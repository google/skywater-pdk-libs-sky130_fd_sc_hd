* File: sky130_fd_sc_hd__inv_8.pxi.spice
* Created: Tue Sep  1 19:10:19 2020
* 
x_PM_SKY130_FD_SC_HD__INV_8%A N_A_c_66_n N_A_M1000_g N_A_M1002_g N_A_c_67_n
+ N_A_M1001_g N_A_M1004_g N_A_c_68_n N_A_M1003_g N_A_M1008_g N_A_c_69_n
+ N_A_M1005_g N_A_M1009_g N_A_c_70_n N_A_M1006_g N_A_M1010_g N_A_c_71_n
+ N_A_M1007_g N_A_M1011_g N_A_c_72_n N_A_M1012_g N_A_M1013_g N_A_c_73_n
+ N_A_M1014_g N_A_M1015_g A A A A A A N_A_c_74_n PM_SKY130_FD_SC_HD__INV_8%A
x_PM_SKY130_FD_SC_HD__INV_8%VPWR N_VPWR_M1002_s N_VPWR_M1004_s N_VPWR_M1009_s
+ N_VPWR_M1011_s N_VPWR_M1015_s N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n
+ N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n VPWR
+ N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_226_n PM_SKY130_FD_SC_HD__INV_8%VPWR
x_PM_SKY130_FD_SC_HD__INV_8%Y N_Y_M1000_d N_Y_M1003_d N_Y_M1006_d N_Y_M1012_d
+ N_Y_M1002_d N_Y_M1008_d N_Y_M1010_d N_Y_M1013_d N_Y_c_290_n N_Y_c_291_n
+ N_Y_c_307_n N_Y_c_302_n N_Y_c_308_n N_Y_c_311_n N_Y_c_292_n N_Y_c_318_n
+ N_Y_c_322_n N_Y_c_326_n N_Y_c_293_n N_Y_c_334_n N_Y_c_338_n N_Y_c_342_n
+ N_Y_c_294_n N_Y_c_350_n N_Y_c_354_n N_Y_c_357_n N_Y_c_295_n N_Y_c_303_n
+ N_Y_c_296_n N_Y_c_368_n N_Y_c_297_n N_Y_c_376_n N_Y_c_298_n N_Y_c_384_n
+ N_Y_c_299_n N_Y_c_392_n Y Y PM_SKY130_FD_SC_HD__INV_8%Y
x_PM_SKY130_FD_SC_HD__INV_8%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1005_s
+ N_VGND_M1007_s N_VGND_M1014_s N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n
+ N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n
+ N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n VGND
+ N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n PM_SKY130_FD_SC_HD__INV_8%VGND
cc_1 VNB N_A_c_66_n 0.0191953f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.995
cc_2 VNB N_A_c_67_n 0.0157981f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_3 VNB N_A_c_68_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=0.995
cc_4 VNB N_A_c_69_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=0.995
cc_5 VNB N_A_c_70_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=0.995
cc_6 VNB N_A_c_71_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.995
cc_7 VNB N_A_c_72_n 0.0157972f $X=-0.19 $Y=-0.24 $X2=3.155 $Y2=0.995
cc_8 VNB N_A_c_73_n 0.0191608f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=0.995
cc_9 VNB N_A_c_74_n 0.13208f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=1.16
cc_10 VNB N_VPWR_c_226_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_290_n 0.00180816f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=1.325
cc_12 VNB N_Y_c_291_n 0.0121685f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=1.985
cc_13 VNB N_Y_c_292_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.56
cc_14 VNB N_Y_c_293_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_Y_c_294_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.105
cc_16 VNB N_Y_c_295_n 0.0115362f $X=-0.19 $Y=-0.24 $X2=0.845 $Y2=1.16
cc_17 VNB N_Y_c_296_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=3.155 $Y2=1.16
cc_18 VNB N_Y_c_297_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=3.365 $Y2=1.16
cc_19 VNB N_Y_c_298_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.845 $Y2=1.2
cc_20 VNB N_Y_c_299_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB Y 0.0229772f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=1.2
cc_22 VNB Y 0.0219886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_464_n 0.0145621f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=0.56
cc_24 VNB N_VGND_c_465_n 0.0166337f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=1.325
cc_25 VNB N_VGND_c_466_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=0.995
cc_26 VNB N_VGND_c_467_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=0.56
cc_27 VNB N_VGND_c_468_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_469_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=1.325
cc_29 VNB N_VGND_c_470_n 0.0121521f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=1.985
cc_30 VNB N_VGND_c_471_n 0.0181978f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.995
cc_31 VNB N_VGND_c_472_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=0.56
cc_32 VNB N_VGND_c_473_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=1.325
cc_33 VNB N_VGND_c_474_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=2.735 $Y2=1.985
cc_34 VNB N_VGND_c_475_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_476_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.575 $Y2=1.325
cc_36 VNB N_VGND_c_477_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.105
cc_37 VNB N_VGND_c_478_n 0.219879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_A_M1002_g 0.0219695f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.985
cc_39 VPB N_A_M1004_g 0.0185026f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.985
cc_40 VPB N_A_M1008_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=1.985
cc_41 VPB N_A_M1009_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=1.985
cc_42 VPB N_A_M1010_g 0.0185065f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.985
cc_43 VPB N_A_M1011_g 0.0185065f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=1.985
cc_44 VPB N_A_M1013_g 0.0185011f $X=-0.19 $Y=1.305 $X2=3.155 $Y2=1.985
cc_45 VPB N_A_M1015_g 0.0219078f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=1.985
cc_46 VPB N_A_c_74_n 0.0227951f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=1.16
cc_47 VPB N_VPWR_c_227_n 0.0152107f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=0.56
cc_48 VPB N_VPWR_c_228_n 0.0294647f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=1.325
cc_49 VPB N_VPWR_c_229_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=0.995
cc_50 VPB N_VPWR_c_230_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=0.56
cc_51 VPB N_VPWR_c_231_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_232_n 0.00358901f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.325
cc_53 VPB N_VPWR_c_233_n 0.012408f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.985
cc_54 VPB N_VPWR_c_234_n 0.0316876f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=0.995
cc_55 VPB N_VPWR_c_235_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=0.56
cc_56 VPB N_VPWR_c_236_n 0.00323736f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=1.325
cc_57 VPB N_VPWR_c_237_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.735 $Y2=1.985
cc_58 VPB N_VPWR_c_238_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_239_n 0.017949f $X=-0.19 $Y=1.305 $X2=3.575 $Y2=1.325
cc_60 VPB N_VPWR_c_240_n 0.00323736f $X=-0.19 $Y=1.305 $X2=2.905 $Y2=1.105
cc_61 VPB N_VPWR_c_226_n 0.0516153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_Y_c_302_n 0.0156116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_Y_c_303_n 0.0109095f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=1.16
cc_64 VPB Y 0.0108936f $X=-0.19 $Y=1.305 $X2=2.53 $Y2=1.2
cc_65 VPB Y 0.0102978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 N_A_M1002_g N_VPWR_c_228_n 0.00321527f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_M1004_g N_VPWR_c_229_n 0.00146448f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_M1008_g N_VPWR_c_229_n 0.00146448f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A_M1008_g N_VPWR_c_230_n 0.00541359f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A_M1009_g N_VPWR_c_230_n 0.00541359f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_M1009_g N_VPWR_c_231_n 0.00146448f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_M1010_g N_VPWR_c_231_n 0.00146448f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A_M1011_g N_VPWR_c_232_n 0.00146448f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_M1013_g N_VPWR_c_232_n 0.00146448f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1015_g N_VPWR_c_234_n 0.0032367f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1002_g N_VPWR_c_235_n 0.00541359f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_M1004_g N_VPWR_c_235_n 0.00541359f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1010_g N_VPWR_c_237_n 0.00541359f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_M1011_g N_VPWR_c_237_n 0.00541359f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_M1013_g N_VPWR_c_239_n 0.00541359f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_M1015_g N_VPWR_c_239_n 0.00541359f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_VPWR_c_226_n 0.0105807f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_M1004_g N_VPWR_c_226_n 0.00950154f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1008_g N_VPWR_c_226_n 0.00950154f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1009_g N_VPWR_c_226_n 0.00950154f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1010_g N_VPWR_c_226_n 0.00950154f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1011_g N_VPWR_c_226_n 0.00950154f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1013_g N_VPWR_c_226_n 0.00950154f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_M1015_g N_VPWR_c_226_n 0.0105352f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_c_66_n N_Y_c_290_n 0.0124304f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_Y_c_307_n 0.0140381f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_c_66_n N_Y_c_308_n 0.0108215f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_67_n N_Y_c_308_n 0.00620543f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_c_68_n N_Y_c_308_n 5.19281e-19 $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_M1002_g N_Y_c_311_n 0.0145598f $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_M1004_g N_Y_c_311_n 0.00975139f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_M1008_g N_Y_c_311_n 6.1949e-19 $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_c_67_n N_Y_c_292_n 0.00890471f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_c_68_n N_Y_c_292_n 0.00890471f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_100 A N_Y_c_292_n 0.0368812f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A_c_74_n N_Y_c_292_n 0.00222429f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_M1004_g N_Y_c_318_n 0.0107189f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_M1008_g N_Y_c_318_n 0.0107189f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_104 A N_Y_c_318_n 0.0320704f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_105 N_A_c_74_n N_Y_c_318_n 0.00201785f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_c_67_n N_Y_c_322_n 5.19281e-19 $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_c_68_n N_Y_c_322_n 0.00620543f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_69_n N_Y_c_322_n 0.00620543f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_c_70_n N_Y_c_322_n 5.19281e-19 $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_M1004_g N_Y_c_326_n 6.1949e-19 $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_M1008_g N_Y_c_326_n 0.00975139f $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_M1009_g N_Y_c_326_n 0.00975139f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_M1010_g N_Y_c_326_n 6.1949e-19 $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_c_69_n N_Y_c_293_n 0.00890471f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_c_70_n N_Y_c_293_n 0.00890471f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_116 A N_Y_c_293_n 0.0368812f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A_c_74_n N_Y_c_293_n 0.00222429f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_M1009_g N_Y_c_334_n 0.0107189f $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_M1010_g N_Y_c_334_n 0.0107189f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_120 A N_Y_c_334_n 0.0320704f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A_c_74_n N_Y_c_334_n 0.00201785f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_c_69_n N_Y_c_338_n 5.19281e-19 $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_70_n N_Y_c_338_n 0.00620543f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_c_71_n N_Y_c_338_n 0.00620543f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_72_n N_Y_c_338_n 5.19281e-19 $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_M1009_g N_Y_c_342_n 6.1949e-19 $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A_M1010_g N_Y_c_342_n 0.00975139f $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_M1011_g N_Y_c_342_n 0.00975139f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_M1013_g N_Y_c_342_n 6.1949e-19 $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_c_71_n N_Y_c_294_n 0.00890471f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_72_n N_Y_c_294_n 0.00890471f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_132 A N_Y_c_294_n 0.0368812f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_133 N_A_c_74_n N_Y_c_294_n 0.00222429f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_M1011_g N_Y_c_350_n 0.0107189f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1013_g N_Y_c_350_n 0.0107189f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_136 A N_Y_c_350_n 0.0320704f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A_c_74_n N_Y_c_350_n 0.00201785f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_71_n N_Y_c_354_n 5.19281e-19 $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_c_72_n N_Y_c_354_n 0.00620543f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_73_n N_Y_c_354_n 0.0108215f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_M1011_g N_Y_c_357_n 6.1949e-19 $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1013_g N_Y_c_357_n 0.00975139f $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1015_g N_Y_c_357_n 0.0145598f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_c_73_n N_Y_c_295_n 0.0121852f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_145 A N_Y_c_295_n 3.17698e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A_M1015_g N_Y_c_303_n 0.0138077f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_147 A N_Y_c_303_n 3.15358e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A_c_66_n N_Y_c_296_n 0.00116017f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_67_n N_Y_c_296_n 0.00116017f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_150 A N_Y_c_296_n 0.0269421f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A_c_74_n N_Y_c_296_n 0.00230339f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_M1002_g N_Y_c_368_n 8.84614e-19 $X=0.635 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_M1004_g N_Y_c_368_n 8.84614e-19 $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_154 A N_Y_c_368_n 0.0213676f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_c_74_n N_Y_c_368_n 0.00209661f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_68_n N_Y_c_297_n 0.00116017f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_69_n N_Y_c_297_n 0.00116017f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_158 A N_Y_c_297_n 0.0269421f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A_c_74_n N_Y_c_297_n 0.00230339f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_M1008_g N_Y_c_376_n 8.84614e-19 $X=1.475 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_M1009_g N_Y_c_376_n 8.84614e-19 $X=1.895 $Y=1.985 $X2=0 $Y2=0
cc_162 A N_Y_c_376_n 0.0213676f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A_c_74_n N_Y_c_376_n 0.00209661f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_c_70_n N_Y_c_298_n 0.00116017f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_71_n N_Y_c_298_n 0.00116017f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_166 A N_Y_c_298_n 0.0269421f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A_c_74_n N_Y_c_298_n 0.00230339f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_M1010_g N_Y_c_384_n 8.84614e-19 $X=2.315 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_M1011_g N_Y_c_384_n 8.84614e-19 $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_170 A N_Y_c_384_n 0.0213676f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A_c_74_n N_Y_c_384_n 0.00209661f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_c_72_n N_Y_c_299_n 0.00116017f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_73_n N_Y_c_299_n 0.00116017f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_174 A N_Y_c_299_n 0.0269421f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_175 N_A_c_74_n N_Y_c_299_n 0.00230339f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_M1013_g N_Y_c_392_n 8.84614e-19 $X=3.155 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_M1015_g N_Y_c_392_n 8.84614e-19 $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_178 A N_Y_c_392_n 0.0213676f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A_c_74_n N_Y_c_392_n 0.00209661f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_c_66_n Y 0.0211079f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_181 A Y 0.015622f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A_c_73_n Y 0.0218736f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_183 A Y 0.0183588f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A_c_66_n N_VGND_c_465_n 0.00321527f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_67_n N_VGND_c_466_n 0.00146448f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_68_n N_VGND_c_466_n 0.00146448f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_68_n N_VGND_c_467_n 0.00422241f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_69_n N_VGND_c_467_n 0.00422241f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_69_n N_VGND_c_468_n 0.00146448f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_70_n N_VGND_c_468_n 0.00146448f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_71_n N_VGND_c_469_n 0.00146448f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_72_n N_VGND_c_469_n 0.00146448f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_73_n N_VGND_c_471_n 0.0032389f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_66_n N_VGND_c_472_n 0.00422241f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_67_n N_VGND_c_472_n 0.00422241f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_70_n N_VGND_c_474_n 0.00422241f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_71_n N_VGND_c_474_n 0.00422241f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_c_72_n N_VGND_c_476_n 0.00422241f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_c_73_n N_VGND_c_476_n 0.00422241f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_66_n N_VGND_c_478_n 0.00677573f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_67_n N_VGND_c_478_n 0.00569656f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_68_n N_VGND_c_478_n 0.00569656f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_69_n N_VGND_c_478_n 0.00569656f $X=1.895 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_70_n N_VGND_c_478_n 0.00569656f $X=2.315 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_c_71_n N_VGND_c_478_n 0.00569656f $X=2.735 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_c_72_n N_VGND_c_478_n 0.00569656f $X=3.155 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_c_73_n N_VGND_c_478_n 0.00673022f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_208 N_VPWR_c_226_n N_Y_M1002_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_209 N_VPWR_c_226_n N_Y_M1008_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_210 N_VPWR_c_226_n N_Y_M1010_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_211 N_VPWR_c_226_n N_Y_M1013_d 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_212 N_VPWR_M1002_s N_Y_c_307_n 0.00209819f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_213 N_VPWR_c_228_n N_Y_c_307_n 0.0059027f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_214 N_VPWR_M1002_s N_Y_c_302_n 0.00218031f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_215 N_VPWR_c_228_n N_Y_c_302_n 0.0157986f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_216 N_VPWR_c_235_n N_Y_c_311_n 0.0189039f $X=1.18 $Y=2.72 $X2=0 $Y2=0
cc_217 N_VPWR_c_226_n N_Y_c_311_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_M1004_s N_Y_c_318_n 0.00311483f $X=1.13 $Y=1.485 $X2=0 $Y2=0
cc_219 N_VPWR_c_229_n N_Y_c_318_n 0.0126919f $X=1.265 $Y=2 $X2=0 $Y2=0
cc_220 N_VPWR_c_230_n N_Y_c_326_n 0.0189039f $X=2.02 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_c_226_n N_Y_c_326_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_M1009_s N_Y_c_334_n 0.00311483f $X=1.97 $Y=1.485 $X2=0 $Y2=0
cc_223 N_VPWR_c_231_n N_Y_c_334_n 0.0126919f $X=2.105 $Y=2 $X2=0 $Y2=0
cc_224 N_VPWR_c_237_n N_Y_c_342_n 0.0189039f $X=2.86 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_226_n N_Y_c_342_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_M1011_s N_Y_c_350_n 0.00311483f $X=2.81 $Y=1.485 $X2=0 $Y2=0
cc_227 N_VPWR_c_232_n N_Y_c_350_n 0.0126919f $X=2.945 $Y=2 $X2=0 $Y2=0
cc_228 N_VPWR_c_239_n N_Y_c_357_n 0.0189039f $X=3.7 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_226_n N_Y_c_357_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_M1015_s N_Y_c_303_n 0.00346511f $X=3.65 $Y=1.485 $X2=0 $Y2=0
cc_231 N_VPWR_c_234_n N_Y_c_303_n 0.0263139f $X=3.785 $Y=2 $X2=0 $Y2=0
cc_232 N_Y_c_290_n N_VGND_M1000_s 7.48374e-19 $X=0.68 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_233 N_Y_c_291_n N_VGND_M1000_s 0.00215453f $X=0.43 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_234 N_Y_c_292_n N_VGND_M1001_s 0.00162148f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_235 N_Y_c_293_n N_VGND_M1005_s 0.00162148f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_236 N_Y_c_294_n N_VGND_M1007_s 0.00162148f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_237 N_Y_c_295_n N_VGND_M1014_s 0.00292039f $X=3.735 $Y=0.81 $X2=0 $Y2=0
cc_238 N_Y_c_291_n N_VGND_c_464_n 0.00295616f $X=0.43 $Y=0.81 $X2=0 $Y2=0
cc_239 N_Y_c_290_n N_VGND_c_465_n 0.00570628f $X=0.68 $Y=0.81 $X2=0 $Y2=0
cc_240 N_Y_c_291_n N_VGND_c_465_n 0.0151569f $X=0.43 $Y=0.81 $X2=0 $Y2=0
cc_241 N_Y_c_292_n N_VGND_c_466_n 0.0122675f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_242 N_Y_c_292_n N_VGND_c_467_n 0.00203746f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_243 N_Y_c_322_n N_VGND_c_467_n 0.0188551f $X=1.685 $Y=0.38 $X2=0 $Y2=0
cc_244 N_Y_c_293_n N_VGND_c_467_n 0.00203746f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_245 N_Y_c_293_n N_VGND_c_468_n 0.0122675f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_246 N_Y_c_294_n N_VGND_c_469_n 0.0122675f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_247 N_Y_c_295_n N_VGND_c_470_n 8.69458e-19 $X=3.735 $Y=0.81 $X2=0 $Y2=0
cc_248 N_Y_c_295_n N_VGND_c_471_n 0.0256874f $X=3.735 $Y=0.81 $X2=0 $Y2=0
cc_249 N_Y_c_290_n N_VGND_c_472_n 0.00203746f $X=0.68 $Y=0.81 $X2=0 $Y2=0
cc_250 N_Y_c_308_n N_VGND_c_472_n 0.0188551f $X=0.845 $Y=0.38 $X2=0 $Y2=0
cc_251 N_Y_c_292_n N_VGND_c_472_n 0.00203746f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_252 N_Y_c_293_n N_VGND_c_474_n 0.00203746f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_253 N_Y_c_338_n N_VGND_c_474_n 0.0188551f $X=2.525 $Y=0.38 $X2=0 $Y2=0
cc_254 N_Y_c_294_n N_VGND_c_474_n 0.00203746f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_255 N_Y_c_294_n N_VGND_c_476_n 0.00203746f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_256 N_Y_c_354_n N_VGND_c_476_n 0.0188551f $X=3.365 $Y=0.38 $X2=0 $Y2=0
cc_257 N_Y_c_295_n N_VGND_c_476_n 0.00203746f $X=3.735 $Y=0.81 $X2=0 $Y2=0
cc_258 N_Y_M1000_d N_VGND_c_478_n 0.00215201f $X=0.71 $Y=0.235 $X2=0 $Y2=0
cc_259 N_Y_M1003_d N_VGND_c_478_n 0.00215201f $X=1.55 $Y=0.235 $X2=0 $Y2=0
cc_260 N_Y_M1006_d N_VGND_c_478_n 0.00215201f $X=2.39 $Y=0.235 $X2=0 $Y2=0
cc_261 N_Y_M1012_d N_VGND_c_478_n 0.00215201f $X=3.23 $Y=0.235 $X2=0 $Y2=0
cc_262 N_Y_c_290_n N_VGND_c_478_n 0.00420836f $X=0.68 $Y=0.81 $X2=0 $Y2=0
cc_263 N_Y_c_291_n N_VGND_c_478_n 0.00562823f $X=0.43 $Y=0.81 $X2=0 $Y2=0
cc_264 N_Y_c_308_n N_VGND_c_478_n 0.0122069f $X=0.845 $Y=0.38 $X2=0 $Y2=0
cc_265 N_Y_c_292_n N_VGND_c_478_n 0.00845923f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_266 N_Y_c_322_n N_VGND_c_478_n 0.0122069f $X=1.685 $Y=0.38 $X2=0 $Y2=0
cc_267 N_Y_c_293_n N_VGND_c_478_n 0.00845923f $X=2.36 $Y=0.81 $X2=0 $Y2=0
cc_268 N_Y_c_338_n N_VGND_c_478_n 0.0122069f $X=2.525 $Y=0.38 $X2=0 $Y2=0
cc_269 N_Y_c_294_n N_VGND_c_478_n 0.00845923f $X=3.2 $Y=0.81 $X2=0 $Y2=0
cc_270 N_Y_c_354_n N_VGND_c_478_n 0.0122069f $X=3.365 $Y=0.38 $X2=0 $Y2=0
cc_271 N_Y_c_295_n N_VGND_c_478_n 0.00667558f $X=3.735 $Y=0.81 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__inv_2.pex.spice
* Created: Tue Sep  1 19:10:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__INV_2%A 1 3 6 8 10 13 15 22
r36 21 22 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.48 $Y=1.16 $X2=0.9
+ $Y2=1.16
r37 18 21 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.27 $Y=1.16
+ $X2=0.48 $Y2=1.16
r38 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r39 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=1.325
+ $X2=0.9 $Y2=1.16
r40 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.9 $Y=1.325 $X2=0.9
+ $Y2=1.985
r41 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=0.995 $X2=0.9
+ $Y2=1.16
r42 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.9 $Y=0.995 $X2=0.9
+ $Y2=0.56
r43 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r44 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.325 $X2=0.48
+ $Y2=1.985
r45 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995 $X2=0.48
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__INV_2%VPWR 1 2 7 9 13 15 19 21 31
r19 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r20 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r21 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r22 22 27 3.83185 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=2.72
+ $X2=0.177 $Y2=2.72
r23 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=2.72
+ $X2=0.69 $Y2=2.72
r24 21 30 3.66464 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=1.202 $Y2=2.72
r25 21 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=0.69 $Y2=2.72
r26 19 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r27 19 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r28 15 18 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=1.13 $Y=1.66
+ $X2=1.13 $Y2=2.34
r29 13 30 3.25055 $w=2.1e-07 $l=1.15521e-07 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.202 $Y2=2.72
r30 13 18 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.13 $Y2=2.34
r31 9 12 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=1.66 $X2=0.24
+ $Y2=2.34
r32 7 27 3.18603 $w=2.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.177 $Y2=2.72
r33 7 12 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.34
r34 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.485 $X2=1.11 $Y2=2.34
r35 2 15 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.485 $X2=1.11 $Y2=1.66
r36 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=2.34
r37 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__INV_2%Y 1 2 9 13 17 18 19 33 36
r22 36 37 2.27618 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.69 $Y=1.53
+ $X2=0.69 $Y2=1.485
r23 33 34 1.92695 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.69 $Y=0.85
+ $X2=0.69 $Y2=0.885
r24 19 36 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=0.69 $Y=1.55 $X2=0.69
+ $Y2=1.53
r25 19 37 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=0.73 $Y=1.465
+ $X2=0.73 $Y2=1.485
r26 18 19 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.73 $Y=1.19
+ $X2=0.73 $Y2=1.465
r27 17 33 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.69 $Y=0.825
+ $X2=0.69 $Y2=0.85
r28 17 18 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.73 $Y=0.91
+ $X2=0.73 $Y2=1.19
r29 17 34 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=0.73 $Y=0.91
+ $X2=0.73 $Y2=0.885
r30 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=1.66
+ $X2=0.69 $Y2=2.34
r31 11 19 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.69 $Y=1.65 $X2=0.69
+ $Y2=1.55
r32 11 13 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.69 $Y=1.65 $X2=0.69
+ $Y2=1.66
r33 7 17 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.69 $Y=0.72
+ $X2=0.69 $Y2=0.825
r34 7 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.69 $Y=0.72 $X2=0.69
+ $Y2=0.38
r35 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.485 $X2=0.69 $Y2=2.34
r36 2 13 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.485 $X2=0.69 $Y2=1.66
r37 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__INV_2%VGND 1 2 7 9 11 13 15 17 27
r20 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r21 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r22 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r23 18 23 3.83185 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r24 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.69
+ $Y2=0
r25 17 26 3.66464 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.202
+ $Y2=0
r26 17 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.69
+ $Y2=0
r27 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r28 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r29 11 26 3.25055 $w=2.1e-07 $l=1.15521e-07 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.202 $Y2=0
r30 11 13 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0.38
r31 7 23 3.18603 $w=2.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.177 $Y2=0
r32 7 9 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r33 2 13 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.975
+ $Y=0.235 $X2=1.11 $Y2=0.38
r34 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends


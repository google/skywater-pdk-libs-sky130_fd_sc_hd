* File: sky130_fd_sc_hd__sdfbbn_1.spice
* Created: Thu Aug 27 14:45:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdfbbn_1.pex.spice"
.subckt sky130_fd_sc_hd__sdfbbn_1  VNB VPB CLK_N SCD SCE D SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* SCE	SCE
* SCD	SCD
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1045 N_VGND_M1045_d N_CLK_N_M1045_g N_A_27_47#_M1045_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_A_193_47#_M1026_d N_A_27_47#_M1026_g N_VGND_M1045_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_381_47# N_SCD_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1013 N_A_453_47#_M1013_d N_SCE_M1013_g A_381_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1239 AS=0.0441 PD=1.43 PS=0.63 NRD=8.568 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1041 N_VGND_M1041_d N_SCE_M1041_g N_A_423_315#_M1041_s VNB NSHORT L=0.15
+ W=0.42 AD=0.05985 AS=0.1092 PD=0.705 PS=1.36 NRD=2.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1042 A_735_47# N_A_423_315#_M1042_g N_VGND_M1041_d VNB NSHORT L=0.15 W=0.42
+ AD=0.05985 AS=0.05985 PD=0.705 PS=0.705 NRD=24.996 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1027 N_A_453_47#_M1027_d N_D_M1027_g A_735_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.05985 PD=0.802308 PS=0.705 NRD=0 NRS=24.996 M=1 R=2.8
+ SA=75001.1 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1014 N_A_917_47#_M1014_d N_A_193_47#_M1014_g N_A_453_47#_M1027_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0747 AS=0.0609231 PD=0.775 PS=0.687692 NRD=0 NRS=16.656 M=1
+ R=2.4 SA=75001.5 SB=75002.7 A=0.054 P=1.02 MULT=1
MM1044 A_1030_47# N_A_27_47#_M1044_g N_A_917_47#_M1014_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0677077 AS=0.0747 PD=0.72 PS=0.775 NRD=44.352 NRS=46.656 M=1 R=2.4
+ SA=75002.1 SB=75002.2 A=0.054 P=1.02 MULT=1
MM1009 N_VGND_M1009_d N_A_1102_21#_M1009_g A_1030_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.08295 AS=0.0789923 PD=0.815 PS=0.84 NRD=34.284 NRS=38.016 M=1 R=2.8
+ SA=75002.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_1241_47#_M1004_d N_SET_B_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0808698 AS=0.08295 PD=0.788491 PS=0.815 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75002.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1040 N_A_1102_21#_M1040_d N_A_917_47#_M1040_g N_A_1241_47#_M1004_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0864 AS=0.12323 PD=0.91 PS=1.20151 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75002.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1032 N_A_1241_47#_M1032_d N_A_1396_21#_M1032_g N_A_1102_21#_M1040_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 A_1614_47# N_A_1102_21#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.64
+ AD=0.12544 AS=0.1664 PD=1.2672 PS=1.8 NRD=26.436 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1010 N_A_1714_47#_M1010_d N_A_27_47#_M1010_g A_1614_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0702 AS=0.07056 PD=0.75 PS=0.7128 NRD=23.328 NRS=46.992 M=1 R=2.4
+ SA=75000.7 SB=75002.6 A=0.054 P=1.02 MULT=1
MM1024 A_1822_47# N_A_193_47#_M1024_g N_A_1714_47#_M1010_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0702 PD=0.687692 PS=0.75 NRD=38.076 NRS=13.332 M=1
+ R=2.4 SA=75001.2 SB=75002.1 A=0.054 P=1.02 MULT=1
MM1003 N_VGND_M1003_d N_A_1887_21#_M1003_g A_1822_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.05985 AS=0.0710769 PD=0.705 PS=0.802308 NRD=2.856 NRS=32.628 M=1 R=2.8
+ SA=75001.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_2004_47#_M1006_d N_SET_B_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.094183 AS=0.05985 PD=0.851887 PS=0.705 NRD=24.276 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_1887_21#_M1020_d N_A_1714_47#_M1020_g N_A_2004_47#_M1006_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0864 AS=0.143517 PD=0.91 PS=1.29811 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75001.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1029 N_A_2004_47#_M1029_d N_A_1396_21#_M1029_g N_A_1887_21#_M1020_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_RESET_B_M1015_g N_A_1396_21#_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_Q_N_M1001_d N_A_1887_21#_M1001_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.121799 PD=1.82 PS=1.19673 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1046 N_VGND_M1046_d N_A_1887_21#_M1046_g N_A_2596_47#_M1046_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_Q_M1018_d N_A_2596_47#_M1018_g N_VGND_M1046_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1025 N_VPWR_M1025_d N_CLK_N_M1025_g N_A_27_47#_M1025_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1033 A_381_363# N_SCD_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1664 PD=0.85 PS=1.8 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.5 A=0.096 P=1.58 MULT=1
MM1038 N_A_453_47#_M1038_d N_A_423_315#_M1038_g A_381_363# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0672 PD=1.8 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_SCE_M1034_g N_A_423_315#_M1034_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75007.8 A=0.063 P=1.14 MULT=1
MM1021 A_752_413# N_SCE_M1021_g N_VPWR_M1034_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=37.5088 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75007.4 A=0.063 P=1.14 MULT=1
MM1017 N_A_453_47#_M1017_d N_D_M1017_g A_752_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07035 AS=0.0567 PD=0.755 PS=0.69 NRD=0 NRS=37.5088 M=1 R=2.8 SA=75001
+ SB=75007 A=0.063 P=1.14 MULT=1
MM1039 N_A_917_47#_M1039_d N_A_27_47#_M1039_g N_A_453_47#_M1017_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.07035 PD=0.69 PS=0.755 NRD=0 NRS=28.1316 M=1
+ R=2.8 SA=75001.5 SB=75006.5 A=0.063 P=1.14 MULT=1
MM1011 A_1017_413# N_A_193_47#_M1011_g N_A_917_47#_M1039_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0945 AS=0.0567 PD=0.87 PS=0.69 NRD=79.7259 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75006.1 A=0.063 P=1.14 MULT=1
MM1035 N_VPWR_M1035_d N_A_1102_21#_M1035_g A_1017_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0945 PD=0.8 PS=0.87 NRD=21.0987 NRS=79.7259 M=1 R=2.8
+ SA=75002.5 SB=75005.5 A=0.063 P=1.14 MULT=1
MM1012 N_A_1102_21#_M1012_d N_SET_B_M1012_g N_VPWR_M1035_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.098 AS=0.0798 PD=0.82 PS=0.8 NRD=53.9386 NRS=25.7873 M=1 R=2.8
+ SA=75003.1 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1036 A_1351_329# N_A_917_47#_M1036_g N_A_1102_21#_M1012_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1134 AS=0.196 PD=1.11 PS=1.64 NRD=18.7544 NRS=0 M=1 R=5.6
+ SA=75001.9 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1030 N_VPWR_M1030_d N_A_1396_21#_M1030_g A_1351_329# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2247 AS=0.1134 PD=1.375 PS=1.11 NRD=5.8509 NRS=18.7544 M=1 R=5.6
+ SA=75002.3 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1047 A_1572_329# N_A_1102_21#_M1047_g N_VPWR_M1030_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2324 AS=0.2247 PD=1.88 PS=1.375 NRD=51.9686 NRS=53.9386 M=1 R=5.6
+ SA=75003 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1031 N_A_1714_47#_M1031_d N_A_193_47#_M1031_g A_1572_329# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.1162 PD=0.69 PS=0.94 NRD=0 NRS=103.957 M=1 R=2.8
+ SA=75005.4 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1019 A_1800_413# N_A_27_47#_M1019_g N_A_1714_47#_M1031_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.0567 PD=0.86 PS=0.69 NRD=77.3816 NRS=0 M=1 R=2.8
+ SA=75005.8 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1043 N_VPWR_M1043_d N_A_1887_21#_M1043_g A_1800_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0924 PD=0.81 PS=0.86 NRD=25.7873 NRS=77.3816 M=1 R=2.8
+ SA=75006.4 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_1887_21#_M1008_d N_SET_B_M1008_g N_VPWR_M1043_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0819 PD=0.78 PS=0.81 NRD=25.7873 NRS=25.7873 M=1 R=2.8
+ SA=75007 SB=75001 A=0.063 P=1.14 MULT=1
MM1023 A_2122_329# N_A_1714_47#_M1023_g N_A_1887_21#_M1008_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.1638 PD=1.05 PS=1.56 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75003.8 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1028 N_VPWR_M1028_d N_A_1396_21#_M1028_g A_2122_329# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2184 AS=0.0882 PD=2.2 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75004.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_RESET_B_M1005_g N_A_1396_21#_M1005_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.120117 AS=0.1664 PD=1.04195 PS=1.8 NRD=40.8381 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1037 N_Q_N_M1037_d N_A_1887_21#_M1037_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.187683 PD=2.52 PS=1.62805 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1022_d N_A_1887_21#_M1022_g N_A_2596_47#_M1022_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=14.6174 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1002 N_Q_M1002_d N_A_2596_47#_M1002_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.181707 PD=2.52 PS=1.61585 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX48_noxref VNB VPB NWDIODE A=23.4972 P=32.49
c_307 VPB 0 2.26019e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__sdfbbn_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o2111ai_2.pex.spice
* Created: Thu Aug 27 14:34:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2111AI_2%D1 1 3 6 8 10 13 15 17 19
c44 8 0 1.49698e-19 $X=0.985 $Y=0.995
r45 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r46 16 17 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.555 $Y=1.16
+ $X2=0.985 $Y2=1.16
r47 15 22 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.48 $Y=1.16
+ $X2=0.26 $Y2=1.16
r48 15 16 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.48 $Y=1.16
+ $X2=0.555 $Y2=1.16
r49 11 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.325
+ $X2=0.985 $Y2=1.16
r50 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.985 $Y=1.325
+ $X2=0.985 $Y2=1.985
r51 8 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=0.995
+ $X2=0.985 $Y2=1.16
r52 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.985 $Y=0.995
+ $X2=0.985 $Y2=0.56
r53 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.325
+ $X2=0.555 $Y2=1.16
r54 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.555 $Y=1.325
+ $X2=0.555 $Y2=1.985
r55 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=1.16
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%C1 3 7 11 15 18 19 20 21 22
c50 18 0 1.52617e-19 $X=1.415 $Y=1.16
c51 3 0 9.02883e-20 $X=1.415 $Y=0.56
r52 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.16 $X2=1.625 $Y2=1.16
r53 21 22 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.61
+ $Y2=1.2
r54 19 26 32.2152 $w=2.7e-07 $l=1.45e-07 $layer=POLY_cond $X=1.77 $Y=1.16
+ $X2=1.625 $Y2=1.16
r55 19 20 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.77 $Y=1.16
+ $X2=1.845 $Y2=1.16
r56 17 26 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.49 $Y=1.16
+ $X2=1.625 $Y2=1.16
r57 17 18 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.49 $Y=1.16
+ $X2=1.415 $Y2=1.16
r58 13 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.845 $Y=1.295
+ $X2=1.845 $Y2=1.16
r59 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.845 $Y=1.295
+ $X2=1.845 $Y2=1.985
r60 9 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.845 $Y=1.025
+ $X2=1.845 $Y2=1.16
r61 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.845 $Y=1.025
+ $X2=1.845 $Y2=0.56
r62 5 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.415 $Y=1.295
+ $X2=1.415 $Y2=1.16
r63 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.415 $Y=1.295
+ $X2=1.415 $Y2=1.985
r64 1 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.415 $Y=1.025
+ $X2=1.415 $Y2=1.16
r65 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.415 $Y=1.025
+ $X2=1.415 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%B1 3 7 11 15 17 18 19 22 23 24
c55 24 0 2.80714e-19 $X=2.99 $Y=1.19
c56 7 0 1.00188e-19 $X=2.705 $Y=1.985
r57 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=1.16 $X2=2.365 $Y2=1.16
r58 24 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.16 $X2=3.02 $Y2=1.16
r59 23 24 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=1.2 $X2=2.99
+ $Y2=1.2
r60 23 29 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=1.2
+ $X2=2.365 $Y2=1.2
r61 22 31 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.185 $Y=1.16
+ $X2=3.02 $Y2=1.16
r62 20 21 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.705 $Y=1.16
+ $X2=2.83 $Y2=1.16
r63 19 28 58.876 $w=2.7e-07 $l=2.65e-07 $layer=POLY_cond $X=2.63 $Y=1.16
+ $X2=2.365 $Y2=1.16
r64 19 20 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.63 $Y=1.16
+ $X2=2.705 $Y2=1.16
r65 18 31 25.55 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=2.905 $Y=1.16
+ $X2=3.02 $Y2=1.16
r66 18 21 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.905 $Y=1.16
+ $X2=2.83 $Y2=1.16
r67 17 28 3.33261 $w=2.7e-07 $l=1.5e-08 $layer=POLY_cond $X=2.35 $Y=1.16
+ $X2=2.365 $Y2=1.16
r68 13 22 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.26 $Y=1.025
+ $X2=3.185 $Y2=1.16
r69 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.26 $Y=1.025
+ $X2=3.26 $Y2=0.56
r70 9 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.83 $Y=1.025
+ $X2=2.83 $Y2=1.16
r71 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.83 $Y=1.025
+ $X2=2.83 $Y2=0.56
r72 5 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.705 $Y=1.295
+ $X2=2.705 $Y2=1.16
r73 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.705 $Y=1.295
+ $X2=2.705 $Y2=1.985
r74 1 17 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.275 $Y=1.295
+ $X2=2.35 $Y2=1.16
r75 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.275 $Y=1.295
+ $X2=2.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%A2 3 7 11 15 18 19 20 21 22 23
c45 23 0 1.00188e-19 $X=4.285 $Y=1.105
c46 20 0 1.45868e-19 $X=4.12 $Y=1.16
c47 18 0 1.49713e-19 $X=3.69 $Y=1.16
c48 7 0 1.31001e-19 $X=3.69 $Y=1.985
r49 22 23 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=1.2 $X2=4.37
+ $Y2=1.2
r50 22 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.915
+ $Y=1.16 $X2=3.915 $Y2=1.16
r51 21 22 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=3.45 $Y=1.2 $X2=3.91
+ $Y2=1.2
r52 19 28 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=3.915 $Y2=1.16
r53 19 20 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=4.12 $Y2=1.16
r54 17 28 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.765 $Y=1.16
+ $X2=3.915 $Y2=1.16
r55 17 18 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.16
+ $X2=3.69 $Y2=1.16
r56 13 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.12 $Y=1.295
+ $X2=4.12 $Y2=1.16
r57 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.12 $Y=1.295
+ $X2=4.12 $Y2=1.985
r58 9 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.12 $Y=1.025
+ $X2=4.12 $Y2=1.16
r59 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.12 $Y=1.025
+ $X2=4.12 $Y2=0.56
r60 5 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.69 $Y=1.295
+ $X2=3.69 $Y2=1.16
r61 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.69 $Y=1.295 $X2=3.69
+ $Y2=1.985
r62 1 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.69 $Y=1.025
+ $X2=3.69 $Y2=1.16
r63 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.69 $Y=1.025
+ $X2=3.69 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%A1 3 7 11 15 18 19 20 21 22
c41 22 0 1.45868e-19 $X=5.29 $Y=1.19
r42 21 22 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=4.8 $Y=1.2 $X2=5.29
+ $Y2=1.2
r43 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=1.16 $X2=4.8 $Y2=1.16
r44 19 26 23.3282 $w=2.7e-07 $l=1.05e-07 $layer=POLY_cond $X=4.905 $Y=1.16
+ $X2=4.8 $Y2=1.16
r45 19 20 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.905 $Y=1.16
+ $X2=4.98 $Y2=1.16
r46 17 26 38.8804 $w=2.7e-07 $l=1.75e-07 $layer=POLY_cond $X=4.625 $Y=1.16
+ $X2=4.8 $Y2=1.16
r47 17 18 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.625 $Y=1.16
+ $X2=4.55 $Y2=1.16
r48 13 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.98 $Y=1.295
+ $X2=4.98 $Y2=1.16
r49 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.98 $Y=1.295
+ $X2=4.98 $Y2=1.985
r50 9 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.98 $Y=1.025
+ $X2=4.98 $Y2=1.16
r51 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.98 $Y=1.025
+ $X2=4.98 $Y2=0.56
r52 5 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.55 $Y=1.295
+ $X2=4.55 $Y2=1.16
r53 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.55 $Y=1.295 $X2=4.55
+ $Y2=1.985
r54 1 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.55 $Y=1.025
+ $X2=4.55 $Y2=1.16
r55 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.55 $Y=1.025
+ $X2=4.55 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%VPWR 1 2 3 4 5 16 18 22 26 30 34 36 38 43
+ 48 53 63 64 70 73 76 79
r84 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r85 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 64 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r89 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r90 61 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.93 $Y=2.72 $X2=4.8
+ $Y2=2.72
r91 61 63 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.93 $Y=2.72
+ $X2=5.29 $Y2=2.72
r92 60 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r93 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r94 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r95 57 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r96 56 59 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r97 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r98 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=2.72
+ $X2=2.92 $Y2=2.72
r99 54 56 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=2.72
+ $X2=3.45 $Y2=2.72
r100 53 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.67 $Y=2.72 $X2=4.8
+ $Y2=2.72
r101 53 59 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.67 $Y=2.72 $X2=4.37
+ $Y2=2.72
r102 52 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r103 52 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r104 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.06 $Y2=2.72
r106 49 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.53 $Y2=2.72
r107 48 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.92 $Y2=2.72
r108 48 51 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.53 $Y2=2.72
r109 47 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 47 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r111 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r112 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r113 44 46 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=2.06 $Y2=2.72
r115 43 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r116 42 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 39 67 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r119 39 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r121 38 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 36 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 32 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.8 $Y=2.635
+ $X2=4.8 $Y2=2.72
r125 32 34 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=4.8 $Y=2.635
+ $X2=4.8 $Y2=2.02
r126 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=2.635
+ $X2=2.92 $Y2=2.72
r127 28 30 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.92 $Y=2.635
+ $X2=2.92 $Y2=2
r128 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=2.635
+ $X2=2.06 $Y2=2.72
r129 24 26 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.06 $Y=2.635
+ $X2=2.06 $Y2=2
r130 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r131 20 22 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r132 16 67 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=2.635
+ $X2=0.212 $Y2=2.72
r133 16 18 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.3 $Y=2.635
+ $X2=0.3 $Y2=1.845
r134 5 34 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=4.625
+ $Y=1.485 $X2=4.765 $Y2=2.02
r135 4 30 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=2.78
+ $Y=1.485 $X2=2.92 $Y2=2
r136 3 26 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.485 $X2=2.06 $Y2=2
r137 2 22 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.485 $X2=1.2 $Y2=2
r138 1 18 300 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_PDIFF $count=2 $X=0.215
+ $Y=1.485 $X2=0.34 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%Y 1 2 3 4 5 16 20 22 26 28 32 34 35 36 37
+ 38 39 40 62 66
c62 62 0 9.02883e-20 $X=0.77 $Y=0.7
c63 36 0 1.52617e-19 $X=0.605 $Y=0.765
r64 66 67 2.47132 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.77 $Y=0.85
+ $X2=0.77 $Y2=0.905
r65 39 40 16.6218 $w=2.58e-07 $l=3.75e-07 $layer=LI1_cond $X=0.735 $Y=1.835
+ $X2=0.735 $Y2=2.21
r66 39 54 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.735 $Y=1.835
+ $X2=0.735 $Y2=1.665
r67 38 49 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=1.58
+ $X2=0.735 $Y2=1.495
r68 38 54 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=1.58
+ $X2=0.735 $Y2=1.665
r69 38 49 1.10812 $w=2.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.735 $Y=1.47
+ $X2=0.735 $Y2=1.495
r70 37 38 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.735 $Y=1.19
+ $X2=0.735 $Y2=1.47
r71 36 66 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.77 $Y=0.835
+ $X2=0.77 $Y2=0.85
r72 36 62 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.77 $Y=0.835
+ $X2=0.77 $Y2=0.7
r73 36 37 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=0.735 $Y=0.92
+ $X2=0.735 $Y2=1.19
r74 36 67 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=0.92
+ $X2=0.735 $Y2=0.905
r75 30 32 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=3.91 $Y=1.665
+ $X2=3.91 $Y2=1.9
r76 29 35 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.575 $Y=1.58 $X2=2.485
+ $Y2=1.58
r77 28 30 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.815 $Y=1.58
+ $X2=3.91 $Y2=1.665
r78 28 29 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.815 $Y=1.58
+ $X2=2.575 $Y2=1.58
r79 24 35 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=1.665
+ $X2=2.485 $Y2=1.58
r80 24 26 11.0909 $w=1.78e-07 $l=1.8e-07 $layer=LI1_cond $X=2.485 $Y=1.665
+ $X2=2.485 $Y2=1.845
r81 23 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=1.58
+ $X2=1.63 $Y2=1.58
r82 22 35 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.395 $Y=1.58 $X2=2.485
+ $Y2=1.58
r83 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.395 $Y=1.58
+ $X2=1.725 $Y2=1.58
r84 18 34 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=1.58
r85 18 20 10.5072 $w=1.88e-07 $l=1.8e-07 $layer=LI1_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=1.845
r86 17 38 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.865 $Y=1.58
+ $X2=0.735 $Y2=1.58
r87 16 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.535 $Y=1.58
+ $X2=1.63 $Y2=1.58
r88 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=1.58
+ $X2=0.865 $Y2=1.58
r89 5 32 600 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_PDIFF $count=1 $X=3.765
+ $Y=1.485 $X2=3.905 $Y2=1.9
r90 4 26 300 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_PDIFF $count=2 $X=2.35
+ $Y=1.485 $X2=2.49 $Y2=1.845
r91 3 20 300 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_PDIFF $count=2 $X=1.49
+ $Y=1.485 $X2=1.63 $Y2=1.845
r92 2 39 300 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=1.485 $X2=0.77 $Y2=1.835
r93 1 62 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.235 $X2=0.77 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%A_664_297# 1 2 3 10 12 14 16 17 18 22
r34 20 22 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.23 $Y=1.685
+ $X2=5.23 $Y2=1.815
r35 19 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.5 $Y=1.6 $X2=4.37
+ $Y2=1.6
r36 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.1 $Y=1.6
+ $X2=5.23 $Y2=1.685
r37 18 19 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.1 $Y=1.6 $X2=4.5
+ $Y2=1.6
r38 17 29 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=4.37 $Y=2.275
+ $X2=4.37 $Y2=2.37
r39 16 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=1.685
+ $X2=4.37 $Y2=1.6
r40 16 17 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=4.37 $Y=1.685
+ $X2=4.37 $Y2=2.275
r41 15 25 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=2.37 $X2=3.44
+ $Y2=2.37
r42 14 29 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=4.24 $Y=2.37 $X2=4.37
+ $Y2=2.37
r43 14 15 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=4.24 $Y=2.37 $X2=3.57
+ $Y2=2.37
r44 10 25 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=3.44 $Y=2.275
+ $X2=3.44 $Y2=2.37
r45 10 12 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.44 $Y=2.275
+ $X2=3.44 $Y2=2
r46 3 22 300 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_PDIFF $count=2 $X=5.055
+ $Y=1.485 $X2=5.195 $Y2=1.815
r47 2 29 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.485 $X2=4.335 $Y2=2.36
r48 2 27 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=4.195
+ $Y=1.485 $X2=4.335 $Y2=1.68
r49 1 25 600 $w=1.7e-07 $l=9.49342e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.485 $X2=3.475 $Y2=2.36
r50 1 12 600 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.485 $X2=3.475 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%A_27_47# 1 2 3 10 12 14 20 21 25
r39 25 27 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.1 $Y=0.705 $X2=2.1
+ $Y2=0.82
r40 20 27 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.925 $Y=0.82 $X2=2.1
+ $Y2=0.82
r41 20 21 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.925 $Y=0.82
+ $X2=1.3 $Y2=0.82
r42 17 21 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=1.207 $Y=0.735
+ $X2=1.3 $Y2=0.82
r43 17 19 6.89435 $w=1.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.207 $Y=0.735
+ $X2=1.207 $Y2=0.62
r44 16 19 10.4914 $w=1.83e-07 $l=1.75e-07 $layer=LI1_cond $X=1.207 $Y=0.445
+ $X2=1.207 $Y2=0.62
r45 15 23 4.12233 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=0.435 $Y=0.352
+ $X2=0.305 $Y2=0.352
r46 14 16 6.81649 $w=1.85e-07 $l=1.31168e-07 $layer=LI1_cond $X=1.115 $Y=0.352
+ $X2=1.207 $Y2=0.445
r47 14 15 40.7666 $w=1.83e-07 $l=6.8e-07 $layer=LI1_cond $X=1.115 $Y=0.352
+ $X2=0.435 $Y2=0.352
r48 10 23 2.94905 $w=2.6e-07 $l=9.3e-08 $layer=LI1_cond $X=0.305 $Y=0.445
+ $X2=0.305 $Y2=0.352
r49 10 12 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.305 $Y=0.445
+ $X2=0.305 $Y2=0.7
r50 3 25 182 $w=1.7e-07 $l=5.48452e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.235 $X2=2.09 $Y2=0.705
r51 2 19 182 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.235 $X2=1.205 $Y2=0.62
r52 1 23 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.34 $Y2=0.36
r53 1 12 182 $w=1.7e-07 $l=5.58167e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.34 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%A_298_47# 1 2 8 12 13
c26 8 0 1.49698e-19 $X=1.775 $Y=0.35
r27 12 13 8.65019 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0.37
+ $X2=2.88 $Y2=0.37
r28 8 10 7.32471 $w=3.08e-07 $l=1.67332e-07 $layer=LI1_cond $X=1.775 $Y=0.35
+ $X2=1.635 $Y2=0.41
r29 8 13 64.5024 $w=1.88e-07 $l=1.105e-06 $layer=LI1_cond $X=1.775 $Y=0.35
+ $X2=2.88 $Y2=0.35
r30 2 12 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.235 $X2=3.045 $Y2=0.36
r31 1 10 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.235 $X2=1.635 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%A_497_47# 1 2 3 4 13 19 21 25 27 29 30 32
r48 28 30 5.22322 $w=1.87e-07 $l=9.5e-08 $layer=LI1_cond $X=4.43 $Y=0.745
+ $X2=4.335 $Y2=0.745
r49 27 32 5.67621 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=5.267 $Y=0.745
+ $X2=5.267 $Y2=0.58
r50 27 28 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=5.1 $Y=0.745 $X2=4.43
+ $Y2=0.745
r51 23 30 1.29491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=4.335 $Y=0.65
+ $X2=4.335 $Y2=0.745
r52 23 25 4.37799 $w=1.88e-07 $l=7.5e-08 $layer=LI1_cond $X=4.335 $Y=0.65
+ $X2=4.335 $Y2=0.575
r53 22 29 5.28167 $w=1.85e-07 $l=9.5e-08 $layer=LI1_cond $X=3.57 $Y=0.747
+ $X2=3.475 $Y2=0.747
r54 21 30 5.22322 $w=1.87e-07 $l=9.59948e-08 $layer=LI1_cond $X=4.24 $Y=0.747
+ $X2=4.335 $Y2=0.745
r55 21 22 40.1671 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=4.24 $Y=0.747
+ $X2=3.57 $Y2=0.747
r56 17 29 1.24671 $w=1.9e-07 $l=9.2e-08 $layer=LI1_cond $X=3.475 $Y=0.655
+ $X2=3.475 $Y2=0.747
r57 17 19 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=3.475 $Y=0.655
+ $X2=3.475 $Y2=0.575
r58 13 29 5.28167 $w=1.85e-07 $l=9.5e-08 $layer=LI1_cond $X=3.38 $Y=0.747
+ $X2=3.475 $Y2=0.747
r59 13 15 45.8624 $w=1.83e-07 $l=7.65e-07 $layer=LI1_cond $X=3.38 $Y=0.747
+ $X2=2.615 $Y2=0.747
r60 4 32 182 $w=1.7e-07 $l=4.33618e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=0.235 $X2=5.255 $Y2=0.58
r61 3 25 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=4.195
+ $Y=0.235 $X2=4.335 $Y2=0.575
r62 2 19 182 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.235 $X2=3.47 $Y2=0.575
r63 1 15 182 $w=1.7e-07 $l=5.66282e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.615 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O2111AI_2%VGND 1 2 9 13 15 17 25 32 33 36 39
r74 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r75 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r76 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r77 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r78 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=4.765
+ $Y2=0
r79 30 32 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=5.29
+ $Y2=0
r80 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r81 29 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r82 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r83 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.905
+ $Y2=0
r84 26 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.37
+ $Y2=0
r85 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.765
+ $Y2=0
r86 25 28 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.37
+ $Y2=0
r87 24 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r88 23 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r89 19 23 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=3.45
+ $Y2=0
r90 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.905
+ $Y2=0
r91 17 23 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.45
+ $Y2=0
r92 15 24 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=3.45
+ $Y2=0
r93 15 19 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r94 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=0.085
+ $X2=4.765 $Y2=0
r95 11 13 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=4.765 $Y=0.085
+ $X2=4.765 $Y2=0.385
r96 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0
r97 7 9 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.905 $Y=0.085 $X2=3.905
+ $Y2=0.385
r98 2 13 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.765 $Y2=0.385
r99 1 9 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.235 $X2=3.905 $Y2=0.385
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__dlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__dlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.435000 2.185000 1.685000 ;
        RECT 1.985000 0.385000 2.185000 1.435000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 0.255000 6.355000 0.595000 ;
        RECT 6.090000 1.495000 6.355000 2.455000 ;
        RECT 6.170000 0.595000 6.355000 1.495000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
      LAYER mcon ;
        RECT 0.145000 1.105000 0.315000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.190000 1.105000 5.510000 1.435000 ;
      LAYER mcon ;
        RECT 5.210000 1.105000 5.380000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085000 1.075000 0.380000 1.120000 ;
        RECT 0.085000 1.120000 5.440000 1.260000 ;
        RECT 0.085000 1.260000 0.380000 1.305000 ;
        RECT 5.150000 1.075000 5.440000 1.120000 ;
        RECT 5.150000 1.260000 5.440000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.260000 0.345000 0.615000 ;
      RECT 0.175000  0.615000 0.780000 0.785000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.785000 0.780000 1.060000 ;
      RECT 0.610000  1.060000 0.840000 1.390000 ;
      RECT 0.610000  1.390000 0.780000 1.795000 ;
      RECT 1.015000  0.260000 1.280000 1.855000 ;
      RECT 1.015000  1.855000 2.590000 2.025000 ;
      RECT 1.015000  2.025000 1.240000 2.465000 ;
      RECT 1.450000  2.195000 1.815000 2.635000 ;
      RECT 1.480000  0.085000 1.810000 0.905000 ;
      RECT 2.390000  0.815000 3.220000 0.985000 ;
      RECT 2.390000  0.985000 2.590000 1.855000 ;
      RECT 2.475000  2.255000 3.225000 2.425000 ;
      RECT 2.790000  0.390000 3.725000 0.560000 ;
      RECT 3.055000  1.155000 4.175000 1.325000 ;
      RECT 3.055000  1.325000 3.225000 2.255000 ;
      RECT 3.395000  2.135000 3.695000 2.635000 ;
      RECT 3.430000  1.535000 4.710000 1.840000 ;
      RECT 3.430000  1.840000 4.130000 1.865000 ;
      RECT 3.555000  0.560000 3.725000 0.995000 ;
      RECT 3.555000  0.995000 4.175000 1.155000 ;
      RECT 3.895000  0.085000 4.145000 0.610000 ;
      RECT 3.910000  1.865000 4.130000 2.435000 ;
      RECT 4.310000  2.010000 4.595000 2.635000 ;
      RECT 4.320000  0.255000 4.580000 0.615000 ;
      RECT 4.345000  0.615000 4.580000 0.995000 ;
      RECT 4.345000  0.995000 4.740000 1.325000 ;
      RECT 4.345000  1.325000 4.710000 1.535000 ;
      RECT 4.840000  0.290000 5.155000 0.620000 ;
      RECT 4.935000  0.620000 5.155000 0.765000 ;
      RECT 4.935000  0.765000 6.000000 0.935000 ;
      RECT 5.005000  1.725000 5.920000 1.895000 ;
      RECT 5.005000  1.895000 5.335000 2.465000 ;
      RECT 5.570000  2.130000 5.920000 2.635000 ;
      RECT 5.670000  0.085000 5.840000 0.545000 ;
      RECT 5.750000  0.935000 6.000000 1.325000 ;
      RECT 5.750000  1.325000 5.920000 1.725000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__dlclkp_1
END LIBRARY

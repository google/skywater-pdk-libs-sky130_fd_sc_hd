* File: sky130_fd_sc_hd__einvp_2.pxi.spice
* Created: Thu Aug 27 14:20:43 2020
* 
x_PM_SKY130_FD_SC_HD__EINVP_2%TE N_TE_M1008_g N_TE_M1004_g N_TE_c_60_n
+ N_TE_c_61_n N_TE_c_62_n N_TE_M1000_g N_TE_c_63_n N_TE_c_64_n N_TE_M1009_g
+ N_TE_c_65_n TE TE PM_SKY130_FD_SC_HD__EINVP_2%TE
x_PM_SKY130_FD_SC_HD__EINVP_2%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1004_s
+ N_A_27_47#_c_110_n N_A_27_47#_M1001_g N_A_27_47#_c_111_n N_A_27_47#_c_112_n
+ N_A_27_47#_c_113_n N_A_27_47#_M1003_g N_A_27_47#_c_114_n N_A_27_47#_c_106_n
+ N_A_27_47#_c_115_n N_A_27_47#_c_116_n N_A_27_47#_c_107_n N_A_27_47#_c_108_n
+ N_A_27_47#_c_109_n PM_SKY130_FD_SC_HD__EINVP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVP_2%A N_A_c_173_n N_A_M1006_g N_A_M1002_g N_A_c_174_n
+ N_A_M1007_g N_A_M1005_g A A A N_A_c_176_n PM_SKY130_FD_SC_HD__EINVP_2%A
x_PM_SKY130_FD_SC_HD__EINVP_2%VPWR N_VPWR_M1004_d N_VPWR_M1001_s N_VPWR_c_213_n
+ N_VPWR_c_214_n VPWR N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n
+ N_VPWR_c_212_n N_VPWR_c_219_n N_VPWR_c_220_n PM_SKY130_FD_SC_HD__EINVP_2%VPWR
x_PM_SKY130_FD_SC_HD__EINVP_2%A_215_309# N_A_215_309#_M1001_d
+ N_A_215_309#_M1003_d N_A_215_309#_M1005_d N_A_215_309#_c_257_n
+ N_A_215_309#_c_265_n N_A_215_309#_c_258_n N_A_215_309#_c_271_n
+ N_A_215_309#_c_259_n N_A_215_309#_c_290_n N_A_215_309#_c_260_n
+ PM_SKY130_FD_SC_HD__EINVP_2%A_215_309#
x_PM_SKY130_FD_SC_HD__EINVP_2%Z N_Z_M1006_s N_Z_M1002_s Z Z Z Z N_Z_c_297_n
+ PM_SKY130_FD_SC_HD__EINVP_2%Z
x_PM_SKY130_FD_SC_HD__EINVP_2%VGND N_VGND_M1008_d N_VGND_M1009_d N_VGND_c_315_n
+ N_VGND_c_316_n VGND N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n
+ N_VGND_c_320_n N_VGND_c_321_n N_VGND_c_322_n PM_SKY130_FD_SC_HD__EINVP_2%VGND
x_PM_SKY130_FD_SC_HD__EINVP_2%A_204_47# N_A_204_47#_M1000_s N_A_204_47#_M1006_d
+ N_A_204_47#_M1007_d N_A_204_47#_c_385_n N_A_204_47#_c_364_n
+ N_A_204_47#_c_369_n N_A_204_47#_c_365_n N_A_204_47#_c_366_n
+ N_A_204_47#_c_367_n PM_SKY130_FD_SC_HD__EINVP_2%A_204_47#
cc_1 VNB N_TE_M1008_g 0.033909f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_TE_c_60_n 0.0185273f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.035
cc_3 VNB N_TE_c_61_n 0.039083f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.035
cc_4 VNB N_TE_c_62_n 0.0141739f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.96
cc_5 VNB N_TE_c_63_n 0.0216364f $X=-0.19 $Y=-0.24 $X2=1.29 $Y2=1.035
cc_6 VNB N_TE_c_64_n 0.0182804f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=0.96
cc_7 VNB N_TE_c_65_n 0.00649751f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.035
cc_8 VNB TE 0.0134128f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_9 VNB N_A_27_47#_c_106_n 0.0155207f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.035
cc_10 VNB N_A_27_47#_c_107_n 0.00998586f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.142
cc_11 VNB N_A_27_47#_c_108_n 0.00709899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_109_n 0.027093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_c_173_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_14 VNB N_A_c_174_n 0.0186926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB A 0.0211887f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=0.96
cc_16 VNB N_A_c_176_n 0.0560577f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_17 VNB N_VPWR_c_212_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_315_n 4.00197e-19 $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.035
cc_19 VNB N_VGND_c_316_n 0.0059279f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.56
cc_20 VNB N_VGND_c_317_n 0.0143218f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=0.56
cc_21 VNB N_VGND_c_318_n 0.0123175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_319_n 0.0360649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_320_n 0.182872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_321_n 0.0047617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_322_n 0.00564938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_204_47#_c_364_n 0.00615837f $X=-0.19 $Y=-0.24 $X2=1.29 $Y2=1.035
cc_27 VNB N_A_204_47#_c_365_n 0.00293188f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.035
cc_28 VNB N_A_204_47#_c_366_n 0.0144618f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_29 VNB N_A_204_47#_c_367_n 0.00165125f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_30 VPB N_TE_M1004_g 0.0539915f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_31 VPB N_TE_c_61_n 0.01029f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.035
cc_32 VPB TE 0.0160305f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_33 VPB N_A_27_47#_c_110_n 0.0174982f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_34 VPB N_A_27_47#_c_111_n 0.00917137f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.035
cc_35 VPB N_A_27_47#_c_112_n 0.0092982f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.96
cc_36 VPB N_A_27_47#_c_113_n 0.0146322f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_37 VPB N_A_27_47#_c_114_n 0.00786149f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=0.96
cc_38 VPB N_A_27_47#_c_115_n 0.0198678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_116_n 0.0214591f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_40 VPB N_A_27_47#_c_108_n 0.0129676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_109_n 0.00100224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_M1002_g 0.0187578f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_43 VPB N_A_M1005_g 0.0211943f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_44 VPB A 0.01327f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=0.96
cc_45 VPB N_A_c_176_n 0.0155642f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_46 VPB N_VPWR_c_213_n 0.00652211f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.035
cc_47 VPB N_VPWR_c_214_n 4.07719e-19 $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_48 VPB N_VPWR_c_215_n 0.0150576f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=0.56
cc_49 VPB N_VPWR_c_216_n 0.0151073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_217_n 0.035677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_212_n 0.050982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_219_n 0.00565587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_220_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_215_309#_c_257_n 0.00737777f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_55 VPB N_A_215_309#_c_258_n 0.00166947f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.035
cc_56 VPB N_A_215_309#_c_259_n 0.00793407f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_57 VPB N_A_215_309#_c_260_n 0.0205972f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.142
cc_58 N_TE_c_63_n N_A_27_47#_c_112_n 0.00686796f $X=1.29 $Y=1.035 $X2=0 $Y2=0
cc_59 N_TE_M1004_g N_A_27_47#_c_116_n 0.0379477f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_60 N_TE_c_60_n N_A_27_47#_c_116_n 5.73392e-19 $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_61 N_TE_c_61_n N_A_27_47#_c_116_n 0.00264156f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_62 TE N_A_27_47#_c_116_n 0.0429593f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_63 N_TE_M1008_g N_A_27_47#_c_107_n 0.0239638f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_64 N_TE_c_60_n N_A_27_47#_c_107_n 0.0151409f $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_65 N_TE_c_61_n N_A_27_47#_c_107_n 0.0173893f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_66 N_TE_c_62_n N_A_27_47#_c_107_n 0.00787261f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_67 N_TE_c_64_n N_A_27_47#_c_107_n 7.19667e-19 $X=1.365 $Y=0.96 $X2=0 $Y2=0
cc_68 N_TE_c_65_n N_A_27_47#_c_107_n 0.00168518f $X=0.945 $Y=1.035 $X2=0 $Y2=0
cc_69 TE N_A_27_47#_c_107_n 0.0471178f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_70 N_TE_c_63_n N_A_27_47#_c_108_n 0.0182405f $X=1.29 $Y=1.035 $X2=0 $Y2=0
cc_71 N_TE_c_65_n N_A_27_47#_c_108_n 0.0111081f $X=0.945 $Y=1.035 $X2=0 $Y2=0
cc_72 N_TE_c_63_n N_A_27_47#_c_109_n 0.00728161f $X=1.29 $Y=1.035 $X2=0 $Y2=0
cc_73 N_TE_M1004_g N_VPWR_c_213_n 0.0113741f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_74 N_TE_M1004_g N_VPWR_c_215_n 0.0046653f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_75 N_TE_M1004_g N_VPWR_c_212_n 0.00523707f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_76 N_TE_M1004_g N_A_215_309#_c_257_n 0.00562299f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_77 N_TE_M1004_g N_A_215_309#_c_258_n 6.77363e-19 $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_78 N_TE_c_63_n N_A_215_309#_c_258_n 0.00116538f $X=1.29 $Y=1.035 $X2=0 $Y2=0
cc_79 N_TE_M1008_g N_VGND_c_315_n 0.00882192f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_80 N_TE_c_60_n N_VGND_c_315_n 5.89318e-19 $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_81 N_TE_c_62_n N_VGND_c_315_n 0.00557165f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_82 N_TE_c_64_n N_VGND_c_315_n 5.32619e-19 $X=1.365 $Y=0.96 $X2=0 $Y2=0
cc_83 N_TE_c_62_n N_VGND_c_316_n 5.66547e-19 $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_84 N_TE_c_64_n N_VGND_c_316_n 0.00807242f $X=1.365 $Y=0.96 $X2=0 $Y2=0
cc_85 N_TE_M1008_g N_VGND_c_317_n 0.00341574f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_86 N_TE_c_62_n N_VGND_c_318_n 0.00564095f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_87 N_TE_c_64_n N_VGND_c_318_n 0.00341689f $X=1.365 $Y=0.96 $X2=0 $Y2=0
cc_88 N_TE_M1008_g N_VGND_c_320_n 0.00501514f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_89 N_TE_c_62_n N_VGND_c_320_n 0.00950335f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_90 N_TE_c_64_n N_VGND_c_320_n 0.0040262f $X=1.365 $Y=0.96 $X2=0 $Y2=0
cc_91 N_TE_c_64_n N_A_204_47#_c_364_n 0.0124477f $X=1.365 $Y=0.96 $X2=0 $Y2=0
cc_92 N_TE_c_63_n N_A_204_47#_c_369_n 0.00186022f $X=1.29 $Y=1.035 $X2=0 $Y2=0
cc_93 N_TE_c_64_n N_A_204_47#_c_365_n 0.00320107f $X=1.365 $Y=0.96 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_114_n N_A_M1002_g 0.0217278f $X=1.655 $Y=1.32 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_108_n N_A_c_176_n 0.00343401f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_109_n N_A_c_176_n 0.0131652f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_116_n N_VPWR_M1004_d 0.00259802f $X=0.687 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_27_47#_c_110_n N_VPWR_c_213_n 0.00199804f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_116_n N_VPWR_c_213_n 0.0238531f $X=0.687 $Y=1.785 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_110_n N_VPWR_c_214_n 0.0109235f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_113_n N_VPWR_c_214_n 0.0120506f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_115_n N_VPWR_c_215_n 0.0176305f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_110_n N_VPWR_c_216_n 0.0046653f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_113_n N_VPWR_c_217_n 0.0046653f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_105 N_A_27_47#_M1004_s N_VPWR_c_212_n 0.00238524f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_110_n N_VPWR_c_212_n 0.00921786f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_113_n N_VPWR_c_212_n 0.00804845f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_115_n N_VPWR_c_212_n 0.00986266f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_116_n N_VPWR_c_212_n 0.00671954f $X=0.687 $Y=1.785 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_c_116_n N_A_215_309#_c_257_n 0.0194181f $X=0.687 $Y=1.785
+ $X2=0 $Y2=0
cc_111 N_A_27_47#_c_110_n N_A_215_309#_c_265_n 0.0156765f $X=1.41 $Y=1.47 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_c_111_n N_A_215_309#_c_265_n 0.00201418f $X=1.655 $Y=1.395
+ $X2=0 $Y2=0
cc_113 N_A_27_47#_c_113_n N_A_215_309#_c_265_n 0.0142044f $X=1.83 $Y=1.47 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_108_n N_A_215_309#_c_265_n 0.0460363f $X=1.79 $Y=1.16 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_116_n N_A_215_309#_c_258_n 0.0151769f $X=0.687 $Y=1.785
+ $X2=0 $Y2=0
cc_116 N_A_27_47#_c_108_n N_A_215_309#_c_258_n 0.0165264f $X=1.79 $Y=1.16 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_113_n N_A_215_309#_c_271_n 0.00463403f $X=1.83 $Y=1.47 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_c_113_n N_Z_c_297_n 2.45355e-19 $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_114_n N_Z_c_297_n 0.00122636f $X=1.655 $Y=1.32 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_108_n N_Z_c_297_n 0.0276571f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_109_n N_Z_c_297_n 2.37454e-19 $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_107_n N_VGND_M1008_d 0.00286332f $X=0.875 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_27_47#_c_107_n N_VGND_c_315_n 0.0227672f $X=0.875 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_106_n N_VGND_c_317_n 0.0177719f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_107_n N_VGND_c_317_n 0.00272678f $X=0.875 $Y=1.16 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_M1008_s N_VGND_c_320_n 0.00228937f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_106_n N_VGND_c_320_n 0.00989054f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_c_107_n N_VGND_c_320_n 0.00593319f $X=0.875 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_112_n N_A_204_47#_c_364_n 7.29275e-19 $X=1.485 $Y=1.395
+ $X2=0 $Y2=0
cc_130 N_A_27_47#_c_108_n N_A_204_47#_c_364_n 0.0688973f $X=1.79 $Y=1.16 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_c_109_n N_A_204_47#_c_364_n 0.00701665f $X=1.79 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_c_108_n N_A_204_47#_c_369_n 0.0141721f $X=1.79 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_M1002_g N_VPWR_c_214_n 0.00102048f $X=2.305 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_M1002_g N_VPWR_c_217_n 0.00357877f $X=2.305 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1005_g N_VPWR_c_217_n 0.00357877f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1002_g N_VPWR_c_212_n 0.00538183f $X=2.305 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_M1005_g N_VPWR_c_212_n 0.00620254f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_138 A N_A_215_309#_M1005_d 0.00347024f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_139 N_A_M1002_g N_A_215_309#_c_265_n 0.00149727f $X=2.305 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_M1002_g N_A_215_309#_c_271_n 0.00463843f $X=2.305 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_M1002_g N_A_215_309#_c_259_n 0.0112878f $X=2.305 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1005_g N_A_215_309#_c_259_n 0.0112437f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_143 A N_A_215_309#_c_260_n 0.0252364f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_144 N_A_c_176_n N_A_215_309#_c_260_n 0.00109684f $X=2.98 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_c_173_n N_Z_c_297_n 0.0115775f $X=2.305 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_Z_c_297_n 0.0129714f $X=2.305 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_c_174_n N_Z_c_297_n 0.0116146f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_Z_c_297_n 0.0165959f $X=2.725 $Y=1.985 $X2=0 $Y2=0
cc_149 A N_Z_c_297_n 0.054832f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_150 N_A_c_176_n N_Z_c_297_n 0.0215591f $X=2.98 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_c_173_n N_VGND_c_316_n 0.00319454f $X=2.305 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_173_n N_VGND_c_319_n 0.00357877f $X=2.305 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_174_n N_VGND_c_319_n 0.00357877f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_173_n N_VGND_c_320_n 0.00664112f $X=2.305 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_174_n N_VGND_c_320_n 0.00620254f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_156 A N_A_204_47#_M1007_d 0.00275832f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_157 N_A_c_173_n N_A_204_47#_c_366_n 0.0129376f $X=2.305 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_174_n N_A_204_47#_c_366_n 0.0112437f $X=2.725 $Y=0.995 $X2=0 $Y2=0
cc_159 A N_A_204_47#_c_366_n 0.0232068f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_160 N_A_c_176_n N_A_204_47#_c_366_n 0.00142902f $X=2.98 $Y=1.16 $X2=0 $Y2=0
cc_161 N_VPWR_c_212_n N_A_215_309#_M1001_d 0.00382897f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_162 N_VPWR_c_212_n N_A_215_309#_M1003_d 0.00533627f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_163 N_VPWR_c_212_n N_A_215_309#_M1005_d 0.00209324f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_213_n N_A_215_309#_c_257_n 0.0278322f $X=0.68 $Y=2.34 $X2=0
+ $Y2=0
cc_165 N_VPWR_c_216_n N_A_215_309#_c_257_n 0.0165671f $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_166 N_VPWR_c_212_n N_A_215_309#_c_257_n 0.0091658f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_167 N_VPWR_M1001_s N_A_215_309#_c_265_n 0.00328966f $X=1.485 $Y=1.545 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_214_n N_A_215_309#_c_265_n 0.0170258f $X=1.62 $Y=2.02 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_214_n N_A_215_309#_c_271_n 0.0260226f $X=1.62 $Y=2.02 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_217_n N_A_215_309#_c_259_n 0.0570633f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_212_n N_A_215_309#_c_259_n 0.0353389f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_214_n N_A_215_309#_c_290_n 0.0123818f $X=1.62 $Y=2.02 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_217_n N_A_215_309#_c_290_n 0.0119545f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_212_n N_A_215_309#_c_290_n 0.006547f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_175 N_VPWR_c_212_n N_Z_M1002_s 0.00216833f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_176 N_A_215_309#_c_259_n N_Z_M1002_s 0.00312348f $X=2.85 $Y=2.38 $X2=0 $Y2=0
cc_177 N_A_215_309#_c_265_n N_Z_c_297_n 0.0126255f $X=1.985 $Y=1.64 $X2=0 $Y2=0
cc_178 N_A_215_309#_c_271_n N_Z_c_297_n 0.0265342f $X=2.07 $Y=1.96 $X2=0 $Y2=0
cc_179 N_A_215_309#_c_259_n N_Z_c_297_n 0.015949f $X=2.85 $Y=2.38 $X2=0 $Y2=0
cc_180 N_Z_M1006_s N_VGND_c_320_n 0.00216833f $X=2.38 $Y=0.235 $X2=0.687
+ $Y2=1.075
cc_181 N_Z_M1006_s N_A_204_47#_c_366_n 0.00303482f $X=2.38 $Y=0.235 $X2=0 $Y2=0
cc_182 N_Z_c_297_n N_A_204_47#_c_366_n 0.015949f $X=2.515 $Y=0.76 $X2=0 $Y2=0
cc_183 N_VGND_c_320_n N_A_204_47#_M1000_s 0.00325955f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_184 N_VGND_c_320_n N_A_204_47#_M1006_d 0.00210127f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_185 N_VGND_c_320_n N_A_204_47#_M1007_d 0.00208521f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_318_n N_A_204_47#_c_385_n 0.0121424f $X=1.41 $Y=0 $X2=0 $Y2=0
cc_187 N_VGND_c_320_n N_A_204_47#_c_385_n 0.00739874f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_188 N_VGND_M1009_d N_A_204_47#_c_364_n 0.0046626f $X=1.44 $Y=0.235 $X2=0
+ $Y2=0
cc_189 N_VGND_c_316_n N_A_204_47#_c_364_n 0.0231246f $X=1.575 $Y=0.38 $X2=0
+ $Y2=0
cc_190 N_VGND_c_318_n N_A_204_47#_c_364_n 0.00232396f $X=1.41 $Y=0 $X2=0 $Y2=0
cc_191 N_VGND_c_319_n N_A_204_47#_c_364_n 0.00296166f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_c_320_n N_A_204_47#_c_364_n 0.0104609f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_c_316_n N_A_204_47#_c_365_n 0.0048719f $X=1.575 $Y=0.38 $X2=0
+ $Y2=0
cc_194 N_VGND_c_319_n N_A_204_47#_c_366_n 0.0547026f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_320_n N_A_204_47#_c_366_n 0.0342286f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_316_n N_A_204_47#_c_367_n 0.0151323f $X=1.575 $Y=0.38 $X2=0
+ $Y2=0
cc_197 N_VGND_c_319_n N_A_204_47#_c_367_n 0.0164632f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_320_n N_A_204_47#_c_367_n 0.0092005f $X=2.99 $Y=0 $X2=0 $Y2=0

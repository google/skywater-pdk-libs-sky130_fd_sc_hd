* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_2.spice
* Created: Thu Aug 27 14:23:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_2.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_2  VNB VPB A KAPWR X VGND VPWR
* 
* VGND	VGND
* X	X
* KAPWR	KAPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_27_47#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.1113 PD=0.745 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_27_47#_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.06825 PD=0.69 PS=0.745 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1003_d N_A_27_47#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_KAPWR_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1625 AS=0.265 PD=1.325 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_27_47#_M1000_g N_KAPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1625 PD=1.27 PS=1.325 NRD=0 NRS=8.8453 M=1 R=6.66667 SA=75000.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1000_d N_A_27_47#_M1005_g N_KAPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=3.5631 P=7.65
c_37 VPB 0 8.20068e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_2.pxi.spice"
*
.ends
*
*

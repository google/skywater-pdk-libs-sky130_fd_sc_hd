* NGSPICE file created from sky130_fd_sc_hd__xor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
M1000 a_470_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=1.33e+12p pd=1.266e+07u as=8.65e+11p ps=7.73e+06u
M1001 X B a_470_47# VNB nshort w=650000u l=150000u
+  ad=3.8675e+11p pd=3.79e+06u as=5.135e+11p ps=5.48e+06u
M1002 VPWR A a_470_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_470_297# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=8.05e+11p ps=7.61e+06u
M1005 VGND A a_470_47# VNB nshort w=650000u l=150000u
+  ad=1.03675e+12p pd=1.099e+07u as=0p ps=0u
M1006 VPWR B a_470_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_112_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_112_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_112_47# B VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=0p ps=0u
M1010 a_470_297# a_112_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1011 VGND A a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_470_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_297# B a_112_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1014 a_112_47# B a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B a_112_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_112_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_112_47# a_470_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_470_47# B X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


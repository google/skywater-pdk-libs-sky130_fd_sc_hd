* File: sky130_fd_sc_hd__and3b_2.spice.pex
* Created: Thu Aug 27 14:08:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND3B_2%A_N 3 7 9 10 16
c26 9 0 1.51555e-19 $X=0.145 $Y=0.765
r27 14 16 29.6615 $w=3.25e-07 $l=2e-07 $layer=POLY_cond $X=0.27 $Y=1.16 $X2=0.47
+ $Y2=1.16
r28 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r29 9 10 13.4814 $w=2.63e-07 $l=3.1e-07 $layer=LI1_cond $X=0.277 $Y=0.85
+ $X2=0.277 $Y2=1.16
r30 5 16 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.16
r31 5 7 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.765
r32 1 16 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=1.16
r33 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_2%A_109_53# 1 2 9 13 17 21 25 28 32
c42 32 0 1.51555e-19 $X=1.43 $Y=1.16
c43 25 0 1.91433e-19 $X=1.22 $Y=1.16
r44 31 32 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.41 $Y=1.16 $X2=1.43
+ $Y2=1.16
r45 26 31 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.22 $Y=1.16
+ $X2=1.41 $Y2=1.16
r46 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.16 $X2=1.22 $Y2=1.16
r47 23 28 1.99325 $w=2.3e-07 $l=1.38e-07 $layer=LI1_cond $X=0.855 $Y=1.13
+ $X2=0.717 $Y2=1.13
r48 23 25 18.2888 $w=2.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.855 $Y=1.13
+ $X2=1.22 $Y2=1.13
r49 19 28 4.44123 $w=2.75e-07 $l=1.15e-07 $layer=LI1_cond $X=0.717 $Y=1.245
+ $X2=0.717 $Y2=1.13
r50 19 21 20.744 $w=2.73e-07 $l=4.95e-07 $layer=LI1_cond $X=0.717 $Y=1.245
+ $X2=0.717 $Y2=1.74
r51 15 28 4.44123 $w=2.75e-07 $l=1.15e-07 $layer=LI1_cond $X=0.717 $Y=1.015
+ $X2=0.717 $Y2=1.13
r52 15 17 22.8393 $w=2.73e-07 $l=5.45e-07 $layer=LI1_cond $X=0.717 $Y=1.015
+ $X2=0.717 $Y2=0.47
r53 11 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.16
r54 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.475
r55 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r56 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.41 $Y=1.325 $X2=1.41
+ $Y2=1.765
r57 2 21 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.555 $X2=0.68 $Y2=1.74
r58 1 17 182 $w=1.7e-07 $l=2.71662e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.265 $X2=0.7 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_2%B 3 8 10 11 14
c38 14 0 1.62801e-19 $X=1.9 $Y=2.3
c39 10 0 3.17214e-19 $X=1.81 $Y=1.2
c40 8 0 3.5796e-20 $X=1.83 $Y=1.765
r41 14 16 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=2.3
+ $X2=1.895 $Y2=2.135
r42 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.9 $Y=2.3
+ $X2=1.9 $Y2=2.3
r43 11 15 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=2.095 $Y=2.295
+ $X2=1.9 $Y2=2.295
r44 9 10 66.5448 $w=1.9e-07 $l=1.85e-07 $layer=POLY_cond $X=1.81 $Y=1.015
+ $X2=1.81 $Y2=1.2
r45 8 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.83 $Y=1.765
+ $X2=1.83 $Y2=2.135
r46 8 10 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.83 $Y=1.765
+ $X2=1.83 $Y2=1.2
r47 3 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.79 $Y=0.475 $X2=1.79
+ $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_2%C 3 7 9 10 15
r46 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.255 $Y2=1.325
r47 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.255 $Y2=0.995
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=1.16 $X2=2.255 $Y2=1.16
r49 10 16 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=2.215 $Y=0.85
+ $X2=2.215 $Y2=1.16
r50 9 10 10.0225 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.115 $Y=0.51
+ $X2=2.115 $Y2=0.765
r51 7 18 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.305 $Y=1.695
+ $X2=2.305 $Y2=1.325
r52 3 17 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.195 $Y=0.475
+ $X2=2.195 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_2%A_215_311# 1 2 3 10 12 15 17 19 22 26 28 32
+ 33 35 38 40 41 44 52
c109 41 0 1.61577e-19 $X=2.2 $Y=1.51
c110 38 0 1.62801e-19 $X=2.095 $Y=1.725
r111 51 52 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.79 $Y=1.16
+ $X2=3.21 $Y2=1.16
r112 45 51 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=2.79 $Y2=1.16
r113 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.735
+ $Y=1.16 $X2=2.735 $Y2=1.16
r114 42 44 13.2781 $w=2.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.705 $Y=1.425
+ $X2=2.705 $Y2=1.16
r115 41 48 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.2 $Y=1.51
+ $X2=2.105 $Y2=1.51
r116 40 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.59 $Y=1.51
+ $X2=2.705 $Y2=1.425
r117 40 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.59 $Y=1.51
+ $X2=2.2 $Y2=1.51
r118 36 48 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=1.595
+ $X2=2.105 $Y2=1.51
r119 36 38 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.105 $Y=1.595
+ $X2=2.105 $Y2=1.725
r120 35 48 25.6396 $w=1.68e-07 $l=3.93e-07 $layer=LI1_cond $X=1.712 $Y=1.51
+ $X2=2.105 $Y2=1.51
r121 34 35 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=1.712 $Y=0.57
+ $X2=1.712 $Y2=1.425
r122 32 35 8.28556 $w=1.68e-07 $l=1.27e-07 $layer=LI1_cond $X=1.585 $Y=1.51
+ $X2=1.712 $Y2=1.51
r123 32 33 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.585 $Y=1.51
+ $X2=1.285 $Y2=1.51
r124 28 34 6.81977 $w=2.65e-07 $l=1.85957e-07 $layer=LI1_cond $X=1.585 $Y=0.437
+ $X2=1.712 $Y2=0.57
r125 28 30 15.8733 $w=2.63e-07 $l=3.65e-07 $layer=LI1_cond $X=1.585 $Y=0.437
+ $X2=1.22 $Y2=0.437
r126 24 33 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=1.167 $Y=1.595
+ $X2=1.285 $Y2=1.51
r127 24 26 8.09162 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.167 $Y=1.595
+ $X2=1.167 $Y2=1.76
r128 20 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r129 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.985
r130 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r131 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=0.56
r132 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.325
+ $X2=2.79 $Y2=1.16
r133 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.79 $Y=1.325
+ $X2=2.79 $Y2=1.985
r134 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=0.995
+ $X2=2.79 $Y2=1.16
r135 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.79 $Y=0.995
+ $X2=2.79 $Y2=0.56
r136 3 38 600 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.555 $X2=2.095 $Y2=1.725
r137 2 26 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.555 $X2=1.2 $Y2=1.76
r138 1 30 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.265 $X2=1.22 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_2%VPWR 1 2 3 4 13 15 19 23 25 27 32 34 36 41
+ 50 57 61
r57 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 54 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 52 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 45 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 45 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r63 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 42 57 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=2.675 $Y=2.72
+ $X2=2.567 $Y2=2.72
r65 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.675 $Y=2.72
+ $X2=2.99 $Y2=2.72
r66 41 60 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=3.505 $Y2=2.72
r67 41 44 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=2.99 $Y2=2.72
r68 40 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 37 47 4.67309 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.2
+ $Y2=2.72
r71 37 39 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.69
+ $Y2=2.72
r72 36 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 36 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 36 50 17.7217 $w=6.13e-07 $l=5.9e-07 $layer=LI1_cond $X=1.337 $Y=2.72
+ $X2=1.337 $Y2=2.13
r75 36 39 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.03 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 34 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 34 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 29 32 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=1.55 $Y=1.86 $X2=1.62
+ $Y2=1.86
r79 25 60 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.462 $Y=2.635
+ $X2=3.505 $Y2=2.72
r80 25 27 29.3547 $w=2.63e-07 $l=6.75e-07 $layer=LI1_cond $X=3.462 $Y=2.635
+ $X2=3.462 $Y2=1.96
r81 21 57 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.567 $Y=2.635
+ $X2=2.567 $Y2=2.72
r82 21 23 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=2.567 $Y=2.635
+ $X2=2.567 $Y2=1.955
r83 20 36 8.47627 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=1.337 $Y2=2.72
r84 19 57 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.46 $Y=2.72
+ $X2=2.567 $Y2=2.72
r85 19 20 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.46 $Y=2.72
+ $X2=1.645 $Y2=2.72
r86 17 29 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.55 $Y=1.955
+ $X2=1.55 $Y2=1.86
r87 17 50 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=1.55 $Y=1.955
+ $X2=1.55 $Y2=2.13
r88 13 47 2.96741 $w=3.15e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.2 $Y2=2.72
r89 13 15 32.744 $w=3.13e-07 $l=8.95e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=1.74
r90 4 27 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.96
r91 3 23 300 $w=1.7e-07 $l=5.61159e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=1.485 $X2=2.58 $Y2=1.955
r92 2 32 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.555 $X2=1.62 $Y2=1.85
r93 1 15 600 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.555 $X2=0.26 $Y2=1.74
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_2%X 1 2 8 11 12 13 14 15 20 23 26
r34 20 23 4.13306 $w=2.45e-07 $l=8.3e-08 $layer=LI1_cond $X=3.037 $Y=0.593
+ $X2=3.037 $Y2=0.51
r35 15 32 8.51056 $w=5.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.445 $Y=1.185
+ $X2=3.075 $Y2=1.185
r36 14 26 10.1091 $w=2.83e-07 $l=2.5e-07 $layer=LI1_cond $X=3.017 $Y=2.21
+ $X2=3.017 $Y2=1.96
r37 13 31 6.78285 $w=2.43e-07 $l=1.21e-07 $layer=LI1_cond $X=3.037 $Y=0.594
+ $X2=3.037 $Y2=0.715
r38 13 20 0.0470385 $w=2.43e-07 $l=1e-09 $layer=LI1_cond $X=3.037 $Y=0.594
+ $X2=3.037 $Y2=0.593
r39 13 23 0.0497959 $w=2.45e-07 $l=1e-09 $layer=LI1_cond $X=3.037 $Y=0.509
+ $X2=3.037 $Y2=0.51
r40 11 26 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=3.017 $Y=1.937
+ $X2=3.017 $Y2=1.96
r41 11 12 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=3.017 $Y=1.937
+ $X2=3.017 $Y2=1.795
r42 9 32 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=3.075 $Y=1.445
+ $X2=3.075 $Y2=1.185
r43 9 12 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.075 $Y=1.445
+ $X2=3.075 $Y2=1.795
r44 8 32 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=3.075 $Y=0.925
+ $X2=3.075 $Y2=1.185
r45 8 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.075 $Y=0.925
+ $X2=3.075 $Y2=0.715
r46 2 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.865
+ $Y=1.485 $X2=3 $Y2=1.96
r47 1 23 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_2%VGND 1 2 3 10 12 16 18 20 22 24 32 41 45
r45 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r46 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r47 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r48 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r49 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r50 33 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.575
+ $Y2=0
r51 33 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.99
+ $Y2=0
r52 32 44 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.505
+ $Y2=0
r53 32 35 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=2.99
+ $Y2=0
r54 31 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r55 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r56 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r57 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r58 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r59 25 38 4.2375 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r60 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.69
+ $Y2=0
r61 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.575
+ $Y2=0
r62 24 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.07
+ $Y2=0
r63 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r64 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r65 18 44 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.462 $Y=0.085
+ $X2=3.505 $Y2=0
r66 18 20 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=3.462 $Y=0.085
+ $X2=3.462 $Y2=0.515
r67 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=0.085
+ $X2=2.575 $Y2=0
r68 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.575 $Y=0.085
+ $X2=2.575 $Y2=0.495
r69 10 38 3.04719 $w=2.7e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.177 $Y2=0
r70 10 12 13.872 $w=2.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.22 $Y2=0.41
r71 3 20 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.515
r72 2 16 182 $w=1.7e-07 $l=4.03949e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.265 $X2=2.575 $Y2=0.495
r73 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.41
.ends


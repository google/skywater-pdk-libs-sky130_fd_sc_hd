* NGSPICE file created from sky130_fd_sc_hd__ebufn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_320_309# VPB phighvt w=940000u l=150000u
+  ad=8.826e+11p pd=7.59e+06u as=1.7987e+12p ps=1.343e+07u
M1001 a_320_309# a_27_47# Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.4e+11p ps=5.08e+06u
M1002 a_214_47# TE_B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1003 VGND a_214_47# a_393_47# VNB nshort w=650000u l=150000u
+  ad=5.9475e+11p pd=5.73e+06u as=9.555e+11p ps=9.44e+06u
M1004 a_393_47# a_214_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_214_47# a_393_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_393_47# a_214_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z a_27_47# a_393_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=0p ps=0u
M1008 a_393_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_320_309# a_27_47# Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_393_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_320_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Z a_27_47# a_320_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1014 a_214_47# TE_B VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1015 Z a_27_47# a_393_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR TE_B a_320_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Z a_27_47# a_320_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1019 a_320_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


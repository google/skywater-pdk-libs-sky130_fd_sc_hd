* File: sky130_fd_sc_hd__xor3_4.pex.spice
* Created: Thu Aug 27 14:50:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XOR3_4%A_79_21# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 38 41 42 43 45 47 49 50 52 54 56 58 59 68
c143 56 0 1.80415e-19 $X=1.932 $Y=1.325
c144 42 0 8.82126e-20 $X=2.375 $Y=1.96
c145 33 0 1.53226e-19 $X=1.83 $Y=1.985
r146 67 68 14.6505 $w=3.29e-07 $l=1e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.83 $Y2=1.16
r147 66 67 46.8815 $w=3.29e-07 $l=3.2e-07 $layer=POLY_cond $X=1.41 $Y=1.16
+ $X2=1.73 $Y2=1.16
r148 65 66 14.6505 $w=3.29e-07 $l=1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.41 $Y2=1.16
r149 64 65 46.8815 $w=3.29e-07 $l=3.2e-07 $layer=POLY_cond $X=0.99 $Y=1.16
+ $X2=1.31 $Y2=1.16
r150 63 64 14.6505 $w=3.29e-07 $l=1e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.99 $Y2=1.16
r151 62 63 46.8815 $w=3.29e-07 $l=3.2e-07 $layer=POLY_cond $X=0.57 $Y=1.16
+ $X2=0.89 $Y2=1.16
r152 61 62 14.6505 $w=3.29e-07 $l=1e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.57 $Y2=1.16
r153 58 59 10.5404 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=3.595 $Y=0.355
+ $X2=3.41 $Y2=0.355
r154 54 55 18.4591 $w=2.3e-07 $l=3.48e-07 $layer=LI1_cond $X=1.932 $Y=0.865
+ $X2=2.28 $Y2=0.865
r155 50 52 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=2.545 $Y=2.32
+ $X2=3.6 $Y2=2.32
r156 49 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=2.235
+ $X2=2.545 $Y2=2.32
r157 48 49 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=2.045
+ $X2=2.46 $Y2=2.235
r158 47 59 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=2.365 $Y=0.34
+ $X2=3.41 $Y2=0.34
r159 45 55 2.50919 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.28 $Y=0.695
+ $X2=2.28 $Y2=0.865
r160 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.28 $Y=0.425
+ $X2=2.365 $Y2=0.34
r161 44 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.28 $Y=0.425
+ $X2=2.28 $Y2=0.695
r162 42 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=1.96
+ $X2=2.46 $Y2=2.045
r163 42 43 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.375 $Y=1.96
+ $X2=2.045 $Y2=1.96
r164 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.96 $Y=1.875
+ $X2=2.045 $Y2=1.96
r165 41 56 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.96 $Y=1.875
+ $X2=1.96 $Y2=1.325
r166 39 68 10.9878 $w=3.29e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.16
+ $X2=1.83 $Y2=1.16
r167 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.905
+ $Y=1.16 $X2=1.905 $Y2=1.16
r168 36 56 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.932 $Y=1.213
+ $X2=1.932 $Y2=1.325
r169 36 38 2.71464 $w=2.23e-07 $l=5.3e-08 $layer=LI1_cond $X=1.932 $Y=1.213
+ $X2=1.932 $Y2=1.16
r170 35 54 0.876693 $w=2.25e-07 $l=2.12e-07 $layer=LI1_cond $X=1.932 $Y=1.077
+ $X2=1.932 $Y2=0.865
r171 35 38 4.25123 $w=2.23e-07 $l=8.3e-08 $layer=LI1_cond $X=1.932 $Y=1.077
+ $X2=1.932 $Y2=1.16
r172 31 68 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.16
r173 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.985
r174 28 67 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r175 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r176 24 66 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r177 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.985
r178 21 65 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r179 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r180 17 64 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.325
+ $X2=0.99 $Y2=1.16
r181 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.99 $Y=1.325
+ $X2=0.99 $Y2=1.985
r182 14 63 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r183 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r184 10 62 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.325
+ $X2=0.57 $Y2=1.16
r185 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.57 $Y=1.325
+ $X2=0.57 $Y2=1.985
r186 7 61 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r187 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r188 2 52 600 $w=1.7e-07 $l=7.79824e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.625 $X2=3.6 $Y2=2.32
r189 1 58 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.46
+ $Y=0.245 $X2=3.595 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%C 1 3 4 6 7 11 13 15 16 17 20 21
c67 7 0 8.82126e-20 $X=3.27 $Y=1.16
r68 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.33
+ $Y=1.16 $X2=3.33 $Y2=1.16
r69 17 21 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.09 $Y=1.16 $X2=3.33
+ $Y2=1.16
r70 13 20 37.0704 $w=1.5e-07 $l=1.19896e-07 $layer=POLY_cond $X=3.385 $Y=0.985
+ $X2=3.27 $Y2=0.995
r71 13 15 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.385 $Y=0.985
+ $X2=3.385 $Y2=0.565
r72 9 20 37.0704 $w=1.5e-07 $l=3.95727e-07 $layer=POLY_cond $X=3.345 $Y=1.355
+ $X2=3.27 $Y2=0.995
r73 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.345 $Y=1.355
+ $X2=3.345 $Y2=2.045
r74 8 16 5.03009 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.49 $Y=1.16 $X2=2.37
+ $Y2=1.16
r75 7 20 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.16
+ $X2=3.27 $Y2=0.995
r76 7 8 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=3.27 $Y=1.16 $X2=2.49
+ $Y2=1.16
r77 4 16 37.0704 $w=1.5e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.415 $Y=0.995
+ $X2=2.37 $Y2=1.16
r78 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.415 $Y=0.995
+ $X2=2.415 $Y2=0.675
r79 1 16 37.0704 $w=1.5e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.325 $Y=1.325
+ $X2=2.37 $Y2=1.16
r80 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.325 $Y=1.325
+ $X2=2.325 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%A_480_297# 1 2 9 13 14 16 18 21 27 28 31
c77 14 0 1.53226e-19 $X=2.625 $Y=1.535
r78 28 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=1.16
+ $X2=3.875 $Y2=0.995
r79 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.875
+ $Y=1.16 $X2=3.875 $Y2=1.16
r80 24 27 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.77 $Y=1.16
+ $X2=3.875 $Y2=1.16
r81 20 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.77 $Y=1.325
+ $X2=3.77 $Y2=1.16
r82 20 21 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.77 $Y=1.325
+ $X2=3.77 $Y2=1.535
r83 19 23 3.40825 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.71 $Y=1.62 $X2=2.54
+ $Y2=1.62
r84 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=1.62
+ $X2=3.77 $Y2=1.535
r85 18 19 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=3.685 $Y=1.62
+ $X2=2.71 $Y2=1.62
r86 14 23 3.40825 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.625 $Y=1.535
+ $X2=2.54 $Y2=1.62
r87 14 16 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.625 $Y=1.535
+ $X2=2.625 $Y2=0.76
r88 13 31 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.935 $Y=0.565
+ $X2=3.935 $Y2=0.995
r89 7 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=1.325
+ $X2=3.875 $Y2=1.16
r90 7 9 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=3.875 $Y=1.325
+ $X2=3.875 $Y2=2.045
r91 2 23 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.485 $X2=2.575 $Y2=1.62
r92 1 16 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.465 $X2=2.625 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%A_1031_297# 1 2 9 13 15 17 19 21 22 23 27 35
+ 37 38 39 40 47 49 50 58
c168 49 0 1.83334e-19 $X=8.15 $Y=0.85
c169 15 0 1.24749e-19 $X=8.325 $Y=1.28
r170 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.27
+ $Y=1.11 $X2=8.27 $Y2=1.11
r171 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.2 $Y=0.85 $X2=8.2
+ $Y2=1.11
r172 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.15 $Y=0.85
+ $X2=8.15 $Y2=0.85
r173 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.77 $Y=0.85
+ $X2=6.77 $Y2=0.85
r174 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.39 $Y=0.85
+ $X2=5.39 $Y2=0.85
r175 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.915 $Y=0.85
+ $X2=6.77 $Y2=0.85
r176 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.005 $Y=0.85
+ $X2=8.15 $Y2=0.85
r177 39 40 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=8.005 $Y=0.85
+ $X2=6.915 $Y2=0.85
r178 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.535 $Y=0.85
+ $X2=5.39 $Y2=0.85
r179 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=0.85
+ $X2=6.77 $Y2=0.85
r180 37 38 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=6.625 $Y=0.85
+ $X2=5.535 $Y2=0.85
r181 35 47 7.77229 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=6.747 $Y=0.995
+ $X2=6.747 $Y2=0.85
r182 31 35 6.36987 $w=2.73e-07 $l=1.52e-07 $layer=LI1_cond $X=6.595 $Y=1.132
+ $X2=6.747 $Y2=1.132
r183 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.595
+ $Y=1.16 $X2=6.595 $Y2=1.16
r184 28 58 34.8134 $w=2.38e-07 $l=7.25e-07 $layer=LI1_cond $X=5.42 $Y=1.445
+ $X2=5.42 $Y2=0.72
r185 27 28 1.42499 $w=2.4e-07 $l=1.35e-07 $layer=LI1_cond $X=5.42 $Y=1.58
+ $X2=5.42 $Y2=1.445
r186 25 27 5.5488 $w=2.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.29 $Y=1.58
+ $X2=5.42 $Y2=1.58
r187 22 32 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.86 $Y=1.16
+ $X2=6.595 $Y2=1.16
r188 22 23 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.86 $Y=1.16
+ $X2=6.935 $Y2=1.16
r189 19 55 38.945 $w=2.68e-07 $l=1.92678e-07 $layer=POLY_cond $X=8.33 $Y=0.945
+ $X2=8.27 $Y2=1.11
r190 19 21 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.33 $Y=0.945
+ $X2=8.33 $Y2=0.535
r191 15 55 39.8442 $w=2.68e-07 $l=1.95576e-07 $layer=POLY_cond $X=8.325 $Y=1.28
+ $X2=8.27 $Y2=1.11
r192 15 17 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=8.325 $Y=1.28
+ $X2=8.325 $Y2=2.065
r193 11 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.935 $Y=1.325
+ $X2=6.935 $Y2=1.16
r194 11 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.935 $Y=1.325
+ $X2=6.935 $Y2=1.805
r195 7 23 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.935 $Y=0.995
+ $X2=6.935 $Y2=1.16
r196 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.935 $Y=0.995
+ $X2=6.935 $Y2=0.455
r197 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.155
+ $Y=1.485 $X2=5.29 $Y2=1.63
r198 1 58 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.235 $X2=5.455 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%B 3 7 9 10 13 18 19 20 23 27 31 34 35 37 38
+ 41
r121 37 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.875 $Y=1.53
+ $X2=8.15 $Y2=1.53
r122 35 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.16
+ $X2=7.79 $Y2=1.325
r123 35 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.16
+ $X2=7.79 $Y2=0.995
r124 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.79
+ $Y=1.16 $X2=7.79 $Y2=1.16
r125 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.79 $Y=1.445
+ $X2=7.875 $Y2=1.53
r126 32 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.79 $Y=1.445
+ $X2=7.79 $Y2=1.16
r127 28 30 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.08 $Y=1.16
+ $X2=5.245 $Y2=1.16
r128 27 42 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.81 $Y=1.965
+ $X2=7.81 $Y2=1.325
r129 25 27 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.81 $Y=2.465
+ $X2=7.81 $Y2=1.965
r130 23 41 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.73 $Y=0.565
+ $X2=7.73 $Y2=0.995
r131 19 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.735 $Y=2.54
+ $X2=7.81 $Y2=2.465
r132 19 20 761.457 $w=1.5e-07 $l=1.485e-06 $layer=POLY_cond $X=7.735 $Y=2.54
+ $X2=6.25 $Y2=2.54
r133 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.175 $Y=2.465
+ $X2=6.25 $Y2=2.54
r134 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.175 $Y=2.465
+ $X2=6.175 $Y2=1.905
r135 15 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.175 $Y=1.235
+ $X2=6.175 $Y2=1.16
r136 15 18 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.175 $Y=1.235
+ $X2=6.175 $Y2=1.905
r137 11 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.175 $Y=1.085
+ $X2=6.175 $Y2=1.16
r138 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.175 $Y=1.085
+ $X2=6.175 $Y2=0.565
r139 10 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.32 $Y=1.16
+ $X2=5.245 $Y2=1.16
r140 9 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.1 $Y=1.16
+ $X2=6.175 $Y2=1.16
r141 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.1 $Y=1.16 $X2=5.32
+ $Y2=1.16
r142 5 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.245 $Y=1.085
+ $X2=5.245 $Y2=1.16
r143 5 7 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.245 $Y=1.085
+ $X2=5.245 $Y2=0.56
r144 1 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.08 $Y=1.235
+ $X2=5.08 $Y2=1.16
r145 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.08 $Y=1.235
+ $X2=5.08 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%A 3 6 8 11 12 13
c43 13 0 1.83334e-19 $X=8.76 $Y=0.995
r44 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=1.16
+ $X2=8.76 $Y2=1.325
r45 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=1.16
+ $X2=8.76 $Y2=0.995
r46 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.75
+ $Y=1.16 $X2=8.75 $Y2=1.16
r47 8 12 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=8.61 $Y=1.2 $X2=8.75
+ $Y2=1.2
r48 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.83 $Y=1.985
+ $X2=8.83 $Y2=1.325
r49 3 13 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.83 $Y=0.555
+ $X2=8.83 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%A_1135_365# 1 2 3 4 15 18 22 24 28 29 30 31
+ 36 37 38 41 44 45 48
c133 36 0 1.98666e-19 $X=9.25 $Y=1.16
c134 31 0 1.06604e-19 $X=9.19 $Y=1.495
c135 30 0 1.15937e-19 $X=9.19 $Y=1.325
r136 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.61 $Y=0.51
+ $X2=8.61 $Y2=0.51
r137 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.85 $Y=0.51
+ $X2=5.85 $Y2=0.51
r138 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.995 $Y=0.51
+ $X2=5.85 $Y2=0.51
r139 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.465 $Y=0.51
+ $X2=8.61 $Y2=0.51
r140 37 38 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=8.465 $Y=0.51
+ $X2=5.995 $Y2=0.51
r141 36 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.16
+ $X2=9.25 $Y2=1.325
r142 36 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.16
+ $X2=9.25 $Y2=0.995
r143 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.25
+ $Y=1.16 $X2=9.25 $Y2=1.16
r144 33 35 20.4335 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=9.22 $Y=0.82
+ $X2=9.22 $Y2=1.16
r145 32 45 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=8.64 $Y=0.735
+ $X2=8.64 $Y2=0.51
r146 30 35 10.2745 $w=2.03e-07 $l=1.79374e-07 $layer=LI1_cond $X=9.19 $Y=1.325
+ $X2=9.22 $Y2=1.16
r147 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.19 $Y=1.325
+ $X2=9.19 $Y2=1.495
r148 29 32 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=8.785 $Y=0.82
+ $X2=8.64 $Y2=0.735
r149 28 33 1.77774 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.105 $Y=0.82
+ $X2=9.22 $Y2=0.82
r150 28 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.105 $Y=0.82
+ $X2=8.785 $Y2=0.82
r151 24 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.105 $Y=1.6
+ $X2=9.19 $Y2=1.495
r152 24 26 25.6147 $w=2.08e-07 $l=4.85e-07 $layer=LI1_cond $X=9.105 $Y=1.6
+ $X2=8.62 $Y2=1.6
r153 20 41 3.61456 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=0.595
+ $X2=5.8 $Y2=0.43
r154 20 22 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.8 $Y=0.595
+ $X2=5.8 $Y2=1.94
r155 18 49 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.29 $Y=1.985
+ $X2=9.29 $Y2=1.325
r156 15 48 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.29 $Y=0.555
+ $X2=9.29 $Y2=0.995
r157 4 26 600 $w=1.7e-07 $l=2.32164e-07 $layer=licon1_PDIFF $count=1 $X=8.4
+ $Y=1.645 $X2=8.62 $Y2=1.62
r158 3 22 600 $w=1.7e-07 $l=1.73205e-07 $layer=licon1_PDIFF $count=1 $X=5.675
+ $Y=1.825 $X2=5.8 $Y2=1.94
r159 2 45 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=8.405
+ $Y=0.235 $X2=8.62 $Y2=0.625
r160 1 41 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.245 $X2=5.965 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 39 44 48
+ 53 61 68 69 72 75 78 81 84 87
c119 5 0 1.06604e-19 $X=8.905 $Y=1.485
r120 84 87 0.000284542 $w=4.8e-07 $l=1e-09 $layer=MET1_cond $X=0.229 $Y=2.72
+ $X2=0.23 $Y2=2.72
r121 81 82 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r122 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r125 69 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=8.97 $Y2=2.72
r126 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r127 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.245 $Y=2.72
+ $X2=9.08 $Y2=2.72
r128 66 68 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=9.245 $Y=2.72
+ $X2=9.89 $Y2=2.72
r129 65 82 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=8.97 $Y2=2.72
r130 65 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r131 64 65 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r132 62 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=2.72
+ $X2=4.87 $Y2=2.72
r133 62 64 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.035 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 61 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.915 $Y=2.72
+ $X2=9.08 $Y2=2.72
r135 61 64 236.497 $w=1.68e-07 $l=3.625e-06 $layer=LI1_cond $X=8.915 $Y=2.72
+ $X2=5.29 $Y2=2.72
r136 60 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r137 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r138 57 60 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.37 $Y2=2.72
r139 57 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r140 56 59 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r142 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.04 $Y2=2.72
r143 54 56 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.53 $Y2=2.72
r144 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=2.72
+ $X2=4.87 $Y2=2.72
r145 53 59 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.705 $Y=2.72
+ $X2=4.37 $Y2=2.72
r146 52 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r147 52 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r149 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r150 49 51 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r151 48 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=2.04 $Y2=2.72
r152 48 51 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=1.61 $Y2=2.72
r153 47 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r154 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r155 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r156 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r157 42 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r158 39 47 0.10528 $w=4.8e-07 $l=3.7e-07 $layer=MET1_cond $X=0.32 $Y=2.72
+ $X2=0.69 $Y2=2.72
r159 39 87 0.0256088 $w=4.8e-07 $l=9e-08 $layer=MET1_cond $X=0.32 $Y=2.72
+ $X2=0.23 $Y2=2.72
r160 37 42 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=0.275 $Y=2.72
+ $X2=0.23 $Y2=2.72
r161 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=2.72
+ $X2=0.36 $Y2=2.72
r162 36 46 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.69 $Y2=2.72
r163 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.36 $Y2=2.72
r164 32 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.08 $Y=2.635
+ $X2=9.08 $Y2=2.72
r165 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.08 $Y=2.635
+ $X2=9.08 $Y2=2.36
r166 28 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=2.635
+ $X2=4.87 $Y2=2.72
r167 28 30 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.87 $Y=2.635
+ $X2=4.87 $Y2=2.32
r168 24 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r169 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.3
r170 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r171 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.3
r172 16 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.36 $Y=2.635
+ $X2=0.36 $Y2=2.72
r173 16 18 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.36 $Y=2.635
+ $X2=0.36 $Y2=2.3
r174 5 34 600 $w=1.7e-07 $l=9.58514e-07 $layer=licon1_PDIFF $count=1 $X=8.905
+ $Y=1.485 $X2=9.08 $Y2=2.36
r175 4 30 600 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.87 $Y2=2.32
r176 3 26 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2.3
r177 2 22 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.485 $X2=1.2 $Y2=2.3
r178 1 18 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.485 $X2=0.36 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%X 1 2 3 4 15 19 21 22 24 27 31 33 34 42
r55 40 42 7.27933 $w=6e-07 $l=3.58e-07 $layer=LI1_cond $X=1.262 $Y=1.742
+ $X2=1.62 $Y2=1.742
r56 34 40 0.244 $w=6e-07 $l=1.2e-08 $layer=LI1_cond $X=1.25 $Y=1.742 $X2=1.262
+ $Y2=1.742
r57 34 37 9.55667 $w=6e-07 $l=4.7e-07 $layer=LI1_cond $X=1.25 $Y=1.742 $X2=0.78
+ $Y2=1.742
r58 29 42 8.31678 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=1.62 $Y=2.045
+ $X2=1.62 $Y2=1.742
r59 29 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.62 $Y=2.045
+ $X2=1.62 $Y2=2.3
r60 25 33 5.55835 $w=2.42e-07 $l=4.15e-07 $layer=LI1_cond $X=1.52 $Y=0.66
+ $X2=1.105 $Y2=0.66
r61 25 27 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.52 $Y=0.66 $X2=1.52
+ $Y2=0.56
r62 24 40 4.52168 $w=3.15e-07 $l=3.02e-07 $layer=LI1_cond $X=1.262 $Y=1.44
+ $X2=1.262 $Y2=1.742
r63 23 33 5.55835 $w=2.42e-07 $l=3.3441e-07 $layer=LI1_cond $X=1.262 $Y=0.925
+ $X2=1.105 $Y2=0.66
r64 23 24 18.8415 $w=3.13e-07 $l=5.15e-07 $layer=LI1_cond $X=1.262 $Y=0.925
+ $X2=1.262 $Y2=1.44
r65 21 33 1.02508 $w=2.65e-07 $l=1.32e-07 $layer=LI1_cond $X=1.105 $Y=0.792
+ $X2=1.105 $Y2=0.66
r66 21 22 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=1.105 $Y=0.792
+ $X2=0.765 $Y2=0.792
r67 17 37 8.31678 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=0.78 $Y=2.045
+ $X2=0.78 $Y2=1.742
r68 17 19 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.78 $Y=2.045
+ $X2=0.78 $Y2=2.3
r69 13 22 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=0.68 $Y=0.66
+ $X2=0.765 $Y2=0.792
r70 13 15 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.68 $Y=0.66 $X2=0.68
+ $Y2=0.56
r71 4 42 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=1.62
r72 4 31 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=2.3
r73 3 37 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=0.645
+ $Y=1.485 $X2=0.78 $Y2=1.62
r74 3 19 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.485 $X2=0.78 $Y2=2.3
r75 2 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.56
r76 1 15 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%A_602_325# 1 2 3 4 13 18 21 23 25 27 30 32 34
+ 35 37 38 44 48
c142 34 0 1.24749e-19 $X=7.95 $Y=0.38
r143 47 48 11.956 $w=2.5e-07 $l=2.45e-07 $layer=LI1_cond $X=4.11 $Y=1.535
+ $X2=4.355 $Y2=1.535
r144 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.77 $Y=1.53
+ $X2=6.77 $Y2=1.53
r145 41 48 5.612 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=4.47 $Y=1.535
+ $X2=4.355 $Y2=1.535
r146 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.47 $Y=1.53
+ $X2=4.47 $Y2=1.53
r147 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.615 $Y=1.53
+ $X2=4.47 $Y2=1.53
r148 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.53
+ $X2=6.77 $Y2=1.53
r149 37 38 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=6.625 $Y=1.53
+ $X2=4.615 $Y2=1.53
r150 34 35 13.3743 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=7.95 $Y=0.36
+ $X2=7.705 $Y2=0.36
r151 32 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.195 $Y=0.34
+ $X2=7.705 $Y2=0.34
r152 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.11 $Y=0.425
+ $X2=7.195 $Y2=0.34
r153 29 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.11 $Y=0.425
+ $X2=7.11 $Y2=1.445
r154 28 45 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=6.83 $Y=1.53
+ $X2=6.622 $Y2=1.53
r155 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.025 $Y=1.53
+ $X2=7.11 $Y2=1.445
r156 27 28 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.025 $Y=1.53
+ $X2=6.83 $Y2=1.53
r157 23 45 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=6.622 $Y=1.615
+ $X2=6.622 $Y2=1.53
r158 23 25 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=6.622 $Y=1.615
+ $X2=6.622 $Y2=1.62
r159 19 48 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.355 $Y=1.375
+ $X2=4.355 $Y2=1.535
r160 19 21 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.355 $Y=1.375
+ $X2=4.355 $Y2=0.76
r161 17 47 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.11 $Y=1.695
+ $X2=4.11 $Y2=1.535
r162 17 18 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.11 $Y=1.695
+ $X2=4.11 $Y2=1.895
r163 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.025 $Y=1.98
+ $X2=4.11 $Y2=1.895
r164 13 15 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.025 $Y=1.98
+ $X2=3.135 $Y2=1.98
r165 4 25 300 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=2 $X=6.25
+ $Y=1.485 $X2=6.59 $Y2=1.62
r166 3 15 600 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.625 $X2=3.135 $Y2=1.98
r167 2 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.805
+ $Y=0.245 $X2=7.95 $Y2=0.38
r168 1 21 182 $w=1.7e-07 $l=6.65507e-07 $layer=licon1_NDIFF $count=1 $X=4.01
+ $Y=0.245 $X2=4.355 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%A_608_49# 1 2 3 4 13 18 19 20 22 23 24 26 28
+ 29 32 33 34 36 39 43 48 50 52 53 55
c179 55 0 1.81066e-19 $X=6.16 $Y=2.36
r180 53 54 13.934 $w=1.97e-07 $l=2.25e-07 $layer=LI1_cond $X=6.16 $Y=0.772
+ $X2=6.385 $Y2=0.772
r181 50 51 8.30177 $w=1.69e-07 $l=1.15e-07 $layer=LI1_cond $X=4.695 $Y=1.12
+ $X2=4.81 $Y2=1.12
r182 46 48 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.335 $Y=2.32
+ $X2=4.45 $Y2=2.32
r183 41 54 1.60063 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=6.385 $Y=0.655
+ $X2=6.385 $Y2=0.772
r184 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.385 $Y=0.655
+ $X2=6.385 $Y2=0.545
r185 37 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=2.36
+ $X2=6.16 $Y2=2.36
r186 37 39 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=6.245 $Y=2.36
+ $X2=8.105 $Y2=2.36
r187 36 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.16 $Y=2.275
+ $X2=6.16 $Y2=2.36
r188 35 53 1.60063 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.16 $Y=0.89
+ $X2=6.16 $Y2=0.772
r189 35 36 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=6.16 $Y=0.89
+ $X2=6.16 $Y2=2.275
r190 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=2.36
+ $X2=6.16 $Y2=2.36
r191 33 34 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.075 $Y=2.36
+ $X2=5.54 $Y2=2.36
r192 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=2.275
+ $X2=5.54 $Y2=2.36
r193 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.455 $Y=2.065
+ $X2=5.455 $Y2=2.275
r194 30 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=1.98
+ $X2=4.81 $Y2=1.98
r195 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.37 $Y=1.98
+ $X2=5.455 $Y2=2.065
r196 29 30 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.37 $Y=1.98
+ $X2=4.895 $Y2=1.98
r197 28 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=1.895
+ $X2=4.81 $Y2=1.98
r198 27 51 0.680474 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=1.205
+ $X2=4.81 $Y2=1.12
r199 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.81 $Y=1.205
+ $X2=4.81 $Y2=1.895
r200 26 50 0.680474 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=1.035
+ $X2=4.695 $Y2=1.12
r201 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.695 $Y=0.425
+ $X2=4.695 $Y2=1.035
r202 23 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.725 $Y=1.98
+ $X2=4.81 $Y2=1.98
r203 23 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.725 $Y=1.98
+ $X2=4.535 $Y2=1.98
r204 22 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=2.235
+ $X2=4.45 $Y2=2.32
r205 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=2.065
+ $X2=4.535 $Y2=1.98
r206 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.45 $Y=2.065
+ $X2=4.45 $Y2=2.235
r207 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.61 $Y=0.34
+ $X2=4.695 $Y2=0.425
r208 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.61 $Y=0.34
+ $X2=4.1 $Y2=0.34
r209 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=0.425
+ $X2=4.1 $Y2=0.34
r210 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.015 $Y=0.425
+ $X2=4.015 $Y2=0.655
r211 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.93 $Y=0.74
+ $X2=4.015 $Y2=0.655
r212 13 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.93 $Y=0.74
+ $X2=3.175 $Y2=0.74
r213 4 39 600 $w=1.7e-07 $l=8.17634e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.645 $X2=8.105 $Y2=2.36
r214 3 46 600 $w=1.7e-07 $l=8.66372e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.625 $X2=4.335 $Y2=2.32
r215 2 43 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=6.25
+ $Y=0.245 $X2=6.385 $Y2=0.545
r216 1 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.04
+ $Y=0.245 $X2=3.175 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%A_1402_49# 1 2 3 4 15 18 23 26 29 31 36
c62 29 0 1.98666e-19 $X=9.19 $Y=1.99
r63 34 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.5 $Y=0.42 $X2=9.59
+ $Y2=0.42
r64 28 29 16.3406 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=9.5 $Y=1.99 $X2=9.19
+ $Y2=1.99
r65 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.59 $Y=1.875
+ $X2=9.59 $Y2=1.99
r66 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.59 $Y=0.585
+ $X2=9.59 $Y2=0.42
r67 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=9.59 $Y=0.585
+ $X2=9.59 $Y2=1.875
r68 21 31 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=9.545 $Y=1.99
+ $X2=9.59 $Y2=1.99
r69 21 28 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=9.545 $Y=1.99
+ $X2=9.5 $Y2=1.99
r70 21 23 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=9.545 $Y=2.105
+ $X2=9.545 $Y2=2.3
r71 20 29 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=7.6 $Y=2.02
+ $X2=9.19 $Y2=2.02
r72 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.535 $Y=2.02
+ $X2=7.6 $Y2=2.02
r73 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.45 $Y=1.935
+ $X2=7.535 $Y2=2.02
r74 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=7.45 $Y=1.935
+ $X2=7.45 $Y2=0.76
r75 4 28 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=9.365
+ $Y=1.485 $X2=9.5 $Y2=1.96
r76 4 23 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.365
+ $Y=1.485 $X2=9.5 $Y2=2.3
r77 3 20 600 $w=1.7e-07 $l=8.14709e-07 $layer=licon1_PDIFF $count=1 $X=7.01
+ $Y=1.485 $X2=7.6 $Y2=2.02
r78 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.365
+ $Y=0.235 $X2=9.5 $Y2=0.42
r79 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=7.01
+ $Y=0.245 $X2=7.45 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__XOR3_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 45 47 69 70 76 79
r133 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r134 73 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r135 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r136 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r137 66 67 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r138 64 67 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.29 $Y=0 $X2=8.97
+ $Y2=0
r139 63 66 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=5.29 $Y=0 $X2=8.97
+ $Y2=0
r140 63 64 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r141 61 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r142 60 61 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r143 58 61 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=4.83 $Y2=0
r144 57 60 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.83
+ $Y2=0
r145 57 58 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r146 55 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r147 55 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r148 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r149 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r150 52 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r151 51 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r152 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r153 48 73 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r154 48 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r155 47 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r156 47 50 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r157 45 51 0.10528 $w=4.8e-07 $l=3.7e-07 $layer=MET1_cond $X=0.32 $Y=0 $X2=0.69
+ $Y2=0
r158 45 79 0.0284542 $w=4.8e-07 $l=1e-07 $layer=MET1_cond $X=0.32 $Y=0 $X2=0.22
+ $Y2=0
r159 43 66 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=8.995 $Y=0 $X2=8.97
+ $Y2=0
r160 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.995 $Y=0 $X2=9.08
+ $Y2=0
r161 42 69 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.165 $Y=0
+ $X2=9.89 $Y2=0
r162 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.165 $Y=0 $X2=9.08
+ $Y2=0
r163 40 60 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.95 $Y=0 $X2=4.83
+ $Y2=0
r164 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=0 $X2=5.035
+ $Y2=0
r165 39 63 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.12 $Y=0 $X2=5.29
+ $Y2=0
r166 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=0 $X2=5.035
+ $Y2=0
r167 37 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r168 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.94
+ $Y2=0
r169 36 57 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.07
+ $Y2=0
r170 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.94
+ $Y2=0
r171 32 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.08 $Y=0.085
+ $X2=9.08 $Y2=0
r172 32 34 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.08 $Y=0.085
+ $X2=9.08 $Y2=0.4
r173 28 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.035 $Y=0.085
+ $X2=5.035 $Y2=0
r174 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.035 $Y=0.085
+ $X2=5.035 $Y2=0.38
r175 24 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r176 24 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.36
r177 20 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r178 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r179 16 73 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r180 16 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r181 5 34 182 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=1 $X=8.905
+ $Y=0.235 $X2=9.08 $Y2=0.4
r182 4 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.235 $X2=5.035 $Y2=0.38
r183 3 26 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.36
r184 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r185 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o2111a_4.pex.spice
* Created: Thu Aug 27 14:33:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2111A_4%D1 1 3 6 8 10 14 16 17
r40 21 23 34.5433 $w=3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.255 $Y=1.16
+ $X2=0.47 $Y2=1.16
r41 16 17 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.16 $X2=0.23
+ $Y2=1.53
r42 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r43 8 23 67.48 $w=3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16 $X2=0.47
+ $Y2=1.16
r44 8 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r45 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r46 4 23 18.9685 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r47 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r48 1 23 18.9685 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%C1 1 3 6 10 14 18 19 21 22 23 30 35 41
c85 41 0 2.31747e-19 $X=2.552 $Y=1.197
c86 19 0 1.47037e-19 $X=1.31 $Y=1.16
c87 14 0 3.95163e-19 $X=2.57 $Y=1.985
r88 34 41 1.50194 $w=2.15e-07 $l=1.23e-07 $layer=LI1_cond $X=2.552 $Y=1.32
+ $X2=2.552 $Y2=1.197
r89 33 41 5.15 $w=2.44e-07 $l=1.03e-07 $layer=LI1_cond $X=2.655 $Y=1.197
+ $X2=2.552 $Y2=1.197
r90 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.16 $X2=2.655 $Y2=1.16
r91 30 32 14.2257 $w=2.88e-07 $l=8.5e-08 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.655 $Y2=1.16
r92 29 30 10.0417 $w=2.88e-07 $l=6e-08 $layer=POLY_cond $X=2.51 $Y=1.16 $X2=2.57
+ $Y2=1.16
r93 23 35 3.07165 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.552 $Y=1.575
+ $X2=2.552 $Y2=1.49
r94 23 35 1.23285 $w=2.13e-07 $l=2.3e-08 $layer=LI1_cond $X=2.552 $Y=1.467
+ $X2=2.552 $Y2=1.49
r95 23 34 7.87949 $w=2.13e-07 $l=1.47e-07 $layer=LI1_cond $X=2.552 $Y=1.467
+ $X2=2.552 $Y2=1.32
r96 22 41 1.1 $w=2.44e-07 $l=2.2e-08 $layer=LI1_cond $X=2.53 $Y=1.197 $X2=2.552
+ $Y2=1.197
r97 21 23 42.2826 $w=2.93e-07 $l=1.05e-06 $layer=LI1_cond $X=1.395 $Y=1.575
+ $X2=2.445 $Y2=1.575
r98 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.16 $X2=1.31 $Y2=1.16
r99 16 21 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=1.272 $Y=1.49
+ $X2=1.395 $Y2=1.575
r100 16 18 15.5227 $w=2.43e-07 $l=3.3e-07 $layer=LI1_cond $X=1.272 $Y=1.49
+ $X2=1.272 $Y2=1.16
r101 12 30 18.0107 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.57 $Y=1.305
+ $X2=2.57 $Y2=1.16
r102 12 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.57 $Y=1.305
+ $X2=2.57 $Y2=1.985
r103 8 29 18.0107 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.51 $Y=1.015
+ $X2=2.51 $Y2=1.16
r104 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.51 $Y=1.015
+ $X2=2.51 $Y2=0.56
r105 4 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r106 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r107 1 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r108 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%B1 3 7 11 15 17 24
c46 15 0 1.65495e-19 $X=2.15 $Y=1.985
r47 22 24 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.94 $Y=1.16
+ $X2=2.15 $Y2=1.16
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=1.16 $X2=1.94 $Y2=1.16
r49 19 22 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.94 $Y2=1.16
r50 17 23 6.115 $w=2.43e-07 $l=1.3e-07 $layer=LI1_cond $X=2.07 $Y=1.197 $X2=1.94
+ $Y2=1.197
r51 13 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r52 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r53 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r54 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r55 5 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r56 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295 $X2=1.73
+ $Y2=1.985
r57 1 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r58 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%A2 3 5 7 8 10 13 15 18 22 25 26 33 37
c84 37 0 1.69571e-19 $X=3.452 $Y=1.49
c85 33 0 1.29832e-19 $X=3.33 $Y=1.127
c86 26 0 1.75007e-19 $X=3.365 $Y=1.445
c87 25 0 5.05851e-20 $X=3.45 $Y=1.19
c88 22 0 1.11734e-19 $X=4.82 $Y=1.16
c89 3 0 6.62528e-20 $X=3.33 $Y=1.985
r90 31 33 5.00346 $w=2.89e-07 $l=3e-08 $layer=POLY_cond $X=3.3 $Y=1.127 $X2=3.33
+ $Y2=1.127
r91 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.3
+ $Y=1.16 $X2=3.3 $Y2=1.16
r92 26 37 2.72785 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.452 $Y=1.575
+ $X2=3.452 $Y2=1.49
r93 26 37 0.898515 $w=2.93e-07 $l=2.3e-08 $layer=LI1_cond $X=3.452 $Y=1.467
+ $X2=3.452 $Y2=1.49
r94 26 36 5.74268 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=3.452 $Y=1.467
+ $X2=3.452 $Y2=1.32
r95 25 36 0.100412 $w=2.43e-07 $l=2e-09 $layer=LI1_cond $X=3.45 $Y=1.197
+ $X2=3.452 $Y2=1.197
r96 25 32 7.53086 $w=2.43e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=1.197
+ $X2=3.3 $Y2=1.197
r97 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.82
+ $Y=1.16 $X2=4.82 $Y2=1.16
r98 19 22 3.76308 $w=2.43e-07 $l=8e-08 $layer=LI1_cond $X=4.74 $Y=1.197 $X2=4.82
+ $Y2=1.197
r99 17 19 2.87745 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4.74 $Y=1.32
+ $X2=4.74 $Y2=1.197
r100 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.74 $Y=1.32
+ $X2=4.74 $Y2=1.49
r101 16 26 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.6 $Y=1.575
+ $X2=3.452 $Y2=1.575
r102 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.655 $Y=1.575
+ $X2=4.74 $Y2=1.49
r103 15 16 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=4.655 $Y=1.575
+ $X2=3.6 $Y2=1.575
r104 11 23 33.6564 $w=2.93e-07 $l=1.74284e-07 $layer=POLY_cond $X=4.89 $Y=1.025
+ $X2=4.8 $Y2=1.16
r105 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.89 $Y=1.025
+ $X2=4.89 $Y2=0.56
r106 8 23 51.752 $w=2.93e-07 $l=2.94915e-07 $layer=POLY_cond $X=4.69 $Y=1.405
+ $X2=4.8 $Y2=1.16
r107 8 10 186.373 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.69 $Y=1.405
+ $X2=4.69 $Y2=1.985
r108 5 33 25.8512 $w=2.89e-07 $l=2.31892e-07 $layer=POLY_cond $X=3.485 $Y=0.96
+ $X2=3.33 $Y2=1.127
r109 5 7 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.485 $Y=0.96 $X2=3.485
+ $Y2=0.56
r110 1 33 18.0918 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=3.33 $Y=1.295
+ $X2=3.33 $Y2=1.127
r111 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.33 $Y=1.295
+ $X2=3.33 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%A1 1 3 4 6 7 9 10 12 13 20
r46 18 20 21.8328 $w=2.87e-07 $l=1.3e-07 $layer=POLY_cond $X=4.055 $Y=1.197
+ $X2=4.185 $Y2=1.197
r47 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.055
+ $Y=1.16 $X2=4.055 $Y2=1.16
r48 16 18 17.6341 $w=2.87e-07 $l=1.05e-07 $layer=POLY_cond $X=3.95 $Y=1.197
+ $X2=4.055 $Y2=1.197
r49 13 19 17.9579 $w=2.14e-07 $l=3.15e-07 $layer=LI1_cond $X=4.37 $Y=1.197
+ $X2=4.055 $Y2=1.197
r50 10 20 31.0697 $w=2.87e-07 $l=2.9011e-07 $layer=POLY_cond $X=4.37 $Y=0.985
+ $X2=4.185 $Y2=1.197
r51 10 12 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.37 $Y=0.985
+ $X2=4.37 $Y2=0.56
r52 7 20 17.9292 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=4.185 $Y=1.41
+ $X2=4.185 $Y2=1.197
r53 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.185 $Y=1.41
+ $X2=4.185 $Y2=1.985
r54 4 16 17.9292 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=3.95 $Y=0.985
+ $X2=3.95 $Y2=1.197
r55 4 6 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.95 $Y=0.985
+ $X2=3.95 $Y2=0.56
r56 1 16 32.7491 $w=2.87e-07 $l=2.94795e-07 $layer=POLY_cond $X=3.755 $Y=1.41
+ $X2=3.95 $Y2=1.197
r57 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.755 $Y=1.41
+ $X2=3.755 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%A_27_297# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 51 55 59 60 63 67 71 74 75 86 93 94 97 98 100 113
c174 86 0 6.66153e-20 $X=6.595 $Y=1.16
c175 75 0 1.45e-19 $X=5.55 $Y=1.197
c176 67 0 1.29832e-19 $X=4.775 $Y=1.917
c177 60 0 1.29227e-19 $X=1.23 $Y=1.917
c178 59 0 1.78096e-20 $X=1.795 $Y=1.917
c179 25 0 1.11734e-19 $X=5.63 $Y=1.985
r180 112 113 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=6.87 $Y=1.16
+ $X2=6.89 $Y2=1.16
r181 109 110 9.99782 $w=2.7e-07 $l=4.5e-08 $layer=POLY_cond $X=6.425 $Y=1.16
+ $X2=6.47 $Y2=1.16
r182 106 107 13.3304 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=5.99 $Y=1.16
+ $X2=6.05 $Y2=1.16
r183 96 98 10.1746 $w=6.33e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=2.147
+ $X2=3.285 $Y2=2.147
r184 96 97 15.0719 $w=6.33e-07 $l=4.25e-07 $layer=LI1_cond $X=3.12 $Y=2.147
+ $X2=2.695 $Y2=2.147
r185 87 112 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=6.595 $Y=1.16
+ $X2=6.87 $Y2=1.16
r186 87 110 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=6.595 $Y=1.16
+ $X2=6.47 $Y2=1.16
r187 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.595
+ $Y=1.16 $X2=6.595 $Y2=1.16
r188 84 109 37.7695 $w=2.7e-07 $l=1.7e-07 $layer=POLY_cond $X=6.255 $Y=1.16
+ $X2=6.425 $Y2=1.16
r189 84 107 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=6.255 $Y=1.16
+ $X2=6.05 $Y2=1.16
r190 83 86 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=6.255 $Y=1.197
+ $X2=6.595 $Y2=1.197
r191 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.255
+ $Y=1.16 $X2=6.255 $Y2=1.16
r192 81 106 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.915 $Y=1.16
+ $X2=5.99 $Y2=1.16
r193 81 104 63.3195 $w=2.7e-07 $l=2.85e-07 $layer=POLY_cond $X=5.915 $Y=1.16
+ $X2=5.63 $Y2=1.16
r194 80 83 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=5.915 $Y=1.197
+ $X2=6.255 $Y2=1.197
r195 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.915
+ $Y=1.16 $X2=5.915 $Y2=1.16
r196 78 104 12.2196 $w=2.7e-07 $l=5.5e-08 $layer=POLY_cond $X=5.575 $Y=1.16
+ $X2=5.63 $Y2=1.16
r197 78 101 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.575 $Y=1.16
+ $X2=5.485 $Y2=1.16
r198 77 80 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=5.575 $Y=1.197
+ $X2=5.915 $Y2=1.197
r199 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.575
+ $Y=1.16 $X2=5.575 $Y2=1.16
r200 75 77 1.17596 $w=2.43e-07 $l=2.5e-08 $layer=LI1_cond $X=5.55 $Y=1.197
+ $X2=5.575 $Y2=1.197
r201 73 75 7.11011 $w=2.45e-07 $l=1.5995e-07 $layer=LI1_cond $X=5.465 $Y=1.32
+ $X2=5.55 $Y2=1.197
r202 73 74 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.465 $Y=1.32
+ $X2=5.465 $Y2=1.83
r203 72 100 7.76722 $w=1.72e-07 $l=1.45997e-07 $layer=LI1_cond $X=5.065 $Y=1.915
+ $X2=4.92 $Y2=1.917
r204 71 74 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.38 $Y=1.915
+ $X2=5.465 $Y2=1.83
r205 71 72 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.38 $Y=1.915
+ $X2=5.065 $Y2=1.915
r206 67 100 7.76722 $w=1.72e-07 $l=1.45e-07 $layer=LI1_cond $X=4.775 $Y=1.917
+ $X2=4.92 $Y2=1.917
r207 67 98 94.4312 $w=1.73e-07 $l=1.49e-06 $layer=LI1_cond $X=4.775 $Y=1.917
+ $X2=3.285 $Y2=1.917
r208 66 94 6.44382 $w=1.75e-07 $l=1.15e-07 $layer=LI1_cond $X=2.025 $Y=1.917
+ $X2=1.91 $Y2=1.917
r209 66 97 42.4623 $w=1.73e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=1.917
+ $X2=2.695 $Y2=1.917
r210 61 94 0.379591 $w=2.3e-07 $l=8.8e-08 $layer=LI1_cond $X=1.91 $Y=2.005
+ $X2=1.91 $Y2=1.917
r211 61 63 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.91 $Y=2.005
+ $X2=1.91 $Y2=2.3
r212 60 93 9.06286 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=1.23 $Y=1.917
+ $X2=1.1 $Y2=1.917
r213 59 94 6.44382 $w=1.75e-07 $l=1.15e-07 $layer=LI1_cond $X=1.795 $Y=1.917
+ $X2=1.91 $Y2=1.917
r214 59 60 35.8078 $w=1.73e-07 $l=5.65e-07 $layer=LI1_cond $X=1.795 $Y=1.917
+ $X2=1.23 $Y2=1.917
r215 53 93 29.1249 $w=1.73e-07 $l=4.13e-07 $layer=LI1_cond $X=0.687 $Y=1.917
+ $X2=1.1 $Y2=1.917
r216 53 55 35.7424 $w=3.43e-07 $l=1.07e-06 $layer=LI1_cond $X=0.687 $Y=1.83
+ $X2=0.687 $Y2=0.76
r217 51 53 33.1445 $w=1.73e-07 $l=4.7e-07 $layer=LI1_cond $X=0.217 $Y=1.917
+ $X2=0.687 $Y2=1.917
r218 47 113 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.89 $Y=1.295
+ $X2=6.89 $Y2=1.16
r219 47 49 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.89 $Y=1.295
+ $X2=6.89 $Y2=1.985
r220 43 112 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.87 $Y=1.025
+ $X2=6.87 $Y2=1.16
r221 43 45 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.87 $Y=1.025
+ $X2=6.87 $Y2=0.56
r222 39 110 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.47 $Y=1.295
+ $X2=6.47 $Y2=1.16
r223 39 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.47 $Y=1.295
+ $X2=6.47 $Y2=1.985
r224 35 109 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.425 $Y=1.025
+ $X2=6.425 $Y2=1.16
r225 35 37 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.425 $Y=1.025
+ $X2=6.425 $Y2=0.56
r226 31 107 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.05 $Y=1.295
+ $X2=6.05 $Y2=1.16
r227 31 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.05 $Y=1.295
+ $X2=6.05 $Y2=1.985
r228 27 106 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.99 $Y=1.025
+ $X2=5.99 $Y2=1.16
r229 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.99 $Y=1.025
+ $X2=5.99 $Y2=0.56
r230 23 104 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.63 $Y=1.295
+ $X2=5.63 $Y2=1.16
r231 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.63 $Y=1.295
+ $X2=5.63 $Y2=1.985
r232 19 101 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.485 $Y=1.025
+ $X2=5.485 $Y2=1.16
r233 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.485 $Y=1.025
+ $X2=5.485 $Y2=0.56
r234 6 100 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.765
+ $Y=1.485 $X2=4.9 $Y2=1.96
r235 5 96 200 $w=1.7e-07 $l=6.71751e-07 $layer=licon1_PDIFF $count=3 $X=2.645
+ $Y=1.485 $X2=3.12 $Y2=1.96
r236 4 63 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.3
r237 3 93 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r238 2 51 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r239 1 55 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 51 52 54 55 56 58 70 77 82 87 93 96 99 102 106
c130 7 0 3.98522e-20 $X=6.965 $Y=1.485
r131 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r132 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r133 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r135 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 91 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r137 91 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r138 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r139 88 102 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.415 $Y=2.72
+ $X2=6.255 $Y2=2.72
r140 88 90 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.415 $Y=2.72
+ $X2=6.67 $Y2=2.72
r141 87 105 4.74443 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=7.152 $Y2=2.72
r142 87 90 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=6.67 $Y2=2.72
r143 86 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r144 86 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r145 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r146 83 99 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.585 $Y=2.72
+ $X2=5.415 $Y2=2.72
r147 83 85 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=2.72
+ $X2=5.75 $Y2=2.72
r148 82 102 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=6.255 $Y2=2.72
r149 82 85 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r150 81 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r151 81 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r152 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r153 78 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=2.72
+ $X2=3.97 $Y2=2.72
r154 78 80 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.135 $Y=2.72
+ $X2=4.37 $Y2=2.72
r155 77 99 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.245 $Y=2.72
+ $X2=5.415 $Y2=2.72
r156 77 80 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=5.245 $Y=2.72
+ $X2=4.37 $Y2=2.72
r157 76 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r158 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r159 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r160 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r161 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r162 70 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.97 $Y2=2.72
r163 70 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.45 $Y2=2.72
r164 69 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r165 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r166 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r167 66 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r168 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r169 63 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r170 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r171 58 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r172 58 60 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r173 56 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r174 56 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r175 54 68 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.07 $Y2=2.72
r176 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.36 $Y2=2.72
r177 53 72 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.53 $Y2=2.72
r178 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.36 $Y2=2.72
r179 51 65 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.4 $Y=2.72
+ $X2=1.15 $Y2=2.72
r180 51 52 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.4 $Y=2.72
+ $X2=1.512 $Y2=2.72
r181 50 68 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=2.07 $Y2=2.72
r182 50 52 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.512 $Y2=2.72
r183 46 105 2.97959 $w=3.25e-07 $l=1.05119e-07 $layer=LI1_cond $X=7.107 $Y=2.635
+ $X2=7.152 $Y2=2.72
r184 46 48 22.517 $w=3.23e-07 $l=6.35e-07 $layer=LI1_cond $X=7.107 $Y=2.635
+ $X2=7.107 $Y2=2
r185 42 102 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=2.635
+ $X2=6.255 $Y2=2.72
r186 42 44 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=6.255 $Y=2.635
+ $X2=6.255 $Y2=2
r187 38 99 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=2.635
+ $X2=5.415 $Y2=2.72
r188 38 40 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=5.415 $Y=2.635
+ $X2=5.415 $Y2=2.34
r189 34 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.72
r190 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.36
r191 30 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r192 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.36
r193 26 52 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.512 $Y=2.635
+ $X2=1.512 $Y2=2.72
r194 26 28 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=1.512 $Y=2.635
+ $X2=1.512 $Y2=2.36
r195 22 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r196 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r197 7 48 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=2
r198 6 44 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.125
+ $Y=1.485 $X2=6.26 $Y2=2
r199 5 40 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=5.295
+ $Y=1.485 $X2=5.42 $Y2=2.34
r200 4 36 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.485 $X2=3.97 $Y2=2.36
r201 3 32 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.36
r202 2 28 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.36
r203 1 24 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35 37
+ 38 39 40 41 47 48
c57 39 0 3.98522e-20 $X=7.13 $Y=0.85
r58 41 48 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=1.58 $X2=7.14
+ $Y2=1.495
r59 41 48 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.14 $Y=1.47
+ $X2=7.14 $Y2=1.495
r60 40 41 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.14 $Y=1.19
+ $X2=7.14 $Y2=1.47
r61 39 47 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=0.78 $X2=7.14
+ $Y2=0.865
r62 39 40 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.14 $Y=0.9 $X2=7.14
+ $Y2=1.19
r63 39 47 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.14 $Y=0.9 $X2=7.14
+ $Y2=0.865
r64 36 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.775 $Y=1.58
+ $X2=6.68 $Y2=1.58
r65 35 41 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.005 $Y=1.58
+ $X2=7.14 $Y2=1.58
r66 35 36 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.005 $Y=1.58
+ $X2=6.775 $Y2=1.58
r67 34 37 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.745 $Y=0.78 $X2=6.645
+ $Y2=0.78
r68 33 39 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.005 $Y=0.78
+ $X2=7.14 $Y2=0.78
r69 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.005 $Y=0.78
+ $X2=6.745 $Y2=0.78
r70 29 38 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.68 $Y=1.665
+ $X2=6.68 $Y2=1.58
r71 29 31 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=6.68 $Y=1.665
+ $X2=6.68 $Y2=1.96
r72 25 37 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=0.695
+ $X2=6.645 $Y2=0.78
r73 25 27 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=6.645 $Y=0.695
+ $X2=6.645 $Y2=0.42
r74 23 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.585 $Y=1.58
+ $X2=6.68 $Y2=1.58
r75 23 24 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.585 $Y=1.58
+ $X2=5.925 $Y2=1.58
r76 21 37 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.545 $Y=0.78 $X2=6.645
+ $Y2=0.78
r77 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.545 $Y=0.78
+ $X2=5.875 $Y2=0.78
r78 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.84 $Y=1.665
+ $X2=5.925 $Y2=1.58
r79 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.84 $Y=1.665
+ $X2=5.84 $Y2=1.96
r80 13 22 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=5.762 $Y=0.695
+ $X2=5.875 $Y2=0.78
r81 13 15 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=5.762 $Y=0.695
+ $X2=5.762 $Y2=0.42
r82 4 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.545
+ $Y=1.485 $X2=6.68 $Y2=1.96
r83 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.705
+ $Y=1.485 $X2=5.84 $Y2=1.96
r84 2 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.5
+ $Y=0.235 $X2=6.64 $Y2=0.42
r85 1 15 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.235 $X2=5.78 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%A_27_47# 1 2 3 16 19
r28 14 16 81.1721 $w=2.28e-07 $l=1.62e-06 $layer=LI1_cond $X=1.1 $Y=0.37
+ $X2=2.72 $Y2=0.37
r29 12 19 3.52738 $w=2.3e-07 $l=1.23e-07 $layer=LI1_cond $X=0.345 $Y=0.37
+ $X2=0.222 $Y2=0.37
r30 12 14 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.345 $Y=0.37
+ $X2=1.1 $Y2=0.37
r31 3 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.235 $X2=2.72 $Y2=0.38
r32 2 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r33 1 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%A_361_47# 1 2 3 10 16 18 20 22 25
r47 20 27 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=4.665 $Y=0.655
+ $X2=4.665 $Y2=0.77
r48 20 22 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=4.665 $Y=0.655
+ $X2=4.665 $Y2=0.42
r49 19 25 4.8823 $w=2.3e-07 $l=1.08e-07 $layer=LI1_cond $X=3.825 $Y=0.77
+ $X2=3.717 $Y2=0.77
r50 18 27 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=4.535 $Y=0.77
+ $X2=4.665 $Y2=0.77
r51 18 19 35.5754 $w=2.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.535 $Y=0.77
+ $X2=3.825 $Y2=0.77
r52 14 25 1.58651 $w=2.15e-07 $l=1.15e-07 $layer=LI1_cond $X=3.717 $Y=0.655
+ $X2=3.717 $Y2=0.77
r53 14 16 12.5965 $w=2.13e-07 $l=2.35e-07 $layer=LI1_cond $X=3.717 $Y=0.655
+ $X2=3.717 $Y2=0.42
r54 10 25 4.8823 $w=2.3e-07 $l=1.07e-07 $layer=LI1_cond $X=3.61 $Y=0.77
+ $X2=3.717 $Y2=0.77
r55 10 12 83.6774 $w=2.28e-07 $l=1.67e-06 $layer=LI1_cond $X=3.61 $Y=0.77
+ $X2=1.94 $Y2=0.77
r56 3 27 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.63 $Y2=0.76
r57 3 22 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.63 $Y2=0.42
r58 2 25 182 $w=1.7e-07 $l=6.08379e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.74 $Y2=0.76
r59 2 16 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.74 $Y2=0.42
r60 1 12 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_4%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 40
+ 41 43 44 45 60 64 70 74
r106 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r107 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r108 68 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r109 68 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r110 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r111 65 70 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.375 $Y=0 $X2=6.225
+ $Y2=0
r112 65 67 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.375 $Y=0 $X2=6.67
+ $Y2=0
r113 64 73 5.10352 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=7.137 $Y2=0
r114 64 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.67
+ $Y2=0
r115 63 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r116 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r117 60 70 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.075 $Y=0 $X2=6.225
+ $Y2=0
r118 60 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=5.75 $Y2=0
r119 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r120 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r121 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r122 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r123 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r124 52 53 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r125 48 52 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.99
+ $Y2=0
r126 45 53 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=2.99 $Y2=0
r127 45 48 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r128 43 58 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.035 $Y=0
+ $X2=4.83 $Y2=0
r129 43 44 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=5.035 $Y=0
+ $X2=5.167 $Y2=0
r130 42 62 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.75
+ $Y2=0
r131 42 44 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.167
+ $Y2=0
r132 40 55 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.91
+ $Y2=0
r133 40 41 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.18
+ $Y2=0
r134 39 58 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.365 $Y=0
+ $X2=4.83 $Y2=0
r135 39 41 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.365 $Y=0 $X2=4.18
+ $Y2=0
r136 37 52 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.11 $Y=0 $X2=2.99
+ $Y2=0
r137 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=0 $X2=3.275
+ $Y2=0
r138 36 55 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.91
+ $Y2=0
r139 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.275
+ $Y2=0
r140 32 73 2.91958 $w=3.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.137 $Y2=0
r141 32 34 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.095 $Y2=0.38
r142 28 70 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.225 $Y2=0
r143 28 30 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.225 $Y2=0.36
r144 24 44 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.167 $Y=0.085
+ $X2=5.167 $Y2=0
r145 24 26 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=5.167 $Y=0.085
+ $X2=5.167 $Y2=0.38
r146 20 41 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=0.085
+ $X2=4.18 $Y2=0
r147 20 22 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.18 $Y=0.085
+ $X2=4.18 $Y2=0.38
r148 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=0.085
+ $X2=3.275 $Y2=0
r149 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.275 $Y=0.085
+ $X2=3.275 $Y2=0.38
r150 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.38
r151 4 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.065
+ $Y=0.235 $X2=6.21 $Y2=0.36
r152 3 26 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.965
+ $Y=0.235 $X2=5.15 $Y2=0.38
r153 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.235 $X2=4.16 $Y2=0.38
r154 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.235 $X2=3.275 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__clkbuf_2.pex.spice
* Created: Tue Sep  1 19:00:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKBUF_2%A 3 5 7 8 9
c28 3 0 5.879e-20 $X=0.475 $Y=0.445
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.16 $X2=0.53 $Y2=1.16
r30 9 14 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.16
r31 8 14 9.92381 $w=3.58e-07 $l=3.1e-07 $layer=LI1_cond $X=0.605 $Y=0.85
+ $X2=0.605 $Y2=1.16
r32 5 13 49.3808 $w=3.11e-07 $l=2.4955e-07 $layer=POLY_cond $X=0.475 $Y=1.395
+ $X2=0.505 $Y2=1.16
r33 5 7 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.475 $Y=1.395
+ $X2=0.475 $Y2=1.985
r34 1 13 53.2554 $w=3.11e-07 $l=2.74591e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.505 $Y2=1.16
r35 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_2%A_27_47# 1 2 7 9 10 12 13 15 16 18 20 23 25
+ 29 30 35 37
c59 29 0 7.4402e-20 $X=1.05 $Y=1.16
r60 32 35 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r61 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r62 27 29 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.09 $Y=1.495
+ $X2=1.09 $Y2=1.16
r63 26 37 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.355 $Y=1.58
+ $X2=0.22 $Y2=1.58
r64 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.965 $Y=1.58
+ $X2=1.09 $Y2=1.495
r65 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.965 $Y=1.58
+ $X2=0.355 $Y2=1.58
r66 21 37 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=1.58
r67 21 23 3.41465 $w=2.68e-07 $l=8e-08 $layer=LI1_cond $X=0.22 $Y=1.665 $X2=0.22
+ $Y2=1.745
r68 20 37 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.17 $Y=1.495
+ $X2=0.22 $Y2=1.58
r69 19 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r70 19 20 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.495
r71 16 30 42.1856 $w=2.85e-07 $l=3.23381e-07 $layer=POLY_cond $X=1.37 $Y=1.395
+ $X2=1.16 $Y2=1.16
r72 16 18 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.37 $Y=1.395
+ $X2=1.37 $Y2=1.985
r73 13 30 72.6277 $w=2.85e-07 $l=5.09289e-07 $layer=POLY_cond $X=1.37 $Y=0.745
+ $X2=1.16 $Y2=1.16
r74 13 15 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.37 $Y=0.745 $X2=1.37
+ $Y2=0.445
r75 10 30 42.1856 $w=2.85e-07 $l=3.23381e-07 $layer=POLY_cond $X=0.95 $Y=1.395
+ $X2=1.16 $Y2=1.16
r76 10 12 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.95 $Y=1.395
+ $X2=0.95 $Y2=1.985
r77 7 30 72.6277 $w=2.85e-07 $l=2.1e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=1.16 $Y2=1.16
r78 7 9 96.4 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=0.95 $Y=1.16 $X2=0.95
+ $Y2=0.445
r79 2 23 300 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.745
r80 1 35 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_2%VPWR 1 2 9 11 13 15 17 22 28 32
r31 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r32 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r35 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.69 $Y2=2.72
r37 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.15 $Y2=2.72
r38 22 31 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.627 $Y2=2.72
r39 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.15 $Y2=2.72
r40 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r42 15 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r44 11 31 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.582 $Y=2.635
+ $X2=1.627 $Y2=2.72
r45 11 13 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.582 $Y=2.635
+ $X2=1.582 $Y2=2.295
r46 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.635 $X2=0.69
+ $Y2=2.72
r47 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=1.94
r48 2 13 600 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=1.485 $X2=1.58 $Y2=2.295
r49 1 9 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.94
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_2%X 1 2 9 13 15 16 17 18 28
c35 15 0 5.879e-20 $X=1.525 $Y=0.765
c36 2 0 7.4402e-20 $X=1.025 $Y=1.485
r37 26 40 25.5408 $w=1.73e-07 $l=4.03e-07 $layer=LI1_cond $X=1.555 $Y=1.942
+ $X2=1.152 $Y2=1.942
r38 25 28 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=1.555 $Y=0.825
+ $X2=1.555 $Y2=0.85
r39 18 26 3.48571 $w=1.73e-07 $l=5.5e-08 $layer=LI1_cond $X=1.61 $Y=1.942
+ $X2=1.555 $Y2=1.942
r40 18 26 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=1.555 $Y=1.82
+ $X2=1.555 $Y2=1.855
r41 17 18 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=1.555 $Y=1.53
+ $X2=1.555 $Y2=1.82
r42 16 17 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.555 $Y=1.19
+ $X2=1.555 $Y2=1.53
r43 15 25 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.61 $Y=0.74
+ $X2=1.555 $Y2=0.74
r44 15 16 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=1.555 $Y=0.88
+ $X2=1.555 $Y2=1.19
r45 15 28 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=1.555 $Y=0.88
+ $X2=1.555 $Y2=0.85
r46 11 40 0.409621 $w=1.85e-07 $l=8.8e-08 $layer=LI1_cond $X=1.152 $Y=2.03
+ $X2=1.152 $Y2=1.942
r47 11 13 14.3882 $w=1.83e-07 $l=2.4e-07 $layer=LI1_cond $X=1.152 $Y=2.03
+ $X2=1.152 $Y2=2.27
r48 7 25 26.9444 $w=1.68e-07 $l=4.13e-07 $layer=LI1_cond $X=1.142 $Y=0.74
+ $X2=1.555 $Y2=0.74
r49 7 9 12.714 $w=2.03e-07 $l=2.35e-07 $layer=LI1_cond $X=1.142 $Y=0.655
+ $X2=1.142 $Y2=0.42
r50 2 13 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.485 $X2=1.16 $Y2=2.27
r51 1 9 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.16 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_2%VGND 1 2 9 11 13 15 17 22 28 32
r30 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r31 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r32 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r33 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r34 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r35 23 28 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.692
+ $Y2=0
r36 23 25 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.15
+ $Y2=0
r37 22 31 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.627
+ $Y2=0
r38 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.15
+ $Y2=0
r39 17 28 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.692
+ $Y2=0
r40 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.23
+ $Y2=0
r41 15 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r42 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r43 11 31 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.582 $Y=0.085
+ $X2=1.627 $Y2=0
r44 11 13 10.8364 $w=3.33e-07 $l=3.15e-07 $layer=LI1_cond $X=1.582 $Y=0.085
+ $X2=1.582 $Y2=0.4
r45 7 28 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r46 7 9 13.2007 $w=2.73e-07 $l=3.15e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.4
r47 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.4
r48 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__einvn_1.spice.pex
* Created: Thu Aug 27 14:20:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVN_1%TE_B 3 5 7 9 11 13 14 15 20
c39 5 0 1.55584e-19 $X=0.47 $Y=1.41
r40 19 21 33.8755 $w=2.49e-07 $l=1.75e-07 $layer=POLY_cond $X=0.407 $Y=1.16
+ $X2=0.407 $Y2=1.335
r41 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.16 $X2=0.405 $Y2=1.16
r42 14 15 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.297 $Y=1.19
+ $X2=0.297 $Y2=1.53
r43 14 20 0.813489 $w=4.23e-07 $l=3e-08 $layer=LI1_cond $X=0.297 $Y=1.19
+ $X2=0.297 $Y2=1.16
r44 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.945 $Y=1.41
+ $X2=0.945 $Y2=1.985
r45 10 21 14.627 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=0.545 $Y=1.335
+ $X2=0.407 $Y2=1.335
r46 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.87 $Y=1.335
+ $X2=0.945 $Y2=1.41
r47 9 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.87 $Y=1.335
+ $X2=0.545 $Y2=1.335
r48 5 21 22.0795 $w=2.49e-07 $l=1.01735e-07 $layer=POLY_cond $X=0.47 $Y=1.41
+ $X2=0.407 $Y2=1.335
r49 5 7 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.47 $Y=1.41 $X2=0.47
+ $Y2=2.165
r50 1 19 39.5011 $w=2.49e-07 $l=1.93959e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.407 $Y2=1.16
r51 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_1%A_27_47# 1 2 9 12 14 17 18 19 20 24 25 27 28
+ 30
c59 28 0 1.65488e-19 $X=1.067 $Y=1.615
c60 17 0 1.55584e-19 $X=0.685 $Y=0.7
r61 27 28 16.7862 $w=1.83e-07 $l=2.8e-07 $layer=LI1_cond $X=0.777 $Y=1.895
+ $X2=0.777 $Y2=1.615
r62 25 30 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=1.387 $Y=1.16
+ $X2=1.387 $Y2=0.995
r63 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.365
+ $Y=1.16 $X2=1.365 $Y2=1.16
r64 22 28 13.9894 $w=7.63e-07 $l=3.82e-07 $layer=LI1_cond $X=1.067 $Y=1.233
+ $X2=1.067 $Y2=1.615
r65 22 24 1.14136 $w=7.63e-07 $l=7.3e-08 $layer=LI1_cond $X=1.067 $Y=1.233
+ $X2=1.067 $Y2=1.16
r66 21 24 5.86313 $w=7.63e-07 $l=3.75e-07 $layer=LI1_cond $X=1.067 $Y=0.785
+ $X2=1.067 $Y2=1.16
r67 19 27 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=0.685 $Y=1.98
+ $X2=0.777 $Y2=1.895
r68 19 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.685 $Y=1.98
+ $X2=0.37 $Y2=1.98
r69 17 21 11.2654 $w=1.7e-07 $l=4.22367e-07 $layer=LI1_cond $X=0.685 $Y=0.7
+ $X2=1.067 $Y2=0.785
r70 17 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.685 $Y=0.7
+ $X2=0.37 $Y2=0.7
r71 14 20 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.227 $Y=2.065
+ $X2=0.37 $Y2=1.98
r72 14 16 4.2807 $w=2.85e-07 $l=1e-07 $layer=LI1_cond $X=0.227 $Y=2.065
+ $X2=0.227 $Y2=2.165
r73 10 18 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.227 $Y=0.615
+ $X2=0.37 $Y2=0.7
r74 10 12 6.87422 $w=2.83e-07 $l=1.7e-07 $layer=LI1_cond $X=0.227 $Y=0.615
+ $X2=0.227 $Y2=0.445
r75 9 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.355 $Y=0.56
+ $X2=1.355 $Y2=0.995
r76 2 16 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.165
r77 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_1%A 1 3 6 8 9 10 17
r28 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.83 $Y=1.16
+ $X2=2.055 $Y2=1.16
r29 9 10 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.092 $Y=1.16
+ $X2=2.092 $Y2=1.53
r30 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.16 $X2=2.055 $Y2=1.16
r31 8 9 14.5819 $w=2.43e-07 $l=3.1e-07 $layer=LI1_cond $X=2.092 $Y=0.85
+ $X2=2.092 $Y2=1.16
r32 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.325 $X2=1.83
+ $Y2=1.985
r34 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.995 $X2=1.83
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_1%VPWR 1 6 8 10 20 21 24
r27 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r28 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 18 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r30 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 17 20 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r33 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=0.705 $Y2=2.72
r34 15 17 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.705 $Y2=2.72
r36 10 12 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r37 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r39 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r40 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.36
r41 1 6 600 $w=1.7e-07 $l=5.89597e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.705 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_1%Z 1 2 7 9 11 12
r34 32 34 5.8045 $w=6.78e-07 $l=3.3e-07 $layer=LI1_cond $X=1.71 $Y=2.125
+ $X2=2.04 $Y2=2.125
r35 22 39 4.46199 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=1.71 $Y=0.595
+ $X2=1.71 $Y2=0.425
r36 12 34 0.439735 $w=6.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.065 $Y=2.125
+ $X2=2.04 $Y2=2.125
r37 11 39 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=2.04 $Y=0.425
+ $X2=1.71 $Y2=0.425
r38 9 32 1.84689 $w=6.78e-07 $l=1.05e-07 $layer=LI1_cond $X=1.605 $Y=2.125
+ $X2=1.71 $Y2=2.125
r39 9 32 8.75737 $w=1.8e-07 $l=3.4e-07 $layer=LI1_cond $X=1.71 $Y=1.785 $X2=1.71
+ $Y2=2.125
r40 9 22 55.7784 $w=2.48e-07 $l=1.19e-06 $layer=LI1_cond $X=1.71 $Y=1.785
+ $X2=1.71 $Y2=0.595
r41 7 9 8.09112 $w=6.78e-07 $l=4.6e-07 $layer=LI1_cond $X=1.145 $Y=2.125
+ $X2=1.605 $Y2=2.125
r42 2 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=1.96
r43 1 11 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_1%VGND 1 4 13 14 19 25
r23 23 25 12.5253 $w=5.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=1.44 $Y2=0.18
r24 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r25 21 23 1.57973 $w=5.28e-07 $l=7e-08 $layer=LI1_cond $X=1.08 $Y=0.18 $X2=1.15
+ $Y2=0.18
r26 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r27 17 21 8.80133 $w=5.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.69 $Y=0.18
+ $X2=1.08 $Y2=0.18
r28 17 19 9.36586 $w=5.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=0.18
+ $X2=0.54 $Y2=0.18
r29 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r30 14 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r31 13 25 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.44
+ $Y2=0
r32 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r33 8 19 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.54
+ $Y2=0
r34 4 18 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r35 4 8 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r36 1 21 91 $w=1.7e-07 $l=5.94222e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=1.08 $Y2=0.36
.ends


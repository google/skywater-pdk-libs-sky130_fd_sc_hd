* File: sky130_fd_sc_hd__or2_0.pxi.spice
* Created: Thu Aug 27 14:42:27 2020
* 
x_PM_SKY130_FD_SC_HD__OR2_0%B N_B_c_40_n N_B_M1003_g N_B_M1005_g B N_B_c_41_n
+ N_B_c_42_n PM_SKY130_FD_SC_HD__OR2_0%B
x_PM_SKY130_FD_SC_HD__OR2_0%A N_A_M1000_g N_A_M1004_g A A N_A_c_66_n N_A_c_67_n
+ PM_SKY130_FD_SC_HD__OR2_0%A
x_PM_SKY130_FD_SC_HD__OR2_0%A_68_355# N_A_68_355#_M1003_d N_A_68_355#_M1005_s
+ N_A_68_355#_M1001_g N_A_68_355#_M1002_g N_A_68_355#_c_97_n N_A_68_355#_c_118_n
+ N_A_68_355#_c_104_n N_A_68_355#_c_98_n N_A_68_355#_c_99_n N_A_68_355#_c_100_n
+ N_A_68_355#_c_101_n PM_SKY130_FD_SC_HD__OR2_0%A_68_355#
x_PM_SKY130_FD_SC_HD__OR2_0%VPWR N_VPWR_M1004_d N_VPWR_c_161_n VPWR
+ N_VPWR_c_162_n N_VPWR_c_163_n N_VPWR_c_160_n N_VPWR_c_165_n
+ PM_SKY130_FD_SC_HD__OR2_0%VPWR
x_PM_SKY130_FD_SC_HD__OR2_0%X N_X_M1001_d N_X_M1002_d N_X_c_183_n N_X_c_185_n X
+ PM_SKY130_FD_SC_HD__OR2_0%X
x_PM_SKY130_FD_SC_HD__OR2_0%VGND N_VGND_M1003_s N_VGND_M1000_d N_VGND_c_204_n
+ N_VGND_c_205_n N_VGND_c_206_n N_VGND_c_207_n N_VGND_c_208_n VGND
+ N_VGND_c_209_n N_VGND_c_210_n PM_SKY130_FD_SC_HD__OR2_0%VGND
cc_1 VNB N_B_c_40_n 0.0194184f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.995
cc_2 VNB N_B_c_41_n 0.0158543f $X=-0.19 $Y=-0.24 $X2=0.415 $Y2=1.16
cc_3 VNB N_B_c_42_n 0.0384897f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.16
cc_4 VNB A 0.00619407f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_5 VNB N_A_c_66_n 0.0206308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_c_67_n 0.0173825f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.16
cc_7 VNB N_A_68_355#_c_97_n 0.00285007f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.16
cc_8 VNB N_A_68_355#_c_98_n 9.29659e-19 $X=-0.19 $Y=-0.24 $X2=0.415 $Y2=1.305
cc_9 VNB N_A_68_355#_c_99_n 0.0280564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_68_355#_c_100_n 0.00287913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_68_355#_c_101_n 0.0216537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_160_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_X_c_183_n 0.0205143f $X=-0.19 $Y=-0.24 $X2=0.415 $Y2=1.16
cc_14 VNB X 0.0277943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_204_n 0.0147919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_205_n 0.0332999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_206_n 0.0159217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_207_n 0.0200192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_208_n 0.00413547f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.305
cc_20 VNB N_VGND_c_209_n 0.0275441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_210_n 0.172303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_B_M1005_g 0.0401273f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.985
cc_23 VPB N_B_c_41_n 0.0218965f $X=-0.19 $Y=1.305 $X2=0.415 $Y2=1.16
cc_24 VPB N_B_c_42_n 0.0121029f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_25 VPB N_A_M1004_g 0.033464f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.985
cc_26 VPB A 0.00416763f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_27 VPB N_A_c_66_n 0.0045414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_68_355#_M1002_g 0.0440153f $X=-0.19 $Y=1.305 $X2=0.415 $Y2=1.16
cc_29 VPB N_A_68_355#_c_97_n 0.00331581f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_30 VPB N_A_68_355#_c_104_n 0.0158375f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.305
cc_31 VPB N_A_68_355#_c_98_n 0.00413395f $X=-0.19 $Y=1.305 $X2=0.415 $Y2=1.305
cc_32 VPB N_A_68_355#_c_99_n 0.00846547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_161_n 0.0114507f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.985
cc_34 VPB N_VPWR_c_162_n 0.036681f $X=-0.19 $Y=1.305 $X2=0.415 $Y2=1.16
cc_35 VPB N_VPWR_c_163_n 0.0227838f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.305
cc_36 VPB N_VPWR_c_160_n 0.0669479f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_165_n 0.00562253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_X_c_185_n 0.0212819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB X 0.0430122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 N_B_M1005_g N_A_M1004_g 0.040374f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_41 N_B_c_42_n A 5.98102e-19 $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_42 N_B_c_42_n N_A_c_66_n 0.040374f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_43 N_B_c_40_n N_A_c_67_n 0.0114906f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_44 N_B_c_40_n N_A_68_355#_c_97_n 0.00770487f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_45 N_B_M1005_g N_A_68_355#_c_97_n 0.0136145f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_46 N_B_c_41_n N_A_68_355#_c_97_n 0.0457832f $X=0.415 $Y=1.16 $X2=0 $Y2=0
cc_47 N_B_c_42_n N_A_68_355#_c_97_n 0.00965871f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_48 N_B_M1005_g N_A_68_355#_c_104_n 0.0138966f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_49 N_B_c_41_n N_A_68_355#_c_104_n 0.0200194f $X=0.415 $Y=1.16 $X2=0 $Y2=0
cc_50 N_B_c_42_n N_A_68_355#_c_104_n 0.00322375f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_51 N_B_c_40_n N_A_68_355#_c_100_n 0.00481232f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_52 N_B_M1005_g N_VPWR_c_162_n 0.0042703f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_53 N_B_M1005_g N_VPWR_c_160_n 0.00495008f $X=0.675 $Y=1.985 $X2=0 $Y2=0
cc_54 N_B_c_40_n N_VGND_c_205_n 0.00455481f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_55 N_B_c_41_n N_VGND_c_205_n 0.0203438f $X=0.415 $Y=1.16 $X2=0 $Y2=0
cc_56 N_B_c_42_n N_VGND_c_205_n 0.00552608f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_57 N_B_c_40_n N_VGND_c_207_n 0.00492879f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_58 N_B_c_40_n N_VGND_c_210_n 0.00512902f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A_M1004_g N_A_68_355#_M1002_g 0.0284977f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_60 A N_A_68_355#_c_97_n 0.0465022f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_61 N_A_c_67_n N_A_68_355#_c_97_n 0.0105666f $X=1.095 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A_M1004_g N_A_68_355#_c_118_n 0.0128723f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_63 A N_A_68_355#_c_118_n 0.0238808f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_64 N_A_c_66_n N_A_68_355#_c_118_n 3.7381e-19 $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_M1004_g N_A_68_355#_c_104_n 9.32062e-19 $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_A_68_355#_c_98_n 0.00112241f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_67 A N_A_68_355#_c_98_n 0.0429878f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_c_66_n N_A_68_355#_c_98_n 3.04326e-19 $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_69 A N_A_68_355#_c_99_n 0.00441772f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_66_n N_A_68_355#_c_99_n 0.0198385f $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_67_n N_A_68_355#_c_100_n 3.54959e-19 $X=1.095 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_c_67_n N_A_68_355#_c_101_n 0.00893741f $X=1.095 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_VPWR_c_161_n 0.00404488f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_M1004_g N_VPWR_c_162_n 0.00472107f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_VPWR_c_160_n 0.00495008f $X=1.035 $Y=1.985 $X2=0 $Y2=0
cc_76 A N_VGND_c_206_n 0.0137474f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A_c_66_n N_VGND_c_206_n 3.87822e-19 $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_c_67_n N_VGND_c_206_n 0.00395206f $X=1.095 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_c_67_n N_VGND_c_207_n 0.00510437f $X=1.095 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_c_67_n N_VGND_c_210_n 0.00512902f $X=1.095 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_68_355#_c_118_n A_150_355# 0.00353666f $X=1.525 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_82 N_A_68_355#_c_104_n A_150_355# 7.13894e-19 $X=0.84 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_68_355#_c_118_n N_VPWR_M1004_d 0.00605639f $X=1.525 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_68_355#_M1002_g N_VPWR_c_161_n 0.00968529f $X=1.52 $Y=2.095 $X2=0
+ $Y2=0
cc_85 N_A_68_355#_c_118_n N_VPWR_c_161_n 0.0195718f $X=1.525 $Y=1.87 $X2=0 $Y2=0
cc_86 N_A_68_355#_c_104_n N_VPWR_c_162_n 0.00739201f $X=0.84 $Y=1.87 $X2=0 $Y2=0
cc_87 N_A_68_355#_M1002_g N_VPWR_c_163_n 0.00412397f $X=1.52 $Y=2.095 $X2=0
+ $Y2=0
cc_88 N_A_68_355#_M1002_g N_VPWR_c_160_n 0.00446972f $X=1.52 $Y=2.095 $X2=0
+ $Y2=0
cc_89 N_A_68_355#_c_118_n N_VPWR_c_160_n 0.0179074f $X=1.525 $Y=1.87 $X2=0 $Y2=0
cc_90 N_A_68_355#_c_104_n N_VPWR_c_160_n 0.0188086f $X=0.84 $Y=1.87 $X2=0 $Y2=0
cc_91 N_A_68_355#_c_118_n N_X_M1002_d 0.00235343f $X=1.525 $Y=1.87 $X2=0 $Y2=0
cc_92 N_A_68_355#_c_98_n N_X_c_183_n 0.00817936f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_68_355#_c_99_n N_X_c_183_n 0.00382537f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_68_355#_c_101_n N_X_c_183_n 0.00401959f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_68_355#_M1002_g N_X_c_185_n 0.00649949f $X=1.52 $Y=2.095 $X2=0 $Y2=0
cc_96 N_A_68_355#_c_118_n N_X_c_185_n 0.00333158f $X=1.525 $Y=1.87 $X2=0 $Y2=0
cc_97 N_A_68_355#_M1002_g X 0.00948915f $X=1.52 $Y=2.095 $X2=0 $Y2=0
cc_98 N_A_68_355#_c_118_n X 0.0144304f $X=1.525 $Y=1.87 $X2=0 $Y2=0
cc_99 N_A_68_355#_c_98_n X 0.0610867f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_68_355#_c_99_n X 0.00826352f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_68_355#_c_101_n X 0.00478275f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_68_355#_c_100_n N_VGND_c_205_n 0.0154652f $X=0.825 $Y=0.66 $X2=0
+ $Y2=0
cc_103 N_A_68_355#_c_100_n N_VGND_c_206_n 0.0133733f $X=0.825 $Y=0.66 $X2=0
+ $Y2=0
cc_104 N_A_68_355#_c_101_n N_VGND_c_206_n 0.00333768f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_105 N_A_68_355#_c_100_n N_VGND_c_207_n 0.00934653f $X=0.825 $Y=0.66 $X2=0
+ $Y2=0
cc_106 N_A_68_355#_c_101_n N_VGND_c_209_n 0.00484683f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_107 N_A_68_355#_c_100_n N_VGND_c_210_n 0.00960978f $X=0.825 $Y=0.66 $X2=0
+ $Y2=0
cc_108 N_A_68_355#_c_101_n N_VGND_c_210_n 0.00512902f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_109 N_VPWR_c_161_n N_X_c_185_n 0.0145243f $X=1.31 $Y=2.21 $X2=0 $Y2=0
cc_110 N_VPWR_c_163_n N_X_c_185_n 0.0360862f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_111 N_VPWR_c_160_n N_X_c_185_n 0.0202188f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_112 N_VPWR_c_161_n X 4.08387e-19 $X=1.31 $Y=2.21 $X2=0 $Y2=0
cc_113 N_X_c_183_n N_VGND_c_209_n 0.0141465f $X=2.022 $Y=0.675 $X2=0 $Y2=0
cc_114 N_X_c_183_n N_VGND_c_210_n 0.0193184f $X=2.022 $Y=0.675 $X2=0 $Y2=0

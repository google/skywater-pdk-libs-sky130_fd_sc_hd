# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__mux4_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 0.995000 1.240000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.495000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.250000 1.055000 5.580000 1.675000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.800000 1.055000 5.045000 1.675000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265000 0.995000 3.565000 1.995000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 0.995000 6.345000 1.675000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315000 0.255000 9.575000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 2.800000  0.085000 3.090000 0.805000 ;
        RECT 5.150000  0.085000 5.320000 0.545000 ;
        RECT 6.010000  0.085000 6.340000 0.465000 ;
        RECT 8.895000  0.085000 9.065000 0.545000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
        RECT 9.345000 -0.085000 9.515000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.515000 2.255000 0.845000 2.635000 ;
        RECT 3.235000 2.255000 3.565000 2.635000 ;
        RECT 5.060000 2.255000 5.390000 2.635000 ;
        RECT 5.980000 2.255000 6.330000 2.635000 ;
        RECT 8.815000 2.255000 9.145000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
        RECT 9.345000 2.635000 9.515000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.260000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 1.185000 0.805000 ;
      RECT 0.175000 1.795000 1.705000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 1.015000 0.255000 2.090000 0.425000 ;
      RECT 1.015000 0.425000 1.185000 0.635000 ;
      RECT 1.015000 2.135000 1.185000 2.295000 ;
      RECT 1.015000 2.295000 2.545000 2.465000 ;
      RECT 1.410000 0.595000 1.750000 0.765000 ;
      RECT 1.410000 0.765000 1.700000 0.935000 ;
      RECT 1.410000 0.935000 1.580000 1.455000 ;
      RECT 1.410000 1.455000 2.045000 1.625000 ;
      RECT 1.535000 1.965000 1.705000 2.125000 ;
      RECT 1.875000 1.625000 2.045000 1.955000 ;
      RECT 1.875000 1.955000 2.205000 2.125000 ;
      RECT 1.920000 0.425000 2.090000 0.760000 ;
      RECT 2.080000 1.105000 2.620000 1.285000 ;
      RECT 2.260000 0.430000 2.620000 1.105000 ;
      RECT 2.260000 1.285000 2.620000 1.395000 ;
      RECT 2.260000 1.395000 3.065000 1.625000 ;
      RECT 2.375000 1.795000 2.545000 2.295000 ;
      RECT 2.715000 1.625000 3.065000 2.465000 ;
      RECT 3.380000 0.255000 4.980000 0.425000 ;
      RECT 3.380000 0.425000 3.550000 0.795000 ;
      RECT 3.720000 0.595000 4.050000 0.845000 ;
      RECT 3.735000 0.845000 4.050000 0.920000 ;
      RECT 3.735000 0.920000 3.905000 1.445000 ;
      RECT 3.735000 1.445000 4.495000 1.615000 ;
      RECT 3.825000 1.785000 3.995000 2.295000 ;
      RECT 3.825000 2.295000 4.835000 2.465000 ;
      RECT 4.075000 1.095000 4.405000 1.105000 ;
      RECT 4.075000 1.105000 4.460000 1.265000 ;
      RECT 4.165000 1.615000 4.495000 2.125000 ;
      RECT 4.220000 0.595000 4.390000 0.715000 ;
      RECT 4.220000 0.715000 5.740000 0.885000 ;
      RECT 4.220000 0.885000 4.390000 0.925000 ;
      RECT 4.290000 1.265000 4.460000 1.275000 ;
      RECT 4.625000 0.425000 4.980000 0.465000 ;
      RECT 4.665000 1.915000 5.730000 2.085000 ;
      RECT 4.665000 2.085000 4.835000 2.295000 ;
      RECT 5.495000 0.295000 5.740000 0.715000 ;
      RECT 5.560000 2.085000 5.730000 2.465000 ;
      RECT 6.500000 2.135000 6.685000 2.465000 ;
      RECT 6.510000 0.325000 6.685000 0.655000 ;
      RECT 6.515000 0.655000 6.685000 1.105000 ;
      RECT 6.515000 1.105000 6.805000 1.275000 ;
      RECT 6.515000 1.275000 6.685000 2.135000 ;
      RECT 6.980000 0.765000 7.220000 0.935000 ;
      RECT 6.980000 0.935000 7.150000 2.135000 ;
      RECT 6.980000 2.135000 7.190000 2.465000 ;
      RECT 7.030000 0.255000 7.200000 0.415000 ;
      RECT 7.030000 0.415000 7.560000 0.585000 ;
      RECT 7.360000 2.255000 7.690000 2.295000 ;
      RECT 7.360000 2.295000 8.645000 2.465000 ;
      RECT 7.390000 0.585000 7.560000 1.755000 ;
      RECT 7.390000 1.755000 8.175000 1.985000 ;
      RECT 7.730000 0.255000 8.725000 0.425000 ;
      RECT 7.730000 0.425000 7.900000 0.585000 ;
      RECT 7.845000 1.985000 8.175000 2.125000 ;
      RECT 7.970000 0.765000 8.385000 0.925000 ;
      RECT 7.970000 0.925000 8.380000 0.935000 ;
      RECT 8.190000 1.105000 8.645000 1.275000 ;
      RECT 8.210000 0.595000 8.385000 0.765000 ;
      RECT 8.475000 1.665000 9.125000 1.835000 ;
      RECT 8.475000 1.835000 8.645000 2.295000 ;
      RECT 8.555000 0.425000 8.725000 0.715000 ;
      RECT 8.555000 0.715000 9.125000 0.885000 ;
      RECT 8.955000 0.885000 9.125000 1.665000 ;
    LAYER mcon ;
      RECT 1.530000 0.765000 1.700000 0.935000 ;
      RECT 2.450000 1.105000 2.620000 1.275000 ;
      RECT 4.290000 1.105000 4.460000 1.275000 ;
      RECT 4.325000 1.785000 4.495000 1.955000 ;
      RECT 6.635000 1.105000 6.805000 1.275000 ;
      RECT 7.050000 0.765000 7.220000 0.935000 ;
      RECT 7.555000 1.785000 7.725000 1.955000 ;
      RECT 8.475000 1.105000 8.645000 1.275000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 8.200000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 2.390000 1.075000 2.680000 1.120000 ;
      RECT 2.390000 1.120000 4.520000 1.260000 ;
      RECT 2.390000 1.260000 2.680000 1.305000 ;
      RECT 4.230000 1.075000 4.520000 1.120000 ;
      RECT 4.230000 1.260000 4.520000 1.305000 ;
      RECT 4.265000 1.755000 4.555000 1.800000 ;
      RECT 4.265000 1.800000 7.785000 1.940000 ;
      RECT 4.265000 1.940000 4.555000 1.985000 ;
      RECT 6.575000 1.075000 6.865000 1.120000 ;
      RECT 6.575000 1.120000 8.705000 1.260000 ;
      RECT 6.575000 1.260000 6.865000 1.305000 ;
      RECT 6.990000 0.735000 7.280000 0.780000 ;
      RECT 6.990000 0.920000 7.280000 0.965000 ;
      RECT 7.495000 1.755000 7.785000 1.800000 ;
      RECT 7.495000 1.940000 7.785000 1.985000 ;
      RECT 7.910000 0.735000 8.200000 0.780000 ;
      RECT 7.910000 0.920000 8.200000 0.965000 ;
      RECT 8.415000 1.075000 8.705000 1.120000 ;
      RECT 8.415000 1.260000 8.705000 1.305000 ;
  END
END sky130_fd_sc_hd__mux4_1

* File: sky130_fd_sc_hd__dlygate4sd3_1.spice.SKY130_FD_SC_HD__DLYGATE4SD3_1.pxi
* Created: Thu Aug 27 14:18:52 2020
* 
x_PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A N_A_M1003_g N_A_M1001_g A A N_A_c_59_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A
x_PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_49_47# N_A_49_47#_M1003_s
+ N_A_49_47#_M1001_s N_A_49_47#_c_88_n N_A_49_47#_c_92_n N_A_49_47#_c_89_n
+ N_A_49_47#_c_90_n N_A_49_47#_c_93_n N_A_49_47#_c_94_n N_A_49_47#_c_107_n
+ N_A_49_47#_M1002_g N_A_49_47#_M1006_g
+ PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_49_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_285_47# N_A_285_47#_M1002_d
+ N_A_285_47#_M1006_d N_A_285_47#_c_146_n N_A_285_47#_M1005_g
+ N_A_285_47#_M1004_g N_A_285_47#_c_148_n N_A_285_47#_c_153_n
+ N_A_285_47#_c_149_n N_A_285_47#_c_150_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_285_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_391_47# N_A_391_47#_M1005_s
+ N_A_391_47#_M1004_s N_A_391_47#_M1000_g N_A_391_47#_M1007_g
+ N_A_391_47#_c_204_n N_A_391_47#_c_211_n N_A_391_47#_c_205_n
+ N_A_391_47#_c_206_n N_A_391_47#_c_212_n N_A_391_47#_c_213_n
+ N_A_391_47#_c_207_n N_A_391_47#_c_214_n N_A_391_47#_c_208_n
+ N_A_391_47#_c_209_n PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_391_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%VPWR N_VPWR_M1001_d N_VPWR_M1004_d
+ N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_276_n VPWR
+ N_VPWR_c_277_n N_VPWR_c_272_n N_VPWR_c_279_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%VPWR
x_PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%X N_X_M1000_d N_X_M1007_d X X X X X X X X
+ PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%X
x_PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%VGND N_VGND_M1003_d N_VGND_M1005_d
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n VGND
+ N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%VGND
cc_1 VNB N_A_M1003_g 0.0353054f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.445
cc_2 VNB A 0.0196429f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_3 VNB N_A_c_59_n 0.0279487f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_4 VNB N_A_49_47#_c_88_n 0.0186011f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_5 VNB N_A_49_47#_c_89_n 0.00890424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_49_47#_c_90_n 0.00988507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_49_47#_M1002_g 0.0920344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_285_47#_c_146_n 0.0415925f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=2.275
cc_9 VNB N_A_285_47#_M1005_g 0.0635286f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_10 VNB N_A_285_47#_c_148_n 0.00952725f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.16
cc_11 VNB N_A_285_47#_c_149_n 0.00815436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_285_47#_c_150_n 0.0011096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_391_47#_c_204_n 0.00509535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_391_47#_c_205_n 3.80283e-19 $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.335
cc_15 VNB N_A_391_47#_c_206_n 0.00376132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_391_47#_c_207_n 6.40166e-19 $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.335
cc_17 VNB N_A_391_47#_c_208_n 0.0227093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_391_47#_c_209_n 0.0193118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_272_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.0257322f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=2.275
cc_21 VNB X 0.0247986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_330_n 0.00527691f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_23 VNB N_VGND_c_331_n 0.00558565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_332_n 0.0475366f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_25 VNB N_VGND_c_333_n 0.00622287f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_26 VNB N_VGND_c_334_n 0.0189062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_335_n 0.213803f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_336_n 0.0248367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A_M1001_g 0.0597844f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=2.275
cc_30 VPB A 0.0246649f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_31 VPB N_A_c_59_n 0.00575535f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_32 VPB N_A_49_47#_c_92_n 0.0186015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_49_47#_c_93_n 0.0091095f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.16
cc_34 VPB N_A_49_47#_c_94_n 0.012349f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_35 VPB N_A_49_47#_M1002_g 0.105104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_285_47#_c_146_n 0.00996844f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=2.275
cc_37 VPB N_A_285_47#_M1004_g 0.10235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_285_47#_c_153_n 0.0103019f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.325
cc_39 VPB N_A_285_47#_c_149_n 0.0118567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_285_47#_c_150_n 0.0013759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_391_47#_M1007_g 0.0237951f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_391_47#_c_211_n 0.00509572f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=0.995
cc_43 VPB N_A_391_47#_c_212_n 0.0010446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_391_47#_c_213_n 0.00469613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_391_47#_c_214_n 0.00121303f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.335
cc_46 VPB N_A_391_47#_c_208_n 0.00475269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_273_n 0.00527691f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_48 VPB N_VPWR_c_274_n 0.00558565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_275_n 0.0475366f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_50 VPB N_VPWR_c_276_n 0.00622287f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_51 VPB N_VPWR_c_277_n 0.0189062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_272_n 0.0579295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_279_n 0.0248367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB X 0.0346962f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_55 VPB X 0.00990325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB X 0.00831449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 N_A_M1003_g N_A_49_47#_c_88_n 0.00372379f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_58 N_A_M1001_g N_A_49_47#_c_92_n 0.00372379f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_A_49_47#_c_89_n 0.0134838f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_60 A N_A_49_47#_c_89_n 0.0226442f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_61 N_A_c_59_n N_A_49_47#_c_89_n 4.78834e-19 $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_62 A N_A_49_47#_c_90_n 0.0254749f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_c_59_n N_A_49_47#_c_90_n 0.00324355f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_M1001_g N_A_49_47#_c_93_n 0.0157889f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_65 A N_A_49_47#_c_93_n 0.0231476f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_66 A N_A_49_47#_c_94_n 0.0262024f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_c_59_n N_A_49_47#_c_94_n 5.46546e-19 $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_M1003_g N_A_49_47#_c_107_n 0.0010616f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_69 N_A_M1001_g N_A_49_47#_c_107_n 0.00103729f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_70 A N_A_49_47#_c_107_n 0.045705f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A_c_59_n N_A_49_47#_c_107_n 5.61125e-19 $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_A_49_47#_M1002_g 0.0897342f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_73 A N_A_49_47#_M1002_g 0.00422688f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_M1003_g N_A_285_47#_c_148_n 6.68187e-19 $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_M1001_g N_A_285_47#_c_153_n 6.87329e-19 $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_VPWR_c_273_n 0.00306527f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_77 N_A_M1001_g N_VPWR_c_272_n 0.00688647f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_VPWR_c_279_n 0.00435702f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_79 N_A_M1003_g N_VGND_c_330_n 0.00306527f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A_M1003_g N_VGND_c_335_n 0.00688647f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_81 N_A_M1003_g N_VGND_c_336_n 0.00435702f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_49_47#_M1002_g N_A_285_47#_c_146_n 0.00601759f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_83 N_A_49_47#_c_89_n N_A_285_47#_c_148_n 0.0137617f $X=0.945 $Y=0.8 $X2=0
+ $Y2=0
cc_84 N_A_49_47#_c_107_n N_A_285_47#_c_148_n 0.0124474f $X=1.06 $Y=1.16 $X2=0
+ $Y2=0
cc_85 N_A_49_47#_M1002_g N_A_285_47#_c_148_n 0.0309284f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_86 N_A_49_47#_c_93_n N_A_285_47#_c_153_n 0.0178092f $X=0.945 $Y=1.895 $X2=0
+ $Y2=0
cc_87 N_A_49_47#_c_107_n N_A_285_47#_c_153_n 0.0124474f $X=1.06 $Y=1.16 $X2=0
+ $Y2=0
cc_88 N_A_49_47#_M1002_g N_A_285_47#_c_153_n 0.0334042f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_89 N_A_49_47#_c_107_n N_A_285_47#_c_150_n 0.0432881f $X=1.06 $Y=1.16 $X2=0
+ $Y2=0
cc_90 N_A_49_47#_M1002_g N_A_285_47#_c_150_n 0.0253227f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_91 N_A_49_47#_M1002_g N_A_391_47#_c_204_n 9.68806e-19 $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_92 N_A_49_47#_M1002_g N_A_391_47#_c_211_n 9.68806e-19 $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_93 N_A_49_47#_M1002_g N_A_391_47#_c_206_n 7.08938e-19 $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_94 N_A_49_47#_M1002_g N_A_391_47#_c_213_n 9.17449e-19 $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_95 N_A_49_47#_c_93_n N_VPWR_c_273_n 0.0166562f $X=0.945 $Y=1.895 $X2=0 $Y2=0
cc_96 N_A_49_47#_M1002_g N_VPWR_c_273_n 0.0031499f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_49_47#_c_93_n N_VPWR_c_275_n 0.00342886f $X=0.945 $Y=1.895 $X2=0 $Y2=0
cc_98 N_A_49_47#_M1002_g N_VPWR_c_275_n 0.015717f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_49_47#_M1001_s N_VPWR_c_272_n 0.00218964f $X=0.245 $Y=2.065 $X2=0
+ $Y2=0
cc_100 N_A_49_47#_c_92_n N_VPWR_c_272_n 0.0108988f $X=0.37 $Y=2.21 $X2=0 $Y2=0
cc_101 N_A_49_47#_c_93_n N_VPWR_c_272_n 0.0101892f $X=0.945 $Y=1.895 $X2=0 $Y2=0
cc_102 N_A_49_47#_M1002_g N_VPWR_c_272_n 0.0225563f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_103 N_A_49_47#_c_92_n N_VPWR_c_279_n 0.018707f $X=0.37 $Y=2.21 $X2=0 $Y2=0
cc_104 N_A_49_47#_c_93_n N_VPWR_c_279_n 0.00238773f $X=0.945 $Y=1.895 $X2=0
+ $Y2=0
cc_105 N_A_49_47#_c_89_n N_VGND_c_330_n 0.0162823f $X=0.945 $Y=0.8 $X2=0 $Y2=0
cc_106 N_A_49_47#_M1002_g N_VGND_c_330_n 0.0031499f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_107 N_A_49_47#_c_89_n N_VGND_c_332_n 0.00342446f $X=0.945 $Y=0.8 $X2=0 $Y2=0
cc_108 N_A_49_47#_M1002_g N_VGND_c_332_n 0.015717f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_49_47#_M1003_s N_VGND_c_335_n 0.00218964f $X=0.245 $Y=0.235 $X2=0
+ $Y2=0
cc_110 N_A_49_47#_c_88_n N_VGND_c_335_n 0.010877f $X=0.37 $Y=0.51 $X2=0 $Y2=0
cc_111 N_A_49_47#_c_89_n N_VGND_c_335_n 0.0101153f $X=0.945 $Y=0.8 $X2=0 $Y2=0
cc_112 N_A_49_47#_M1002_g N_VGND_c_335_n 0.0225563f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_113 N_A_49_47#_c_88_n N_VGND_c_336_n 0.0186092f $X=0.37 $Y=0.51 $X2=0 $Y2=0
cc_114 N_A_49_47#_c_89_n N_VGND_c_336_n 0.00234724f $X=0.945 $Y=0.8 $X2=0 $Y2=0
cc_115 N_A_285_47#_M1004_g N_A_391_47#_M1007_g 0.0349265f $X=2.465 $Y=2.275
+ $X2=0 $Y2=0
cc_116 N_A_285_47#_M1005_g N_A_391_47#_c_204_n 0.0044735f $X=2.465 $Y=0.445
+ $X2=0 $Y2=0
cc_117 N_A_285_47#_c_148_n N_A_391_47#_c_204_n 0.0354712f $X=1.56 $Y=0.51 $X2=0
+ $Y2=0
cc_118 N_A_285_47#_M1004_g N_A_391_47#_c_211_n 0.0044735f $X=2.465 $Y=2.275
+ $X2=0 $Y2=0
cc_119 N_A_285_47#_c_153_n N_A_391_47#_c_211_n 0.0354712f $X=1.56 $Y=2.21 $X2=0
+ $Y2=0
cc_120 N_A_285_47#_c_146_n N_A_391_47#_c_205_n 4.78834e-19 $X=2.465 $Y=0.995
+ $X2=0 $Y2=0
cc_121 N_A_285_47#_M1005_g N_A_391_47#_c_205_n 0.0289622f $X=2.465 $Y=0.445
+ $X2=0 $Y2=0
cc_122 N_A_285_47#_c_149_n N_A_391_47#_c_205_n 0.016816f $X=2.08 $Y=1.16 $X2=0
+ $Y2=0
cc_123 N_A_285_47#_c_146_n N_A_391_47#_c_206_n 0.00623751f $X=2.465 $Y=0.995
+ $X2=0 $Y2=0
cc_124 N_A_285_47#_c_148_n N_A_391_47#_c_206_n 0.0140938f $X=1.56 $Y=0.51 $X2=0
+ $Y2=0
cc_125 N_A_285_47#_c_149_n N_A_391_47#_c_206_n 0.0244854f $X=2.08 $Y=1.16 $X2=0
+ $Y2=0
cc_126 N_A_285_47#_M1004_g N_A_391_47#_c_212_n 0.0406621f $X=2.465 $Y=2.275
+ $X2=0 $Y2=0
cc_127 N_A_285_47#_c_149_n N_A_391_47#_c_212_n 0.0172142f $X=2.08 $Y=1.16 $X2=0
+ $Y2=0
cc_128 N_A_285_47#_c_146_n N_A_391_47#_c_213_n 0.00105103f $X=2.465 $Y=0.995
+ $X2=0 $Y2=0
cc_129 N_A_285_47#_c_153_n N_A_391_47#_c_213_n 0.0182391f $X=1.56 $Y=2.21 $X2=0
+ $Y2=0
cc_130 N_A_285_47#_c_149_n N_A_391_47#_c_213_n 0.0257425f $X=2.08 $Y=1.16 $X2=0
+ $Y2=0
cc_131 N_A_285_47#_c_146_n N_A_391_47#_c_207_n 0.0137387f $X=2.465 $Y=0.995
+ $X2=0 $Y2=0
cc_132 N_A_285_47#_M1005_g N_A_391_47#_c_207_n 0.0151228f $X=2.465 $Y=0.445
+ $X2=0 $Y2=0
cc_133 N_A_285_47#_c_149_n N_A_391_47#_c_207_n 0.0224245f $X=2.08 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_285_47#_M1004_g N_A_391_47#_c_214_n 0.0225833f $X=2.465 $Y=2.275
+ $X2=0 $Y2=0
cc_135 N_A_285_47#_c_149_n N_A_391_47#_c_214_n 0.0235171f $X=2.08 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_285_47#_c_146_n N_A_391_47#_c_208_n 0.0214767f $X=2.465 $Y=0.995
+ $X2=0 $Y2=0
cc_137 N_A_285_47#_M1005_g N_A_391_47#_c_209_n 0.0220837f $X=2.465 $Y=0.445
+ $X2=0 $Y2=0
cc_138 N_A_285_47#_c_153_n N_VPWR_c_273_n 0.0120708f $X=1.56 $Y=2.21 $X2=0 $Y2=0
cc_139 N_A_285_47#_M1004_g N_VPWR_c_274_n 0.00331596f $X=2.465 $Y=2.275 $X2=0
+ $Y2=0
cc_140 N_A_285_47#_M1004_g N_VPWR_c_275_n 0.0145406f $X=2.465 $Y=2.275 $X2=0
+ $Y2=0
cc_141 N_A_285_47#_c_153_n N_VPWR_c_275_n 0.0258435f $X=1.56 $Y=2.21 $X2=0 $Y2=0
cc_142 N_A_285_47#_M1006_d N_VPWR_c_272_n 0.00210122f $X=1.425 $Y=2.065 $X2=0
+ $Y2=0
cc_143 N_A_285_47#_M1004_g N_VPWR_c_272_n 0.0178211f $X=2.465 $Y=2.275 $X2=0
+ $Y2=0
cc_144 N_A_285_47#_c_153_n N_VPWR_c_272_n 0.0148749f $X=1.56 $Y=2.21 $X2=0 $Y2=0
cc_145 N_A_285_47#_c_148_n N_VGND_c_330_n 0.0120708f $X=1.56 $Y=0.51 $X2=0 $Y2=0
cc_146 N_A_285_47#_M1005_g N_VGND_c_331_n 0.00331596f $X=2.465 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_285_47#_M1005_g N_VGND_c_332_n 0.0145406f $X=2.465 $Y=0.445 $X2=0
+ $Y2=0
cc_148 N_A_285_47#_c_148_n N_VGND_c_332_n 0.0258435f $X=1.56 $Y=0.51 $X2=0 $Y2=0
cc_149 N_A_285_47#_M1002_d N_VGND_c_335_n 0.00210122f $X=1.425 $Y=0.235 $X2=0
+ $Y2=0
cc_150 N_A_285_47#_M1005_g N_VGND_c_335_n 0.0178211f $X=2.465 $Y=0.445 $X2=0
+ $Y2=0
cc_151 N_A_285_47#_c_148_n N_VGND_c_335_n 0.0148749f $X=1.56 $Y=0.51 $X2=0 $Y2=0
cc_152 N_A_391_47#_c_212_n N_VPWR_M1004_d 0.00315266f $X=2.59 $Y=1.895 $X2=0
+ $Y2=0
cc_153 N_A_391_47#_c_214_n N_VPWR_M1004_d 0.00135896f $X=2.815 $Y=1.785 $X2=0
+ $Y2=0
cc_154 N_A_391_47#_M1007_g N_VPWR_c_274_n 0.00321658f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_391_47#_c_212_n N_VPWR_c_274_n 0.0206549f $X=2.59 $Y=1.895 $X2=0
+ $Y2=0
cc_156 N_A_391_47#_c_211_n N_VPWR_c_275_n 0.0183485f $X=2.08 $Y=2.21 $X2=0 $Y2=0
cc_157 N_A_391_47#_c_212_n N_VPWR_c_275_n 0.00739553f $X=2.59 $Y=1.895 $X2=0
+ $Y2=0
cc_158 N_A_391_47#_M1007_g N_VPWR_c_277_n 0.00583607f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_391_47#_M1004_s N_VPWR_c_272_n 0.00218964f $X=1.955 $Y=2.065 $X2=0
+ $Y2=0
cc_160 N_A_391_47#_M1007_g N_VPWR_c_272_n 0.0117105f $X=3.115 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_391_47#_c_211_n N_VPWR_c_272_n 0.0107063f $X=2.08 $Y=2.21 $X2=0 $Y2=0
cc_162 N_A_391_47#_c_212_n N_VPWR_c_272_n 0.0130675f $X=2.59 $Y=1.895 $X2=0
+ $Y2=0
cc_163 N_A_391_47#_M1007_g X 0.00261074f $X=3.115 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_391_47#_c_207_n X 0.0336214f $X=2.815 $Y=1.325 $X2=0 $Y2=0
cc_165 N_A_391_47#_c_214_n X 0.00719162f $X=2.815 $Y=1.785 $X2=0 $Y2=0
cc_166 N_A_391_47#_c_208_n X 0.00762512f $X=3.06 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_391_47#_c_209_n X 0.00260914f $X=3.06 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_391_47#_c_207_n N_VGND_M1005_d 0.00256816f $X=2.815 $Y=1.325 $X2=0
+ $Y2=0
cc_169 N_A_391_47#_c_207_n N_VGND_c_331_n 0.0206549f $X=2.815 $Y=1.325 $X2=0
+ $Y2=0
cc_170 N_A_391_47#_c_208_n N_VGND_c_331_n 3.85782e-19 $X=3.06 $Y=1.16 $X2=0
+ $Y2=0
cc_171 N_A_391_47#_c_209_n N_VGND_c_331_n 0.00321658f $X=3.06 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_391_47#_c_204_n N_VGND_c_332_n 0.0182527f $X=2.08 $Y=0.51 $X2=0 $Y2=0
cc_173 N_A_391_47#_c_205_n N_VGND_c_332_n 0.00542751f $X=2.59 $Y=0.8 $X2=0 $Y2=0
cc_174 N_A_391_47#_c_207_n N_VGND_c_332_n 0.00187568f $X=2.815 $Y=1.325 $X2=0
+ $Y2=0
cc_175 N_A_391_47#_c_209_n N_VGND_c_334_n 0.00583607f $X=3.06 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_391_47#_M1005_s N_VGND_c_335_n 0.00218964f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_177 N_A_391_47#_c_204_n N_VGND_c_335_n 0.0106848f $X=2.08 $Y=0.51 $X2=0 $Y2=0
cc_178 N_A_391_47#_c_205_n N_VGND_c_335_n 0.00864014f $X=2.59 $Y=0.8 $X2=0 $Y2=0
cc_179 N_A_391_47#_c_207_n N_VGND_c_335_n 0.00432656f $X=2.815 $Y=1.325 $X2=0
+ $Y2=0
cc_180 N_A_391_47#_c_209_n N_VGND_c_335_n 0.0117105f $X=3.06 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_272_n N_X_M1007_d 0.00283025f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_182 N_VPWR_c_277_n X 0.0258765f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_183 N_VPWR_c_272_n X 0.01475f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_184 X N_VGND_c_334_n 0.0258153f $X=3.385 $Y=0.425 $X2=0 $Y2=0
cc_185 N_X_M1000_d N_VGND_c_335_n 0.00283025f $X=3.19 $Y=0.235 $X2=0 $Y2=0
cc_186 X N_VGND_c_335_n 0.0147317f $X=3.385 $Y=0.425 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o32ai_1.pxi.spice
* Created: Tue Sep  1 19:26:01 2020
* 
x_PM_SKY130_FD_SC_HD__O32AI_1%B1 N_B1_c_48_n N_B1_M1008_g N_B1_M1005_g B1 B1
+ N_B1_c_51_n PM_SKY130_FD_SC_HD__O32AI_1%B1
x_PM_SKY130_FD_SC_HD__O32AI_1%B2 N_B2_c_77_n N_B2_M1002_g N_B2_c_78_n
+ N_B2_M1009_g B2 PM_SKY130_FD_SC_HD__O32AI_1%B2
x_PM_SKY130_FD_SC_HD__O32AI_1%A3 N_A3_c_114_n N_A3_M1003_g N_A3_M1007_g A3
+ N_A3_c_116_n PM_SKY130_FD_SC_HD__O32AI_1%A3
x_PM_SKY130_FD_SC_HD__O32AI_1%A2 N_A2_M1004_g N_A2_M1001_g A2 A2 A2 A2
+ N_A2_c_152_n N_A2_c_153_n PM_SKY130_FD_SC_HD__O32AI_1%A2
x_PM_SKY130_FD_SC_HD__O32AI_1%A1 N_A1_M1006_g N_A1_M1000_g A1 N_A1_c_188_n
+ N_A1_c_189_n PM_SKY130_FD_SC_HD__O32AI_1%A1
x_PM_SKY130_FD_SC_HD__O32AI_1%VPWR N_VPWR_M1005_s N_VPWR_M1000_d N_VPWR_c_211_n
+ N_VPWR_c_212_n N_VPWR_c_213_n N_VPWR_c_214_n VPWR N_VPWR_c_215_n
+ N_VPWR_c_210_n PM_SKY130_FD_SC_HD__O32AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O32AI_1%Y N_Y_M1008_d N_Y_M1002_d N_Y_c_249_n Y Y
+ N_Y_c_260_n PM_SKY130_FD_SC_HD__O32AI_1%Y
x_PM_SKY130_FD_SC_HD__O32AI_1%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1009_d
+ N_A_27_47#_M1004_d N_A_27_47#_c_281_n N_A_27_47#_c_294_n N_A_27_47#_c_286_n
+ N_A_27_47#_c_296_n N_A_27_47#_c_291_n N_A_27_47#_c_307_p
+ PM_SKY130_FD_SC_HD__O32AI_1%A_27_47#
x_PM_SKY130_FD_SC_HD__O32AI_1%VGND N_VGND_M1003_d N_VGND_M1006_d N_VGND_c_319_n
+ N_VGND_c_320_n VGND N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n
+ N_VGND_c_324_n PM_SKY130_FD_SC_HD__O32AI_1%VGND
cc_1 VNB N_B1_c_48_n 0.0192677f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB B1 0.0124125f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB B1 0.0114803f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_B1_c_51_n 0.0346233f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_5 VNB N_B2_c_77_n 0.0257716f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B2_c_78_n 0.0173227f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_7 VNB B2 0.00294533f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_8 VNB N_A3_c_114_n 0.0196684f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_9 VNB A3 0.00255055f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_10 VNB N_A3_c_116_n 0.025377f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_11 VNB A2 0.00426905f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_12 VNB N_A2_c_152_n 0.0263868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_153_n 0.0189338f $X=-0.19 $Y=-0.24 $X2=0.217 $Y2=0.85
cc_14 VNB A1 0.0175497f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_15 VNB N_A1_c_188_n 0.0280291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_189_n 0.0213312f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_17 VNB N_VPWR_c_210_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB Y 0.00284436f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_19 VNB N_A_27_47#_c_281_n 0.0103631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_319_n 0.0121329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_320_n 0.0275124f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB N_VGND_c_321_n 0.0120821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_322_n 0.0374298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_323_n 0.0161873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_324_n 0.179907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_B1_M1005_g 0.0246012f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_27 VPB B1 0.0032255f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_28 VPB N_B1_c_51_n 0.010654f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_29 VPB N_B2_c_77_n 0.00745045f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_30 VPB N_B2_M1002_g 0.0202802f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_31 VPB B2 0.00114193f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_32 VPB N_A3_M1007_g 0.02214f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB A3 0.00253463f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_34 VPB N_A3_c_116_n 0.00690727f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_35 VPB N_A2_M1001_g 0.0202784f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB A2 0.00126071f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_37 VPB N_A2_c_152_n 0.00649864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A1_M1000_g 0.0254041f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB A1 0.00307229f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_40 VPB N_A1_c_188_n 0.00583657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_211_n 0.0102356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_212_n 0.043052f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_43 VPB N_VPWR_c_213_n 0.012107f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_44 VPB N_VPWR_c_214_n 0.0474273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_215_n 0.0604155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_210_n 0.0429311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB Y 0.00103429f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_48 N_B1_c_51_n N_B2_c_77_n 0.0520212f $X=0.47 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_49 N_B1_M1005_g N_B2_M1002_g 0.0484651f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_50 N_B1_c_48_n N_B2_c_78_n 0.0209421f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_51 N_B1_c_51_n B2 4.89155e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_52 N_B1_M1005_g N_VPWR_c_212_n 0.00463875f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_53 B1 N_VPWR_c_212_n 0.0224803f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_54 N_B1_c_51_n N_VPWR_c_212_n 0.00190713f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_55 N_B1_M1005_g N_VPWR_c_215_n 0.00562613f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_56 N_B1_M1005_g N_VPWR_c_210_n 0.0108402f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_57 N_B1_c_48_n N_Y_c_249_n 0.00394766f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_58 N_B1_c_48_n Y 0.00272122f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_59 N_B1_M1005_g Y 0.0253044f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_60 B1 Y 0.00942316f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_61 B1 Y 0.0231913f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_62 N_B1_c_51_n Y 0.00690825f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_63 B1 N_A_27_47#_M1008_s 0.00377188f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_64 N_B1_c_48_n N_A_27_47#_c_281_n 0.0133506f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_65 B1 N_A_27_47#_c_281_n 0.0170233f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_66 N_B1_c_51_n N_A_27_47#_c_281_n 8.56211e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B1_c_48_n N_A_27_47#_c_286_n 5.36508e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_68 N_B1_c_48_n N_VGND_c_322_n 0.00357877f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B1_c_48_n N_VGND_c_324_n 0.00634206f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_70 N_B2_c_78_n N_A3_c_114_n 0.0104997f $X=0.945 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_71 N_B2_M1002_g N_A3_M1007_g 0.0107268f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_72 B2 N_A3_M1007_g 9.8795e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_73 N_B2_c_77_n A3 2.86966e-19 $X=0.83 $Y=1.325 $X2=0 $Y2=0
cc_74 N_B2_M1002_g A3 5.85235e-19 $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_75 B2 A3 0.0501598f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_76 N_B2_c_77_n N_A3_c_116_n 0.0204609f $X=0.83 $Y=1.325 $X2=0 $Y2=0
cc_77 B2 N_A3_c_116_n 0.00220465f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_78 N_B2_M1002_g N_VPWR_c_215_n 0.00357877f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B2_M1002_g N_VPWR_c_210_n 0.00574497f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_80 B2 N_Y_M1002_d 0.00516282f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_81 N_B2_c_77_n N_Y_c_249_n 0.00307547f $X=0.83 $Y=1.325 $X2=0 $Y2=0
cc_82 N_B2_c_77_n Y 0.00417395f $X=0.83 $Y=1.325 $X2=0 $Y2=0
cc_83 N_B2_c_78_n Y 0.00336315f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_84 B2 Y 0.0421293f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_85 N_B2_c_77_n N_Y_c_260_n 7.98464e-19 $X=0.83 $Y=1.325 $X2=0 $Y2=0
cc_86 N_B2_M1002_g N_Y_c_260_n 0.0237178f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_87 B2 N_Y_c_260_n 0.0275775f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_88 N_B2_c_77_n N_A_27_47#_c_281_n 4.5205e-19 $X=0.83 $Y=1.325 $X2=0 $Y2=0
cc_89 N_B2_c_78_n N_A_27_47#_c_281_n 0.0109882f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_90 B2 N_A_27_47#_c_281_n 0.00452809f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_91 N_B2_c_78_n N_A_27_47#_c_286_n 0.00293147f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B2_c_77_n N_A_27_47#_c_291_n 0.00214908f $X=0.83 $Y=1.325 $X2=0 $Y2=0
cc_93 N_B2_c_78_n N_A_27_47#_c_291_n 0.001483f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_94 B2 N_A_27_47#_c_291_n 0.0171683f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B2_c_78_n N_VGND_c_322_n 0.0035787f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B2_c_78_n N_VGND_c_324_n 0.00547417f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A3_M1007_g N_A2_M1001_g 0.0251635f $X=1.59 $Y=1.985 $X2=0 $Y2=0
cc_98 A3 N_A2_M1001_g 4.96216e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_99 N_A3_M1007_g A2 0.00985913f $X=1.59 $Y=1.985 $X2=0 $Y2=0
cc_100 A3 A2 0.0365235f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A3_c_116_n A2 0.00224623f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_102 A3 N_A2_c_152_n 0.00111538f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A3_c_116_n N_A2_c_152_n 0.0130878f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A3_c_114_n N_A2_c_153_n 0.0112299f $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A3_M1007_g N_VPWR_c_215_n 0.00539883f $X=1.59 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A3_M1007_g N_VPWR_c_210_n 0.0108116f $X=1.59 $Y=1.985 $X2=0 $Y2=0
cc_107 A3 N_Y_M1002_d 0.00177033f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A3_M1007_g N_Y_c_260_n 0.0117878f $X=1.59 $Y=1.985 $X2=0 $Y2=0
cc_109 A3 N_Y_c_260_n 0.00675541f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_110 N_A3_c_116_n N_Y_c_260_n 0.00316808f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A3_c_114_n N_A_27_47#_c_294_n 0.00240691f $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A3_c_114_n N_A_27_47#_c_286_n 0.00714468f $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A3_c_114_n N_A_27_47#_c_296_n 0.0123148f $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_114 A3 N_A_27_47#_c_296_n 0.0204534f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A3_c_116_n N_A_27_47#_c_296_n 0.00451082f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A3_c_114_n N_A_27_47#_c_291_n 8.93991e-19 $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A3_c_114_n N_VGND_c_322_n 0.00420986f $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A3_c_114_n N_VGND_c_323_n 0.00596003f $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A3_c_114_n N_VGND_c_324_n 0.00654428f $X=1.405 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A2_M1001_g N_A1_M1000_g 0.0318511f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_121 A2 A1 0.014292f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A2_c_152_n A1 0.00131363f $X=2.14 $Y=1.16 $X2=0 $Y2=0
cc_123 A2 N_A1_c_188_n 0.00431955f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A2_c_152_n N_A1_c_188_n 0.0318511f $X=2.14 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A2_c_153_n N_A1_c_189_n 0.0318511f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A2_M1001_g N_VPWR_c_214_n 0.00395305f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_127 A2 N_VPWR_c_214_n 0.032307f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_128 N_A2_M1001_g N_VPWR_c_215_n 0.00480635f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_129 A2 N_VPWR_c_215_n 0.0184704f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A2_M1001_g N_VPWR_c_210_n 0.00878191f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_131 A2 N_VPWR_c_210_n 0.0109684f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A2_M1001_g N_Y_c_260_n 5.52454e-19 $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_133 A2 N_Y_c_260_n 0.0294328f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_134 A2 A_333_297# 0.0159751f $X=1.99 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_135 A2 N_A_27_47#_c_296_n 0.0209826f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A2_c_152_n N_A_27_47#_c_296_n 0.00114453f $X=2.14 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A2_c_153_n N_A_27_47#_c_296_n 0.0142853f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A2_c_153_n N_VGND_c_320_n 9.51265e-19 $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_c_153_n N_VGND_c_321_n 0.00341689f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A2_c_153_n N_VGND_c_323_n 0.00883082f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A2_c_153_n N_VGND_c_324_n 0.0040385f $X=2.14 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_VPWR_c_214_n 0.0231747f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_143 A1 N_VPWR_c_214_n 0.0346598f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A1_c_188_n N_VPWR_c_214_n 0.00401953f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A1_M1000_g N_VPWR_c_215_n 0.0046653f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1000_g N_VPWR_c_210_n 0.00799591f $X=2.65 $Y=1.985 $X2=0 $Y2=0
cc_147 A1 N_VGND_c_320_n 0.0345181f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A1_c_188_n N_VGND_c_320_n 0.00401953f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A1_c_189_n N_VGND_c_320_n 0.0125086f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A1_c_189_n N_VGND_c_321_n 0.0046653f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_189_n N_VGND_c_323_n 8.21686e-19 $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A1_c_189_n N_VGND_c_324_n 0.00799591f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_153 N_VPWR_c_210_n A_109_297# 0.00168633f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_154 N_VPWR_c_210_n N_Y_M1002_d 0.00492478f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_215_n Y 0.00983417f $X=2.695 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_c_210_n Y 0.00646331f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_215_n N_Y_c_260_n 0.0527352f $X=2.695 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_c_210_n N_Y_c_260_n 0.031551f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_159 N_VPWR_c_210_n A_333_297# 0.0131909f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_160 N_VPWR_c_210_n A_461_297# 0.0115413f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_161 A_109_297# Y 9.38831e-19 $X=0.545 $Y=1.485 $X2=0.26 $Y2=2.34
cc_162 N_Y_M1008_d N_A_27_47#_c_281_n 0.00420893f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_163 N_Y_c_249_n N_A_27_47#_c_281_n 0.0169039f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_164 N_Y_M1008_d N_VGND_c_324_n 0.00261003f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_296_n N_VGND_M1003_d 0.0203053f $X=2.355 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_27_47#_c_296_n N_VGND_c_321_n 0.00232396f $X=2.355 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_307_p N_VGND_c_321_n 0.0062327f $X=2.44 $Y=0.54 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_281_n N_VGND_c_322_n 0.0542362f $X=1.015 $Y=0.37 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_294_n N_VGND_c_322_n 0.0189339f $X=1.18 $Y=0.485 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_296_n N_VGND_c_322_n 0.00241908f $X=2.355 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_296_n N_VGND_c_323_n 0.0449411f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1008_s N_VGND_c_324_n 0.00209344f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1009_d N_VGND_c_324_n 0.00247321f $X=1.02 $Y=0.235 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_M1004_d N_VGND_c_324_n 0.00421763f $X=2.305 $Y=0.235 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_281_n N_VGND_c_324_n 0.03326f $X=1.015 $Y=0.37 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_294_n N_VGND_c_324_n 0.0124151f $X=1.18 $Y=0.485 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_296_n N_VGND_c_324_n 0.0110354f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_307_p N_VGND_c_324_n 0.00596842f $X=2.44 $Y=0.54 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a21oi_2.spice.pex
* Created: Thu Aug 27 14:01:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21OI_2%A2 1 3 7 11 14 16 19 21 22 25 29 31
c80 22 0 2.65731e-19 $X=1.77 $Y=1.16
c81 19 0 2.22276e-19 $X=1.767 $Y=1.495
r82 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.4
+ $Y=1.16 $X2=0.4 $Y2=1.16
r83 25 36 1.31569 $w=4.98e-07 $l=5.5e-08 $layer=LI1_cond $X=0.395 $Y=1.53
+ $X2=0.395 $Y2=1.585
r84 25 29 8.85098 $w=4.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.395 $Y=1.53
+ $X2=0.395 $Y2=1.16
r85 22 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.16
+ $X2=1.77 $Y2=0.995
r86 21 24 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=1.16
+ $X2=1.77 $Y2=1.245
r87 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.16 $X2=1.77 $Y2=1.16
r88 19 24 8.86495 $w=3.23e-07 $l=2.5e-07 $layer=LI1_cond $X=1.767 $Y=1.495
+ $X2=1.767 $Y2=1.245
r89 17 36 6.79934 $w=1.8e-07 $l=2.5e-07 $layer=LI1_cond $X=0.645 $Y=1.585
+ $X2=0.395 $Y2=1.585
r90 16 19 7.57412 $w=1.8e-07 $l=2.02049e-07 $layer=LI1_cond $X=1.605 $Y=1.585
+ $X2=1.767 $Y2=1.495
r91 16 17 59.1515 $w=1.78e-07 $l=9.6e-07 $layer=LI1_cond $X=1.605 $Y=1.585
+ $X2=0.645 $Y2=1.585
r92 12 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=1.16
r93 12 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=1.985
r94 11 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.71 $Y=0.56
+ $X2=1.71 $Y2=0.995
r95 5 28 35.7425 $w=3.34e-07 $l=1.85769e-07 $layer=POLY_cond $X=0.495 $Y=1.015
+ $X2=0.402 $Y2=1.16
r96 5 7 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=1.015
+ $X2=0.495 $Y2=0.56
r97 1 28 35.7425 $w=3.34e-07 $l=1.83807e-07 $layer=POLY_cond $X=0.49 $Y=1.305
+ $X2=0.402 $Y2=1.16
r98 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.49 $Y=1.305 $X2=0.49
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_2%A1 1 3 6 8 10 13 15 21 22
r51 20 22 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.29 $Y=1.16 $X2=1.35
+ $Y2=1.16
r52 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.29
+ $Y=1.16 $X2=1.29 $Y2=1.16
r53 17 20 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=1.29 $Y2=1.16
r54 15 21 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.29 $Y2=1.16
r55 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=1.16
r56 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=1.985
r57 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=1.16
r58 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=0.56
r59 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=1.16
r60 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.92 $Y=1.325 $X2=0.92
+ $Y2=1.985
r61 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=0.995
+ $X2=0.92 $Y2=1.16
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.92 $Y=0.995 $X2=0.92
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_2%B1 3 7 11 15 17 21 22 26
r47 21 22 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.937 $Y=1.16
+ $X2=2.937 $Y2=1.53
r48 21 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r49 18 20 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=2.19 $Y=1.16
+ $X2=2.61 $Y2=1.16
r50 17 26 54.8156 $w=2.9e-07 $l=2.65e-07 $layer=POLY_cond $X=2.685 $Y=1.16
+ $X2=2.95 $Y2=1.16
r51 17 20 15.5139 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=2.685 $Y=1.16
+ $X2=2.61 $Y2=1.16
r52 13 20 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.61 $Y=1.305
+ $X2=2.61 $Y2=1.16
r53 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.61 $Y=1.305
+ $X2=2.61 $Y2=1.985
r54 9 20 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.61 $Y=1.015
+ $X2=2.61 $Y2=1.16
r55 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.61 $Y=1.015
+ $X2=2.61 $Y2=0.56
r56 5 18 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.19 $Y=1.305
+ $X2=2.19 $Y2=1.16
r57 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.19 $Y=1.305 $X2=2.19
+ $Y2=1.985
r58 1 18 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.19 $Y=1.015
+ $X2=2.19 $Y2=1.16
r59 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.19 $Y=1.015
+ $X2=2.19 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_2%A_27_297# 1 2 3 4 13 15 17 21 23 25 26 27 28
+ 31 36
c57 25 0 1.34834e-19 $X=1.98 $Y=2.025
c58 23 0 1.30898e-19 $X=1.815 $Y=1.94
c59 3 0 1.08624e-19 $X=1.845 $Y=1.485
r60 29 31 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=2.937 $Y=2.285
+ $X2=2.937 $Y2=1.96
r61 27 29 7.42255 $w=1.8e-07 $l=1.91792e-07 $layer=LI1_cond $X=2.785 $Y=2.375
+ $X2=2.937 $Y2=2.285
r62 27 28 39.4343 $w=1.78e-07 $l=6.4e-07 $layer=LI1_cond $X=2.785 $Y=2.375
+ $X2=2.145 $Y2=2.375
r63 26 28 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.98 $Y=2.285
+ $X2=2.145 $Y2=2.375
r64 25 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.025 $X2=1.98
+ $Y2=1.94
r65 25 26 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.98 $Y=2.025
+ $X2=1.98 $Y2=2.285
r66 24 36 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.22 $Y=1.94
+ $X2=1.135 $Y2=1.98
r67 23 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=1.94
+ $X2=1.98 $Y2=1.94
r68 23 24 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.815 $Y=1.94
+ $X2=1.22 $Y2=1.94
r69 19 36 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.135 $Y=2.105
+ $X2=1.135 $Y2=1.98
r70 19 21 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.135 $Y=2.105
+ $X2=1.135 $Y2=2.3
r71 18 34 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=0.37 $Y=1.98 $X2=0.24
+ $Y2=1.98
r72 17 36 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=1.98 $X2=1.135
+ $Y2=1.98
r73 17 18 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.05 $Y=1.98
+ $X2=0.37 $Y2=1.98
r74 13 34 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.105
+ $X2=0.24 $Y2=1.98
r75 13 15 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=0.24 $Y=2.105
+ $X2=0.24 $Y2=2.3
r76 4 31 300 $w=1.7e-07 $l=5.80732e-07 $layer=licon1_PDIFF $count=2 $X=2.685
+ $Y=1.485 $X2=2.92 $Y2=1.96
r77 3 38 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=1.485 $X2=1.98 $Y2=2.02
r78 2 36 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.135 $Y2=1.94
r79 2 21 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.135 $Y2=2.3
r80 1 34 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.96
r81 1 15 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_2%VPWR 1 2 9 13 15 17 22 29 30 33 36
c52 2 0 1.13651e-19 $X=1.425 $Y=1.485
r53 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 30 37 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=1.56 $Y2=2.72
r58 27 29 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=0.705 $Y2=2.72
r63 23 25 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.56 $Y2=2.72
r65 22 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.705 $Y2=2.72
r67 17 19 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 11 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=2.635
+ $X2=1.56 $Y2=2.72
r71 11 13 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.56 $Y=2.635
+ $X2=1.56 $Y2=2.36
r72 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r73 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.36
r74 2 13 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.485 $X2=1.56 $Y2=2.36
r75 1 9 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.705 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_2%Y 1 2 3 12 14 15 18 22 23 26
r48 23 26 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=2.455 $Y=0.51
+ $X2=2.455 $Y2=0.42
r49 20 23 3.78145 $w=3.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.455 $Y=0.615
+ $X2=2.455 $Y2=0.51
r50 20 22 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0.615
+ $X2=2.455 $Y2=0.7
r51 16 22 3.05675 $w=3.1e-07 $l=8.9861e-08 $layer=LI1_cond $X=2.465 $Y=0.785
+ $X2=2.455 $Y2=0.7
r52 16 18 31.6922 $w=2.98e-07 $l=8.25e-07 $layer=LI1_cond $X=2.465 $Y=0.785
+ $X2=2.465 $Y2=1.61
r53 14 22 3.57226 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.295 $Y=0.7
+ $X2=2.455 $Y2=0.7
r54 14 15 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=2.295 $Y=0.7
+ $X2=1.3 $Y2=0.7
r55 10 15 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=1.127 $Y=0.615
+ $X2=1.3 $Y2=0.7
r56 10 12 8.51806 $w=3.43e-07 $l=2.55e-07 $layer=LI1_cond $X=1.127 $Y=0.615
+ $X2=1.127 $Y2=0.36
r57 3 18 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.485 $X2=2.4 $Y2=1.61
r58 2 26 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.42
r59 2 22 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.76
r60 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.235 $X2=1.135 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21OI_2%VGND 1 2 3 10 12 16 18 20 23 24 25 34 43
r47 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r48 37 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r49 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 34 42 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.007
+ $Y2=0
r51 34 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.53
+ $Y2=0
r52 33 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r53 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r54 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r55 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r56 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 27 39 4.4461 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r58 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r59 25 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r60 25 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r61 23 32 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.76 $Y=0 $X2=1.61
+ $Y2=0
r62 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.76 $Y=0 $X2=1.925
+ $Y2=0
r63 22 36 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.53
+ $Y2=0
r64 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.925
+ $Y2=0
r65 18 42 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=3.007 $Y2=0
r66 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=2.96 $Y2=0.38
r67 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.925 $Y=0.085
+ $X2=1.925 $Y2=0
r68 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.925 $Y=0.085
+ $X2=1.925 $Y2=0.36
r69 10 39 3.03143 $w=2.95e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.247 $Y=0.085
+ $X2=0.197 $Y2=0
r70 10 12 10.7431 $w=2.93e-07 $l=2.75e-07 $layer=LI1_cond $X=0.247 $Y=0.085
+ $X2=0.247 $Y2=0.36
r71 3 20 91 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=2 $X=2.685
+ $Y=0.235 $X2=2.96 $Y2=0.38
r72 2 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.235 $X2=1.925 $Y2=0.36
r73 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends


* NGSPICE file created from sky130_fd_sc_hd__dlrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=1.0568e+12p ps=9.48e+06u
M1001 a_664_425# a_193_47# a_560_425# VPB phighvt w=360000u l=150000u
+  ad=1.644e+11p pd=1.67e+06u as=1.332e+11p ps=1.46e+06u
M1002 a_711_21# a_560_425# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.3e+11p pd=2.66e+06u as=0p ps=0u
M1003 VGND D a_299_47# VNB nshort w=420000u l=150000u
+  ad=5.375e+11p pd=6.04e+06u as=1.092e+11p ps=1.36e+06u
M1004 a_560_425# a_27_47# a_465_369# VPB phighvt w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1005 a_929_47# a_560_425# a_711_21# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=1.69e+11p ps=1.82e+06u
M1006 a_465_47# a_299_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
M1007 a_560_425# a_193_47# a_465_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1008 VGND RESET_B a_929_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR GATE a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1010 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1011 Q a_711_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1012 a_465_369# a_299_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR RESET_B a_711_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR D a_299_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1015 a_654_47# a_27_47# a_560_425# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1016 VGND a_711_21# a_654_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q a_711_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1018 VPWR a_711_21# a_664_425# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND GATE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends


* File: sky130_fd_sc_hd__a2111oi_2.spice.pex
* Created: Thu Aug 27 13:59:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2111OI_2%C1 1 3 6 10 14 17 20 25 26 28 34 37 39 42
c84 37 0 1.9492e-19 $X=1.81 $Y=0.995
c85 28 0 1.67185e-19 $X=1.525 $Y=1.445
c86 26 0 1.44232e-19 $X=1.78 $Y=1.16
c87 10 0 1.65935e-19 $X=1.79 $Y=1.985
r88 39 42 0.245201 $w=2.33e-07 $l=5e-09 $layer=LI1_cond $X=1.615 $Y=1.562
+ $X2=1.61 $Y2=1.562
r89 28 39 3.0562 $w=2.35e-07 $l=9.2e-08 $layer=LI1_cond $X=1.707 $Y=1.562
+ $X2=1.615 $Y2=1.562
r90 28 42 1.96161 $w=2.33e-07 $l=4e-08 $layer=LI1_cond $X=1.57 $Y=1.562 $X2=1.61
+ $Y2=1.562
r91 26 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.16
+ $X2=1.81 $Y2=1.325
r92 26 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.16
+ $X2=1.81 $Y2=0.995
r93 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=1.16 $X2=1.78 $Y2=1.16
r94 22 28 8.45579 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=1.707 $Y=1.275
+ $X2=1.707 $Y2=1.445
r95 21 25 3.43381 $w=2.43e-07 $l=7.3e-08 $layer=LI1_cond $X=1.707 $Y=1.152
+ $X2=1.78 $Y2=1.152
r96 21 22 2.40932 $w=1.85e-07 $l=1.23e-07 $layer=LI1_cond $X=1.707 $Y=1.152
+ $X2=1.707 $Y2=1.275
r97 20 28 54.6797 $w=2.33e-07 $l=1.115e-06 $layer=LI1_cond $X=0.455 $Y=1.562
+ $X2=1.57 $Y2=1.562
r98 18 34 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.29 $Y=1.16 $X2=0.5
+ $Y2=1.16
r99 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.16 $X2=0.29 $Y2=1.16
r100 15 20 7.07017 $w=2.35e-07 $l=2.15708e-07 $layer=LI1_cond $X=0.29 $Y=1.445
+ $X2=0.455 $Y2=1.562
r101 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.29 $Y=1.445
+ $X2=0.29 $Y2=1.16
r102 14 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.56 $X2=1.9
+ $Y2=0.995
r103 10 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.79 $Y=1.985
+ $X2=1.79 $Y2=1.325
r104 4 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.325
+ $X2=0.5 $Y2=1.16
r105 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.5 $Y=1.325 $X2=0.5
+ $Y2=1.985
r106 1 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=0.995
+ $X2=0.5 $Y2=1.16
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.5 $Y=0.995 $X2=0.5
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%D1 1 3 6 8 10 13 15 21 22
r51 20 22 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.26 $Y=1.16 $X2=1.36
+ $Y2=1.16
r52 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.26
+ $Y=1.16 $X2=1.26 $Y2=1.16
r53 17 20 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=1.26 $Y2=1.16
r54 15 21 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=1.15 $Y=1.175 $X2=1.26
+ $Y2=1.175
r55 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.16
r56 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.985
r57 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=0.995
+ $X2=1.36 $Y2=1.16
r58 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.36 $Y=0.995
+ $X2=1.36 $Y2=0.56
r59 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.16
r60 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.93 $Y=1.325 $X2=0.93
+ $Y2=1.985
r61 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.16
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.93 $Y=0.995 $X2=0.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%B1 3 5 7 10 12 14 15 22 23
c49 3 0 1.67185e-19 $X=2.26 $Y=1.985
r50 21 23 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.915 $Y2=1.16
r51 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.69
+ $Y=1.16 $X2=2.69 $Y2=1.16
r52 19 21 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.375 $Y=1.16
+ $X2=2.69 $Y2=1.16
r53 17 19 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.375 $Y2=1.16
r54 15 22 0.535558 $w=6.68e-07 $l=3e-08 $layer=LI1_cond $X=2.52 $Y=1.19 $X2=2.52
+ $Y2=1.16
r55 12 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.995
+ $X2=2.915 $Y2=1.16
r56 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.915 $Y=0.995
+ $X2=2.915 $Y2=0.56
r57 8 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.16
r58 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.985
r59 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=0.995
+ $X2=2.375 $Y2=1.16
r60 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.375 $Y=0.995
+ $X2=2.375 $Y2=0.56
r61 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.325
+ $X2=2.26 $Y2=1.16
r62 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.26 $Y=1.325 $X2=2.26
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%A1 1 3 6 10 13 17 22 23 25 26 27 32 35
r75 26 27 49.3546 $w=2.28e-07 $l=9.85e-07 $layer=LI1_cond $X=4.895 $Y=1.56
+ $X2=3.91 $Y2=1.56
r76 25 27 9.77071 $w=2.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.715 $Y=1.56
+ $X2=3.91 $Y2=1.56
r77 23 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=1.16
+ $X2=5.06 $Y2=1.325
r78 23 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=1.16
+ $X2=5.06 $Y2=0.995
r79 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.06
+ $Y=1.16 $X2=5.06 $Y2=1.16
r80 20 26 7.45331 $w=2.3e-07 $l=2.47919e-07 $layer=LI1_cond $X=5.092 $Y=1.445
+ $X2=4.895 $Y2=1.56
r81 20 22 8.31509 $w=3.93e-07 $l=2.85e-07 $layer=LI1_cond $X=5.092 $Y=1.445
+ $X2=5.092 $Y2=1.16
r82 18 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.55 $Y=1.16 $X2=3.64
+ $Y2=1.16
r83 18 29 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.55 $Y=1.16
+ $X2=3.345 $Y2=1.16
r84 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.16 $X2=3.55 $Y2=1.16
r85 15 25 6.8319 $w=2.3e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.59 $Y=1.445
+ $X2=3.715 $Y2=1.56
r86 15 17 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=3.59 $Y=1.445
+ $X2=3.59 $Y2=1.16
r87 13 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.97 $Y=1.985
+ $X2=4.97 $Y2=1.325
r88 10 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.97 $Y=0.56
+ $X2=4.97 $Y2=0.995
r89 4 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.325
+ $X2=3.64 $Y2=1.16
r90 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.64 $Y=1.325 $X2=3.64
+ $Y2=1.985
r91 1 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=0.995
+ $X2=3.345 $Y2=1.16
r92 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.345 $Y=0.995
+ $X2=3.345 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%A2 1 3 6 10 12 14 15 23
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=1.16 $X2=4.52 $Y2=1.16
r46 20 22 3.44503 $w=3.35e-07 $l=2e-08 $layer=POLY_cond $X=4.5 $Y=1.157 $X2=4.52
+ $Y2=1.157
r47 19 20 74.0681 $w=3.35e-07 $l=4.3e-07 $layer=POLY_cond $X=4.07 $Y=1.157
+ $X2=4.5 $Y2=1.157
r48 15 23 0.475263 $w=7.53e-07 $l=3e-08 $layer=LI1_cond $X=4.347 $Y=1.19
+ $X2=4.347 $Y2=1.16
r49 12 22 3.44503 $w=3.35e-07 $l=2e-08 $layer=POLY_cond $X=4.54 $Y=1.157
+ $X2=4.52 $Y2=1.157
r50 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.54 $Y=0.99
+ $X2=4.54 $Y2=0.56
r51 8 20 21.5811 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=4.5 $Y=1.325 $X2=4.5
+ $Y2=1.157
r52 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.5 $Y=1.325 $X2=4.5
+ $Y2=1.985
r53 4 19 21.5811 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=4.07 $Y=1.325
+ $X2=4.07 $Y2=1.157
r54 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.07 $Y=1.325 $X2=4.07
+ $Y2=1.985
r55 1 19 4.30629 $w=3.35e-07 $l=2.5e-08 $layer=POLY_cond $X=4.045 $Y=1.157
+ $X2=4.07 $Y2=1.157
r56 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.045 $Y=0.99
+ $X2=4.045 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%A_28_297# 1 2 3 12 14 15 18 22
r40 18 22 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.815 $Y=2.38
+ $X2=2.9 $Y2=2.3
r41 18 20 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.815 $Y=2.38
+ $X2=2.185 $Y2=2.38
r42 15 17 90.1866 $w=1.88e-07 $l=1.545e-06 $layer=LI1_cond $X=0.46 $Y=2.37
+ $X2=2.005 $Y2=2.37
r43 14 20 5.69365 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=2.09 $Y=2.37
+ $X2=2.185 $Y2=2.37
r44 14 17 4.96172 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=2.37
+ $X2=2.005 $Y2=2.37
r45 10 15 7.69972 $w=1.9e-07 $l=2.22486e-07 $layer=LI1_cond $X=0.28 $Y=2.275
+ $X2=0.46 $Y2=2.37
r46 10 12 8.16314 $w=3.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.28 $Y=2.275
+ $X2=0.28 $Y2=2.02
r47 3 22 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.485 $X2=2.9 $Y2=2.3
r48 2 17 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.485 $X2=2.005 $Y2=2.36
r49 1 12 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.485 $X2=0.285 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%Y 1 2 3 4 5 6 19 21 23 25 31 33 37 40 41
+ 45 47 52 54 55 57 59 63 67 70
c131 55 0 1.44232e-19 $X=2.14 $Y=1.535
c132 54 0 1.9492e-19 $X=2.13 $Y=0.74
r133 67 70 2.15657 $w=1.78e-07 $l=3.5e-08 $layer=LI1_cond $X=3.025 $Y=1.535
+ $X2=2.99 $Y2=1.535
r134 63 67 3.89832 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=3.14 $Y=1.535
+ $X2=3.025 $Y2=1.535
r135 63 70 1.5404 $w=1.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.965 $Y=1.535
+ $X2=2.99 $Y2=1.535
r136 56 63 25.0968 $w=2.78e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=0.845
+ $X2=3.14 $Y2=1.445
r137 56 57 2.22146 $w=2.3e-07 $l=3.05205e-07 $layer=LI1_cond $X=3.14 $Y=0.845
+ $X2=2.965 $Y2=0.615
r138 55 63 50.8333 $w=1.78e-07 $l=8.25e-07 $layer=LI1_cond $X=2.14 $Y=1.535
+ $X2=2.965 $Y2=1.535
r139 48 57 3.9698 $w=1.9e-07 $l=3.745e-07 $layer=LI1_cond $X=3.295 $Y=0.71
+ $X2=2.965 $Y2=0.615
r140 47 59 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=5.187 $Y=0.71
+ $X2=5.187 $Y2=0.38
r141 47 48 100.694 $w=1.88e-07 $l=1.725e-06 $layer=LI1_cond $X=5.02 $Y=0.71
+ $X2=3.295 $Y2=0.71
r142 43 57 2.22146 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=0.615
+ $X2=2.965 $Y2=0.615
r143 43 45 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.13 $Y=0.615
+ $X2=3.13 $Y2=0.375
r144 42 54 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0.73
+ $X2=2.13 $Y2=0.73
r145 41 57 3.9698 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=2.965 $Y=0.73
+ $X2=2.965 $Y2=0.615
r146 41 42 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.965 $Y=0.73
+ $X2=2.295 $Y2=0.73
r147 39 55 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.055 $Y=1.625
+ $X2=2.14 $Y2=1.535
r148 39 40 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.055 $Y=1.625
+ $X2=2.055 $Y2=1.85
r149 35 54 0.0811015 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=2.13 $Y=0.615
+ $X2=2.13 $Y2=0.73
r150 35 37 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.13 $Y=0.615
+ $X2=2.13 $Y2=0.4
r151 34 52 5.44316 $w=2.3e-07 $l=1.23e-07 $layer=LI1_cond $X=1.295 $Y=0.73
+ $X2=1.172 $Y2=0.73
r152 33 54 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=0.73
+ $X2=2.13 $Y2=0.73
r153 33 34 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.965 $Y=0.73
+ $X2=1.295 $Y2=0.73
r154 29 52 1.11607 $w=2.45e-07 $l=1.15e-07 $layer=LI1_cond $X=1.172 $Y=0.615
+ $X2=1.172 $Y2=0.73
r155 29 31 9.17251 $w=2.43e-07 $l=1.95e-07 $layer=LI1_cond $X=1.172 $Y=0.615
+ $X2=1.172 $Y2=0.42
r156 25 40 7.17723 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.97 $Y=1.977
+ $X2=2.055 $Y2=1.85
r157 25 27 37.2849 $w=2.53e-07 $l=8.25e-07 $layer=LI1_cond $X=1.97 $Y=1.977
+ $X2=1.145 $Y2=1.977
r158 24 50 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=0.38 $Y=0.73
+ $X2=0.25 $Y2=0.73
r159 23 52 5.44316 $w=2.3e-07 $l=1.22e-07 $layer=LI1_cond $X=1.05 $Y=0.73
+ $X2=1.172 $Y2=0.73
r160 23 24 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.05 $Y=0.73
+ $X2=0.38 $Y2=0.73
r161 19 50 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=0.25 $Y=0.615
+ $X2=0.25 $Y2=0.73
r162 19 21 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=0.25 $Y=0.615
+ $X2=0.25 $Y2=0.42
r163 6 27 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.485 $X2=1.145 $Y2=1.98
r164 5 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.045
+ $Y=0.235 $X2=5.185 $Y2=0.38
r165 4 45 91 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=2 $X=2.99
+ $Y=0.235 $X2=3.13 $Y2=0.375
r166 3 54 182 $w=1.7e-07 $l=5.77321e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.13 $Y2=0.74
r167 3 37 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.13 $Y2=0.4
r168 2 52 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.145 $Y2=0.76
r169 2 31 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.145 $Y2=0.42
r170 1 50 182 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.285 $Y2=0.76
r171 1 21 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.285 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%A_467_297# 1 2 3 4 13 17 19 23 25 27 29 31
+ 37 39
c58 31 0 1.65935e-19 $X=2.475 $Y=1.88
r59 31 34 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.475 $Y=1.88
+ $X2=2.475 $Y2=1.975
r60 27 41 3.0592 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=5.235 $Y=2.105
+ $X2=5.235 $Y2=1.975
r61 27 29 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.235 $Y=2.105
+ $X2=5.235 $Y2=2.36
r62 26 39 4.38255 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=4.4 $Y=1.975
+ $X2=4.295 $Y2=1.975
r63 25 41 3.88283 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=1.975
+ $X2=5.235 $Y2=1.975
r64 25 26 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=5.07 $Y=1.975
+ $X2=4.4 $Y2=1.975
r65 21 39 2.05017 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=4.295 $Y=2.105
+ $X2=4.295 $Y2=1.975
r66 21 23 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=4.295 $Y=2.105
+ $X2=4.295 $Y2=2.3
r67 20 37 7.95815 $w=2.1e-07 $l=4.43959e-07 $layer=LI1_cond $X=3.52 $Y=1.97
+ $X2=3.155 $Y2=1.795
r68 19 39 4.38255 $w=2.55e-07 $l=1.07471e-07 $layer=LI1_cond $X=4.19 $Y=1.97
+ $X2=4.295 $Y2=1.975
r69 19 20 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=4.19 $Y=1.97
+ $X2=3.52 $Y2=1.97
r70 15 37 0.549021 $w=3.65e-07 $l=3.80263e-07 $layer=LI1_cond $X=3.337 $Y=2.095
+ $X2=3.155 $Y2=1.795
r71 15 17 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=3.337 $Y=2.095
+ $X2=3.337 $Y2=2.3
r72 14 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=1.88
+ $X2=2.475 $Y2=1.88
r73 13 37 7.95815 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=1.88
+ $X2=3.155 $Y2=1.795
r74 13 14 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=3.155 $Y=1.88
+ $X2=2.64 $Y2=1.88
r75 4 41 600 $w=1.7e-07 $l=6.22796e-07 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=1.485 $X2=5.235 $Y2=2.02
r76 4 29 600 $w=1.7e-07 $l=9.65337e-07 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=1.485 $X2=5.235 $Y2=2.36
r77 3 39 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=1.485 $X2=4.285 $Y2=1.96
r78 3 23 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=1.485 $X2=4.285 $Y2=2.3
r79 2 37 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.485 $X2=3.43 $Y2=1.96
r80 2 17 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.485 $X2=3.43 $Y2=2.3
r81 1 34 600 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.475 $Y2=1.975
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r71 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r72 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r73 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r74 31 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r76 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=2.72
+ $X2=3.855 $Y2=2.72
r77 28 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.02 $Y=2.72
+ $X2=4.37 $Y2=2.72
r78 27 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 26 27 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r80 22 26 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=2.72
+ $X2=3.855 $Y2=2.72
r82 20 26 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.69 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 18 27 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.45 $Y2=2.72
r84 18 22 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 16 30 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.57 $Y=2.72 $X2=4.37
+ $Y2=2.72
r86 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.57 $Y=2.72
+ $X2=4.735 $Y2=2.72
r87 15 33 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.9 $Y=2.72 $X2=5.29
+ $Y2=2.72
r88 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=2.72
+ $X2=4.735 $Y2=2.72
r89 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.735 $Y=2.635
+ $X2=4.735 $Y2=2.72
r90 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.735 $Y=2.635
+ $X2=4.735 $Y2=2.36
r91 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=2.635
+ $X2=3.855 $Y2=2.72
r92 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.855 $Y=2.635
+ $X2=3.855 $Y2=2.36
r93 2 13 600 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=4.575
+ $Y=1.485 $X2=4.735 $Y2=2.36
r94 1 9 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=1.485 $X2=3.855 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_2%VGND 1 2 3 4 15 19 21 25 29 31 33 38 43 53
+ 54 57 60 63 66
r80 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r81 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r82 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r83 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r84 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r85 54 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r86 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r87 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.29
+ $Y2=0
r88 51 53 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=5.29
+ $Y2=0
r89 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r90 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r91 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r92 47 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r93 46 49 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r94 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r95 44 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.63
+ $Y2=0
r96 44 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.99
+ $Y2=0
r97 43 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.29
+ $Y2=0
r98 43 49 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.125 $Y=0 $X2=3.91
+ $Y2=0
r99 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r100 42 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r101 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r102 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.715
+ $Y2=0
r103 39 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.15
+ $Y2=0
r104 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.63
+ $Y2=0
r105 38 41 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.15 $Y2=0
r106 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.715
+ $Y2=0
r107 33 35 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.23
+ $Y2=0
r108 31 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r109 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r110 27 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=0.085
+ $X2=4.29 $Y2=0
r111 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.29 $Y=0.085
+ $X2=4.29 $Y2=0.36
r112 23 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r113 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.36
r114 22 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.63
+ $Y2=0
r115 21 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.63
+ $Y2=0
r116 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=1.795 $Y2=0
r117 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0
r118 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0.36
r119 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r120 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.36
r121 4 29 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=4.12
+ $Y=0.235 $X2=4.29 $Y2=0.36
r122 3 25 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.235 $X2=2.63 $Y2=0.36
r123 2 19 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.63 $Y2=0.36
r124 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.36
.ends


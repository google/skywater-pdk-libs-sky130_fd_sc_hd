* File: sky130_fd_sc_hd__a2111o_4.spice
* Created: Thu Aug 27 13:58:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2111o_4.pex.spice"
.subckt sky130_fd_sc_hd__a2111o_4  VNB VPB D1 C1 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_D1_M1000_g N_A_44_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1000_d N_D1_M1001_g N_A_44_47#_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_C1_M1015_g N_A_44_47#_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.102375 AS=0.091 PD=0.965 PS=0.93 NRD=7.38 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1015_d N_C1_M1016_g N_A_44_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.102375 AS=0.108875 PD=0.965 PS=0.985 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1008 N_A_44_47#_M1016_s N_B1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.2665 PD=0.985 PS=1.47 NRD=10.152 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1019 N_A_44_47#_M1019_d N_B1_M1019_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.2665 PD=0.935 PS=1.47 NRD=0.912 NRS=3.684 M=1 R=4.33333
+ SA=75003 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_A_770_47#_M1010_d N_A1_M1010_g N_A_44_47#_M1019_d VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.092625 PD=0.93 PS=0.935 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.4 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1026 N_A_770_47#_M1010_d N_A1_M1026_g N_A_44_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.182 PD=0.93 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A2_M1011_g N_A_770_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.091 PD=1.86 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_A2_M1022_g N_A_770_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1009_d N_A_44_47#_M1009_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1012 N_X_M1009_d N_A_44_47#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1020 N_X_M1020_d N_A_44_47#_M1020_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1021 N_X_M1020_d N_A_44_47#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_44_47#_M1005_d N_D1_M1005_g N_A_30_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1018 N_A_44_47#_M1005_d N_D1_M1018_g N_A_30_297#_M1018_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1006 N_A_285_297#_M1006_d N_C1_M1006_g N_A_30_297#_M1018_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1024 N_A_285_297#_M1006_d N_C1_M1024_g N_A_30_297#_M1024_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.26 PD=1.28 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_477_297#_M1004_d N_B1_M1004_g N_A_285_297#_M1004_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1014 N_A_477_297#_M1014_d N_B1_M1014_g N_A_285_297#_M1004_s VPB PHIGHVT L=0.15
+ W=1 AD=0.2575 AS=0.14 PD=1.515 PS=1.28 NRD=23.6203 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_477_297#_M1014_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.2575 PD=1.28 PS=1.515 NRD=0 NRS=22.6353 M=1 R=6.66667 SA=75001.3
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1002_d N_A1_M1017_g N_A_477_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.26 PD=1.28 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_477_297#_M1003_d N_A2_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.26 PD=1.28 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1023 N_A_477_297#_M1003_d N_A2_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_44_47#_M1007_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1013 N_X_M1007_d N_A_44_47#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1025 N_X_M1025_d N_A_44_47#_M1025_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1027 N_X_M1025_d N_A_44_47#_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hd__a2111o_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nor3_4.pxi.spice
* Created: Tue Sep  1 19:18:30 2020
* 
x_PM_SKY130_FD_SC_HD__NOR3_4%A N_A_c_96_n N_A_M1003_g N_A_M1002_g N_A_c_97_n
+ N_A_M1005_g N_A_M1012_g N_A_c_98_n N_A_M1009_g N_A_M1015_g N_A_c_99_n
+ N_A_M1010_g N_A_M1022_g A N_A_c_100_n N_A_c_101_n PM_SKY130_FD_SC_HD__NOR3_4%A
x_PM_SKY130_FD_SC_HD__NOR3_4%B N_B_c_170_n N_B_M1011_g N_B_M1000_g N_B_c_171_n
+ N_B_M1013_g N_B_M1007_g N_B_c_172_n N_B_M1017_g N_B_M1016_g N_B_M1020_g
+ N_B_M1018_g N_B_c_182_n N_B_c_183_n N_B_c_184_n N_B_c_185_n N_B_c_173_n
+ N_B_c_174_n N_B_c_175_n B N_B_c_176_n N_B_c_177_n PM_SKY130_FD_SC_HD__NOR3_4%B
x_PM_SKY130_FD_SC_HD__NOR3_4%C N_C_c_304_n N_C_M1006_g N_C_M1001_g N_C_c_305_n
+ N_C_M1014_g N_C_M1004_g N_C_c_306_n N_C_M1019_g N_C_M1008_g N_C_c_307_n
+ N_C_M1021_g N_C_M1023_g C N_C_c_325_n N_C_c_308_n PM_SKY130_FD_SC_HD__NOR3_4%C
x_PM_SKY130_FD_SC_HD__NOR3_4%A_27_297# N_A_27_297#_M1002_s N_A_27_297#_M1012_s
+ N_A_27_297#_M1022_s N_A_27_297#_M1007_d N_A_27_297#_M1018_d
+ N_A_27_297#_c_393_n N_A_27_297#_c_428_p N_A_27_297#_c_394_n
+ N_A_27_297#_c_429_p N_A_27_297#_c_395_n N_A_27_297#_c_396_n
+ N_A_27_297#_c_430_p N_A_27_297#_c_431_p N_A_27_297#_c_456_p
+ N_A_27_297#_c_397_n N_A_27_297#_c_410_n N_A_27_297#_c_412_n
+ N_A_27_297#_c_414_n N_A_27_297#_c_435_p N_A_27_297#_c_415_n
+ PM_SKY130_FD_SC_HD__NOR3_4%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR3_4%VPWR N_VPWR_M1002_d N_VPWR_M1015_d N_VPWR_c_487_n
+ N_VPWR_c_488_n VPWR N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n
+ N_VPWR_c_486_n N_VPWR_c_493_n N_VPWR_c_494_n PM_SKY130_FD_SC_HD__NOR3_4%VPWR
x_PM_SKY130_FD_SC_HD__NOR3_4%A_449_297# N_A_449_297#_M1000_s
+ N_A_449_297#_M1016_s N_A_449_297#_M1004_s N_A_449_297#_M1023_s
+ N_A_449_297#_c_569_n N_A_449_297#_c_570_n N_A_449_297#_c_597_n
+ N_A_449_297#_c_584_n N_A_449_297#_c_586_n N_A_449_297#_c_571_n
+ N_A_449_297#_c_605_n N_A_449_297#_c_606_n
+ PM_SKY130_FD_SC_HD__NOR3_4%A_449_297#
x_PM_SKY130_FD_SC_HD__NOR3_4%Y N_Y_M1003_d N_Y_M1009_d N_Y_M1011_d N_Y_M1017_d
+ N_Y_M1014_s N_Y_M1021_s N_Y_M1001_d N_Y_M1008_d N_Y_c_651_n N_Y_c_634_n
+ N_Y_c_635_n N_Y_c_662_n N_Y_c_636_n N_Y_c_667_n N_Y_c_637_n N_Y_c_685_n
+ N_Y_c_638_n N_Y_c_689_n N_Y_c_727_n N_Y_c_639_n N_Y_c_648_n N_Y_c_694_n
+ N_Y_c_640_n N_Y_c_641_n N_Y_c_642_n N_Y_c_643_n N_Y_c_704_n N_Y_c_644_n
+ N_Y_c_706_n N_Y_c_645_n N_Y_c_646_n N_Y_c_649_n Y PM_SKY130_FD_SC_HD__NOR3_4%Y
x_PM_SKY130_FD_SC_HD__NOR3_4%VGND N_VGND_M1003_s N_VGND_M1005_s N_VGND_M1010_s
+ N_VGND_M1013_s N_VGND_M1006_d N_VGND_M1019_d N_VGND_M1020_s N_VGND_c_828_n
+ N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n
+ N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n
+ N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n N_VGND_c_843_n
+ N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n VGND N_VGND_c_847_n
+ N_VGND_c_848_n N_VGND_c_849_n PM_SKY130_FD_SC_HD__NOR3_4%VGND
cc_1 VNB N_A_c_96_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_97_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_A_c_98_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_A_c_99_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB N_A_c_100_n 0.0200187f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_6 VNB N_A_c_101_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_7 VNB N_B_c_170_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B_c_171_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_9 VNB N_B_c_172_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_10 VNB N_B_c_173_n 0.00679719f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_11 VNB N_B_c_174_n 0.00562963f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_12 VNB N_B_c_175_n 0.0277563f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_13 VNB N_B_c_176_n 0.0461096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B_c_177_n 0.0198341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_C_c_304_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_16 VNB N_C_c_305_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_17 VNB N_C_c_306_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_18 VNB N_C_c_307_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_19 VNB N_C_c_308_n 0.0628802f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_20 VNB N_VPWR_c_486_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_634_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_22 VNB N_Y_c_635_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_636_n 0.00429924f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_24 VNB N_Y_c_637_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_25 VNB N_Y_c_638_n 0.00270792f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.18
cc_26 VNB N_Y_c_639_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_640_n 0.0115223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_641_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_642_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_643_n 0.00253348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_644_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_645_n 0.00379732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_646_n 0.0373197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB Y 0.0224851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_828_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_36 VNB N_VGND_c_829_n 0.0329389f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_37 VNB N_VGND_c_830_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_831_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_832_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_40 VNB N_VGND_c_833_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_41 VNB N_VGND_c_834_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_835_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_836_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_837_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_838_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_839_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_840_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_841_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_842_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_843_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_844_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_845_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_846_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_847_n 0.0169798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_848_n 0.298095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_849_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VPB N_A_M1002_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_58 VPB N_A_M1012_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_59 VPB N_A_M1015_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_60 VPB N_A_M1022_g 0.0185045f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_61 VPB N_A_c_101_n 0.0108808f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_62 VPB N_B_M1000_g 0.018818f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_63 VPB N_B_M1007_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_64 VPB N_B_M1016_g 0.0184964f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_65 VPB N_B_M1018_g 0.0220961f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_66 VPB N_B_c_182_n 0.00216655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_B_c_183_n 0.0091446f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_68 VPB N_B_c_184_n 2.71549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_B_c_185_n 0.00119459f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_70 VPB N_B_c_175_n 0.00685079f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.16
cc_71 VPB N_B_c_176_n 0.00714529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_C_M1001_g 0.0187789f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_73 VPB N_C_M1004_g 0.0180879f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_74 VPB N_C_M1008_g 0.0180987f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_75 VPB N_C_M1023_g 0.0183623f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_76 VPB N_C_c_308_n 0.0105278f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.16
cc_77 VPB N_A_27_297#_c_393_n 0.00371072f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_78 VPB N_A_27_297#_c_394_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_79 VPB N_A_27_297#_c_395_n 0.00240493f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_80 VPB N_A_27_297#_c_396_n 0.00414042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_297#_c_397_n 0.00204609f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.16
cc_82 VPB N_VPWR_c_487_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_83 VPB N_VPWR_c_488_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_84 VPB N_VPWR_c_489_n 0.0180608f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_85 VPB N_VPWR_c_490_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.995
cc_86 VPB N_VPWR_c_491_n 0.105302f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_87 VPB N_VPWR_c_486_n 0.0497918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_493_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_89 VPB N_VPWR_c_494_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_90 VPB N_A_449_297#_c_569_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.995
cc_91 VPB N_A_449_297#_c_570_n 0.00257184f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_92 VPB N_A_449_297#_c_571_n 0.00223882f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_93 VPB N_Y_c_648_n 0.00902013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Y_c_649_n 0.0385079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB Y 0.027853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 N_A_c_99_n N_B_c_170_n 0.0195974f $X=1.75 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_97 N_A_M1022_g N_B_M1000_g 0.0195974f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_c_100_n N_B_c_173_n 0.0121231f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_c_101_n N_B_c_173_n 2.62535e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_c_100_n N_B_c_176_n 2.62535e-19 $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_c_101_n N_B_c_176_n 0.0195974f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_c_100_n N_A_27_297#_c_393_n 0.021852f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_M1002_g N_A_27_297#_c_394_n 0.0134951f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_M1012_g N_A_27_297#_c_394_n 0.0132273f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_c_100_n N_A_27_297#_c_394_n 0.041703f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_c_101_n N_A_27_297#_c_394_n 0.00211509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_M1015_g N_A_27_297#_c_395_n 0.0132273f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_M1022_g N_A_27_297#_c_395_n 0.0132131f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_c_100_n N_A_27_297#_c_395_n 0.0409754f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_c_101_n N_A_27_297#_c_395_n 0.00211509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_c_100_n N_A_27_297#_c_397_n 0.0204549f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_c_101_n N_A_27_297#_c_397_n 0.00220041f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_M1002_g N_VPWR_c_487_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_M1012_g N_VPWR_c_487_n 0.00157837f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_M1015_g N_VPWR_c_488_n 0.00157837f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_M1022_g N_VPWR_c_488_n 0.00302074f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_M1002_g N_VPWR_c_489_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_M1012_g N_VPWR_c_490_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_M1015_g N_VPWR_c_490_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_M1022_g N_VPWR_c_491_n 0.00585385f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_M1002_g N_VPWR_c_486_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_M1012_g N_VPWR_c_486_n 0.0104367f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_M1015_g N_VPWR_c_486_n 0.0104367f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_M1022_g N_VPWR_c_486_n 0.010464f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_c_96_n N_Y_c_651_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_97_n N_Y_c_651_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_98_n N_Y_c_651_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_97_n N_Y_c_634_n 0.00870364f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_98_n N_Y_c_634_n 0.00870364f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_100_n N_Y_c_634_n 0.0362443f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_101_n N_Y_c_634_n 0.00222133f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_c_96_n N_Y_c_635_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_97_n N_Y_c_635_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_100_n N_Y_c_635_n 0.0266272f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_101_n N_Y_c_635_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_97_n N_Y_c_662_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_98_n N_Y_c_662_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_c_99_n N_Y_c_662_n 0.00630972f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_c_99_n N_Y_c_636_n 0.00865686f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_100_n N_Y_c_636_n 0.00826974f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_c_99_n N_Y_c_667_n 5.22228e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_98_n N_Y_c_641_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_c_99_n N_Y_c_641_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_100_n N_Y_c_641_n 0.0266272f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_c_101_n N_Y_c_641_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_c_96_n N_VGND_c_829_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_100_n N_VGND_c_829_n 0.0233945f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_c_97_n N_VGND_c_830_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_98_n N_VGND_c_830_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_99_n N_VGND_c_831_n 0.00146448f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_96_n N_VGND_c_837_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_97_n N_VGND_c_837_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_98_n N_VGND_c_839_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_99_n N_VGND_c_839_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_96_n N_VGND_c_848_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_c_97_n N_VGND_c_848_n 0.0057163f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_98_n N_VGND_c_848_n 0.0057163f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_99_n N_VGND_c_848_n 0.0057435f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B_c_172_n N_C_c_304_n 0.0148255f $X=3.01 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_160 N_B_M1016_g N_C_M1001_g 0.0148255f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_161 N_B_c_182_n N_C_M1001_g 0.0029914f $X=3.6 $Y=1.445 $X2=0 $Y2=0
cc_162 N_B_c_184_n N_C_M1001_g 0.00117404f $X=3.685 $Y=1.53 $X2=0 $Y2=0
cc_163 N_B_c_182_n N_C_M1004_g 0.00270232f $X=3.6 $Y=1.445 $X2=0 $Y2=0
cc_164 N_B_c_183_n N_C_M1004_g 0.0109874f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_165 N_B_c_183_n N_C_M1008_g 0.0103077f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_166 N_B_c_177_n N_C_c_307_n 0.0124239f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B_M1018_g N_C_M1023_g 0.043976f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_168 N_B_c_183_n N_C_M1023_g 0.010294f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_169 N_B_c_185_n N_C_M1023_g 0.00227715f $X=5.08 $Y=1.445 $X2=0 $Y2=0
cc_170 N_B_c_183_n N_C_c_325_n 0.0646929f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_171 N_B_c_173_n N_C_c_325_n 0.0168497f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_172 N_B_c_174_n N_C_c_325_n 0.0126856f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B_c_175_n N_C_c_325_n 2.51215e-19 $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B_c_182_n N_C_c_308_n 0.00472016f $X=3.6 $Y=1.445 $X2=0 $Y2=0
cc_175 N_B_c_183_n N_C_c_308_n 0.00427825f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_176 N_B_c_185_n N_C_c_308_n 3.07103e-19 $X=5.08 $Y=1.445 $X2=0 $Y2=0
cc_177 N_B_c_173_n N_C_c_308_n 0.0235052f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_178 N_B_c_174_n N_C_c_308_n 9.04748e-19 $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B_c_175_n N_C_c_308_n 0.0209639f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B_c_176_n N_C_c_308_n 0.0148255f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B_M1000_g N_A_27_297#_c_396_n 2.57315e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B_M1000_g N_A_27_297#_c_410_n 0.0180937f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B_M1007_g N_A_27_297#_c_410_n 0.0133705f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B_M1000_g N_A_27_297#_c_412_n 3.26991e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B_M1007_g N_A_27_297#_c_412_n 0.00199018f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B_M1018_g N_A_27_297#_c_414_n 0.00248744f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B_M1016_g N_A_27_297#_c_415_n 0.00303361f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B_M1018_g N_A_27_297#_c_415_n 0.00173656f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B_c_183_n N_A_27_297#_c_415_n 0.0012671f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_190 N_B_c_184_n N_A_27_297#_c_415_n 3.67354e-19 $X=3.685 $Y=1.53 $X2=0 $Y2=0
cc_191 N_B_M1000_g N_VPWR_c_491_n 0.00357877f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B_M1007_g N_VPWR_c_491_n 0.00357877f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B_M1016_g N_VPWR_c_491_n 0.00585385f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B_M1018_g N_VPWR_c_491_n 0.00585385f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B_M1000_g N_VPWR_c_486_n 0.00525237f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B_M1007_g N_VPWR_c_486_n 0.00463869f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B_M1016_g N_VPWR_c_486_n 0.0053842f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B_M1018_g N_VPWR_c_486_n 0.00634478f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B_c_183_n N_A_449_297#_M1004_s 0.00162946f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_200 N_B_c_183_n N_A_449_297#_M1023_s 0.00162946f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_201 N_B_M1007_g N_A_449_297#_c_569_n 0.0100078f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B_M1016_g N_A_449_297#_c_569_n 0.00991964f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B_c_173_n N_A_449_297#_c_569_n 0.041703f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_204 N_B_c_176_n N_A_449_297#_c_569_n 0.00211509f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B_c_184_n N_A_449_297#_c_570_n 0.00271526f $X=3.685 $Y=1.53 $X2=0 $Y2=0
cc_206 N_B_c_173_n N_A_449_297#_c_570_n 0.0214236f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_207 N_B_M1000_g N_A_449_297#_c_571_n 2.57315e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B_c_173_n N_A_449_297#_c_571_n 0.0197947f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_209 N_B_c_176_n N_A_449_297#_c_571_n 0.00217153f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B_c_183_n N_Y_M1001_d 3.33457e-19 $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_211 N_B_c_184_n N_Y_M1001_d 0.00152582f $X=3.685 $Y=1.53 $X2=0 $Y2=0
cc_212 N_B_c_183_n N_Y_M1008_d 0.0016256f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_213 N_B_c_170_n N_Y_c_662_n 5.22228e-19 $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B_c_170_n N_Y_c_636_n 0.00865686f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B_c_173_n N_Y_c_636_n 0.00826974f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_216 N_B_c_170_n N_Y_c_667_n 0.00630972f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B_c_171_n N_Y_c_667_n 0.00630972f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B_c_172_n N_Y_c_667_n 5.22228e-19 $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B_c_171_n N_Y_c_637_n 0.00870364f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B_c_172_n N_Y_c_637_n 0.00870364f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B_c_173_n N_Y_c_637_n 0.0362443f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_222 N_B_c_176_n N_Y_c_637_n 0.00222133f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B_c_171_n N_Y_c_685_n 5.22228e-19 $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B_c_172_n N_Y_c_685_n 0.00630972f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B_c_183_n N_Y_c_638_n 0.0051766f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_226 N_B_c_173_n N_Y_c_638_n 0.0223602f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_227 N_B_c_183_n N_Y_c_689_n 0.0307122f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_228 N_B_M1018_g N_Y_c_648_n 0.0127965f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B_c_183_n N_Y_c_648_n 0.0297391f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_230 N_B_c_174_n N_Y_c_648_n 0.00711886f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B_c_175_n N_Y_c_648_n 0.00236763f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B_c_177_n N_Y_c_694_n 0.0069263f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B_c_174_n N_Y_c_640_n 0.0254021f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B_c_175_n N_Y_c_640_n 0.00345541f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B_c_177_n N_Y_c_640_n 0.0108868f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B_c_170_n N_Y_c_642_n 0.00113286f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B_c_171_n N_Y_c_642_n 0.00113286f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B_c_173_n N_Y_c_642_n 0.0266272f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_239 N_B_c_176_n N_Y_c_642_n 0.00230339f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_240 N_B_c_172_n N_Y_c_643_n 0.00112787f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B_c_173_n N_Y_c_643_n 0.0276736f $X=3.515 $Y=1.18 $X2=0 $Y2=0
cc_242 N_B_c_183_n N_Y_c_704_n 0.00242944f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_243 N_B_c_184_n N_Y_c_704_n 0.0100253f $X=3.685 $Y=1.53 $X2=0 $Y2=0
cc_244 N_B_c_183_n N_Y_c_706_n 0.0116461f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_245 N_B_c_183_n N_Y_c_645_n 0.00867576f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_246 N_B_c_174_n N_Y_c_645_n 0.00557001f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_247 N_B_c_175_n N_Y_c_645_n 0.00102373f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B_c_177_n N_Y_c_645_n 0.00112787f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B_c_177_n N_Y_c_646_n 0.00309584f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B_M1018_g N_Y_c_649_n 0.00476503f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B_M1018_g Y 0.00956267f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_252 N_B_c_183_n Y 0.00690775f $X=4.995 $Y=1.53 $X2=0 $Y2=0
cc_253 N_B_c_185_n Y 0.00586153f $X=5.08 $Y=1.445 $X2=0 $Y2=0
cc_254 N_B_c_174_n Y 0.0162231f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B_c_175_n Y 0.00501066f $X=5.16 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B_c_177_n Y 0.0024947f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B_c_170_n N_VGND_c_831_n 0.00146448f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B_c_171_n N_VGND_c_832_n 0.00146448f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_259 N_B_c_172_n N_VGND_c_832_n 0.00146448f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B_c_177_n N_VGND_c_835_n 0.00423334f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_261 N_B_c_177_n N_VGND_c_836_n 0.00316354f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_262 N_B_c_170_n N_VGND_c_841_n 0.00423334f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_263 N_B_c_171_n N_VGND_c_841_n 0.00423334f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_264 N_B_c_172_n N_VGND_c_843_n 0.00423334f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_265 N_B_c_170_n N_VGND_c_848_n 0.0057435f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_266 N_B_c_171_n N_VGND_c_848_n 0.0057163f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B_c_172_n N_VGND_c_848_n 0.0057435f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B_c_177_n N_VGND_c_848_n 0.00706957f $X=5.16 $Y=0.995 $X2=0 $Y2=0
cc_269 N_C_M1023_g N_A_27_297#_c_414_n 2.77803e-19 $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_270 N_C_M1001_g N_A_27_297#_c_415_n 0.00804291f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_271 N_C_M1004_g N_A_27_297#_c_415_n 0.00329221f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_272 N_C_M1008_g N_A_27_297#_c_415_n 0.00329221f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_273 N_C_M1023_g N_A_27_297#_c_415_n 0.00330658f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_274 N_C_M1001_g N_VPWR_c_491_n 0.00357877f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_275 N_C_M1004_g N_VPWR_c_491_n 0.00357877f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_276 N_C_M1008_g N_VPWR_c_491_n 0.00357877f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_277 N_C_M1023_g N_VPWR_c_491_n 0.00357877f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_278 N_C_M1001_g N_VPWR_c_486_n 0.00475717f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_279 N_C_M1004_g N_VPWR_c_486_n 0.00472997f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_280 N_C_M1008_g N_VPWR_c_486_n 0.00472997f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_281 N_C_M1023_g N_VPWR_c_486_n 0.00475717f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_282 N_C_M1001_g N_A_449_297#_c_570_n 2.57315e-19 $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_283 N_C_M1001_g N_A_449_297#_c_584_n 0.00766643f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_284 N_C_M1004_g N_A_449_297#_c_584_n 0.00822051f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_285 N_C_M1008_g N_A_449_297#_c_586_n 0.00822051f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_286 N_C_M1023_g N_A_449_297#_c_586_n 0.0082601f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_287 N_C_c_304_n N_Y_c_685_n 0.00630972f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_288 N_C_c_305_n N_Y_c_685_n 5.22228e-19 $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_289 N_C_c_304_n N_Y_c_638_n 0.00870364f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_290 N_C_c_305_n N_Y_c_638_n 0.00968707f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_291 N_C_c_325_n N_Y_c_638_n 0.00266908f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_292 N_C_c_308_n N_Y_c_638_n 0.00222006f $X=4.69 $Y=1.16 $X2=0 $Y2=0
cc_293 N_C_M1004_g N_Y_c_689_n 0.00930781f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_294 N_C_M1008_g N_Y_c_689_n 0.00930781f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_295 N_C_c_304_n N_Y_c_727_n 5.22228e-19 $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_296 N_C_c_305_n N_Y_c_727_n 0.00630972f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_297 N_C_c_306_n N_Y_c_727_n 0.00630972f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_298 N_C_c_307_n N_Y_c_727_n 5.22228e-19 $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_299 N_C_c_306_n N_Y_c_639_n 0.00869873f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_300 N_C_c_307_n N_Y_c_639_n 0.00869873f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_301 N_C_c_325_n N_Y_c_639_n 0.0363039f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_302 N_C_c_308_n N_Y_c_639_n 0.00222006f $X=4.69 $Y=1.16 $X2=0 $Y2=0
cc_303 N_C_M1023_g N_Y_c_648_n 0.0090766f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_304 N_C_c_306_n N_Y_c_694_n 5.22228e-19 $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_305 N_C_c_307_n N_Y_c_694_n 0.00630972f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_306 N_C_c_304_n N_Y_c_643_n 0.00112787f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_307 N_C_c_308_n N_Y_c_704_n 3.50616e-19 $X=4.69 $Y=1.16 $X2=0 $Y2=0
cc_308 N_C_c_305_n N_Y_c_644_n 0.00113159f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_309 N_C_c_306_n N_Y_c_644_n 0.00113159f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_310 N_C_c_325_n N_Y_c_644_n 0.0266779f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_311 N_C_c_308_n N_Y_c_644_n 0.00230167f $X=4.69 $Y=1.16 $X2=0 $Y2=0
cc_312 N_C_c_307_n N_Y_c_645_n 0.00111217f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_313 N_C_c_325_n N_Y_c_645_n 0.00223821f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_314 N_C_c_304_n N_VGND_c_833_n 0.00146448f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_315 N_C_c_305_n N_VGND_c_833_n 0.00146448f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_316 N_C_c_306_n N_VGND_c_834_n 0.00146448f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_317 N_C_c_307_n N_VGND_c_834_n 0.00146448f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_318 N_C_c_307_n N_VGND_c_835_n 0.00423334f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_319 N_C_c_304_n N_VGND_c_843_n 0.00423334f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_320 N_C_c_305_n N_VGND_c_845_n 0.00423334f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_321 N_C_c_306_n N_VGND_c_845_n 0.00423334f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_322 N_C_c_304_n N_VGND_c_848_n 0.0057435f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_323 N_C_c_305_n N_VGND_c_848_n 0.0057163f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_324 N_C_c_306_n N_VGND_c_848_n 0.0057163f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_325 N_C_c_307_n N_VGND_c_848_n 0.0057435f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_27_297#_c_394_n N_VPWR_M1002_d 0.00165831f $X=0.995 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_327 N_A_27_297#_c_395_n N_VPWR_M1015_d 0.00165831f $X=1.835 $Y=1.54 $X2=0
+ $Y2=0
cc_328 N_A_27_297#_c_394_n N_VPWR_c_487_n 0.0126919f $X=0.995 $Y=1.54 $X2=0
+ $Y2=0
cc_329 N_A_27_297#_c_395_n N_VPWR_c_488_n 0.0126919f $X=1.835 $Y=1.54 $X2=0
+ $Y2=0
cc_330 N_A_27_297#_c_428_p N_VPWR_c_489_n 0.0161885f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_331 N_A_27_297#_c_429_p N_VPWR_c_490_n 0.0142343f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_332 N_A_27_297#_c_430_p N_VPWR_c_491_n 0.0143053f $X=1.96 $Y=2.085 $X2=0
+ $Y2=0
cc_333 N_A_27_297#_c_431_p N_VPWR_c_491_n 0.0142933f $X=2.8 $Y=2.085 $X2=0 $Y2=0
cc_334 N_A_27_297#_c_410_n N_VPWR_c_491_n 0.0346052f $X=2.675 $Y=2.275 $X2=0
+ $Y2=0
cc_335 N_A_27_297#_c_412_n N_VPWR_c_491_n 2.00309e-19 $X=2.68 $Y=2.2 $X2=0 $Y2=0
cc_336 N_A_27_297#_c_414_n N_VPWR_c_491_n 4.20246e-19 $X=5.29 $Y=2.21 $X2=0
+ $Y2=0
cc_337 N_A_27_297#_c_435_p N_VPWR_c_491_n 0.0151494f $X=5.29 $Y=2.21 $X2=0 $Y2=0
cc_338 N_A_27_297#_c_415_n N_VPWR_c_491_n 0.00206198f $X=5.145 $Y=2.2 $X2=0
+ $Y2=0
cc_339 N_A_27_297#_M1002_s N_VPWR_c_486_n 0.00315976f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_340 N_A_27_297#_M1012_s N_VPWR_c_486_n 0.00284632f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_341 N_A_27_297#_M1022_s N_VPWR_c_486_n 0.00246446f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_342 N_A_27_297#_M1007_d N_VPWR_c_486_n 0.00125036f $X=2.665 $Y=1.485 $X2=0
+ $Y2=0
cc_343 N_A_27_297#_M1018_d N_VPWR_c_486_n 0.00107794f $X=5.185 $Y=1.485 $X2=0
+ $Y2=0
cc_344 N_A_27_297#_c_428_p N_VPWR_c_486_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_345 N_A_27_297#_c_429_p N_VPWR_c_486_n 0.00955092f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_346 N_A_27_297#_c_430_p N_VPWR_c_486_n 0.00962794f $X=1.96 $Y=2.085 $X2=0
+ $Y2=0
cc_347 N_A_27_297#_c_431_p N_VPWR_c_486_n 0.00270511f $X=2.8 $Y=2.085 $X2=0
+ $Y2=0
cc_348 N_A_27_297#_c_410_n N_VPWR_c_486_n 0.0130024f $X=2.675 $Y=2.275 $X2=0
+ $Y2=0
cc_349 N_A_27_297#_c_412_n N_VPWR_c_486_n 0.029679f $X=2.68 $Y=2.2 $X2=0 $Y2=0
cc_350 N_A_27_297#_c_414_n N_VPWR_c_486_n 0.0298605f $X=5.29 $Y=2.21 $X2=0 $Y2=0
cc_351 N_A_27_297#_c_435_p N_VPWR_c_486_n 0.00228824f $X=5.29 $Y=2.21 $X2=0
+ $Y2=0
cc_352 N_A_27_297#_c_415_n N_VPWR_c_486_n 0.211701f $X=5.145 $Y=2.2 $X2=0 $Y2=0
cc_353 N_A_27_297#_c_410_n N_A_449_297#_M1000_s 0.00275102f $X=2.675 $Y=2.275
+ $X2=-0.19 $Y2=1.305
cc_354 N_A_27_297#_c_412_n N_A_449_297#_M1000_s 0.00129367f $X=2.68 $Y=2.2
+ $X2=-0.19 $Y2=1.305
cc_355 N_A_27_297#_c_415_n N_A_449_297#_M1016_s 4.81483e-19 $X=5.145 $Y=2.2
+ $X2=0 $Y2=0
cc_356 N_A_27_297#_c_415_n N_A_449_297#_M1023_s 2.09851e-19 $X=5.145 $Y=2.2
+ $X2=0 $Y2=0
cc_357 N_A_27_297#_M1007_d N_A_449_297#_c_569_n 0.00162384f $X=2.665 $Y=1.485
+ $X2=0 $Y2=0
cc_358 N_A_27_297#_c_456_p N_A_449_297#_c_569_n 0.0123012f $X=2.8 $Y=1.96 $X2=0
+ $Y2=0
cc_359 N_A_27_297#_c_410_n N_A_449_297#_c_569_n 0.00282963f $X=2.675 $Y=2.275
+ $X2=0 $Y2=0
cc_360 N_A_27_297#_c_412_n N_A_449_297#_c_569_n 0.0033396f $X=2.68 $Y=2.2 $X2=0
+ $Y2=0
cc_361 N_A_27_297#_c_415_n N_A_449_297#_c_569_n 0.00533813f $X=5.145 $Y=2.2
+ $X2=0 $Y2=0
cc_362 N_A_27_297#_c_431_p N_A_449_297#_c_597_n 0.00510852f $X=2.8 $Y=2.085
+ $X2=0 $Y2=0
cc_363 N_A_27_297#_c_412_n N_A_449_297#_c_597_n 6.00101e-19 $X=2.68 $Y=2.2 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_c_415_n N_A_449_297#_c_597_n 0.0248323f $X=5.145 $Y=2.2 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_c_415_n N_A_449_297#_c_584_n 0.00844892f $X=5.145 $Y=2.2
+ $X2=0 $Y2=0
cc_366 N_A_27_297#_c_415_n N_A_449_297#_c_586_n 0.00557315f $X=5.145 $Y=2.2
+ $X2=0 $Y2=0
cc_367 N_A_27_297#_c_396_n N_A_449_297#_c_571_n 0.00271526f $X=1.96 $Y=1.625
+ $X2=0 $Y2=0
cc_368 N_A_27_297#_c_410_n N_A_449_297#_c_571_n 0.01263f $X=2.675 $Y=2.275 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_412_n N_A_449_297#_c_571_n 0.00351885f $X=2.68 $Y=2.2 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_415_n N_A_449_297#_c_605_n 0.0161944f $X=5.145 $Y=2.2 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_414_n N_A_449_297#_c_606_n 0.00160175f $X=5.29 $Y=2.21
+ $X2=0 $Y2=0
cc_372 N_A_27_297#_c_435_p N_A_449_297#_c_606_n 0.0060695f $X=5.29 $Y=2.21 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_415_n N_A_449_297#_c_606_n 0.0142278f $X=5.145 $Y=2.2 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_c_415_n N_Y_M1001_d 0.00339819f $X=5.145 $Y=2.2 $X2=0 $Y2=0
cc_375 N_A_27_297#_c_415_n N_Y_M1008_d 0.00312809f $X=5.145 $Y=2.2 $X2=0 $Y2=0
cc_376 N_A_27_297#_c_395_n N_Y_c_636_n 3.18413e-19 $X=1.835 $Y=1.54 $X2=0 $Y2=0
cc_377 N_A_27_297#_c_396_n N_Y_c_636_n 0.00936521f $X=1.96 $Y=1.625 $X2=0 $Y2=0
cc_378 N_A_27_297#_c_415_n N_Y_c_689_n 0.00970393f $X=5.145 $Y=2.2 $X2=0 $Y2=0
cc_379 N_A_27_297#_M1018_d N_Y_c_648_n 0.0066394f $X=5.185 $Y=1.485 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_414_n N_Y_c_648_n 0.00969021f $X=5.29 $Y=2.21 $X2=0 $Y2=0
cc_381 N_A_27_297#_c_435_p N_Y_c_648_n 0.0138081f $X=5.29 $Y=2.21 $X2=0 $Y2=0
cc_382 N_A_27_297#_c_415_n N_Y_c_648_n 0.010254f $X=5.145 $Y=2.2 $X2=0 $Y2=0
cc_383 N_A_27_297#_c_415_n N_Y_c_704_n 0.00762843f $X=5.145 $Y=2.2 $X2=0 $Y2=0
cc_384 N_A_27_297#_c_414_n N_Y_c_706_n 0.00192199f $X=5.29 $Y=2.21 $X2=0 $Y2=0
cc_385 N_A_27_297#_c_415_n N_Y_c_706_n 0.00762843f $X=5.145 $Y=2.2 $X2=0 $Y2=0
cc_386 N_A_27_297#_c_414_n N_Y_c_649_n 0.00465658f $X=5.29 $Y=2.21 $X2=0 $Y2=0
cc_387 N_A_27_297#_c_435_p N_Y_c_649_n 0.0252914f $X=5.29 $Y=2.21 $X2=0 $Y2=0
cc_388 N_VPWR_c_486_n N_A_449_297#_M1000_s 0.00165992f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_389 N_VPWR_c_486_n N_A_449_297#_M1016_s 0.00125614f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_486_n N_A_449_297#_M1004_s 0.00120563f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_486_n N_A_449_297#_M1023_s 0.00123032f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_491_n N_A_449_297#_c_597_n 0.0143053f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_486_n N_A_449_297#_c_597_n 0.00271607f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_491_n N_A_449_297#_c_584_n 0.0330174f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_486_n N_A_449_297#_c_584_n 0.00526545f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_491_n N_A_449_297#_c_586_n 0.0330174f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_486_n N_A_449_297#_c_586_n 0.00526944f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_491_n N_A_449_297#_c_605_n 0.0136817f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_486_n N_A_449_297#_c_605_n 0.00252432f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_491_n N_A_449_297#_c_606_n 0.0136817f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_486_n N_A_449_297#_c_606_n 0.00252432f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_486_n N_Y_M1001_d 0.00121934f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_c_486_n N_Y_M1008_d 0.0012148f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_486_n N_Y_c_648_n 0.00618566f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_c_491_n N_Y_c_649_n 0.0199313f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_c_486_n N_Y_c_649_n 0.0111033f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_407 N_A_449_297#_c_584_n N_Y_M1001_d 0.00292711f $X=3.935 $Y=2.38 $X2=0 $Y2=0
cc_408 N_A_449_297#_c_586_n N_Y_M1008_d 0.00292711f $X=4.775 $Y=2.38 $X2=0 $Y2=0
cc_409 N_A_449_297#_M1004_s N_Y_c_689_n 0.00305775f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_410 N_A_449_297#_c_584_n N_Y_c_689_n 0.00333267f $X=3.935 $Y=2.38 $X2=0 $Y2=0
cc_411 N_A_449_297#_c_586_n N_Y_c_689_n 0.00333267f $X=4.775 $Y=2.38 $X2=0 $Y2=0
cc_412 N_A_449_297#_c_605_n N_Y_c_689_n 0.0109639f $X=4.06 $Y=2.3 $X2=0 $Y2=0
cc_413 N_A_449_297#_M1023_s N_Y_c_648_n 0.00320832f $X=4.765 $Y=1.485 $X2=0
+ $Y2=0
cc_414 N_A_449_297#_c_586_n N_Y_c_648_n 0.00318888f $X=4.775 $Y=2.38 $X2=0 $Y2=0
cc_415 N_A_449_297#_c_606_n N_Y_c_648_n 0.0103896f $X=4.9 $Y=2.3 $X2=0 $Y2=0
cc_416 N_A_449_297#_c_584_n N_Y_c_704_n 0.00932136f $X=3.935 $Y=2.38 $X2=0 $Y2=0
cc_417 N_A_449_297#_c_586_n N_Y_c_706_n 0.00932136f $X=4.775 $Y=2.38 $X2=0 $Y2=0
cc_418 N_Y_c_634_n N_VGND_M1005_s 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_419 N_Y_c_636_n N_VGND_M1010_s 0.00162089f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_420 N_Y_c_637_n N_VGND_M1013_s 0.00162089f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_421 N_Y_c_638_n N_VGND_M1006_d 0.00162089f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_422 N_Y_c_639_n N_VGND_M1019_d 0.00162089f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_423 N_Y_c_640_n N_VGND_M1020_s 0.00315681f $X=5.605 $Y=0.815 $X2=0 $Y2=0
cc_424 N_Y_c_635_n N_VGND_c_829_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_425 N_Y_c_634_n N_VGND_c_830_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_426 N_Y_c_636_n N_VGND_c_831_n 0.0122559f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_427 N_Y_c_637_n N_VGND_c_832_n 0.0122559f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_428 N_Y_c_638_n N_VGND_c_833_n 0.0122559f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_429 N_Y_c_639_n N_VGND_c_834_n 0.0122559f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_430 N_Y_c_639_n N_VGND_c_835_n 0.00198695f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_431 N_Y_c_694_n N_VGND_c_835_n 0.0188551f $X=4.9 $Y=0.39 $X2=0 $Y2=0
cc_432 N_Y_c_640_n N_VGND_c_835_n 0.00198695f $X=5.605 $Y=0.815 $X2=0 $Y2=0
cc_433 N_Y_c_640_n N_VGND_c_836_n 0.0127273f $X=5.605 $Y=0.815 $X2=0 $Y2=0
cc_434 N_Y_c_646_n N_VGND_c_836_n 0.0205861f $X=5.75 $Y=0.815 $X2=0 $Y2=0
cc_435 N_Y_c_651_n N_VGND_c_837_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_436 N_Y_c_634_n N_VGND_c_837_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_437 N_Y_c_634_n N_VGND_c_839_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_438 N_Y_c_662_n N_VGND_c_839_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_439 N_Y_c_636_n N_VGND_c_839_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_440 N_Y_c_636_n N_VGND_c_841_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_441 N_Y_c_667_n N_VGND_c_841_n 0.0188551f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_442 N_Y_c_637_n N_VGND_c_841_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_443 N_Y_c_637_n N_VGND_c_843_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_444 N_Y_c_685_n N_VGND_c_843_n 0.0188551f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_445 N_Y_c_638_n N_VGND_c_843_n 0.00198695f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_446 N_Y_c_638_n N_VGND_c_845_n 0.00198695f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_447 N_Y_c_727_n N_VGND_c_845_n 0.0188551f $X=4.06 $Y=0.39 $X2=0 $Y2=0
cc_448 N_Y_c_639_n N_VGND_c_845_n 0.00198695f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_449 N_Y_c_640_n N_VGND_c_847_n 0.00301521f $X=5.605 $Y=0.815 $X2=0 $Y2=0
cc_450 N_Y_c_646_n N_VGND_c_847_n 0.0206482f $X=5.75 $Y=0.815 $X2=0 $Y2=0
cc_451 N_Y_M1003_d N_VGND_c_848_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_452 N_Y_M1009_d N_VGND_c_848_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_453 N_Y_M1011_d N_VGND_c_848_n 0.00215201f $X=2.245 $Y=0.235 $X2=0 $Y2=0
cc_454 N_Y_M1017_d N_VGND_c_848_n 0.00215201f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_455 N_Y_M1014_s N_VGND_c_848_n 0.00215201f $X=3.925 $Y=0.235 $X2=0 $Y2=0
cc_456 N_Y_M1021_s N_VGND_c_848_n 0.00215201f $X=4.765 $Y=0.235 $X2=0 $Y2=0
cc_457 N_Y_c_651_n N_VGND_c_848_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_458 N_Y_c_634_n N_VGND_c_848_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_459 N_Y_c_662_n N_VGND_c_848_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_460 N_Y_c_636_n N_VGND_c_848_n 0.00835832f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_461 N_Y_c_667_n N_VGND_c_848_n 0.0122069f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_462 N_Y_c_637_n N_VGND_c_848_n 0.00835832f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_463 N_Y_c_685_n N_VGND_c_848_n 0.0122069f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_464 N_Y_c_638_n N_VGND_c_848_n 0.00835832f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_465 N_Y_c_727_n N_VGND_c_848_n 0.0122069f $X=4.06 $Y=0.39 $X2=0 $Y2=0
cc_466 N_Y_c_639_n N_VGND_c_848_n 0.00835832f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_467 N_Y_c_694_n N_VGND_c_848_n 0.0122069f $X=4.9 $Y=0.39 $X2=0 $Y2=0
cc_468 N_Y_c_640_n N_VGND_c_848_n 0.00983014f $X=5.605 $Y=0.815 $X2=0 $Y2=0
cc_469 N_Y_c_646_n N_VGND_c_848_n 0.0110914f $X=5.75 $Y=0.815 $X2=0 $Y2=0

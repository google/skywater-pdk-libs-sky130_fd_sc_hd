# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o22ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 1.415000 1.275000 ;
        RECT 1.150000 1.275000 1.415000 1.445000 ;
        RECT 1.150000 1.445000 3.575000 1.615000 ;
        RECT 3.275000 1.075000 3.605000 1.245000 ;
        RECT 3.275000 1.245000 3.575000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.685000 1.075000 3.095000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295000 0.995000 4.940000 1.445000 ;
        RECT 4.295000 1.445000 6.935000 1.615000 ;
        RECT 6.715000 0.995000 6.935000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.110000 1.075000 6.460000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 1.785000 3.915000 1.955000 ;
        RECT 1.845000 1.955000 2.095000 2.125000 ;
        RECT 2.685000 1.955000 2.935000 2.125000 ;
        RECT 3.745000 1.445000 4.125000 1.615000 ;
        RECT 3.745000 1.615000 3.915000 1.785000 ;
        RECT 3.955000 0.645000 7.275000 0.820000 ;
        RECT 3.955000 0.820000 4.125000 1.445000 ;
        RECT 5.255000 1.785000 7.275000 1.955000 ;
        RECT 5.255000 1.955000 5.505000 2.125000 ;
        RECT 6.095000 1.955000 6.345000 2.125000 ;
        RECT 7.105000 0.820000 7.275000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.360000 0.085000 ;
        RECT 0.625000  0.085000 0.795000 0.555000 ;
        RECT 1.465000  0.085000 1.635000 0.555000 ;
        RECT 2.305000  0.085000 2.475000 0.555000 ;
        RECT 3.145000  0.085000 3.315000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.165000 1.445000 0.415000 2.635000 ;
        RECT 1.005000 2.125000 1.255000 2.635000 ;
        RECT 3.565000 2.125000 3.785000 2.635000 ;
        RECT 4.425000 2.125000 4.665000 2.635000 ;
        RECT 6.935000 2.125000 7.215000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.125000 0.255000 0.455000 0.725000 ;
      RECT 0.125000 0.725000 1.295000 0.735000 ;
      RECT 0.125000 0.735000 3.785000 0.905000 ;
      RECT 0.585000 1.445000 0.835000 1.785000 ;
      RECT 0.585000 1.785000 1.675000 1.955000 ;
      RECT 0.585000 1.955000 0.835000 2.465000 ;
      RECT 0.965000 0.255000 1.295000 0.725000 ;
      RECT 1.425000 1.955000 1.675000 2.295000 ;
      RECT 1.425000 2.295000 3.395000 2.465000 ;
      RECT 1.805000 0.255000 2.135000 0.725000 ;
      RECT 1.805000 0.725000 2.975000 0.735000 ;
      RECT 2.265000 2.125000 2.515000 2.295000 ;
      RECT 2.645000 0.255000 2.975000 0.725000 ;
      RECT 3.105000 2.125000 3.395000 2.295000 ;
      RECT 3.485000 0.255000 7.245000 0.475000 ;
      RECT 3.485000 0.475000 3.785000 0.735000 ;
      RECT 3.955000 2.125000 4.255000 2.465000 ;
      RECT 4.085000 1.785000 5.085000 1.955000 ;
      RECT 4.085000 1.955000 4.255000 2.125000 ;
      RECT 4.835000 1.955000 5.085000 2.295000 ;
      RECT 4.835000 2.295000 6.765000 2.465000 ;
      RECT 5.675000 2.125000 5.925000 2.295000 ;
      RECT 6.515000 2.135000 6.765000 2.295000 ;
  END
END sky130_fd_sc_hd__o22ai_4
END LIBRARY

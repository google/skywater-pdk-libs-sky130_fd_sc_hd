* File: sky130_fd_sc_hd__o21a_1.pxi.spice
* Created: Tue Sep  1 19:21:06 2020
* 
x_PM_SKY130_FD_SC_HD__O21A_1%A_79_21# N_A_79_21#_M1001_s N_A_79_21#_M1002_d
+ N_A_79_21#_c_52_n N_A_79_21#_M1007_g N_A_79_21#_M1000_g N_A_79_21#_c_53_n
+ N_A_79_21#_c_54_n N_A_79_21#_c_59_n N_A_79_21#_c_86_p N_A_79_21#_c_60_n
+ N_A_79_21#_c_94_p N_A_79_21#_c_55_n PM_SKY130_FD_SC_HD__O21A_1%A_79_21#
x_PM_SKY130_FD_SC_HD__O21A_1%B1 N_B1_M1002_g N_B1_M1001_g B1 N_B1_c_109_n
+ N_B1_c_110_n N_B1_c_111_n PM_SKY130_FD_SC_HD__O21A_1%B1
x_PM_SKY130_FD_SC_HD__O21A_1%A2 N_A2_M1004_g N_A2_c_142_n N_A2_M1005_g A2
+ N_A2_c_144_n PM_SKY130_FD_SC_HD__O21A_1%A2
x_PM_SKY130_FD_SC_HD__O21A_1%A1 N_A1_c_181_n N_A1_M1003_g N_A1_M1006_g
+ N_A1_c_182_n N_A1_c_183_n A1 PM_SKY130_FD_SC_HD__O21A_1%A1
x_PM_SKY130_FD_SC_HD__O21A_1%X N_X_M1007_s N_X_M1000_s N_X_c_209_n N_X_c_210_n X
+ N_X_c_211_n PM_SKY130_FD_SC_HD__O21A_1%X
x_PM_SKY130_FD_SC_HD__O21A_1%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_231_n VPWR N_VPWR_c_232_n N_VPWR_c_233_n
+ N_VPWR_c_234_n N_VPWR_c_228_n PM_SKY130_FD_SC_HD__O21A_1%VPWR
x_PM_SKY130_FD_SC_HD__O21A_1%VGND N_VGND_M1007_d N_VGND_M1005_d N_VGND_c_270_n
+ N_VGND_c_271_n N_VGND_c_272_n VGND N_VGND_c_273_n N_VGND_c_274_n
+ N_VGND_c_275_n N_VGND_c_276_n N_VGND_c_277_n PM_SKY130_FD_SC_HD__O21A_1%VGND
x_PM_SKY130_FD_SC_HD__O21A_1%A_297_47# N_A_297_47#_M1001_d N_A_297_47#_M1003_d
+ N_A_297_47#_c_310_n N_A_297_47#_c_311_n N_A_297_47#_c_312_n
+ PM_SKY130_FD_SC_HD__O21A_1%A_297_47#
cc_1 VNB N_A_79_21#_c_52_n 0.0230987f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_53_n 0.00419194f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_3 VNB N_A_79_21#_c_54_n 0.0357061f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_4 VNB N_A_79_21#_c_55_n 0.0148524f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.4
cc_5 VNB N_B1_c_109_n 0.0231136f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_6 VNB N_B1_c_110_n 0.00636433f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_7 VNB N_B1_c_111_n 0.0203098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A2_c_142_n 0.0165981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB A2 0.00551734f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A2_c_144_n 0.0195258f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_11 VNB N_A1_c_181_n 0.021688f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=0.235
cc_12 VNB N_A1_c_182_n 0.00772443f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_13 VNB N_A1_c_183_n 0.0365712f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_14 VNB A1 0.00103399f $X=-0.19 $Y=-0.24 $X2=0.737 $Y2=0.905
cc_15 VNB N_X_c_209_n 0.0240441f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_X_c_210_n 0.00831783f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_17 VNB N_X_c_211_n 0.0135933f $X=-0.19 $Y=-0.24 $X2=0.737 $Y2=1.16
cc_18 VNB N_VPWR_c_228_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_270_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_VGND_c_271_n 0.0325477f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_21 VNB N_VGND_c_272_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.737 $Y2=1.475
cc_22 VNB N_VGND_c_273_n 0.0177718f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=1.582
cc_23 VNB N_VGND_c_274_n 0.0171188f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.485
cc_24 VNB N_VGND_c_275_n 0.164518f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.4
cc_25 VNB N_VGND_c_276_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=1.66
cc_26 VNB N_VGND_c_277_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_27 VNB N_A_297_47#_c_310_n 0.0138983f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_28 VNB N_A_297_47#_c_311_n 0.0183573f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_29 VNB N_A_297_47#_c_312_n 0.00377637f $X=-0.19 $Y=-0.24 $X2=0.737 $Y2=1.16
cc_30 VPB N_A_79_21#_M1000_g 0.0248065f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_31 VPB N_A_79_21#_c_53_n 0.00294623f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_32 VPB N_A_79_21#_c_54_n 0.0100537f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_33 VPB N_A_79_21#_c_59_n 0.00422752f $X=-0.19 $Y=1.305 $X2=1.415 $Y2=1.582
cc_34 VPB N_A_79_21#_c_60_n 0.00398386f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=1.69
cc_35 VPB N_B1_M1002_g 0.0230031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_B1_c_109_n 0.00488313f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_37 VPB N_A2_M1004_g 0.0207348f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB A2 0.00269279f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_39 VPB N_A2_c_144_n 0.00564698f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_40 VPB N_A1_M1006_g 0.0205232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A1_c_183_n 0.0120094f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_42 VPB A1 0.0130423f $X=-0.19 $Y=1.305 $X2=0.737 $Y2=0.905
cc_43 VPB N_X_c_211_n 0.047502f $X=-0.19 $Y=1.305 $X2=0.737 $Y2=1.16
cc_44 VPB N_VPWR_c_229_n 0.00211789f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_45 VPB N_VPWR_c_230_n 0.0103102f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_46 VPB N_VPWR_c_231_n 0.0251685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_232_n 0.0155059f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_48 VPB N_VPWR_c_233_n 0.0276998f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=2.34
cc_49 VPB N_VPWR_c_234_n 0.0111749f $X=-0.19 $Y=1.305 $X2=1.2 $Y2=0.74
cc_50 VPB N_VPWR_c_228_n 0.0432594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 N_A_79_21#_M1000_g N_B1_M1002_g 0.00779362f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_52 N_A_79_21#_c_59_n N_B1_M1002_g 0.0182983f $X=1.415 $Y=1.582 $X2=0 $Y2=0
cc_53 N_A_79_21#_c_53_n N_B1_c_109_n 0.00584643f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_54 N_A_79_21#_c_54_n N_B1_c_109_n 0.00894747f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_79_21#_c_59_n N_B1_c_109_n 0.00121736f $X=1.415 $Y=1.582 $X2=0 $Y2=0
cc_56 N_A_79_21#_c_60_n N_B1_c_109_n 0.00242985f $X=1.58 $Y=1.69 $X2=0 $Y2=0
cc_57 N_A_79_21#_c_55_n N_B1_c_109_n 0.00254116f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_58 N_A_79_21#_c_53_n N_B1_c_110_n 0.0182545f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_79_21#_c_54_n N_B1_c_110_n 8.06426e-19 $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_79_21#_c_59_n N_B1_c_110_n 0.0260672f $X=1.415 $Y=1.582 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_60_n N_B1_c_110_n 0.00999421f $X=1.58 $Y=1.69 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_55_n N_B1_c_110_n 0.0211872f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_53_n N_B1_c_111_n 0.00240138f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_55_n N_B1_c_111_n 0.00720802f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_55_n N_A2_c_142_n 8.41953e-19 $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_60_n A2 0.00372259f $X=1.58 $Y=1.69 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_60_n N_A2_c_144_n 2.43595e-19 $X=1.58 $Y=1.69 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_52_n N_X_c_209_n 0.00855649f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_55_n N_X_c_209_n 0.0133645f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_52_n N_X_c_210_n 0.00367098f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_53_n N_X_c_210_n 0.00957984f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_54_n N_X_c_210_n 0.00270383f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_79_21#_M1000_g N_X_c_211_n 0.00372063f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_53_n N_X_c_211_n 0.0279843f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_54_n N_X_c_211_n 0.00861623f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_86_p N_X_c_211_n 6.35484e-19 $X=0.88 $Y=1.582 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_59_n N_VPWR_M1000_d 0.00468864f $X=1.415 $Y=1.582 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_79_21#_c_86_p N_VPWR_M1000_d 0.00542943f $X=0.88 $Y=1.582 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_79_21#_M1000_g N_VPWR_c_229_n 0.0149022f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_54_n N_VPWR_c_229_n 7.70146e-19 $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_59_n N_VPWR_c_229_n 0.0251727f $X=1.415 $Y=1.582 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_86_p N_VPWR_c_229_n 0.0232617f $X=0.88 $Y=1.582 $X2=0 $Y2=0
cc_83 N_A_79_21#_M1000_g N_VPWR_c_232_n 0.0046653f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_94_p N_VPWR_c_233_n 0.0212535f $X=1.58 $Y=2.34 $X2=0 $Y2=0
cc_85 N_A_79_21#_M1002_d N_VPWR_c_228_n 0.00524128f $X=1.37 $Y=1.485 $X2=0 $Y2=0
cc_86 N_A_79_21#_M1000_g N_VPWR_c_228_n 0.00886468f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_94_p N_VPWR_c_228_n 0.0126319f $X=1.58 $Y=2.34 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_55_n N_VGND_M1007_d 0.00365741f $X=1.2 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_79_21#_c_52_n N_VGND_c_270_n 0.00438629f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_54_n N_VGND_c_270_n 7.01852e-19 $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_55_n N_VGND_c_270_n 0.0318141f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_55_n N_VGND_c_271_n 0.0270574f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_52_n N_VGND_c_273_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_79_21#_M1001_s N_VGND_c_275_n 0.00209319f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_c_52_n N_VGND_c_275_n 0.0117818f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_55_n N_VGND_c_275_n 0.0209875f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_60_n N_A_297_47#_c_312_n 0.00638412f $X=1.58 $Y=1.69 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_55_n N_A_297_47#_c_312_n 0.0015618f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_99 N_B1_M1002_g N_A2_M1004_g 0.021201f $X=1.295 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B1_c_111_n N_A2_c_142_n 0.0213706f $X=1.362 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_c_109_n A2 6.49952e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B1_c_110_n A2 0.0187037f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B1_c_109_n N_A2_c_144_n 0.01981f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B1_c_110_n N_A2_c_144_n 9.25913e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B1_M1002_g N_VPWR_c_229_n 0.0128132f $X=1.295 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B1_M1002_g N_VPWR_c_233_n 0.00486043f $X=1.295 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B1_M1002_g N_VPWR_c_228_n 0.00857998f $X=1.295 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B1_c_111_n N_VGND_c_270_n 0.00194637f $X=1.362 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B1_c_111_n N_VGND_c_271_n 0.00539841f $X=1.362 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B1_c_111_n N_VGND_c_275_n 0.0111166f $X=1.362 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B1_c_109_n N_A_297_47#_c_312_n 2.49375e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B1_c_110_n N_A_297_47#_c_312_n 0.00315292f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A2_c_142_n N_A1_c_181_n 0.0266571f $X=1.87 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_114 A2 N_A1_c_182_n 0.0145078f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A2_M1004_g N_A1_c_183_n 0.042447f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_116 A2 N_A1_c_183_n 0.0158285f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A2_c_144_n N_A1_c_183_n 0.0217242f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_118 A2 A1 0.0177041f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_119 N_A2_M1004_g N_VPWR_c_229_n 0.00110024f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A2_M1004_g N_VPWR_c_231_n 0.00145653f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_121 A2 N_VPWR_c_231_n 0.0342467f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A2_M1004_g N_VPWR_c_233_n 0.00585385f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_123 A2 N_VPWR_c_233_n 0.00952185f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A2_M1004_g N_VPWR_c_228_n 0.011145f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_125 A2 N_VPWR_c_228_n 0.00795591f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_126 A2 A_382_297# 0.0200344f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_127 N_A2_c_142_n N_VGND_c_271_n 0.00434208f $X=1.87 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A2_c_142_n N_VGND_c_272_n 0.00268723f $X=1.87 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_142_n N_VGND_c_275_n 0.00602168f $X=1.87 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A2_c_142_n N_A_297_47#_c_310_n 0.00885038f $X=1.87 $Y=0.995 $X2=0 $Y2=0
cc_131 A2 N_A_297_47#_c_310_n 0.00850238f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A2_c_144_n N_A_297_47#_c_310_n 0.001482f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A2_c_142_n N_A_297_47#_c_311_n 7.01622e-19 $X=1.87 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A2_c_142_n N_A_297_47#_c_312_n 0.00317768f $X=1.87 $Y=0.995 $X2=0 $Y2=0
cc_135 A2 N_A_297_47#_c_312_n 0.0240965f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A2_c_144_n N_A_297_47#_c_312_n 0.00164575f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_137 A1 N_VPWR_M1006_d 0.00478094f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_138 N_A1_M1006_g N_VPWR_c_231_n 0.0139319f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_c_182_n N_VPWR_c_231_n 0.00177857f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A1_c_183_n N_VPWR_c_231_n 0.0021218f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_141 A1 N_VPWR_c_231_n 0.0128236f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_142 N_A1_M1006_g N_VPWR_c_233_n 0.0046653f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A1_M1006_g N_VPWR_c_228_n 0.00808301f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A1_c_181_n N_VGND_c_272_n 0.00268723f $X=2.29 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A1_c_181_n N_VGND_c_274_n 0.00422241f $X=2.29 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A1_c_181_n N_VGND_c_275_n 0.00667797f $X=2.29 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A1_c_181_n N_A_297_47#_c_310_n 0.0142466f $X=2.29 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A1_c_182_n N_A_297_47#_c_310_n 0.0281343f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A1_c_183_n N_A_297_47#_c_310_n 0.00724435f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A1_c_181_n N_A_297_47#_c_311_n 0.00630897f $X=2.29 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_181_n N_A_297_47#_c_312_n 2.32235e-19 $X=2.29 $Y=0.995 $X2=0 $Y2=0
cc_152 N_X_c_211_n N_VPWR_c_232_n 0.0194075f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_153 N_X_M1000_s N_VPWR_c_228_n 0.00399293f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_154 N_X_c_211_n N_VPWR_c_228_n 0.0107063f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_155 N_X_c_209_n N_VGND_c_273_n 0.0217551f $X=0.26 $Y=0.395 $X2=0 $Y2=0
cc_156 N_X_M1007_s N_VGND_c_275_n 0.00209319f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_157 N_X_c_209_n N_VGND_c_275_n 0.0128119f $X=0.26 $Y=0.395 $X2=0 $Y2=0
cc_158 N_VPWR_c_228_n A_382_297# 0.00562644f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_159 N_VGND_c_275_n N_A_297_47#_M1001_d 0.00393089f $X=2.53 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_160 N_VGND_c_275_n N_A_297_47#_M1003_d 0.00209319f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_161 N_VGND_M1005_d N_A_297_47#_c_310_n 0.00162148f $X=1.945 $Y=0.235 $X2=0
+ $Y2=0
cc_162 N_VGND_c_271_n N_A_297_47#_c_310_n 0.00203746f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_163 N_VGND_c_272_n N_A_297_47#_c_310_n 0.0122675f $X=2.08 $Y=0.38 $X2=0 $Y2=0
cc_164 N_VGND_c_274_n N_A_297_47#_c_310_n 0.00203746f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_165 N_VGND_c_275_n N_A_297_47#_c_310_n 0.00845923f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_166 N_VGND_c_274_n N_A_297_47#_c_311_n 0.0216897f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_167 N_VGND_c_275_n N_A_297_47#_c_311_n 0.0127966f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_168 N_VGND_c_271_n N_A_297_47#_c_312_n 0.00505518f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_169 N_VGND_c_275_n N_A_297_47#_c_312_n 0.00936078f $X=2.53 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nor2_8.spice
* Created: Thu Aug 27 14:31:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor2_8.pex.spice"
.subckt sky130_fd_sc_hd__nor2_8  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_Y_M1004_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75006.5 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1004_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75006.1 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75005.6 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1008_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75005.2 A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1012_d N_A_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1021 N_Y_M1017_d N_A_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1007_d N_B_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1018_d N_B_M1018_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1018_d N_B_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.8
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1024 N_Y_M1024_d N_B_M1024_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1025 N_Y_M1024_d N_B_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1026 N_Y_M1026_d N_B_M1026_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1028 N_Y_M1026_d N_B_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_297#_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75006.5 A=0.15 P=2.3 MULT=1
MM1003 N_A_27_297#_M1003_d N_A_M1003_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75006.1 A=0.15 P=2.3 MULT=1
MM1009 N_A_27_297#_M1003_d N_A_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75005.7 A=0.15 P=2.3 MULT=1
MM1010 N_A_27_297#_M1010_d N_A_M1010_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1014 N_A_27_297#_M1010_d N_A_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1019 N_A_27_297#_M1019_d N_A_M1019_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1020 N_A_27_297#_M1019_d N_A_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1029 N_A_27_297#_M1029_d N_A_M1029_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_A_27_297#_M1029_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1000_d N_B_M1002_g N_A_27_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1005_d N_B_M1005_g N_A_27_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1016 N_Y_M1005_d N_B_M1016_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.8
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1022 N_Y_M1022_d N_B_M1022_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1027 N_Y_M1022_d N_B_M1027_g N_A_27_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.7
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1030 N_Y_M1030_d N_B_M1030_g N_A_27_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1031 N_Y_M1030_d N_B_M1031_g N_A_27_297#_M1031_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=12.4227 P=18.69
*
.include "sky130_fd_sc_hd__nor2_8.pxi.spice"
*
.ends
*
*

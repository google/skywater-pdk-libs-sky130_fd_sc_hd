* File: sky130_fd_sc_hd__einvp_4.spice
* Created: Thu Aug 27 14:20:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__einvp_4.spice.pex"
.subckt sky130_fd_sc_hd__einvp_4  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_TE_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1015_d N_TE_M1003_g N_A_193_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.09425 PD=0.92 PS=0.94 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75000.6
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_TE_M1007_g N_A_193_47#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.09425 PD=0.92 PS=0.94 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1007_d N_TE_M1009_g N_A_193_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_TE_M1010_g N_A_193_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_Z_M1013_d N_A_M1013_g N_A_193_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1014 N_Z_M1013_d N_A_M1014_g N_A_193_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1016 N_Z_M1016_d N_A_M1016_g N_A_193_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_Z_M1016_d N_A_M1017_g N_A_193_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_TE_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_215_309#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.2444 AS=0.1269 PD=2.4 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667 SA=75000.2
+ SB=75003.2 A=0.141 P=2.18 MULT=1
MM1001 N_A_215_309#_M1001_d N_A_27_47#_M1001_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75000.6 SB=75002.8 A=0.141 P=2.18 MULT=1
MM1002 N_A_215_309#_M1001_d N_A_27_47#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667 SA=75001
+ SB=75002.3 A=0.141 P=2.18 MULT=1
MM1006 N_A_215_309#_M1006_d N_A_27_47#_M1006_g N_VPWR_M1002_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.155294 AS=0.1269 PD=1.28402 PS=1.21 NRD=5.2205 NRS=0 M=1 R=6.26667
+ SA=75001.4 SB=75001.9 A=0.141 P=2.18 MULT=1
MM1004 N_Z_M1004_d N_A_M1004_g N_A_215_309#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.165206 PD=1.27 PS=1.36598 NRD=0 NRS=3.9203 M=1 R=6.66667
+ SA=75001.8 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1005 N_Z_M1004_d N_A_M1005_g N_A_215_309#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1008 N_Z_M1008_d N_A_M1008_g N_A_215_309#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_Z_M1008_d N_A_M1012_g N_A_215_309#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=8.7312 P=14.09
c_44 VNB 0 8.32198e-20 $X=0.15 $Y=-0.085
c_82 VPB 0 1.1096e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__einvp_4.spice.SKY130_FD_SC_HD__EINVP_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__ebufn_4.spice
* Created: Thu Aug 27 14:19:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__ebufn_4.spice.pex"
.subckt sky130_fd_sc_hd__ebufn_4  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_27_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121875 AS=0.169 PD=1.025 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_A_214_47#_M1014_d N_TE_B_M1014_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.121875 PD=1.82 PS=1.025 NRD=0 NRS=18.456 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_214_47#_M1003_g N_A_393_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1003_d N_A_214_47#_M1004_g N_A_393_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_214_47#_M1005_g N_A_393_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1005_d N_A_214_47#_M1006_g N_A_393_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75001.4 SB=75002 A=0.0975 P=1.6 MULT=1
MM1007 N_Z_M1007_d N_A_27_47#_M1007_g N_A_393_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75002 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1008 N_Z_M1007_d N_A_27_47#_M1008_g N_A_393_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.4 SB=75001 A=0.0975 P=1.6 MULT=1
MM1010 N_Z_M1010_d N_A_27_47#_M1010_g N_A_393_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.8 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_Z_M1010_d N_A_27_47#_M1015_g N_A_393_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_27_47#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1875 AS=0.26 PD=1.375 PS=2.52 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1002 N_A_214_47#_M1002_d N_TE_B_M1002_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1875 PD=2.52 PS=1.375 NRD=0 NRS=11.8003 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_TE_B_M1000_g N_A_320_309#_M1000_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.2444 PD=1.21 PS=2.4 NRD=0 NRS=0 M=1 R=6.26667 SA=75000.2
+ SB=75003.6 A=0.141 P=2.18 MULT=1
MM1011 N_VPWR_M1000_d N_TE_B_M1011_g N_A_320_309#_M1011_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75000.6 SB=75003.2 A=0.141 P=2.18 MULT=1
MM1016 N_VPWR_M1016_d N_TE_B_M1016_g N_A_320_309#_M1011_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667 SA=75001
+ SB=75002.8 A=0.141 P=2.18 MULT=1
MM1019 N_VPWR_M1016_d N_TE_B_M1019_g N_A_320_309#_M1019_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.363644 PD=1.21 PS=1.70072 NRD=0 NRS=17.8088 M=1
+ R=6.26667 SA=75001.4 SB=75002.4 A=0.141 P=2.18 MULT=1
MM1001 N_A_320_309#_M1019_s N_A_27_47#_M1001_g N_Z_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.386856 AS=0.135 PD=1.80928 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75002.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1009 N_A_320_309#_M1009_d N_A_27_47#_M1009_g N_Z_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1012 N_A_320_309#_M1009_d N_A_27_47#_M1012_g N_Z_M1012_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_A_320_309#_M1017_d N_A_27_47#_M1017_g N_Z_M1012_s VPB PHIGHVT L=0.15
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_54 VNB 0 1.48146e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__ebufn_4.spice.SKY130_FD_SC_HD__EBUFN_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__buf_4.pex.spice
* Created: Tue Sep  1 18:59:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUF_4%A 3 7 9 15
c31 9 0 1.40316e-19 $X=0.235 $Y=1.19
r32 12 15 34.1305 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.16
+ $X2=0.47 $Y2=1.16
r33 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.305
+ $Y=1.16 $X2=0.305 $Y2=1.16
r34 5 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r35 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=1.985
r36 1 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r37 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 39 41 45
+ 47 48 49 52 54 57 62 68
c106 68 0 1.40316e-19 $X=2.15 $Y=1.16
r107 67 68 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=2.15 $Y2=1.16
r108 66 67 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r109 58 66 74.4282 $w=2.7e-07 $l=3.35e-07 $layer=POLY_cond $X=0.975 $Y=1.16
+ $X2=1.31 $Y2=1.16
r110 58 63 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=0.975 $Y=1.16
+ $X2=0.89 $Y2=1.16
r111 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.16 $X2=0.975 $Y2=1.16
r112 55 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=1.16
+ $X2=0.725 $Y2=1.16
r113 55 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=1.16
+ $X2=0.975 $Y2=1.16
r114 53 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.245
+ $X2=0.725 $Y2=1.16
r115 53 54 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.725 $Y=1.245
+ $X2=0.725 $Y2=1.485
r116 52 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.075
+ $X2=0.725 $Y2=1.16
r117 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.725 $Y=0.905
+ $X2=0.725 $Y2=1.075
r118 50 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.57
+ $X2=0.26 $Y2=1.57
r119 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.64 $Y=1.57
+ $X2=0.725 $Y2=1.485
r120 49 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.64 $Y=1.57
+ $X2=0.425 $Y2=1.57
r121 47 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.64 $Y=0.82
+ $X2=0.725 $Y2=0.905
r122 47 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.64 $Y=0.82
+ $X2=0.345 $Y2=0.82
r123 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.345 $Y2=0.82
r124 43 45 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.56
r125 39 61 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.655
+ $X2=0.26 $Y2=1.57
r126 39 41 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.26 $Y=1.655
+ $X2=0.26 $Y2=2.31
r127 35 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r128 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r129 31 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r130 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r131 27 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r132 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r133 23 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r134 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r135 19 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r136 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r137 15 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r138 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r139 11 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r140 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r141 7 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.16
r142 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r143 2 61 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r144 2 41 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r145 1 45 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_4%VPWR 1 2 3 12 16 18 20 25 26 27 29 31 41 46 50
r46 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 41 49 4.52492 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.477 $Y2=2.72
r51 41 43 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 40 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 40 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 37 46 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=0.715 $Y2=2.72
r56 37 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 31 46 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.715 $Y2=2.72
r58 29 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 27 31 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.595 $Y2=2.72
r60 27 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r61 25 39 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.52 $Y2=2.72
r63 24 43 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=2.07 $Y2=2.72
r64 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.52 $Y2=2.72
r65 20 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.36 $Y=1.66
+ $X2=2.36 $Y2=2.34
r66 18 49 3.24126 $w=3.3e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.477 $Y2=2.72
r67 18 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.34
r68 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r69 14 16 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2
r70 10 46 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.72
r71 10 12 30.4917 $w=2.38e-07 $l=6.35e-07 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2
r72 3 23 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.34
r73 3 20 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.66
r74 2 16 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2
r75 1 12 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_4%X 1 2 3 4 15 19 23 27 29 30 31 32 33
r44 32 33 5.39369 $w=6.63e-07 $l=2.55e-07 $layer=LI1_cond $X=1.777 $Y=1.19
+ $X2=1.777 $Y2=1.445
r45 31 41 2.86771 $w=3.32e-07 $l=8.5e-08 $layer=LI1_cond $X=1.777 $Y=0.82
+ $X2=1.777 $Y2=0.905
r46 31 32 6.52406 $w=4.93e-07 $l=2.7e-07 $layer=LI1_cond $X=1.777 $Y=0.92
+ $X2=1.777 $Y2=1.19
r47 31 41 0.362448 $w=4.93e-07 $l=1.5e-08 $layer=LI1_cond $X=1.777 $Y=0.92
+ $X2=1.777 $Y2=0.905
r48 30 33 13.1335 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=1.185 $Y=1.53
+ $X2=1.53 $Y2=1.53
r49 29 31 14.1322 $w=3.08e-07 $l=3.45e-07 $layer=LI1_cond $X=1.185 $Y=0.82
+ $X2=1.53 $Y2=0.82
r50 25 33 2.86771 $w=3.32e-07 $l=2.01057e-07 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=1.777 $Y2=1.53
r51 25 27 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=1.94 $Y2=1.755
r52 21 31 2.86771 $w=3.32e-07 $l=2.01057e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.777 $Y2=0.82
r53 21 23 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.56
r54 17 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.1 $Y=1.615
+ $X2=1.185 $Y2=1.53
r55 17 19 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.1 $Y=1.615 $X2=1.1
+ $Y2=1.755
r56 13 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.185 $Y2=0.82
r57 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.1 $Y2=0.56
r58 4 27 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.755
r59 3 19 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.755
r60 2 23 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.56
r61 1 15 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_4%VGND 1 2 3 12 16 18 20 23 24 26 27 28 30 40 46
r48 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r49 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r50 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r51 40 45 4.52492 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.477
+ $Y2=0
r52 40 42 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.07
+ $Y2=0
r53 39 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r54 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r55 30 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r56 28 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r57 26 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.15
+ $Y2=0
r58 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.52
+ $Y2=0
r59 25 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=2.07
+ $Y2=0
r60 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.52
+ $Y2=0
r61 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.23
+ $Y2=0
r62 23 24 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.645
+ $Y2=0
r63 22 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=1.15
+ $Y2=0
r64 22 24 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.645
+ $Y2=0
r65 18 45 3.24126 $w=3.3e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.477 $Y2=0
r66 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.38
r67 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r68 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.4
r69 10 24 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=0.085
+ $X2=0.645 $Y2=0
r70 10 12 15.1258 $w=2.38e-07 $l=3.15e-07 $layer=LI1_cond $X=0.645 $Y=0.085
+ $X2=0.645 $Y2=0.4
r71 3 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.38
r72 2 16 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r73 1 12 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends


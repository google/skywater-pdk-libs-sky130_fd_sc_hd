* File: sky130_fd_sc_hd__dlrtn_4.pex.spice
* Created: Tue Sep  1 19:05:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRTN_4%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%A_27_47# 1 2 9 13 17 20 24 28 29 30 38 42 45
+ 47 52 54 56 57 60 63 64 68 71 75 79
c167 20 0 1.41946e-19 $X=3.34 $Y=2.275
c168 13 0 2.6965e-20 $X=0.89 $Y=2.135
c169 9 0 2.6965e-20 $X=0.89 $Y=0.445
r170 64 79 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.1 $Y=1.53
+ $X2=3.1 $Y2=1.415
r171 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.02 $Y=1.53
+ $X2=3.02 $Y2=1.53
r172 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r173 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.875 $Y=1.53
+ $X2=3.02 $Y2=1.53
r175 56 57 2.51856 $w=1.4e-07 $l=2.035e-06 $layer=MET1_cond $X=2.875 $Y=1.53
+ $X2=0.84 $Y2=1.53
r176 52 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=0.87
+ $X2=2.805 $Y2=0.705
r177 51 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.805 $Y=0.87
+ $X2=3.015 $Y2=0.87
r178 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=0.87 $X2=2.805 $Y2=0.87
r179 49 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r180 48 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r181 46 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r182 45 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r183 45 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r184 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r185 39 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=3.185 $Y=1.74
+ $X2=3.34 $Y2=1.74
r186 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.74 $X2=3.185 $Y2=1.74
r187 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.1 $Y=1.585
+ $X2=3.1 $Y2=1.53
r188 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.1 $Y=1.585
+ $X2=3.1 $Y2=1.74
r189 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=1.035
+ $X2=3.015 $Y2=0.87
r190 34 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.015 $Y=1.035
+ $X2=3.015 $Y2=1.415
r191 32 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r192 31 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r193 30 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r194 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r195 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r196 28 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r197 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r198 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r199 18 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.34 $Y=1.875
+ $X2=3.34 $Y2=1.74
r200 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.34 $Y=1.875
+ $X2=3.34 $Y2=2.275
r201 17 71 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.795 $Y=0.415
+ $X2=2.795 $Y2=0.705
r202 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r203 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r204 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r205 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r206 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r207 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.63 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.63 $Y=1.04
+ $X2=1.835 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.04 $X2=1.63 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.63 $Y=1.19 $X2=1.63
+ $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.205
+ $X2=1.835 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.835 $Y=1.205
+ $X2=1.835 $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=0.875
+ $X2=1.835 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.835 $Y=0.875
+ $X2=1.835 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%A_300_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c83 32 0 1.12109e-19 $X=2.26 $Y=0.93
c84 18 0 7.13094e-20 $X=1.975 $Y=0.7
r85 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=0.93
+ $X2=2.26 $Y2=1.095
r86 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=0.93
+ $X2=2.26 $Y2=0.765
r87 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=0.93 $X2=2.26 $Y2=0.93
r88 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.625 $Y=0.51
+ $X2=1.625 $Y2=0.7
r89 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.06 $Y=1.095
+ $X2=2.16 $Y2=0.93
r90 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.06 $Y=1.095 $X2=2.06
+ $Y2=1.495
r91 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.975 $Y=1.58
+ $X2=2.06 $Y2=1.495
r92 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.975 $Y=1.58
+ $X2=1.79 $Y2=1.58
r93 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.7
+ $X2=1.625 $Y2=0.7
r94 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.975 $Y=0.7
+ $X2=2.16 $Y2=0.93
r95 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.975 $Y=0.7
+ $X2=1.71 $Y2=0.7
r96 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=1.79 $Y2=1.58
r97 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=1.625 $Y2=1.99
r98 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.255 $Y=2.165
+ $X2=2.255 $Y2=1.095
r99 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.255 $Y=0.445
+ $X2=2.255 $Y2=0.765
r100 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.845 $X2=1.625 $Y2=1.99
r101 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.235 $X2=1.625 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%A_193_47# 1 2 9 11 12 15 19 22 24 26 27 30
+ 33 37 38
c113 38 0 1.41946e-19 $X=2.675 $Y=1.52
r114 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.52 $X2=2.675 $Y2=1.52
r115 34 38 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.617 $Y=1.87
+ $X2=2.617 $Y2=1.52
r116 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.56 $Y=1.87
+ $X2=2.56 $Y2=1.87
r117 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r118 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r119 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.415 $Y=1.87
+ $X2=2.56 $Y2=1.87
r120 26 27 1.37995 $w=1.4e-07 $l=1.115e-06 $layer=MET1_cond $X=2.415 $Y=1.87
+ $X2=1.3 $Y2=1.87
r121 24 30 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r122 24 25 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r123 22 25 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r124 18 37 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.675 $Y=1.55
+ $X2=2.675 $Y2=1.52
r125 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.675 $Y=1.55
+ $X2=2.675 $Y2=1.685
r126 17 37 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.675 $Y=1.395
+ $X2=2.675 $Y2=1.52
r127 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.225 $Y=1.245
+ $X2=3.225 $Y2=0.415
r128 12 17 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.81 $Y=1.32
+ $X2=2.675 $Y2=1.395
r129 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.15 $Y=1.32
+ $X2=3.225 $Y2=1.245
r130 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.15 $Y=1.32
+ $X2=2.81 $Y2=1.32
r131 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.685
r132 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r133 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%A_725_21# 1 2 9 13 15 17 20 22 24 27 29 31
+ 34 36 38 41 43 46 50 52 53 56 58 63 66 75
c153 75 0 1.81835e-20 $X=6.89 $Y=1.16
r154 74 75 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=6.43 $Y=1.16
+ $X2=6.89 $Y2=1.16
r155 73 74 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=5.995 $Y=1.16
+ $X2=6.43 $Y2=1.16
r156 64 73 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=5.54 $Y=1.16
+ $X2=5.995 $Y2=1.16
r157 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.54
+ $Y=1.16 $X2=5.54 $Y2=1.16
r158 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.54 $Y=1.535
+ $X2=5.54 $Y2=1.16
r159 60 63 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.54 $Y=0.825
+ $X2=5.54 $Y2=1.16
r160 59 66 4.08801 $w=2.5e-07 $l=1.28938e-07 $layer=LI1_cond $X=4.945 $Y=1.62
+ $X2=4.85 $Y2=1.7
r161 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=1.62
+ $X2=5.54 $Y2=1.535
r162 58 59 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.455 $Y=1.62
+ $X2=4.945 $Y2=1.62
r163 54 66 2.34704 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=1.865
+ $X2=4.85 $Y2=1.7
r164 54 56 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=4.85 $Y=1.865
+ $X2=4.85 $Y2=2.27
r165 52 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=0.74
+ $X2=5.54 $Y2=0.825
r166 52 53 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.455 $Y=0.74
+ $X2=4.595 $Y2=0.74
r167 48 53 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=4.42 $Y=0.655
+ $X2=4.595 $Y2=0.74
r168 48 50 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.42 $Y=0.655
+ $X2=4.42 $Y2=0.4
r169 46 67 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.93 $Y=1.7 $X2=3.7
+ $Y2=1.7
r170 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.7 $X2=3.93 $Y2=1.7
r171 43 66 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.755 $Y=1.7
+ $X2=4.85 $Y2=1.7
r172 43 45 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.755 $Y=1.7
+ $X2=3.93 $Y2=1.7
r173 39 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.16
r174 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.985
r175 36 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=1.16
r176 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=0.56
r177 32 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.16
r178 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.985
r179 29 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=1.16
r180 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=0.56
r181 25 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.16
r182 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.985
r183 22 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=1.16
r184 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=0.56
r185 18 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=1.325
+ $X2=5.54 $Y2=1.16
r186 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.54 $Y=1.325
+ $X2=5.54 $Y2=1.985
r187 15 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=0.995
+ $X2=5.54 $Y2=1.16
r188 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.54 $Y=0.995
+ $X2=5.54 $Y2=0.56
r189 11 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.7 $Y=1.865
+ $X2=3.7 $Y2=1.7
r190 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.7 $Y=1.865
+ $X2=3.7 $Y2=2.275
r191 7 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.7 $Y=1.535
+ $X2=3.7 $Y2=1.7
r192 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.7 $Y=1.535 $X2=3.7
+ $Y2=0.445
r193 2 66 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=1.485 $X2=4.85 $Y2=1.755
r194 2 56 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=1.485 $X2=4.85 $Y2=2.27
r195 1 50 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.235 $X2=4.43 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%A_562_413# 1 2 9 13 15 16 17 21 26 28 29 31
c86 31 0 1.0585e-19 $X=4.15 $Y=1.16
c87 29 0 1.65126e-19 $X=3.655 $Y=1.175
r88 34 35 6.98473 $w=2.62e-07 $l=1.5e-07 $layer=LI1_cond $X=3.42 $Y=1.175
+ $X2=3.57 $Y2=1.175
r89 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.15
+ $Y=1.16 $X2=4.15 $Y2=1.16
r90 29 35 3.68445 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=1.175 $X2=3.57
+ $Y2=1.175
r91 29 31 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=3.655 $Y=1.175
+ $X2=4.15 $Y2=1.175
r92 27 35 3.26844 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=1.175
r93 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=2.255
r94 26 34 3.26844 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.42 $Y=1.025
+ $X2=3.42 $Y2=1.175
r95 25 26 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.42 $Y=0.535
+ $X2=3.42 $Y2=1.025
r96 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.485 $Y=2.34
+ $X2=3.57 $Y2=2.255
r97 21 23 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.485 $Y=2.34
+ $X2=3.07 $Y2=2.34
r98 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.45
+ $X2=3.42 $Y2=0.535
r99 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.335 $Y=0.45
+ $X2=3.01 $Y2=0.45
r100 15 32 92.2021 $w=2.7e-07 $l=4.15e-07 $layer=POLY_cond $X=4.565 $Y=1.16
+ $X2=4.15 $Y2=1.16
r101 15 16 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.565 $Y=1.16
+ $X2=4.64 $Y2=1.16
r102 11 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.64 $Y=1.295
+ $X2=4.64 $Y2=1.16
r103 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.64 $Y=1.295
+ $X2=4.64 $Y2=1.985
r104 7 16 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.64 $Y=1.025
+ $X2=4.64 $Y2=1.16
r105 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.64 $Y=1.025
+ $X2=4.64 $Y2=0.56
r106 2 23 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.065 $X2=3.07 $Y2=2.34
r107 1 19 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.235 $X2=3.01 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%RESET_B 1 3 6 8 11 12
c40 11 0 1.0585e-19 $X=5.06 $Y=1.16
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.06
+ $Y=1.16 $X2=5.06 $Y2=1.16
r42 8 12 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.88 $Y=1.16 $X2=5.06
+ $Y2=1.16
r43 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=1.325
+ $X2=5.06 $Y2=1.16
r44 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.06 $Y=1.325 $X2=5.06
+ $Y2=1.985
r45 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=0.995
+ $X2=5.06 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.06 $Y=0.995 $X2=5.06
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%VPWR 1 2 3 4 5 6 7 24 28 32 34 38 42 44 48
+ 52 54 58 60 65 70 78 83 89 92 95 98 101 104 108
c122 42 0 1.81835e-20 $X=5.3 $Y=2.02
r123 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r124 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r125 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r126 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r127 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r128 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r129 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r130 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r131 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r132 87 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r133 87 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r134 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r135 84 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.405 $Y=2.72
+ $X2=6.27 $Y2=2.72
r136 84 86 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.405 $Y=2.72
+ $X2=6.67 $Y2=2.72
r137 83 107 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=7.152 $Y2=2.72
r138 83 86 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=6.67 $Y2=2.72
r139 82 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r140 82 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r142 79 98 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.585 $Y=2.72
+ $X2=4.445 $Y2=2.72
r143 79 81 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.585 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 78 101 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.115 $Y=2.72
+ $X2=5.3 $Y2=2.72
r145 78 81 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.115 $Y=2.72
+ $X2=4.83 $Y2=2.72
r146 77 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r147 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r148 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r149 74 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r150 73 76 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r151 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r152 71 92 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.117 $Y2=2.72
r153 71 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.53 $Y2=2.72
r154 70 95 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.97 $Y2=2.72
r155 70 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.45 $Y2=2.72
r156 69 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r157 69 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r158 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r159 66 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r160 66 68 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r161 65 92 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.96 $Y=2.72
+ $X2=2.117 $Y2=2.72
r162 65 68 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.96 $Y=2.72
+ $X2=1.61 $Y2=2.72
r163 60 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r164 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r165 58 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r166 58 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r167 54 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.11 $Y=1.66
+ $X2=7.11 $Y2=2.34
r168 52 107 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=7.11 $Y=2.635
+ $X2=7.152 $Y2=2.72
r169 52 57 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.11 $Y=2.635
+ $X2=7.11 $Y2=2.34
r170 48 51 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.27 $Y=1.66
+ $X2=6.27 $Y2=2.34
r171 46 104 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=2.635
+ $X2=6.27 $Y2=2.72
r172 46 51 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.27 $Y=2.635
+ $X2=6.27 $Y2=2.34
r173 45 101 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.3 $Y2=2.72
r174 44 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.135 $Y=2.72
+ $X2=6.27 $Y2=2.72
r175 44 45 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.135 $Y=2.72
+ $X2=5.485 $Y2=2.72
r176 40 101 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.72
r177 40 42 19.1555 $w=3.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.02
r178 36 98 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.445 $Y=2.635
+ $X2=4.445 $Y2=2.72
r179 36 38 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.445 $Y=2.635
+ $X2=4.445 $Y2=2.34
r180 35 95 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.115 $Y=2.72
+ $X2=3.97 $Y2=2.72
r181 34 98 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.445 $Y2=2.72
r182 34 35 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.115 $Y2=2.72
r183 30 95 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.72
r184 30 32 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=3.97 $Y=2.635
+ $X2=3.97 $Y2=2.3
r185 26 92 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.117 $Y=2.635
+ $X2=2.117 $Y2=2.72
r186 26 28 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.117 $Y=2.635
+ $X2=2.117 $Y2=2
r187 22 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r188 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r189 7 57 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=2.34
r190 7 54 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=1.66
r191 6 51 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.485 $X2=6.22 $Y2=2.34
r192 6 48 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.485 $X2=6.22 $Y2=1.66
r193 5 42 300 $w=1.7e-07 $l=6.11964e-07 $layer=licon1_PDIFF $count=2 $X=5.135
+ $Y=1.485 $X2=5.3 $Y2=2.02
r194 4 38 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.485 $X2=4.43 $Y2=2.34
r195 3 32 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.775
+ $Y=2.065 $X2=3.91 $Y2=2.3
r196 2 28 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.91
+ $Y=1.845 $X2=2.045 $Y2=2
r197 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%Q 1 2 3 4 14 19 24 26 27 29 30 31 33 35 50
+ 56
r60 50 59 2.13585 $w=5.58e-07 $l=1e-07 $layer=LI1_cond $X=6.575 $Y=1.045
+ $X2=6.675 $Y2=1.045
r61 33 35 9.82493 $w=5.58e-07 $l=4.6e-07 $layer=LI1_cond $X=6.72 $Y=1.045
+ $X2=7.18 $Y2=1.045
r62 33 59 0.961134 $w=5.58e-07 $l=4.5e-08 $layer=LI1_cond $X=6.72 $Y=1.045
+ $X2=6.675 $Y2=1.045
r63 33 59 6.84897 $w=2e-07 $l=2.8e-07 $layer=LI1_cond $X=6.675 $Y=0.765
+ $X2=6.675 $Y2=1.045
r64 33 56 11.2591 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=6.675 $Y=0.765
+ $X2=6.675 $Y2=0.49
r65 31 50 6.72794 $w=5.58e-07 $l=3.15e-07 $layer=LI1_cond $X=6.26 $Y=1.045
+ $X2=6.575 $Y2=1.045
r66 30 48 3.63929 $w=2.83e-07 $l=9e-08 $layer=LI1_cond $X=5.822 $Y=2.21
+ $X2=5.822 $Y2=2.3
r67 28 31 6.30077 $w=5.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.965 $Y=1.045
+ $X2=6.26 $Y2=1.045
r68 28 29 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=1.045
+ $X2=5.88 $Y2=1.045
r69 26 30 7.80426 $w=2.83e-07 $l=1.93e-07 $layer=LI1_cond $X=5.822 $Y=2.017
+ $X2=5.822 $Y2=2.21
r70 26 27 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=5.822 $Y=2.017
+ $X2=5.822 $Y2=1.875
r71 22 24 5.26115 $w=2.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.775 $Y=0.37
+ $X2=5.88 $Y2=0.37
r72 17 59 6.84897 $w=2e-07 $l=2.8e-07 $layer=LI1_cond $X=6.675 $Y=1.325
+ $X2=6.675 $Y2=1.045
r73 17 19 35.2136 $w=1.98e-07 $l=6.35e-07 $layer=LI1_cond $X=6.675 $Y=1.325
+ $X2=6.675 $Y2=1.96
r74 15 29 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=5.88 $Y=1.325
+ $X2=5.88 $Y2=1.045
r75 15 27 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.88 $Y=1.325
+ $X2=5.88 $Y2=1.875
r76 14 29 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=5.88 $Y=0.765
+ $X2=5.88 $Y2=1.045
r77 13 24 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.88 $Y=0.485
+ $X2=5.88 $Y2=0.37
r78 13 14 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.88 $Y=0.485
+ $X2=5.88 $Y2=0.765
r79 4 19 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=6.505
+ $Y=1.485 $X2=6.66 $Y2=1.96
r80 3 48 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.615
+ $Y=1.485 $X2=5.765 $Y2=2.3
r81 2 56 182 $w=1.7e-07 $l=3.23342e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.66 $Y2=0.49
r82 1 22 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=5.615
+ $Y=0.235 $X2=5.775 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DLRTN_4%VGND 1 2 3 4 5 6 21 25 29 33 35 39 41 43 45
+ 47 52 57 65 70 76 79 82 85 88 92
c126 92 0 2.71124e-20 $X=7.13 $Y=0
c127 2 0 7.13094e-20 $X=1.91 $Y=0.235
r128 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r129 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r130 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r131 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r132 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r133 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r134 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r135 74 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r136 74 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r137 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r138 71 88 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=6.27
+ $Y2=0
r139 71 73 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.405 $Y=0
+ $X2=6.67 $Y2=0
r140 70 91 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=7.152 $Y2=0
r141 70 73 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=6.67 $Y2=0
r142 69 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r143 69 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r144 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r145 66 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=0 $X2=3.91
+ $Y2=0
r146 66 68 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.075 $Y=0
+ $X2=4.83 $Y2=0
r147 65 85 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=5.27
+ $Y2=0
r148 65 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=4.83
+ $Y2=0
r149 64 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r150 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r151 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r152 61 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r153 60 63 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r154 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r155 58 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.045
+ $Y2=0
r156 58 60 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.53
+ $Y2=0
r157 57 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.91
+ $Y2=0
r158 57 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.45
+ $Y2=0
r159 56 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r160 56 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r161 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r162 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r163 53 55 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r164 52 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.045
+ $Y2=0
r165 52 55 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.61
+ $Y2=0
r166 47 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r167 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r168 45 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r169 45 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r170 41 91 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=7.11 $Y=0.085
+ $X2=7.152 $Y2=0
r171 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.11 $Y=0.085
+ $X2=7.11 $Y2=0.38
r172 37 88 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0
r173 37 39 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0.38
r174 36 85 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.27
+ $Y2=0
r175 35 88 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.135 $Y=0 $X2=6.27
+ $Y2=0
r176 35 36 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.135 $Y=0
+ $X2=5.44 $Y2=0
r177 31 85 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=0.085
+ $X2=5.27 $Y2=0
r178 31 33 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=5.27 $Y=0.085
+ $X2=5.27 $Y2=0.36
r179 27 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=0.085
+ $X2=3.91 $Y2=0
r180 27 29 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.91 $Y=0.085
+ $X2=3.91 $Y2=0.445
r181 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0
r182 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0.36
r183 19 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r184 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r185 6 43 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.965
+ $Y=0.235 $X2=7.1 $Y2=0.38
r186 5 39 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=6.07
+ $Y=0.235 $X2=6.22 $Y2=0.38
r187 4 33 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.135
+ $Y=0.235 $X2=5.275 $Y2=0.36
r188 3 29 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.775
+ $Y=0.235 $X2=3.91 $Y2=0.445
r189 2 25 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.235 $X2=2.045 $Y2=0.36
r190 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o211a_2.pex.spice
* Created: Thu Aug 27 14:34:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O211A_2%C1 3 6 7 10 12 13 15
c25 12 0 1.45172e-19 $X=0.327 $Y=0.995
r26 10 13 52.4268 $w=4.45e-07 $l=2.1e-07 $layer=POLY_cond $X=0.327 $Y=1.16
+ $X2=0.327 $Y2=1.37
r27 10 12 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.327 $Y=1.16
+ $X2=0.327 $Y2=0.995
r28 7 15 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.16 $X2=0.23
+ $Y2=1.16
r29 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r30 6 13 197.62 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.37
r31 3 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%B1 3 6 8 11 13
r33 11 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=0.93 $Y2=1.325
r34 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=0.93 $Y2=0.995
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.16 $X2=0.965 $Y2=1.16
r36 8 12 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=0.965 $Y2=1.16
r37 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.985
+ $X2=0.905 $Y2=1.325
r38 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.835 $Y=0.56
+ $X2=0.835 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%A2 3 6 7 10 12 13
r28 10 13 54.0123 $w=3.9e-07 $l=2.25e-07 $layer=POLY_cond $X=1.67 $Y=1.16
+ $X2=1.67 $Y2=1.385
r29 10 12 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.16
+ $X2=1.67 $Y2=0.995
r30 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.685
+ $Y=1.16 $X2=1.685 $Y2=1.16
r31 6 13 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.79 $Y=1.985 $X2=1.79
+ $Y2=1.385
r32 3 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.77 $Y=0.56 $X2=1.77
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%A1 3 7 8 11 12 13
r35 11 14 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=1.325
r36 11 13 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r38 8 12 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=1.16
+ $X2=2.24 $Y2=1.16
r39 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.2 $Y=0.56 $X2=2.2
+ $Y2=0.995
r40 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.985
+ $X2=2.15 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%A_27_47# 1 2 3 10 12 15 17 19 22 26 28 29 30
+ 31 34 36 39 40 42 50 56
c101 40 0 1.13771e-19 $X=2.665 $Y=1.16
r102 43 53 71.0206 $w=3.25e-07 $l=4e-07 $layer=POLY_cond $X=3.09 $Y=1.157
+ $X2=2.69 $Y2=1.157
r103 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.16 $X2=3.09 $Y2=1.16
r104 40 42 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.665 $Y=1.16
+ $X2=3.09 $Y2=1.16
r105 38 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.58 $Y=1.325
+ $X2=2.665 $Y2=1.16
r106 38 39 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.58 $Y=1.325
+ $X2=2.58 $Y2=1.51
r107 37 50 10.5328 $w=2.55e-07 $l=3.35e-07 $layer=LI1_cond $X=1.695 $Y=1.637
+ $X2=1.36 $Y2=1.637
r108 36 39 7.17723 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.495 $Y=1.637
+ $X2=2.58 $Y2=1.51
r109 36 37 36.1551 $w=2.53e-07 $l=8e-07 $layer=LI1_cond $X=2.495 $Y=1.637
+ $X2=1.695 $Y2=1.637
r110 32 50 1.77602 $w=6.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.36 $Y=1.765
+ $X2=1.36 $Y2=1.637
r111 32 34 2.23149 $w=6.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.36 $Y=1.765
+ $X2=1.36 $Y2=1.89
r112 30 50 10.5328 $w=2.55e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=1.637
+ $X2=1.36 $Y2=1.637
r113 30 31 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.025 $Y=1.637
+ $X2=0.71 $Y2=1.637
r114 29 31 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=0.62 $Y=1.637
+ $X2=0.71 $Y2=1.637
r115 29 45 17.9872 $w=2.53e-07 $l=3.98e-07 $layer=LI1_cond $X=0.62 $Y=1.637
+ $X2=0.222 $Y2=1.637
r116 28 49 15.927 $w=5.31e-07 $l=5.43171e-07 $layer=LI1_cond $X=0.62 $Y=0.825
+ $X2=0.402 $Y2=0.38
r117 28 29 42.2071 $w=1.78e-07 $l=6.85e-07 $layer=LI1_cond $X=0.62 $Y=0.825
+ $X2=0.62 $Y2=1.51
r118 24 45 0.504477 $w=2.65e-07 $l=1.28e-07 $layer=LI1_cond $X=0.222 $Y=1.765
+ $X2=0.222 $Y2=1.637
r119 24 26 2.39186 $w=2.63e-07 $l=5.5e-08 $layer=LI1_cond $X=0.222 $Y=1.765
+ $X2=0.222 $Y2=1.82
r120 20 56 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=3.12 $Y=1.32
+ $X2=3.12 $Y2=1.157
r121 20 22 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.12 $Y=1.32
+ $X2=3.12 $Y2=1.985
r122 17 56 3.55103 $w=3.25e-07 $l=2e-08 $layer=POLY_cond $X=3.1 $Y=1.157
+ $X2=3.12 $Y2=1.157
r123 17 43 1.77551 $w=3.25e-07 $l=1e-08 $layer=POLY_cond $X=3.1 $Y=1.157
+ $X2=3.09 $Y2=1.157
r124 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.1 $Y=0.995
+ $X2=3.1 $Y2=0.56
r125 13 53 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=2.69 $Y=1.32
+ $X2=2.69 $Y2=1.157
r126 13 15 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.69 $Y=1.32
+ $X2=2.69 $Y2=1.985
r127 10 53 3.55103 $w=3.25e-07 $l=2e-08 $layer=POLY_cond $X=2.67 $Y=1.157
+ $X2=2.69 $Y2=1.157
r128 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=0.56
r129 3 34 150 $w=1.7e-07 $l=7.24741e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=1.485 $X2=1.53 $Y2=1.89
r130 2 26 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.82
r131 1 49 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%VPWR 1 2 3 12 16 18 20 22 24 29 37 43 46 50
r54 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 41 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 41 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 38 46 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.63 $Y=2.72
+ $X2=2.415 $Y2=2.72
r61 38 40 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.63 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 37 49 4.60552 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=3.425 $Y2=2.72
r63 37 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 36 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 32 35 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r69 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 29 46 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.415 $Y2=2.72
r73 29 35 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.2 $Y=2.72 $X2=2.07
+ $Y2=2.72
r74 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 24 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 22 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 18 49 3.16065 $w=3.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.335 $Y=2.635
+ $X2=3.425 $Y2=2.72
r79 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.335 $Y=2.635
+ $X2=3.335 $Y2=2.34
r80 14 46 1.67165 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.72
r81 14 16 16.4826 $w=4.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.02
r82 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=2.72
r83 10 12 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=2.02
r84 3 20 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.485 $X2=3.335 $Y2=2.34
r85 2 16 300 $w=1.7e-07 $l=6.22796e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.415 $Y2=2.02
r86 1 12 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%X 1 2 9 13 15 16 17 18 20 23 25
r45 23 25 3.69697 $w=1.93e-07 $l=6.5e-08 $layer=LI1_cond $X=3.442 $Y=0.785
+ $X2=3.442 $Y2=0.85
r46 20 23 3.20299 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.442 $Y=0.7
+ $X2=3.442 $Y2=0.785
r47 20 25 0.568765 $w=1.93e-07 $l=1e-08 $layer=LI1_cond $X=3.442 $Y=0.86
+ $X2=3.442 $Y2=0.85
r48 19 20 59.4359 $w=1.93e-07 $l=1.045e-06 $layer=LI1_cond $X=3.442 $Y=1.905
+ $X2=3.442 $Y2=0.86
r49 17 20 3.65518 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.345 $Y=0.7
+ $X2=3.442 $Y2=0.7
r50 17 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.345 $Y=0.7
+ $X2=3.05 $Y2=0.7
r51 15 19 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=3.345 $Y=1.99
+ $X2=3.442 $Y2=1.905
r52 15 16 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.345 $Y=1.99 $X2=3
+ $Y2=1.99
r53 11 16 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.905 $Y=2.075
+ $X2=3 $Y2=1.99
r54 11 13 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=2.905 $Y=2.075
+ $X2=2.905 $Y2=2.3
r55 7 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.885 $Y=0.615
+ $X2=3.05 $Y2=0.7
r56 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.885 $Y=0.615
+ $X2=2.885 $Y2=0.36
r57 2 13 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.485 $X2=2.905 $Y2=2.3
r58 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.745
+ $Y=0.235 $X2=2.885 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%A_182_47# 1 2 11
c18 11 0 1.45172e-19 $X=1.985 $Y=0.73
r19 8 11 54.8708 $w=1.88e-07 $l=9.4e-07 $layer=LI1_cond $X=1.045 $Y=0.73
+ $X2=1.985 $Y2=0.73
r20 2 11 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=1.985 $Y2=0.73
r21 1 8 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.045 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_2%VGND 1 2 3 12 16 18 20 23 24 25 27 39 44 48
r53 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r54 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r56 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r57 39 47 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.45
+ $Y2=0
r58 39 41 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=2.99
+ $Y2=0
r59 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r60 38 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r61 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r62 35 44 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.557
+ $Y2=0
r63 35 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=2.07
+ $Y2=0
r64 34 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r65 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r66 29 33 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r67 27 44 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.557
+ $Y2=0
r68 27 33 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.15
+ $Y2=0
r69 25 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r70 25 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 23 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.07
+ $Y2=0
r72 23 24 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.432
+ $Y2=0
r73 22 41 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.99
+ $Y2=0
r74 22 24 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.432
+ $Y2=0
r75 18 47 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.385 $Y=0.085
+ $X2=3.45 $Y2=0
r76 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.385 $Y=0.085
+ $X2=3.385 $Y2=0.36
r77 14 24 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.432 $Y=0.085
+ $X2=2.432 $Y2=0
r78 14 16 13.486 $w=2.33e-07 $l=2.75e-07 $layer=LI1_cond $X=2.432 $Y=0.085
+ $X2=2.432 $Y2=0.36
r79 10 44 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.557 $Y=0.085
+ $X2=1.557 $Y2=0
r80 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=1.557 $Y=0.085
+ $X2=1.557 $Y2=0.38
r81 3 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.385 $Y2=0.36
r82 2 16 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.435 $Y2=0.36
r83 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.56 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a211o_2.pex.spice
* Created: Thu Aug 27 13:59:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A211O_2%A_79_21# 1 2 3 10 12 15 19 21 23 27 29 30 31
+ 32 35 37 41 45 47 50
c105 27 0 1.22295e-19 $X=1.085 $Y=1.16
r106 49 50 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=0.89 $Y=1.16 $X2=0.9
+ $Y2=1.16
r107 43 45 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.42 $Y=1.66
+ $X2=3.42 $Y2=1.755
r108 39 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.42 $Y=0.695
+ $X2=3.42 $Y2=0.4
r109 38 47 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0.785
+ $X2=2.44 $Y2=0.785
r110 37 39 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.255 $Y=0.785
+ $X2=3.42 $Y2=0.695
r111 37 38 40.0505 $w=1.78e-07 $l=6.5e-07 $layer=LI1_cond $X=3.255 $Y=0.785
+ $X2=2.605 $Y2=0.785
r112 33 47 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.44 $Y=0.695
+ $X2=2.44 $Y2=0.785
r113 33 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.44 $Y=0.695
+ $X2=2.44 $Y2=0.36
r114 31 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.255 $Y=1.575
+ $X2=3.42 $Y2=1.66
r115 31 32 126.893 $w=1.68e-07 $l=1.945e-06 $layer=LI1_cond $X=3.255 $Y=1.575
+ $X2=1.31 $Y2=1.575
r116 29 47 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0.785
+ $X2=2.44 $Y2=0.785
r117 29 30 59.4596 $w=1.78e-07 $l=9.65e-07 $layer=LI1_cond $X=2.275 $Y=0.785
+ $X2=1.31 $Y2=0.785
r118 28 50 27.2691 $w=3.27e-07 $l=1.85e-07 $layer=POLY_cond $X=1.085 $Y=1.16
+ $X2=0.9 $Y2=1.16
r119 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.16 $X2=1.085 $Y2=1.16
r120 25 32 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=1.155 $Y=1.49
+ $X2=1.31 $Y2=1.575
r121 25 27 12.2679 $w=3.08e-07 $l=3.3e-07 $layer=LI1_cond $X=1.155 $Y=1.49
+ $X2=1.155 $Y2=1.16
r122 24 30 7.45983 $w=1.8e-07 $l=1.94872e-07 $layer=LI1_cond $X=1.155 $Y=0.875
+ $X2=1.31 $Y2=0.785
r123 24 27 10.595 $w=3.08e-07 $l=2.85e-07 $layer=LI1_cond $X=1.155 $Y=0.875
+ $X2=1.155 $Y2=1.16
r124 21 50 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=0.995
+ $X2=0.9 $Y2=1.16
r125 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.9 $Y=0.995
+ $X2=0.9 $Y2=0.56
r126 17 49 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r127 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r128 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r129 10 49 61.9083 $w=3.27e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r130 10 13 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.47 $Y2=1.325
r131 10 12 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.47 $Y=1 $X2=0.47
+ $Y2=0.56
r132 3 45 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.755
r133 2 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.4
r134 1 35 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.235 $X2=2.44 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%A2 1 3 6 8 13
c31 8 0 1.85193e-19 $X=1.605 $Y=1.19
r32 13 14 23.8829 $w=3.33e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.157
+ $X2=1.83 $Y2=1.157
r33 11 13 2.89489 $w=3.33e-07 $l=2e-08 $layer=POLY_cond $X=1.645 $Y=1.157
+ $X2=1.665 $Y2=1.157
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.16 $X2=1.645 $Y2=1.16
r35 4 14 21.4384 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.157
r36 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.325 $X2=1.83
+ $Y2=1.985
r37 1 13 21.4384 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=1.665 $Y=0.99
+ $X2=1.665 $Y2=1.157
r38 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.665 $Y=0.99
+ $X2=1.665 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%A1 3 6 8 11 12 13
c33 11 0 1.85193e-19 $X=2.285 $Y=1.16
r34 11 14 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.297 $Y=1.16
+ $X2=2.297 $Y2=1.325
r35 11 13 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.297 $Y=1.16
+ $X2=2.297 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.285
+ $Y=1.16 $X2=2.285 $Y2=1.16
r37 8 12 11.0234 $w=2.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.065 $Y=1.16
+ $X2=2.285 $Y2=1.16
r38 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.37 $Y=1.985
+ $X2=2.37 $Y2=1.325
r39 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.225 $Y=0.56
+ $X2=2.225 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%B1 3 6 8 11 13
c30 11 0 1.82012e-19 $X=2.79 $Y=1.16
r31 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.16
+ $X2=2.79 $Y2=1.325
r32 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.16
+ $X2=2.79 $Y2=0.995
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.16 $X2=2.79 $Y2=1.16
r34 8 12 9.77071 $w=2.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.985 $Y=1.16
+ $X2=2.79 $Y2=1.16
r35 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.85 $Y=1.985
+ $X2=2.85 $Y2=1.325
r36 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.73 $Y=0.56 $X2=2.73
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%C1 1 3 6 8 13
c24 8 0 1.82012e-19 $X=3.45 $Y=1.19
r25 10 13 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.21 $Y=1.16
+ $X2=3.43 $Y2=1.16
r26 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.16 $X2=3.43 $Y2=1.16
r27 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.325 $X2=3.21
+ $Y2=1.985
r29 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.995 $X2=3.21
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%VPWR 1 2 3 10 12 18 22 24 26 31 41 42 48 51
r52 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 39 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 36 51 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2.23 $Y=2.72
+ $X2=2.092 $Y2=2.72
r60 36 38 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r61 35 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 32 48 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=1.127 $Y2=2.72
r65 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.255 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 31 51 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.092 $Y2=2.72
r67 31 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 30 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 27 45 4.46799 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r71 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 26 48 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=1.127
+ $Y2=2.72
r73 26 29 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=0.69
+ $Y2=2.72
r74 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 24 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 20 51 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.092 $Y=2.635
+ $X2=2.092 $Y2=2.72
r77 20 22 11.734 $w=2.73e-07 $l=2.8e-07 $layer=LI1_cond $X=2.092 $Y=2.635
+ $X2=2.092 $Y2=2.355
r78 16 48 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.127 $Y=2.635
+ $X2=1.127 $Y2=2.72
r79 16 18 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=1.127 $Y=2.635
+ $X2=1.127 $Y2=2
r80 12 15 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.237 $Y=1.655
+ $X2=0.237 $Y2=2.335
r81 10 45 3.00953 $w=2.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.192 $Y2=2.72
r82 10 15 11.7198 $w=2.93e-07 $l=3e-07 $layer=LI1_cond $X=0.237 $Y=2.635
+ $X2=0.237 $Y2=2.335
r83 3 22 600 $w=1.7e-07 $l=9.64832e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.105 $Y2=2.355
r84 2 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r85 1 15 400 $w=1.7e-07 $l=9.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.335
r86 1 12 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.655
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%X 1 2 9 11 13 16
r16 16 18 43.3419 $w=2.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.67 $Y=0.76
+ $X2=0.67 $Y2=1.625
r17 13 18 29.3121 $w=2.28e-07 $l=5.85e-07 $layer=LI1_cond $X=0.67 $Y=2.21
+ $X2=0.67 $Y2=1.625
r18 11 16 0.501062 $w=2.28e-07 $l=1e-08 $layer=LI1_cond $X=0.67 $Y=0.75 $X2=0.67
+ $Y2=0.76
r19 11 12 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.67 $Y=0.75
+ $X2=0.67 $Y2=0.635
r20 9 12 11.2625 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=0.665 $Y=0.42
+ $X2=0.665 $Y2=0.635
r21 2 18 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.625
r22 1 16 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.685 $Y2=0.76
r23 1 9 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%A_299_297# 1 2 9 14 16
r25 10 14 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=1.93
+ $X2=1.62 $Y2=1.93
r26 9 16 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=1.93
+ $X2=2.63 $Y2=1.93
r27 9 10 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.465 $Y=1.93
+ $X2=1.785 $Y2=1.93
r28 2 16 300 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=2 $X=2.445
+ $Y=1.485 $X2=2.63 $Y2=2
r29 1 14 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.485 $X2=1.62 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_2%VGND 1 2 3 10 12 16 18 25 32 33 41 47 49
c52 2 0 1.22295e-19 $X=0.975 $Y=0.235
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r54 45 47 10.1557 $w=5.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.61 $Y=0.18
+ $X2=1.795 $Y2=0.18
r55 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r56 43 45 3.49797 $w=5.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.455 $Y=0.18
+ $X2=1.61 $Y2=0.18
r57 40 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r58 39 43 6.88309 $w=5.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=1.455 $Y2=0.18
r59 39 41 10.6071 $w=5.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=0.945 $Y2=0.18
r60 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 33 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r63 30 49 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=2.947
+ $Y2=0
r64 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.45
+ $Y2=0
r65 29 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r66 29 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r67 28 47 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=1.795
+ $Y2=0
r68 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r69 25 49 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.947
+ $Y2=0
r70 25 28 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.53
+ $Y2=0
r71 24 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r72 23 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=0.945
+ $Y2=0
r73 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r74 21 36 4.46799 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r75 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.69
+ $Y2=0
r76 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r77 18 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r78 14 49 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.947 $Y=0.085
+ $X2=2.947 $Y2=0
r79 14 16 11.5244 $w=2.73e-07 $l=2.75e-07 $layer=LI1_cond $X=2.947 $Y=0.085
+ $X2=2.947 $Y2=0.36
r80 10 36 3.00953 $w=2.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.192 $Y2=0
r81 10 12 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.237 $Y2=0.38
r82 3 16 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.235 $X2=2.97 $Y2=0.36
r83 2 43 91 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=2 $X=0.975
+ $Y=0.235 $X2=1.455 $Y2=0.36
r84 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


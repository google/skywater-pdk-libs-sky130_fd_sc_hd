* File: sky130_fd_sc_hd__or4bb_2.pxi.spice
* Created: Thu Aug 27 14:44:49 2020
* 
x_PM_SKY130_FD_SC_HD__OR4BB_2%C_N N_C_N_M1013_g N_C_N_M1003_g C_N C_N
+ N_C_N_c_96_n N_C_N_c_97_n N_C_N_c_98_n PM_SKY130_FD_SC_HD__OR4BB_2%C_N
x_PM_SKY130_FD_SC_HD__OR4BB_2%D_N N_D_N_M1005_g N_D_N_M1015_g D_N N_D_N_c_129_n
+ N_D_N_c_130_n PM_SKY130_FD_SC_HD__OR4BB_2%D_N
x_PM_SKY130_FD_SC_HD__OR4BB_2%A_206_93# N_A_206_93#_M1005_d N_A_206_93#_M1015_d
+ N_A_206_93#_M1000_g N_A_206_93#_M1014_g N_A_206_93#_c_172_n
+ N_A_206_93#_c_166_n N_A_206_93#_c_167_n N_A_206_93#_c_168_n
+ N_A_206_93#_c_169_n N_A_206_93#_c_170_n PM_SKY130_FD_SC_HD__OR4BB_2%A_206_93#
x_PM_SKY130_FD_SC_HD__OR4BB_2%A_27_410# N_A_27_410#_M1003_s N_A_27_410#_M1013_s
+ N_A_27_410#_M1012_g N_A_27_410#_M1010_g N_A_27_410#_c_237_n
+ N_A_27_410#_c_243_n N_A_27_410#_c_244_n N_A_27_410#_c_245_n
+ N_A_27_410#_c_246_n N_A_27_410#_c_247_n N_A_27_410#_c_238_n
+ N_A_27_410#_c_239_n N_A_27_410#_c_240_n N_A_27_410#_c_250_n
+ PM_SKY130_FD_SC_HD__OR4BB_2%A_27_410#
x_PM_SKY130_FD_SC_HD__OR4BB_2%B N_B_M1011_g N_B_M1002_g N_B_c_325_n N_B_c_326_n
+ B N_B_c_329_n PM_SKY130_FD_SC_HD__OR4BB_2%B
x_PM_SKY130_FD_SC_HD__OR4BB_2%A N_A_M1001_g N_A_M1004_g A N_A_c_368_n
+ N_A_c_369_n PM_SKY130_FD_SC_HD__OR4BB_2%A
x_PM_SKY130_FD_SC_HD__OR4BB_2%A_316_413# N_A_316_413#_M1000_d
+ N_A_316_413#_M1002_d N_A_316_413#_M1014_s N_A_316_413#_c_409_n
+ N_A_316_413#_M1006_g N_A_316_413#_M1007_g N_A_316_413#_c_410_n
+ N_A_316_413#_M1008_g N_A_316_413#_M1009_g N_A_316_413#_c_420_n
+ N_A_316_413#_c_514_p N_A_316_413#_c_421_n N_A_316_413#_c_411_n
+ N_A_316_413#_c_412_n N_A_316_413#_c_422_n N_A_316_413#_c_430_n
+ N_A_316_413#_c_524_p N_A_316_413#_c_413_n N_A_316_413#_c_465_n
+ N_A_316_413#_c_423_n N_A_316_413#_c_414_n N_A_316_413#_c_424_n
+ N_A_316_413#_c_415_n N_A_316_413#_c_416_n N_A_316_413#_c_417_n
+ PM_SKY130_FD_SC_HD__OR4BB_2%A_316_413#
x_PM_SKY130_FD_SC_HD__OR4BB_2%VPWR N_VPWR_M1013_d N_VPWR_M1004_d N_VPWR_M1009_d
+ N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n VPWR
+ N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n
+ N_VPWR_c_537_n PM_SKY130_FD_SC_HD__OR4BB_2%VPWR
x_PM_SKY130_FD_SC_HD__OR4BB_2%X N_X_M1006_d N_X_M1007_s N_X_c_605_n N_X_c_607_n
+ N_X_c_603_n X PM_SKY130_FD_SC_HD__OR4BB_2%X
x_PM_SKY130_FD_SC_HD__OR4BB_2%VGND N_VGND_M1003_d N_VGND_M1000_s N_VGND_M1012_d
+ N_VGND_M1001_d N_VGND_M1008_s N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n
+ N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n VGND N_VGND_c_634_n
+ N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n
+ N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n VGND
+ PM_SKY130_FD_SC_HD__OR4BB_2%VGND
cc_1 VNB N_C_N_c_96_n 0.023255f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_2 VNB N_C_N_c_97_n 0.00602296f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_3 VNB N_C_N_c_98_n 0.0208027f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_4 VNB D_N 0.0023514f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_5 VNB N_D_N_c_129_n 0.0268087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_D_N_c_130_n 0.0189069f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_7 VNB N_A_206_93#_M1000_g 0.0325332f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_8 VNB N_A_206_93#_c_166_n 0.00451126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_206_93#_c_167_n 7.21544e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_206_93#_c_168_n 0.012688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_206_93#_c_169_n 0.00175f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_206_93#_c_170_n 0.0346299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_410#_M1012_g 0.0270012f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_14 VNB N_A_27_410#_c_237_n 0.0224435f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.325
cc_15 VNB N_A_27_410#_c_238_n 2.24825e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_410#_c_239_n 0.0221854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_410#_c_240_n 0.0187765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_M1011_g 0.0157284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B_c_325_n 0.0147133f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_20 VNB N_B_c_326_n 0.00821622f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_21 VNB N_A_M1001_g 0.0277171f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.26
cc_22 VNB N_A_c_368_n 0.0200358f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_23 VNB N_A_c_369_n 0.00432763f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_24 VNB N_A_316_413#_c_409_n 0.0160502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_316_413#_c_410_n 0.0187042f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.16
cc_26 VNB N_A_316_413#_c_411_n 0.0116364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_316_413#_c_412_n 0.00452568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_316_413#_c_413_n 0.00233469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_316_413#_c_414_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_316_413#_c_415_n 0.00185649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_316_413#_c_416_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_316_413#_c_417_n 0.0455382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_537_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_603_n 7.68963e-19 $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_35 VNB N_VGND_c_628_n 0.0126821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_629_n 0.00646225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_630_n 3.08095e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_631_n 3.22528e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_632_n 0.0112126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_633_n 0.0129123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_634_n 0.0189629f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_635_n 0.01289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_636_n 0.0111699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_637_n 0.0171221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_638_n 0.0243657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_639_n 0.0055533f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_640_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_641_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_642_n 0.259422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_C_N_M1013_g 0.0562707f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.26
cc_51 VPB N_C_N_c_96_n 0.00470919f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_52 VPB N_C_N_c_97_n 0.00234555f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_53 VPB N_D_N_M1015_g 0.0229539f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_54 VPB D_N 5.16049e-19 $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_55 VPB N_D_N_c_129_n 0.00583034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_206_93#_M1014_g 0.0635781f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_57 VPB N_A_206_93#_c_172_n 0.00893839f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_58 VPB N_A_206_93#_c_167_n 0.00403233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_206_93#_c_170_n 0.010455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_410#_M1010_g 0.0190829f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_61 VPB N_A_27_410#_c_237_n 0.0263492f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.325
cc_62 VPB N_A_27_410#_c_243_n 0.016454f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.19
cc_63 VPB N_A_27_410#_c_244_n 0.0206891f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.53
cc_64 VPB N_A_27_410#_c_245_n 0.00680513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_410#_c_246_n 0.00561423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_410#_c_247_n 0.00201079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_410#_c_238_n 9.16196e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_410#_c_239_n 0.00435359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_410#_c_250_n 0.0111036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B_M1011_g 0.0267766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB B 0.0122602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_B_c_329_n 0.0353878f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_73 VPB N_A_M1004_g 0.0209374f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.675
cc_74 VPB N_A_c_368_n 0.00399502f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_75 VPB N_A_c_369_n 0.0033301f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_76 VPB N_A_316_413#_M1007_g 0.0209283f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_77 VPB N_A_316_413#_M1009_g 0.0241426f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_316_413#_c_420_n 0.00969822f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_316_413#_c_421_n 0.00241773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_316_413#_c_422_n 0.003558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_316_413#_c_423_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_316_413#_c_424_n 0.00130727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_316_413#_c_417_n 0.00736414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_538_n 0.0141254f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_85 VPB N_VPWR_c_539_n 0.0103523f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.325
cc_86 VPB N_VPWR_c_540_n 0.0111834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_541_n 0.00851481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_542_n 0.0145108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_543_n 0.0640044f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_544_n 0.018077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_545_n 0.00519112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_546_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_537_n 0.0691573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_X_c_603_n 0.00111849f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_95 N_C_N_M1013_g N_D_N_M1015_g 0.0243255f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_96 N_C_N_c_97_n N_D_N_M1015_g 0.00414707f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_97 N_C_N_c_96_n D_N 2.85663e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_98 N_C_N_c_97_n D_N 0.0259635f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_99 N_C_N_c_96_n N_D_N_c_129_n 0.019221f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_100 N_C_N_c_97_n N_D_N_c_129_n 0.00225922f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_101 N_C_N_c_98_n N_D_N_c_130_n 0.0104665f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_102 N_C_N_c_97_n N_A_206_93#_c_172_n 0.011488f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_103 N_C_N_c_97_n N_A_206_93#_c_167_n 0.00632897f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_104 N_C_N_M1013_g N_A_27_410#_c_237_n 0.0134005f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_105 N_C_N_c_96_n N_A_27_410#_c_237_n 0.00753785f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_106 N_C_N_c_97_n N_A_27_410#_c_237_n 0.0529229f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_107 N_C_N_c_98_n N_A_27_410#_c_237_n 0.00528758f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_108 N_C_N_M1013_g N_A_27_410#_c_243_n 0.00143901f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_109 N_C_N_M1013_g N_A_27_410#_c_244_n 0.0144867f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_110 N_C_N_c_96_n N_A_27_410#_c_244_n 7.20998e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_111 N_C_N_c_97_n N_A_27_410#_c_244_n 0.0280218f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C_N_c_98_n N_A_27_410#_c_240_n 3.39406e-19 $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_113 N_C_N_c_97_n N_VPWR_M1013_d 0.00442525f $X=0.515 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_114 N_C_N_M1013_g N_VPWR_c_538_n 0.0100087f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_115 N_C_N_M1013_g N_VPWR_c_542_n 0.00334979f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_116 N_C_N_M1013_g N_VPWR_c_537_n 0.0048928f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_117 N_C_N_c_97_n N_VGND_c_628_n 0.0108718f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C_N_c_98_n N_VGND_c_628_n 0.00422719f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_119 N_C_N_c_98_n N_VGND_c_638_n 0.00510437f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_120 N_C_N_c_98_n N_VGND_c_642_n 0.00512902f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_121 N_D_N_M1015_g N_A_206_93#_c_172_n 0.00298359f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_122 D_N N_A_206_93#_c_172_n 0.0141771f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_123 N_D_N_c_129_n N_A_206_93#_c_172_n 0.00360045f $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_124 D_N N_A_206_93#_c_166_n 0.00627858f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_125 N_D_N_c_129_n N_A_206_93#_c_166_n 2.39293e-19 $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_126 N_D_N_c_130_n N_A_206_93#_c_166_n 0.00428594f $X=1.035 $Y=0.995 $X2=0
+ $Y2=0
cc_127 N_D_N_M1015_g N_A_206_93#_c_167_n 0.00310772f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_128 D_N N_A_206_93#_c_167_n 0.00627858f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_129 N_D_N_c_129_n N_A_206_93#_c_167_n 2.39293e-19 $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_130 D_N N_A_206_93#_c_168_n 0.012483f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_131 N_D_N_c_129_n N_A_206_93#_c_168_n 0.00272654f $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_D_N_c_130_n N_A_206_93#_c_168_n 3.44947e-19 $X=1.035 $Y=0.995 $X2=0
+ $Y2=0
cc_133 D_N N_A_206_93#_c_169_n 0.0143051f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_134 N_D_N_c_129_n N_A_206_93#_c_169_n 5.83479e-19 $X=1.035 $Y=1.16 $X2=0
+ $Y2=0
cc_135 D_N N_A_206_93#_c_170_n 8.65104e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_136 N_D_N_c_129_n N_A_206_93#_c_170_n 0.0118962f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_137 N_D_N_M1015_g N_A_27_410#_c_244_n 0.0156302f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_138 D_N N_A_27_410#_c_244_n 0.00124584f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_139 N_D_N_M1015_g N_VPWR_c_543_n 0.00259183f $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_140 N_D_N_M1015_g N_VPWR_c_537_n 0.00417489f $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_141 N_D_N_c_130_n N_VGND_c_628_n 0.00165256f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_142 N_D_N_c_130_n N_VGND_c_629_n 0.00207743f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_143 N_D_N_c_130_n N_VGND_c_634_n 0.00510437f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_144 N_D_N_c_130_n N_VGND_c_642_n 0.00512902f $X=1.035 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_206_93#_M1000_g N_A_27_410#_M1012_g 0.0209129f $X=1.895 $Y=0.445
+ $X2=0 $Y2=0
cc_146 N_A_206_93#_M1014_g N_A_27_410#_M1010_g 0.0243913f $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_147 N_A_206_93#_M1015_d N_A_27_410#_c_244_n 0.00247126f $X=1.03 $Y=1.485
+ $X2=0 $Y2=0
cc_148 N_A_206_93#_M1014_g N_A_27_410#_c_244_n 0.00812129f $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_149 N_A_206_93#_c_172_n N_A_27_410#_c_244_n 0.041501f $X=1.41 $Y=1.61 $X2=0
+ $Y2=0
cc_150 N_A_206_93#_c_169_n N_A_27_410#_c_244_n 0.0045774f $X=1.67 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_206_93#_c_170_n N_A_27_410#_c_244_n 0.00315934f $X=1.915 $Y=1.16
+ $X2=0 $Y2=0
cc_152 N_A_206_93#_M1014_g N_A_27_410#_c_245_n 0.010188f $X=1.915 $Y=2.275 $X2=0
+ $Y2=0
cc_153 N_A_206_93#_c_172_n N_A_27_410#_c_245_n 0.00916297f $X=1.41 $Y=1.61 $X2=0
+ $Y2=0
cc_154 N_A_206_93#_M1014_g N_A_27_410#_c_246_n 0.0064787f $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_155 N_A_206_93#_M1014_g N_A_27_410#_c_247_n 0.00882292f $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_156 N_A_206_93#_c_172_n N_A_27_410#_c_247_n 0.00555401f $X=1.41 $Y=1.61 $X2=0
+ $Y2=0
cc_157 N_A_206_93#_c_167_n N_A_27_410#_c_247_n 0.00928736f $X=1.505 $Y=1.525
+ $X2=0 $Y2=0
cc_158 N_A_206_93#_c_169_n N_A_27_410#_c_247_n 0.00673601f $X=1.67 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_206_93#_c_170_n N_A_27_410#_c_247_n 0.00187495f $X=1.915 $Y=1.16
+ $X2=0 $Y2=0
cc_160 N_A_206_93#_M1014_g N_A_27_410#_c_238_n 8.16443e-19 $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_161 N_A_206_93#_c_166_n N_A_27_410#_c_238_n 0.00178546f $X=1.505 $Y=1.075
+ $X2=0 $Y2=0
cc_162 N_A_206_93#_c_167_n N_A_27_410#_c_238_n 0.00442275f $X=1.505 $Y=1.525
+ $X2=0 $Y2=0
cc_163 N_A_206_93#_c_169_n N_A_27_410#_c_238_n 0.0062484f $X=1.67 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A_206_93#_c_170_n N_A_27_410#_c_238_n 0.00131394f $X=1.915 $Y=1.16
+ $X2=0 $Y2=0
cc_165 N_A_206_93#_c_169_n N_A_27_410#_c_239_n 4.74955e-19 $X=1.67 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_206_93#_c_170_n N_A_27_410#_c_239_n 0.0213915f $X=1.915 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_206_93#_M1014_g N_B_M1011_g 0.00153736f $X=1.915 $Y=2.275 $X2=0 $Y2=0
cc_168 N_A_206_93#_M1014_g B 0.00223393f $X=1.915 $Y=2.275 $X2=0 $Y2=0
cc_169 N_A_206_93#_M1014_g N_B_c_329_n 0.00325164f $X=1.915 $Y=2.275 $X2=0 $Y2=0
cc_170 N_A_206_93#_M1014_g N_A_316_413#_c_420_n 0.00971256f $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_171 N_A_206_93#_M1014_g N_A_316_413#_c_421_n 0.00494253f $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_172 N_A_206_93#_M1000_g N_A_316_413#_c_412_n 0.00222847f $X=1.895 $Y=0.445
+ $X2=0 $Y2=0
cc_173 N_A_206_93#_c_168_n N_A_316_413#_c_412_n 0.00818093f $X=1.165 $Y=0.66
+ $X2=0 $Y2=0
cc_174 N_A_206_93#_M1014_g N_A_316_413#_c_430_n 0.00129708f $X=1.915 $Y=2.275
+ $X2=0 $Y2=0
cc_175 N_A_206_93#_M1014_g N_VPWR_c_543_n 0.00375986f $X=1.915 $Y=2.275 $X2=0
+ $Y2=0
cc_176 N_A_206_93#_M1014_g N_VPWR_c_537_n 0.00798404f $X=1.915 $Y=2.275 $X2=0
+ $Y2=0
cc_177 N_A_206_93#_c_168_n N_VGND_M1000_s 4.10598e-19 $X=1.165 $Y=0.66 $X2=0
+ $Y2=0
cc_178 N_A_206_93#_c_168_n N_VGND_c_628_n 8.07382e-19 $X=1.165 $Y=0.66 $X2=0
+ $Y2=0
cc_179 N_A_206_93#_M1000_g N_VGND_c_629_n 0.00890499f $X=1.895 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_206_93#_c_168_n N_VGND_c_629_n 0.0108733f $X=1.165 $Y=0.66 $X2=0
+ $Y2=0
cc_181 N_A_206_93#_c_169_n N_VGND_c_629_n 0.00625028f $X=1.67 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_A_206_93#_c_170_n N_VGND_c_629_n 0.00414886f $X=1.915 $Y=1.16 $X2=0
+ $Y2=0
cc_183 N_A_206_93#_M1000_g N_VGND_c_630_n 6.24366e-19 $X=1.895 $Y=0.445 $X2=0
+ $Y2=0
cc_184 N_A_206_93#_c_168_n N_VGND_c_634_n 0.0095527f $X=1.165 $Y=0.66 $X2=0
+ $Y2=0
cc_185 N_A_206_93#_M1000_g N_VGND_c_635_n 0.0046653f $X=1.895 $Y=0.445 $X2=0
+ $Y2=0
cc_186 N_A_206_93#_M1000_g N_VGND_c_642_n 0.00808301f $X=1.895 $Y=0.445 $X2=0
+ $Y2=0
cc_187 N_A_206_93#_c_168_n N_VGND_c_642_n 0.0131649f $X=1.165 $Y=0.66 $X2=0
+ $Y2=0
cc_188 N_A_27_410#_c_246_n N_B_M1011_g 7.72856e-19 $X=2.25 $Y=1.5 $X2=0 $Y2=0
cc_189 N_A_27_410#_c_238_n N_B_M1011_g 8.95596e-19 $X=2.335 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_27_410#_c_239_n N_B_M1011_g 0.0641534f $X=2.335 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_27_410#_M1012_g N_B_c_325_n 0.0136904f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A_27_410#_M1012_g N_B_c_326_n 0.0126742f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A_27_410#_c_238_n N_A_c_369_n 0.0217601f $X=2.335 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_27_410#_c_239_n N_A_c_369_n 0.00220685f $X=2.335 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_27_410#_c_244_n N_A_316_413#_c_420_n 0.0272384f $X=1.77 $Y=1.95 $X2=0
+ $Y2=0
cc_196 N_A_27_410#_c_246_n N_A_316_413#_c_420_n 0.00376842f $X=2.25 $Y=1.5 $X2=0
+ $Y2=0
cc_197 N_A_27_410#_M1010_g N_A_316_413#_c_421_n 0.00197943f $X=2.395 $Y=1.695
+ $X2=0 $Y2=0
cc_198 N_A_27_410#_c_244_n N_A_316_413#_c_421_n 0.00625142f $X=1.77 $Y=1.95
+ $X2=0 $Y2=0
cc_199 N_A_27_410#_M1012_g N_A_316_413#_c_411_n 0.0113758f $X=2.35 $Y=0.445
+ $X2=0 $Y2=0
cc_200 N_A_27_410#_c_246_n N_A_316_413#_c_411_n 0.00169186f $X=2.25 $Y=1.5 $X2=0
+ $Y2=0
cc_201 N_A_27_410#_c_238_n N_A_316_413#_c_411_n 0.012736f $X=2.335 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_27_410#_c_239_n N_A_316_413#_c_411_n 0.00340859f $X=2.335 $Y=1.16
+ $X2=0 $Y2=0
cc_203 N_A_27_410#_c_246_n N_A_316_413#_c_412_n 0.00590033f $X=2.25 $Y=1.5 $X2=0
+ $Y2=0
cc_204 N_A_27_410#_M1010_g N_A_316_413#_c_422_n 0.0121016f $X=2.395 $Y=1.695
+ $X2=0 $Y2=0
cc_205 N_A_27_410#_c_246_n N_A_316_413#_c_422_n 0.00656826f $X=2.25 $Y=1.5 $X2=0
+ $Y2=0
cc_206 N_A_27_410#_c_244_n N_A_316_413#_c_430_n 0.00786633f $X=1.77 $Y=1.95
+ $X2=0 $Y2=0
cc_207 N_A_27_410#_c_245_n N_A_316_413#_c_430_n 0.00628038f $X=1.855 $Y=1.865
+ $X2=0 $Y2=0
cc_208 N_A_27_410#_c_246_n N_A_316_413#_c_430_n 0.0109594f $X=2.25 $Y=1.5 $X2=0
+ $Y2=0
cc_209 N_A_27_410#_c_239_n N_A_316_413#_c_430_n 2.10144e-19 $X=2.335 $Y=1.16
+ $X2=0 $Y2=0
cc_210 N_A_27_410#_c_246_n N_A_316_413#_c_424_n 0.00276731f $X=2.25 $Y=1.5 $X2=0
+ $Y2=0
cc_211 N_A_27_410#_c_244_n N_VPWR_M1013_d 0.00524517f $X=1.77 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_212 N_A_27_410#_c_244_n N_VPWR_c_538_n 0.0229102f $X=1.77 $Y=1.95 $X2=0 $Y2=0
cc_213 N_A_27_410#_c_243_n N_VPWR_c_542_n 0.0168666f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_214 N_A_27_410#_c_244_n N_VPWR_c_542_n 0.00256078f $X=1.77 $Y=1.95 $X2=0
+ $Y2=0
cc_215 N_A_27_410#_M1010_g N_VPWR_c_543_n 0.00327927f $X=2.395 $Y=1.695 $X2=0
+ $Y2=0
cc_216 N_A_27_410#_c_244_n N_VPWR_c_543_n 0.0110846f $X=1.77 $Y=1.95 $X2=0 $Y2=0
cc_217 N_A_27_410#_M1010_g N_VPWR_c_537_n 0.00417489f $X=2.395 $Y=1.695 $X2=0
+ $Y2=0
cc_218 N_A_27_410#_c_243_n N_VPWR_c_537_n 0.00987673f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_219 N_A_27_410#_c_244_n N_VPWR_c_537_n 0.0244843f $X=1.77 $Y=1.95 $X2=0 $Y2=0
cc_220 N_A_27_410#_c_246_n A_398_413# 0.00263772f $X=2.25 $Y=1.5 $X2=-0.19
+ $Y2=-0.24
cc_221 N_A_27_410#_c_240_n N_VGND_c_628_n 0.0105001f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_222 N_A_27_410#_M1012_g N_VGND_c_629_n 6.19205e-19 $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_27_410#_M1012_g N_VGND_c_630_n 0.00742769f $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_27_410#_M1012_g N_VGND_c_635_n 0.00341689f $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_225 N_A_27_410#_c_240_n N_VGND_c_638_n 0.00972557f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_226 N_A_27_410#_M1012_g N_VGND_c_642_n 0.00414154f $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_227 N_A_27_410#_c_240_n N_VGND_c_642_n 0.0107261f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_228 N_B_M1011_g N_A_M1001_g 0.00392288f $X=2.755 $Y=1.695 $X2=0 $Y2=0
cc_229 N_B_c_325_n N_A_M1001_g 0.0207641f $X=2.762 $Y=0.76 $X2=0 $Y2=0
cc_230 N_B_M1011_g N_A_M1004_g 0.0299871f $X=2.755 $Y=1.695 $X2=0 $Y2=0
cc_231 B N_A_M1004_g 8.99686e-19 $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_232 N_B_M1011_g N_A_c_368_n 0.0213087f $X=2.755 $Y=1.695 $X2=0 $Y2=0
cc_233 N_B_M1011_g N_A_c_369_n 0.0141584f $X=2.755 $Y=1.695 $X2=0 $Y2=0
cc_234 N_B_c_326_n N_A_c_369_n 4.43208e-19 $X=2.762 $Y=0.91 $X2=0 $Y2=0
cc_235 B N_A_316_413#_c_420_n 0.0130053f $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_236 N_B_c_329_n N_A_316_413#_c_420_n 6.32819e-19 $X=2.815 $Y=2.335 $X2=0
+ $Y2=0
cc_237 N_B_M1011_g N_A_316_413#_c_421_n 0.00201096f $X=2.755 $Y=1.695 $X2=0
+ $Y2=0
cc_238 B N_A_316_413#_c_421_n 0.00542028f $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_239 N_B_c_325_n N_A_316_413#_c_411_n 0.00699162f $X=2.762 $Y=0.76 $X2=0 $Y2=0
cc_240 N_B_c_326_n N_A_316_413#_c_411_n 0.00481812f $X=2.762 $Y=0.91 $X2=0 $Y2=0
cc_241 N_B_M1011_g N_A_316_413#_c_422_n 0.0107156f $X=2.755 $Y=1.695 $X2=0 $Y2=0
cc_242 B N_A_316_413#_c_422_n 0.0349748f $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_243 N_B_c_329_n N_A_316_413#_c_422_n 0.00101546f $X=2.815 $Y=2.335 $X2=0
+ $Y2=0
cc_244 N_B_M1011_g N_A_316_413#_c_424_n 0.00538706f $X=2.755 $Y=1.695 $X2=0
+ $Y2=0
cc_245 B N_A_316_413#_c_424_n 0.0138251f $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_246 N_B_M1011_g N_VPWR_c_539_n 0.00280623f $X=2.755 $Y=1.695 $X2=0 $Y2=0
cc_247 B N_VPWR_c_539_n 0.0285382f $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_248 N_B_c_329_n N_VPWR_c_539_n 0.00108286f $X=2.815 $Y=2.335 $X2=0 $Y2=0
cc_249 B N_VPWR_c_543_n 0.0396304f $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_250 N_B_c_329_n N_VPWR_c_543_n 0.00774997f $X=2.815 $Y=2.335 $X2=0 $Y2=0
cc_251 B N_VPWR_c_537_n 0.0238619f $X=2.93 $Y=2.125 $X2=0 $Y2=0
cc_252 N_B_c_329_n N_VPWR_c_537_n 0.0109691f $X=2.815 $Y=2.335 $X2=0 $Y2=0
cc_253 N_B_c_325_n N_VGND_c_630_n 0.00716819f $X=2.762 $Y=0.76 $X2=0 $Y2=0
cc_254 N_B_c_325_n N_VGND_c_631_n 6.24658e-19 $X=2.762 $Y=0.76 $X2=0 $Y2=0
cc_255 N_B_c_325_n N_VGND_c_636_n 0.00341689f $X=2.762 $Y=0.76 $X2=0 $Y2=0
cc_256 N_B_c_325_n N_VGND_c_642_n 0.00405445f $X=2.762 $Y=0.76 $X2=0 $Y2=0
cc_257 N_A_M1001_g N_A_316_413#_c_409_n 0.0177679f $X=3.19 $Y=0.445 $X2=0 $Y2=0
cc_258 N_A_M1004_g N_A_316_413#_M1007_g 0.0189405f $X=3.19 $Y=1.695 $X2=0 $Y2=0
cc_259 N_A_c_369_n N_A_316_413#_c_411_n 0.0189424f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A_c_369_n N_A_316_413#_c_422_n 0.0101811f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_M1001_g N_A_316_413#_c_413_n 0.011795f $X=3.19 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_c_368_n N_A_316_413#_c_413_n 0.00220162f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_c_369_n N_A_316_413#_c_413_n 0.0166868f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_M1004_g N_A_316_413#_c_465_n 0.0112137f $X=3.19 $Y=1.695 $X2=0 $Y2=0
cc_265 N_A_c_369_n N_A_316_413#_c_465_n 0.00969518f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_M1004_g N_A_316_413#_c_423_n 0.0034529f $X=3.19 $Y=1.695 $X2=0 $Y2=0
cc_267 N_A_c_368_n N_A_316_413#_c_414_n 5.77159e-19 $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_c_369_n N_A_316_413#_c_414_n 0.0146254f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_M1004_g N_A_316_413#_c_424_n 0.00964298f $X=3.19 $Y=1.695 $X2=0 $Y2=0
cc_270 N_A_c_368_n N_A_316_413#_c_424_n 0.00156816f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_c_369_n N_A_316_413#_c_424_n 0.0112207f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_c_368_n N_A_316_413#_c_415_n 0.00186332f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_c_369_n N_A_316_413#_c_415_n 0.027072f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_M1001_g N_A_316_413#_c_416_n 0.0034529f $X=3.19 $Y=0.445 $X2=0 $Y2=0
cc_275 N_A_c_368_n N_A_316_413#_c_417_n 0.0203649f $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_c_369_n N_A_316_413#_c_417_n 3.52022e-19 $X=3.175 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_M1004_g N_VPWR_c_539_n 0.00293484f $X=3.19 $Y=1.695 $X2=0 $Y2=0
cc_278 N_A_M1004_g N_VPWR_c_543_n 0.00264181f $X=3.19 $Y=1.695 $X2=0 $Y2=0
cc_279 N_A_M1004_g N_VPWR_c_537_n 0.00333991f $X=3.19 $Y=1.695 $X2=0 $Y2=0
cc_280 N_A_M1001_g N_VGND_c_630_n 6.21849e-19 $X=3.19 $Y=0.445 $X2=0 $Y2=0
cc_281 N_A_M1001_g N_VGND_c_631_n 0.00746702f $X=3.19 $Y=0.445 $X2=0 $Y2=0
cc_282 N_A_M1001_g N_VGND_c_636_n 0.00341689f $X=3.19 $Y=0.445 $X2=0 $Y2=0
cc_283 N_A_M1001_g N_VGND_c_642_n 0.00405445f $X=3.19 $Y=0.445 $X2=0 $Y2=0
cc_284 N_A_316_413#_c_465_n N_VPWR_M1004_d 0.00526233f $X=3.465 $Y=1.58 $X2=0
+ $Y2=0
cc_285 N_A_316_413#_M1007_g N_VPWR_c_539_n 0.00348231f $X=3.68 $Y=1.985 $X2=0
+ $Y2=0
cc_286 N_A_316_413#_c_465_n N_VPWR_c_539_n 0.0190361f $X=3.465 $Y=1.58 $X2=0
+ $Y2=0
cc_287 N_A_316_413#_c_424_n N_VPWR_c_539_n 0.00605542f $X=3.06 $Y=1.58 $X2=0
+ $Y2=0
cc_288 N_A_316_413#_c_417_n N_VPWR_c_539_n 2.11345e-19 $X=4.1 $Y=1.16 $X2=0
+ $Y2=0
cc_289 N_A_316_413#_M1009_g N_VPWR_c_541_n 0.00671263f $X=4.1 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_A_316_413#_c_420_n N_VPWR_c_543_n 0.0285048f $X=2.11 $Y=2.29 $X2=0
+ $Y2=0
cc_291 N_A_316_413#_M1007_g N_VPWR_c_544_n 0.00585385f $X=3.68 $Y=1.985 $X2=0
+ $Y2=0
cc_292 N_A_316_413#_M1009_g N_VPWR_c_544_n 0.00503406f $X=4.1 $Y=1.985 $X2=0
+ $Y2=0
cc_293 N_A_316_413#_M1014_s N_VPWR_c_537_n 0.00217968f $X=1.58 $Y=2.065 $X2=0
+ $Y2=0
cc_294 N_A_316_413#_M1007_g N_VPWR_c_537_n 0.0118387f $X=3.68 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_A_316_413#_M1009_g N_VPWR_c_537_n 0.00966033f $X=4.1 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_316_413#_c_420_n N_VPWR_c_537_n 0.0256417f $X=2.11 $Y=2.29 $X2=0
+ $Y2=0
cc_297 N_A_316_413#_c_422_n N_VPWR_c_537_n 0.00841166f $X=2.975 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_316_413#_c_420_n A_398_413# 0.0042428f $X=2.11 $Y=2.29 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_316_413#_c_421_n A_398_413# 0.00292122f $X=2.195 $Y=2.205 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_316_413#_c_430_n A_398_413# 0.00335245f $X=2.28 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_301 N_A_316_413#_c_422_n A_494_297# 0.00366293f $X=2.975 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_302 N_A_316_413#_c_422_n A_566_297# 0.00180544f $X=2.975 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_303 N_A_316_413#_c_424_n A_566_297# 0.00465932f $X=3.06 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_304 N_A_316_413#_c_410_n N_X_c_605_n 0.00536146f $X=4.1 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_316_413#_c_417_n N_X_c_605_n 0.00259703f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_316_413#_M1009_g N_X_c_607_n 0.00294462f $X=4.1 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A_316_413#_c_417_n N_X_c_607_n 0.00288868f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A_316_413#_c_409_n N_X_c_603_n 0.00151661f $X=3.68 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_316_413#_M1007_g N_X_c_603_n 0.00115345f $X=3.68 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_316_413#_c_410_n N_X_c_603_n 0.00462154f $X=4.1 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A_316_413#_M1009_g N_X_c_603_n 0.006621f $X=4.1 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A_316_413#_c_413_n N_X_c_603_n 0.00352178f $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A_316_413#_c_423_n N_X_c_603_n 0.00841218f $X=3.55 $Y=1.495 $X2=0 $Y2=0
cc_314 N_A_316_413#_c_415_n N_X_c_603_n 0.0232251f $X=3.655 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_316_413#_c_416_n N_X_c_603_n 0.00836616f $X=3.602 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_316_413#_c_417_n N_X_c_603_n 0.0221596f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_316_413#_M1009_g X 0.0119134f $X=4.1 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A_316_413#_c_413_n N_VGND_M1001_d 0.00464421f $X=3.465 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_316_413#_c_416_n N_VGND_M1001_d 6.98847e-19 $X=3.602 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_A_316_413#_c_514_p N_VGND_c_630_n 0.0117247f $X=2.11 $Y=0.47 $X2=0
+ $Y2=0
cc_321 N_A_316_413#_c_411_n N_VGND_c_630_n 0.020154f $X=2.895 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_316_413#_c_409_n N_VGND_c_631_n 0.00768198f $X=3.68 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_316_413#_c_410_n N_VGND_c_631_n 9.49203e-19 $X=4.1 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_316_413#_c_413_n N_VGND_c_631_n 0.022675f $X=3.465 $Y=0.74 $X2=0
+ $Y2=0
cc_325 N_A_316_413#_c_417_n N_VGND_c_631_n 2.33671e-19 $X=4.1 $Y=1.16 $X2=0
+ $Y2=0
cc_326 N_A_316_413#_c_410_n N_VGND_c_633_n 0.00888029f $X=4.1 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_316_413#_c_514_p N_VGND_c_635_n 0.00873683f $X=2.11 $Y=0.47 $X2=0
+ $Y2=0
cc_328 N_A_316_413#_c_411_n N_VGND_c_635_n 0.00325972f $X=2.895 $Y=0.74 $X2=0
+ $Y2=0
cc_329 N_A_316_413#_c_411_n N_VGND_c_636_n 0.00273399f $X=2.895 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_316_413#_c_524_p N_VGND_c_636_n 0.00846569f $X=2.98 $Y=0.47 $X2=0
+ $Y2=0
cc_331 N_A_316_413#_c_413_n N_VGND_c_636_n 0.00273399f $X=3.465 $Y=0.74 $X2=0
+ $Y2=0
cc_332 N_A_316_413#_c_409_n N_VGND_c_637_n 0.00524631f $X=3.68 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A_316_413#_c_410_n N_VGND_c_637_n 0.00513402f $X=4.1 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_316_413#_c_413_n N_VGND_c_637_n 3.34073e-19 $X=3.465 $Y=0.74 $X2=0
+ $Y2=0
cc_335 N_A_316_413#_M1000_d N_VGND_c_642_n 0.00472095f $X=1.97 $Y=0.235 $X2=0
+ $Y2=0
cc_336 N_A_316_413#_M1002_d N_VGND_c_642_n 0.00256656f $X=2.845 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_A_316_413#_c_409_n N_VGND_c_642_n 0.00851181f $X=3.68 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A_316_413#_c_410_n N_VGND_c_642_n 0.00966829f $X=4.1 $Y=0.995 $X2=0
+ $Y2=0
cc_339 N_A_316_413#_c_514_p N_VGND_c_642_n 0.00625157f $X=2.11 $Y=0.47 $X2=0
+ $Y2=0
cc_340 N_A_316_413#_c_411_n N_VGND_c_642_n 0.0105623f $X=2.895 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_316_413#_c_524_p N_VGND_c_642_n 0.00625722f $X=2.98 $Y=0.47 $X2=0
+ $Y2=0
cc_342 N_A_316_413#_c_413_n N_VGND_c_642_n 0.00638906f $X=3.465 $Y=0.74 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_537_n A_398_413# 0.00214454f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_344 N_VPWR_c_537_n N_X_M1007_s 0.00393857f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_345 N_VPWR_c_541_n N_X_c_603_n 0.0744686f $X=4.335 $Y=1.66 $X2=0 $Y2=0
cc_346 N_VPWR_c_544_n X 0.0168871f $X=4.25 $Y=2.72 $X2=0 $Y2=0
cc_347 N_VPWR_c_537_n X 0.0102668f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_348 N_VPWR_c_541_n N_VGND_c_633_n 0.00845515f $X=4.335 $Y=1.66 $X2=0 $Y2=0
cc_349 N_X_c_605_n N_VGND_c_633_n 0.0250997f $X=3.995 $Y=0.587 $X2=0 $Y2=0
cc_350 N_X_c_603_n N_VGND_c_633_n 0.0187538f $X=3.942 $Y=1.495 $X2=0 $Y2=0
cc_351 N_X_c_605_n N_VGND_c_637_n 0.00796253f $X=3.995 $Y=0.587 $X2=0 $Y2=0
cc_352 N_X_M1006_d N_VGND_c_642_n 0.00409985f $X=3.755 $Y=0.235 $X2=0 $Y2=0
cc_353 N_X_c_605_n N_VGND_c_642_n 0.00913686f $X=3.995 $Y=0.587 $X2=0 $Y2=0

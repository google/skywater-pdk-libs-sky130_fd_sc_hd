* File: sky130_fd_sc_hd__o2bb2ai_2.spice.pex
* Created: Thu Aug 27 14:38:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%A1_N 3 6 10 13 15 19 20 22 25 26 27 30
c77 27 0 1.20878e-19 $X=0.46 $Y=0.995
c78 20 0 1.20678e-19 $X=1.78 $Y=1.16
r79 25 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.16
+ $X2=0.46 $Y2=1.325
r80 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.16
+ $X2=0.46 $Y2=0.995
r81 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=1.16 $X2=0.46 $Y2=1.16
r82 22 36 7.60125 $w=5.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.357 $Y=1.19
+ $X2=0.357 $Y2=1.53
r83 22 26 0.670698 $w=5.33e-07 $l=3e-08 $layer=LI1_cond $X=0.357 $Y=1.19
+ $X2=0.357 $Y2=1.16
r84 20 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.16
+ $X2=1.78 $Y2=1.325
r85 20 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.16
+ $X2=1.78 $Y2=0.995
r86 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=1.16 $X2=1.78 $Y2=1.16
r87 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.78 $Y=1.445
+ $X2=1.78 $Y2=1.16
r88 16 36 7.58357 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.625 $Y=1.53
+ $X2=0.357 $Y2=1.53
r89 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.615 $Y=1.53
+ $X2=1.78 $Y2=1.445
r90 15 16 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.615 $Y=1.53
+ $X2=0.625 $Y2=1.53
r91 13 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.985
+ $X2=1.75 $Y2=1.325
r92 10 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.56
+ $X2=1.75 $Y2=0.995
r93 6 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.985
+ $X2=0.49 $Y2=1.325
r94 3 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.56 $X2=0.49
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%A2_N 1 3 6 8 10 13 15 22
c45 1 0 6.86556e-20 $X=0.91 $Y=0.995
r46 20 22 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.115 $Y=1.16
+ $X2=1.33 $Y2=1.16
r47 17 20 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.115 $Y2=1.16
r48 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.16 $X2=1.115 $Y2=1.16
r49 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r50 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r51 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r52 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r53 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r54 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325 $X2=0.91
+ $Y2=1.985
r55 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995 $X2=0.91
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%A_113_297# 1 2 3 10 12 15 17 19 22 26 28
+ 30 32 33 35 39 40 52
c104 40 0 1.20678e-19 $X=1.54 $Y=1.875
c105 39 0 1.20878e-19 $X=1.285 $Y=0.775
c106 17 0 1.65973e-19 $X=3.12 $Y=0.995
r107 51 52 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.7 $Y=1.16
+ $X2=3.12 $Y2=1.16
r108 48 51 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.49 $Y=1.16
+ $X2=2.7 $Y2=1.16
r109 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.16 $X2=2.49 $Y2=1.16
r110 40 43 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.875
+ $X2=1.54 $Y2=1.96
r111 37 39 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=0.775
+ $X2=1.285 $Y2=0.775
r112 32 47 8.95764 $w=3.29e-07 $l=2.26164e-07 $layer=LI1_cond $X=2.2 $Y=1.325
+ $X2=2.345 $Y2=1.16
r113 32 33 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.2 $Y=1.325
+ $X2=2.2 $Y2=1.785
r114 31 40 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=1.875
+ $X2=1.54 $Y2=1.875
r115 30 33 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.115 $Y=1.875
+ $X2=2.2 $Y2=1.785
r116 30 31 27.7273 $w=1.78e-07 $l=4.5e-07 $layer=LI1_cond $X=2.115 $Y=1.875
+ $X2=1.665 $Y2=1.875
r117 28 47 12.7933 $w=3.29e-07 $l=4.45393e-07 $layer=LI1_cond $X=2.115 $Y=0.815
+ $X2=2.345 $Y2=1.16
r118 28 39 51.1414 $w=1.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.115 $Y=0.815
+ $X2=1.285 $Y2=0.815
r119 27 35 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=1.875
+ $X2=0.7 $Y2=1.875
r120 26 40 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=1.875
+ $X2=1.54 $Y2=1.875
r121 26 27 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=1.415 $Y=1.875
+ $X2=0.825 $Y2=1.875
r122 20 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.325
+ $X2=3.12 $Y2=1.16
r123 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.12 $Y=1.325
+ $X2=3.12 $Y2=1.985
r124 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=1.16
r125 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=0.56
r126 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.16
r127 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.985
r128 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=1.16
r129 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=0.56
r130 3 43 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.96
r131 2 35 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
r132 1 37 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%B1 1 3 6 10 13 17 18 21 22 26 28 31
c83 1 0 2.9244e-20 $X=3.575 $Y=0.995
r84 27 31 9.76796 $w=5.38e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=1.345
+ $X2=4.73 $Y2=1.345
r85 26 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=1.16
+ $X2=4.895 $Y2=1.325
r86 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=1.16
+ $X2=4.895 $Y2=0.995
r87 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.895
+ $Y=1.16 $X2=4.895 $Y2=1.16
r88 22 27 8.74909 $w=5.38e-07 $l=3.95e-07 $layer=LI1_cond $X=5.29 $Y=1.345
+ $X2=4.895 $Y2=1.345
r89 21 31 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=3.74 $Y=1.53
+ $X2=4.73 $Y2=1.53
r90 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.575
+ $Y=1.16 $X2=3.575 $Y2=1.16
r91 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.575 $Y=1.445
+ $X2=3.74 $Y2=1.53
r92 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.575 $Y=1.445
+ $X2=3.575 $Y2=1.16
r93 13 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.835 $Y=1.985
+ $X2=4.835 $Y2=1.325
r94 10 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.835 $Y=0.56
+ $X2=4.835 $Y2=0.995
r95 4 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.325
+ $X2=3.575 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.575 $Y=1.325
+ $X2=3.575 $Y2=1.985
r97 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%B2 1 3 6 8 10 13 15 22
r48 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.205 $Y=1.16
+ $X2=4.415 $Y2=1.16
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.205
+ $Y=1.16 $X2=4.205 $Y2=1.16
r50 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.995 $Y=1.16
+ $X2=4.205 $Y2=1.16
r51 15 21 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.205 $Y2=1.175
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.325
+ $X2=4.415 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.415 $Y=1.325
+ $X2=4.415 $Y2=1.985
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=0.995
+ $X2=4.415 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.415 $Y=0.995
+ $X2=4.415 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.325
+ $X2=3.995 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.995 $Y=1.325
+ $X2=3.995 $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=0.995
+ $X2=3.995 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.995 $Y=0.995
+ $X2=3.995 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%VPWR 1 2 3 4 5 16 18 22 26 30 33 34 35 37
+ 47 57 58 64 69 72 74
r83 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r84 71 72 9.18355 $w=6.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=2.47
+ $X2=2.575 $Y2=2.47
r85 67 71 7.49781 $w=6.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.07 $Y=2.47
+ $X2=2.49 $Y2=2.47
r86 67 69 11.8613 $w=6.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.07 $Y=2.47
+ $X2=1.835 $Y2=2.47
r87 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r90 55 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r91 55 75 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.45 $Y2=2.72
r92 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r93 52 74 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.49 $Y=2.72
+ $X2=3.347 $Y2=2.72
r94 52 54 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=3.49 $Y=2.72
+ $X2=4.83 $Y2=2.72
r95 51 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r96 51 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r97 50 72 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.575 $Y2=2.72
r98 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r99 47 74 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=3.347 $Y2=2.72
r100 47 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=2.99 $Y2=2.72
r101 46 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r102 46 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r103 45 69 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.835 $Y2=2.72
r104 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r105 43 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.12 $Y2=2.72
r106 43 45 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 41 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r108 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r109 38 61 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.2
+ $Y2=2.72
r110 38 40 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.4 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 37 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=1.12 $Y2=2.72
r112 37 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 35 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r115 33 54 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=4.83 $Y2=2.72
r116 33 34 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=5.067 $Y2=2.72
r117 32 57 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.17 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 32 34 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=5.17 $Y=2.72
+ $X2=5.067 $Y2=2.72
r119 28 34 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.067 $Y=2.635
+ $X2=5.067 $Y2=2.72
r120 28 30 36.5188 $w=2.03e-07 $l=6.75e-07 $layer=LI1_cond $X=5.067 $Y=2.635
+ $X2=5.067 $Y2=1.96
r121 24 74 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.347 $Y=2.635
+ $X2=3.347 $Y2=2.72
r122 24 26 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=3.347 $Y=2.635
+ $X2=3.347 $Y2=2.3
r123 20 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r124 20 22 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.3
r125 16 61 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.2 $Y2=2.72
r126 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.275 $Y2=1.96
r127 5 30 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=4.91
+ $Y=1.485 $X2=5.05 $Y2=1.96
r128 4 26 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.485 $X2=3.33 $Y2=2.3
r129 3 71 300 $w=1.7e-07 $l=1.09827e-06 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=2.49 $Y2=2.3
r130 2 22 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r131 1 18 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%Y 1 2 3 12 16 18 20 23 24 29
c47 20 0 3.27631e-20 $X=2.98 $Y=1.31
r48 29 34 2.29036 $w=4.68e-07 $l=9e-08 $layer=LI1_cond $X=2.98 $Y=1.53 $X2=2.98
+ $Y2=1.62
r49 24 27 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.205 $Y=1.87
+ $X2=4.205 $Y2=1.96
r50 22 34 4.199 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.98 $Y=1.785
+ $X2=2.98 $Y2=1.62
r51 22 23 2.53623 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=1.785
+ $X2=2.98 $Y2=1.87
r52 20 29 5.59866 $w=4.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.98 $Y=1.31
+ $X2=2.98 $Y2=1.53
r53 20 21 7.05581 $w=4.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.98 $Y=1.31
+ $X2=2.98 $Y2=1.075
r54 19 23 4.34722 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.215 $Y=1.87
+ $X2=2.98 $Y2=1.87
r55 18 24 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.08 $Y=1.87
+ $X2=4.205 $Y2=1.87
r56 18 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=4.08 $Y=1.87
+ $X2=3.215 $Y2=1.87
r57 14 23 2.53623 $w=3.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.89 $Y=1.955
+ $X2=2.98 $Y2=1.87
r58 14 16 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=2.89 $Y=1.955
+ $X2=2.89 $Y2=1.96
r59 12 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.91 $Y=0.73
+ $X2=2.91 $Y2=1.075
r60 3 27 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.07
+ $Y=1.485 $X2=4.205 $Y2=1.96
r61 2 34 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.485 $X2=2.91 $Y2=1.62
r62 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.775
+ $Y=1.485 $X2=2.91 $Y2=1.96
r63 1 12 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.235 $X2=2.91 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%A_730_297# 1 2 7 11 14
r17 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.785 $Y=2.3 $X2=3.785
+ $Y2=2.38
r18 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.625 $Y=2.295
+ $X2=4.625 $Y2=1.96
r19 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.91 $Y=2.38
+ $X2=3.785 $Y2=2.38
r20 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.5 $Y=2.38
+ $X2=4.625 $Y2=2.295
r21 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.5 $Y=2.38 $X2=3.91
+ $Y2=2.38
r22 2 11 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.485 $X2=4.625 $Y2=1.96
r23 1 14 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=1.485 $X2=3.785 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%VGND 1 2 3 4 13 15 19 23 27 30 31 33 34 36
+ 37 38 57 58
r81 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r82 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r83 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r84 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r85 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r86 49 52 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r87 48 51 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r88 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r89 46 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r90 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r91 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r92 42 45 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r93 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r94 40 61 3.40825 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r95 40 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r96 38 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r97 38 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r98 36 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.37
+ $Y2=0
r99 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.625
+ $Y2=0
r100 35 57 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.71 $Y=0 $X2=5.29
+ $Y2=0
r101 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.71 $Y=0 $X2=4.625
+ $Y2=0
r102 33 51 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.45
+ $Y2=0
r103 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.785
+ $Y2=0
r104 32 54 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=4.37
+ $Y2=0
r105 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0 $X2=3.785
+ $Y2=0
r106 30 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r107 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r108 29 48 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.07
+ $Y2=0
r109 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r110 25 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0
r111 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0.39
r112 21 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0
r113 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0.39
r114 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r115 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r116 13 61 3.40825 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.182 $Y2=0
r117 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.39
r118 4 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.235 $X2=4.625 $Y2=0.39
r119 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.785 $Y2=0.39
r120 2 19 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r121 1 15 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%A_113_47# 1 2 7 9 13
c22 9 0 6.86556e-20 $X=0.7 $Y=0.73
r23 11 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.785 $Y=0.39
+ $X2=0.66 $Y2=0.39
r24 11 13 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.785 $Y=0.39
+ $X2=1.54 $Y2=0.39
r25 7 16 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=0.475 $X2=0.66
+ $Y2=0.39
r26 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.66 $Y=0.475
+ $X2=0.66 $Y2=0.73
r27 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r28 1 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
r29 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_2%A_471_47# 1 2 3 4 13 15 18 19 20 23 25 29
+ 34 37
c66 37 0 2.9244e-20 $X=4.205 $Y=0.815
c67 20 0 1.65973e-19 $X=3.53 $Y=0.82
r68 32 34 4.10683 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.405
+ $X2=2.575 $Y2=0.405
r69 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.045 $Y=0.725
+ $X2=5.045 $Y2=0.39
r70 26 37 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=4.37 $Y=0.815
+ $X2=4.205 $Y2=0.815
r71 25 27 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.88 $Y=0.815
+ $X2=5.045 $Y2=0.725
r72 25 26 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.88 $Y=0.815
+ $X2=4.37 $Y2=0.815
r73 21 37 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.205 $Y=0.725
+ $X2=4.205 $Y2=0.815
r74 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.205 $Y=0.725
+ $X2=4.205 $Y2=0.39
r75 19 37 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.04 $Y=0.82
+ $X2=4.205 $Y2=0.815
r76 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.04 $Y=0.82
+ $X2=3.53 $Y2=0.82
r77 16 20 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.387 $Y=0.735
+ $X2=3.53 $Y2=0.82
r78 16 18 0.202183 $w=2.83e-07 $l=5e-09 $layer=LI1_cond $X=3.387 $Y=0.735
+ $X2=3.387 $Y2=0.73
r79 15 36 3.04002 $w=2.85e-07 $l=1.1e-07 $layer=LI1_cond $X=3.387 $Y=0.475
+ $X2=3.387 $Y2=0.365
r80 15 18 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.387 $Y=0.475
+ $X2=3.387 $Y2=0.73
r81 13 36 3.92439 $w=2.2e-07 $l=1.42e-07 $layer=LI1_cond $X=3.245 $Y=0.365
+ $X2=3.387 $Y2=0.365
r82 13 34 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=3.245 $Y=0.365
+ $X2=2.575 $Y2=0.365
r83 4 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.235 $X2=5.045 $Y2=0.39
r84 3 23 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.07
+ $Y=0.235 $X2=4.205 $Y2=0.39
r85 2 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.235 $X2=3.33 $Y2=0.39
r86 2 18 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.235 $X2=3.33 $Y2=0.73
r87 1 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.49 $Y2=0.39
.ends


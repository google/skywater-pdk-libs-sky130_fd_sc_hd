* NGSPICE file created from sky130_fd_sc_hd__a21boi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR A1 a_217_297# VPB phighvt w=1e+06u l=150000u
+  ad=6.613e+11p pd=6.47e+06u as=1.095e+12p ps=1.019e+07u
M1001 VGND B1_N a_61_47# VNB nshort w=420000u l=150000u
+  ad=7.66e+11p pd=6.31e+06u as=1.26e+11p ps=1.44e+06u
M1002 a_217_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_637_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=3.575e+11p ps=3.7e+06u
M1004 VGND A2 a_637_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_217_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A2 a_217_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_61_47# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_61_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_217_297# a_61_47# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1010 Y A1 a_479_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.365e+11p ps=1.72e+06u
M1011 a_61_47# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1012 Y a_61_47# a_217_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_479_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__bufbuf_16.pxi.spice
* Created: Thu Aug 27 14:10:12 2020
* 
x_PM_SKY130_FD_SC_HD__BUFBUF_16%A N_A_c_241_n N_A_M1049_g N_A_M1032_g A
+ N_A_c_243_n PM_SKY130_FD_SC_HD__BUFBUF_16%A
x_PM_SKY130_FD_SC_HD__BUFBUF_16%A_109_47# N_A_109_47#_M1049_d
+ N_A_109_47#_M1032_d N_A_109_47#_M1006_g N_A_109_47#_M1003_g
+ N_A_109_47#_M1007_g N_A_109_47#_M1034_g N_A_109_47#_M1011_g
+ N_A_109_47#_M1044_g N_A_109_47#_c_272_n N_A_109_47#_c_282_n
+ N_A_109_47#_c_283_n N_A_109_47#_c_273_n N_A_109_47#_c_274_n
+ N_A_109_47#_c_275_n N_A_109_47#_c_276_n N_A_109_47#_c_277_n
+ N_A_109_47#_c_278_n PM_SKY130_FD_SC_HD__BUFBUF_16%A_109_47#
x_PM_SKY130_FD_SC_HD__BUFBUF_16%A_215_47# N_A_215_47#_M1006_d
+ N_A_215_47#_M1007_d N_A_215_47#_M1003_s N_A_215_47#_M1034_s
+ N_A_215_47#_M1010_g N_A_215_47#_M1013_g N_A_215_47#_M1012_g
+ N_A_215_47#_M1014_g N_A_215_47#_M1020_g N_A_215_47#_M1019_g
+ N_A_215_47#_M1021_g N_A_215_47#_M1024_g N_A_215_47#_M1023_g
+ N_A_215_47#_M1025_g N_A_215_47#_M1033_g N_A_215_47#_M1045_g
+ N_A_215_47#_c_372_n N_A_215_47#_c_387_n N_A_215_47#_c_373_n
+ N_A_215_47#_c_374_n N_A_215_47#_c_388_n N_A_215_47#_c_389_n
+ N_A_215_47#_c_416_n N_A_215_47#_c_419_n N_A_215_47#_c_375_n
+ N_A_215_47#_c_376_n N_A_215_47#_c_377_n N_A_215_47#_c_378_n
+ N_A_215_47#_c_391_n N_A_215_47#_c_379_n N_A_215_47#_c_380_n
+ PM_SKY130_FD_SC_HD__BUFBUF_16%A_215_47#
x_PM_SKY130_FD_SC_HD__BUFBUF_16%A_549_47# N_A_549_47#_M1010_s
+ N_A_549_47#_M1020_s N_A_549_47#_M1023_s N_A_549_47#_M1013_s
+ N_A_549_47#_M1019_s N_A_549_47#_M1025_s N_A_549_47#_M1000_g
+ N_A_549_47#_M1001_g N_A_549_47#_M1009_g N_A_549_47#_M1002_g
+ N_A_549_47#_M1017_g N_A_549_47#_M1004_g N_A_549_47#_M1018_g
+ N_A_549_47#_M1005_g N_A_549_47#_M1026_g N_A_549_47#_M1008_g
+ N_A_549_47#_M1027_g N_A_549_47#_M1015_g N_A_549_47#_M1028_g
+ N_A_549_47#_M1016_g N_A_549_47#_M1029_g N_A_549_47#_M1022_g
+ N_A_549_47#_M1035_g N_A_549_47#_M1030_g N_A_549_47#_M1038_g
+ N_A_549_47#_M1031_g N_A_549_47#_M1040_g N_A_549_47#_M1036_g
+ N_A_549_47#_M1041_g N_A_549_47#_M1037_g N_A_549_47#_M1042_g
+ N_A_549_47#_M1039_g N_A_549_47#_M1043_g N_A_549_47#_M1047_g
+ N_A_549_47#_M1046_g N_A_549_47#_M1048_g N_A_549_47#_M1051_g
+ N_A_549_47#_M1050_g N_A_549_47#_c_628_n N_A_549_47#_c_629_n
+ N_A_549_47#_c_596_n N_A_549_47#_c_597_n N_A_549_47#_c_622_n
+ N_A_549_47#_c_623_n N_A_549_47#_c_658_n N_A_549_47#_c_662_n
+ N_A_549_47#_c_598_n N_A_549_47#_c_624_n N_A_549_47#_c_674_n
+ N_A_549_47#_c_677_n N_A_549_47#_c_599_n N_A_549_47#_c_600_n
+ N_A_549_47#_c_601_n N_A_549_47#_c_602_n N_A_549_47#_c_626_n
+ N_A_549_47#_c_603_n N_A_549_47#_c_627_n N_A_549_47#_c_604_n
+ N_A_549_47#_c_605_n PM_SKY130_FD_SC_HD__BUFBUF_16%A_549_47#
x_PM_SKY130_FD_SC_HD__BUFBUF_16%VPWR N_VPWR_M1032_s N_VPWR_M1003_d
+ N_VPWR_M1044_d N_VPWR_M1014_d N_VPWR_M1024_d N_VPWR_M1045_d N_VPWR_M1002_s
+ N_VPWR_M1005_s N_VPWR_M1015_s N_VPWR_M1022_s N_VPWR_M1031_s N_VPWR_M1037_s
+ N_VPWR_M1047_s N_VPWR_M1050_s N_VPWR_c_1029_n N_VPWR_c_1030_n N_VPWR_c_1031_n
+ N_VPWR_c_1032_n N_VPWR_c_1033_n N_VPWR_c_1034_n N_VPWR_c_1035_n
+ N_VPWR_c_1036_n N_VPWR_c_1037_n N_VPWR_c_1038_n N_VPWR_c_1039_n
+ N_VPWR_c_1040_n N_VPWR_c_1041_n N_VPWR_c_1042_n N_VPWR_c_1043_n
+ N_VPWR_c_1044_n N_VPWR_c_1045_n N_VPWR_c_1046_n N_VPWR_c_1047_n
+ N_VPWR_c_1048_n N_VPWR_c_1049_n N_VPWR_c_1050_n N_VPWR_c_1051_n
+ N_VPWR_c_1052_n N_VPWR_c_1053_n N_VPWR_c_1054_n N_VPWR_c_1055_n
+ N_VPWR_c_1056_n N_VPWR_c_1057_n N_VPWR_c_1058_n N_VPWR_c_1059_n
+ N_VPWR_c_1060_n N_VPWR_c_1061_n N_VPWR_c_1062_n N_VPWR_c_1063_n
+ N_VPWR_c_1064_n VPWR N_VPWR_c_1065_n N_VPWR_c_1066_n N_VPWR_c_1067_n
+ N_VPWR_c_1068_n N_VPWR_c_1069_n N_VPWR_c_1028_n VPWR
+ PM_SKY130_FD_SC_HD__BUFBUF_16%VPWR
x_PM_SKY130_FD_SC_HD__BUFBUF_16%X N_X_M1000_s N_X_M1017_s N_X_M1026_s
+ N_X_M1028_s N_X_M1035_s N_X_M1040_s N_X_M1042_s N_X_M1046_s N_X_M1001_d
+ N_X_M1004_d N_X_M1008_d N_X_M1016_d N_X_M1030_d N_X_M1036_d N_X_M1039_d
+ N_X_M1048_d N_X_c_1257_n N_X_c_1255_n N_X_c_1256_n N_X_c_1220_n N_X_c_1221_n
+ N_X_c_1237_n N_X_c_1238_n N_X_c_1285_n N_X_c_1287_n N_X_c_1291_n N_X_c_1222_n
+ N_X_c_1239_n N_X_c_1303_n N_X_c_1305_n N_X_c_1309_n N_X_c_1223_n N_X_c_1240_n
+ N_X_c_1321_n N_X_c_1325_n N_X_c_1224_n N_X_c_1241_n N_X_c_1337_n N_X_c_1341_n
+ N_X_c_1225_n N_X_c_1242_n N_X_c_1353_n N_X_c_1357_n N_X_c_1226_n N_X_c_1243_n
+ N_X_c_1369_n N_X_c_1373_n N_X_c_1227_n N_X_c_1244_n N_X_c_1385_n N_X_c_1388_n
+ N_X_c_1228_n N_X_c_1245_n N_X_c_1229_n N_X_c_1246_n N_X_c_1230_n N_X_c_1247_n
+ N_X_c_1231_n N_X_c_1248_n N_X_c_1232_n N_X_c_1249_n N_X_c_1233_n N_X_c_1250_n
+ N_X_c_1234_n N_X_c_1251_n N_X_c_1235_n N_X_c_1252_n X X
+ PM_SKY130_FD_SC_HD__BUFBUF_16%X
x_PM_SKY130_FD_SC_HD__BUFBUF_16%VGND N_VGND_M1049_s N_VGND_M1006_s
+ N_VGND_M1011_s N_VGND_M1012_d N_VGND_M1021_d N_VGND_M1033_d N_VGND_M1009_d
+ N_VGND_M1018_d N_VGND_M1027_d N_VGND_M1029_d N_VGND_M1038_d N_VGND_M1041_d
+ N_VGND_M1043_d N_VGND_M1051_d N_VGND_c_1557_n N_VGND_c_1558_n N_VGND_c_1559_n
+ N_VGND_c_1560_n N_VGND_c_1561_n N_VGND_c_1562_n N_VGND_c_1563_n
+ N_VGND_c_1564_n N_VGND_c_1565_n N_VGND_c_1566_n N_VGND_c_1567_n
+ N_VGND_c_1568_n N_VGND_c_1569_n N_VGND_c_1570_n N_VGND_c_1571_n
+ N_VGND_c_1572_n N_VGND_c_1573_n N_VGND_c_1574_n N_VGND_c_1575_n
+ N_VGND_c_1576_n N_VGND_c_1577_n N_VGND_c_1578_n N_VGND_c_1579_n
+ N_VGND_c_1580_n N_VGND_c_1581_n N_VGND_c_1582_n N_VGND_c_1583_n
+ N_VGND_c_1584_n N_VGND_c_1585_n N_VGND_c_1586_n N_VGND_c_1587_n
+ N_VGND_c_1588_n N_VGND_c_1589_n N_VGND_c_1590_n N_VGND_c_1591_n
+ N_VGND_c_1592_n VGND N_VGND_c_1593_n N_VGND_c_1594_n N_VGND_c_1595_n
+ N_VGND_c_1596_n N_VGND_c_1597_n N_VGND_c_1598_n VGND
+ PM_SKY130_FD_SC_HD__BUFBUF_16%VGND
cc_1 VNB N_A_c_241_n 0.024747f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_243_n 0.0430997f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_109_47#_M1006_g 0.0216102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_109_47#_M1003_g 5.49071e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_109_47#_M1007_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_109_47#_M1034_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_109_47#_M1011_g 0.0175122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_109_47#_M1044_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_109_47#_c_272_n 0.00452528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_109_47#_c_273_n 0.00455418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_109_47#_c_274_n 0.0210275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_109_47#_c_275_n 0.00238606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_109_47#_c_276_n 7.86138e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_109_47#_c_277_n 0.00275841f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_109_47#_c_278_n 0.0499058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_215_47#_M1010_g 0.0176384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_215_47#_M1013_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_215_47#_M1012_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_215_47#_M1014_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_215_47#_M1020_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_215_47#_M1019_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_215_47#_M1021_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_215_47#_M1024_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_215_47#_M1023_g 0.0172827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_215_47#_M1025_g 4.49807e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_215_47#_M1033_g 0.017512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_215_47#_M1045_g 4.62853e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_215_47#_c_372_n 0.00451034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_215_47#_c_373_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_215_47#_c_374_n 0.004399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_215_47#_c_375_n 0.00354558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_215_47#_c_376_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_215_47#_c_377_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_215_47#_c_378_n 0.00345692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_215_47#_c_379_n 0.0013705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_215_47#_c_380_n 0.0945106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_549_47#_M1000_g 0.0176384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_549_47#_M1001_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_549_47#_M1009_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_549_47#_M1002_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_549_47#_M1017_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_549_47#_M1004_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_549_47#_M1018_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_549_47#_M1005_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_549_47#_M1026_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_549_47#_M1008_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_549_47#_M1027_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_549_47#_M1015_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_549_47#_M1028_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_549_47#_M1016_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_549_47#_M1029_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_549_47#_M1022_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_549_47#_M1035_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_549_47#_M1030_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_549_47#_M1038_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_549_47#_M1031_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_549_47#_M1040_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_549_47#_M1036_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_549_47#_M1041_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_549_47#_M1037_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_549_47#_M1042_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_549_47#_M1039_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_549_47#_M1043_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_549_47#_M1047_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_549_47#_M1046_g 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_549_47#_M1048_g 4.49834e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_549_47#_M1051_g 0.0207727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_549_47#_M1050_g 4.88213e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_549_47#_c_596_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_549_47#_c_597_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_549_47#_c_598_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_549_47#_c_599_n 0.00356912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_549_47#_c_600_n 5.27693e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_549_47#_c_601_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_549_47#_c_602_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_549_47#_c_603_n 0.00344553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_549_47#_c_604_n 0.00154098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_549_47#_c_605_n 0.258232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VPWR_c_1028_n 0.497461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_X_c_1220_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_X_c_1221_n 0.00223017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_X_c_1222_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_X_c_1223_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_X_c_1224_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_X_c_1225_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_X_c_1226_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_X_c_1227_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_X_c_1228_n 0.00875768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_X_c_1229_n 0.00223011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_X_c_1230_n 0.00223011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_X_c_1231_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_X_c_1232_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_X_c_1233_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_X_c_1234_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_X_c_1235_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB X 0.0201563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1557_n 0.0110515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1558_n 0.00654843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1559_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1560_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1561_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1562_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1563_n 0.00358349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1564_n 0.0173761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1565_n 0.00357798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1566_n 0.00357798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1567_n 0.00358349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1568_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1569_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1570_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1571_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1572_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1573_n 0.0106959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1574_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1575_n 0.0168651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1576_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1577_n 0.0174747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1578_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1579_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1580_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1581_n 0.0168651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1582_n 0.00323787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1583_n 0.0168382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1584_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1585_n 0.0168382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1586_n 0.00323972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1587_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1588_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1589_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1590_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1591_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1592_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1593_n 0.0309534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1594_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1595_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1596_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1597_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1598_n 0.552462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VPB N_A_M1032_g 0.0285932f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_141 VPB N_A_c_243_n 0.0123768f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_142 VPB N_A_109_47#_M1003_g 0.0240397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_109_47#_M1034_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_109_47#_M1044_g 0.0194268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_109_47#_c_282_n 0.00244524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_109_47#_c_283_n 0.00786457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_109_47#_c_276_n 0.00376804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_215_47#_M1013_g 0.0196632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_215_47#_M1014_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_215_47#_M1019_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_215_47#_M1024_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_215_47#_M1025_g 0.0191652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_215_47#_M1045_g 0.0194265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_215_47#_c_387_n 0.00784989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_215_47#_c_388_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_215_47#_c_389_n 0.00447011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_215_47#_c_376_n 0.00301948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_215_47#_c_391_n 0.00360324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_549_47#_M1001_g 0.0196632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_549_47#_M1002_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_549_47#_M1004_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_549_47#_M1005_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_549_47#_M1008_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_549_47#_M1015_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_549_47#_M1016_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_549_47#_M1022_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_549_47#_M1030_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_549_47#_M1031_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_549_47#_M1036_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_549_47#_M1037_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_549_47#_M1039_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_549_47#_M1047_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_549_47#_M1048_g 0.0191785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_549_47#_M1050_g 0.0230602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_549_47#_c_622_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_549_47#_c_623_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_549_47#_c_624_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_549_47#_c_600_n 0.00304142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_549_47#_c_626_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_549_47#_c_627_n 0.00359185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1029_n 0.0110239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1030_n 0.00747885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1031_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1032_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1033_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1034_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1035_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1036_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1037_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1038_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1039_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1040_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1041_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1042_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1043_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1044_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1045_n 0.0110239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1046_n 0.00416524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1047_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1048_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1049_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1050_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1051_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1052_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1053_n 0.0178722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1054_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1055_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1056_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1057_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1058_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1059_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1060_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1061_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1062_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1063_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1064_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1065_n 0.0313815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1066_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1067_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1068_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1069_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1028_n 0.0564248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_X_c_1237_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_X_c_1238_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_X_c_1239_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_X_c_1240_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_X_c_1241_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_X_c_1242_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_X_c_1243_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_X_c_1244_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_X_c_1245_n 7.14981e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_X_c_1246_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_X_c_1247_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_X_c_1248_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_X_c_1249_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_X_c_1250_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_X_c_1251_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_X_c_1252_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB X 0.00700926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB X 0.00935206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 N_A_c_241_n N_A_109_47#_c_272_n 0.00551285f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_M1032_g N_A_109_47#_c_282_n 0.00332847f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_M1032_g N_A_109_47#_c_283_n 0.00962957f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A_c_241_n N_A_109_47#_c_273_n 0.0071377f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_c_241_n N_A_109_47#_c_275_n 0.00292436f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_c_243_n N_A_109_47#_c_276_n 0.00698145f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_247 A N_A_109_47#_c_277_n 0.0167772f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_248 N_A_c_243_n N_A_109_47#_c_277_n 0.00563457f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A_c_241_n N_A_215_47#_c_374_n 3.65437e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_M1032_g N_A_215_47#_c_389_n 4.12832e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A_M1032_g N_VPWR_c_1030_n 0.00526624f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_252 A N_VPWR_c_1030_n 0.0136987f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_253 N_A_c_243_n N_VPWR_c_1030_n 0.00415776f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_M1032_g N_VPWR_c_1065_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A_M1032_g N_VPWR_c_1028_n 0.0117818f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A_c_241_n N_VGND_c_1558_n 0.00482486f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_257 A N_VGND_c_1558_n 0.0136981f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_258 N_A_c_243_n N_VGND_c_1558_n 0.00431355f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_c_241_n N_VGND_c_1593_n 0.00541562f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_c_241_n N_VGND_c_1598_n 0.011782f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_109_47#_M1011_g N_A_215_47#_M1010_g 0.021435f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_262 N_A_109_47#_M1044_g N_A_215_47#_M1013_g 0.021435f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_263 N_A_109_47#_M1006_g N_A_215_47#_c_372_n 0.00636826f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_264 N_A_109_47#_M1007_g N_A_215_47#_c_372_n 5.23702e-19 $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_265 N_A_109_47#_c_272_n N_A_215_47#_c_372_n 0.0365376f $X=0.68 $Y=0.4 $X2=0
+ $Y2=0
cc_266 N_A_109_47#_M1003_g N_A_215_47#_c_387_n 0.0102729f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_A_109_47#_M1034_g N_A_215_47#_c_387_n 6.98608e-19 $X=1.83 $Y=1.985
+ $X2=0 $Y2=0
cc_268 N_A_109_47#_c_283_n N_A_215_47#_c_387_n 0.0654134f $X=0.68 $Y=1.63 $X2=0
+ $Y2=0
cc_269 N_A_109_47#_M1006_g N_A_215_47#_c_373_n 0.00850187f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_270 N_A_109_47#_M1007_g N_A_215_47#_c_373_n 0.00850187f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_271 N_A_109_47#_c_274_n N_A_215_47#_c_373_n 0.0596152f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_272 N_A_109_47#_c_278_n N_A_215_47#_c_373_n 0.00205431f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_273 N_A_109_47#_M1006_g N_A_215_47#_c_374_n 0.00126794f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_274 N_A_109_47#_c_272_n N_A_215_47#_c_374_n 0.0138613f $X=0.68 $Y=0.4 $X2=0
+ $Y2=0
cc_275 N_A_109_47#_c_274_n N_A_215_47#_c_374_n 0.0278128f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_276 N_A_109_47#_M1003_g N_A_215_47#_c_388_n 0.0107189f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_277 N_A_109_47#_M1034_g N_A_215_47#_c_388_n 0.0107189f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_278 N_A_109_47#_c_274_n N_A_215_47#_c_388_n 0.0596157f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_279 N_A_109_47#_c_278_n N_A_215_47#_c_388_n 0.00198252f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_280 N_A_109_47#_M1003_g N_A_215_47#_c_389_n 0.00168781f $X=1.41 $Y=1.985
+ $X2=0 $Y2=0
cc_281 N_A_109_47#_c_282_n N_A_215_47#_c_389_n 0.0138613f $X=0.68 $Y=1.61 $X2=0
+ $Y2=0
cc_282 N_A_109_47#_c_274_n N_A_215_47#_c_389_n 0.0279329f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_283 N_A_109_47#_M1006_g N_A_215_47#_c_416_n 5.24491e-19 $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_284 N_A_109_47#_M1007_g N_A_215_47#_c_416_n 0.00647394f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_285 N_A_109_47#_M1011_g N_A_215_47#_c_416_n 0.00647394f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_286 N_A_109_47#_M1003_g N_A_215_47#_c_419_n 6.99397e-19 $X=1.41 $Y=1.985
+ $X2=0 $Y2=0
cc_287 N_A_109_47#_M1034_g N_A_215_47#_c_419_n 0.0103785f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_109_47#_M1044_g N_A_215_47#_c_419_n 0.0103785f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_A_109_47#_M1011_g N_A_215_47#_c_375_n 0.00412488f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_290 N_A_109_47#_c_278_n N_A_215_47#_c_376_n 0.00407173f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_291 N_A_109_47#_M1007_g N_A_215_47#_c_378_n 0.00123754f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_292 N_A_109_47#_M1011_g N_A_215_47#_c_378_n 0.0107176f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_293 N_A_109_47#_c_278_n N_A_215_47#_c_378_n 0.00205431f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_294 N_A_109_47#_M1034_g N_A_215_47#_c_391_n 0.00139111f $X=1.83 $Y=1.985
+ $X2=0 $Y2=0
cc_295 N_A_109_47#_M1044_g N_A_215_47#_c_391_n 0.0131306f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_109_47#_c_278_n N_A_215_47#_c_391_n 0.00198252f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_297 N_A_109_47#_c_274_n N_A_215_47#_c_379_n 0.0176501f $X=1.96 $Y=1.16 $X2=0
+ $Y2=0
cc_298 N_A_109_47#_c_278_n N_A_215_47#_c_379_n 0.00200384f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_299 N_A_109_47#_c_278_n N_A_215_47#_c_380_n 0.021435f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_300 N_A_109_47#_M1011_g N_A_549_47#_c_628_n 5.23702e-19 $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_301 N_A_109_47#_M1044_g N_A_549_47#_c_629_n 6.98608e-19 $X=2.25 $Y=1.985
+ $X2=0 $Y2=0
cc_302 N_A_109_47#_c_282_n N_VPWR_c_1030_n 0.0397026f $X=0.68 $Y=1.61 $X2=0
+ $Y2=0
cc_303 N_A_109_47#_M1003_g N_VPWR_c_1031_n 0.0027696f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_A_109_47#_M1034_g N_VPWR_c_1031_n 0.00154685f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_A_109_47#_M1044_g N_VPWR_c_1032_n 0.00154685f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_306 N_A_109_47#_M1034_g N_VPWR_c_1047_n 0.00541359f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_A_109_47#_M1044_g N_VPWR_c_1047_n 0.00541359f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_308 N_A_109_47#_M1003_g N_VPWR_c_1065_n 0.00541359f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_109_47#_c_283_n N_VPWR_c_1065_n 0.0210382f $X=0.68 $Y=1.63 $X2=0
+ $Y2=0
cc_310 N_A_109_47#_M1032_d N_VPWR_c_1028_n 0.00209319f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_311 N_A_109_47#_M1003_g N_VPWR_c_1028_n 0.0108276f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A_109_47#_M1034_g N_VPWR_c_1028_n 0.00950154f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A_109_47#_M1044_g N_VPWR_c_1028_n 0.00952874f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_109_47#_c_283_n N_VPWR_c_1028_n 0.0124268f $X=0.68 $Y=1.63 $X2=0
+ $Y2=0
cc_315 N_A_109_47#_c_272_n N_VGND_c_1558_n 0.0248793f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_316 N_A_109_47#_M1006_g N_VGND_c_1559_n 0.00268723f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_317 N_A_109_47#_M1007_g N_VGND_c_1559_n 0.00146448f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_318 N_A_109_47#_M1011_g N_VGND_c_1560_n 0.00146448f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_319 N_A_109_47#_M1007_g N_VGND_c_1575_n 0.00423644f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_320 N_A_109_47#_M1011_g N_VGND_c_1575_n 0.00423644f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_321 N_A_109_47#_M1006_g N_VGND_c_1593_n 0.00424619f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_322 N_A_109_47#_c_272_n N_VGND_c_1593_n 0.02038f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_323 N_A_109_47#_M1049_d N_VGND_c_1598_n 0.0020946f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_A_109_47#_M1006_g N_VGND_c_1598_n 0.00706231f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_325 N_A_109_47#_M1007_g N_VGND_c_1598_n 0.00575105f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_326 N_A_109_47#_M1011_g N_VGND_c_1598_n 0.00577825f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_327 N_A_109_47#_c_272_n N_VGND_c_1598_n 0.0123919f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_328 N_A_215_47#_M1033_g N_A_549_47#_M1000_g 0.0214679f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_329 N_A_215_47#_M1045_g N_A_549_47#_M1001_g 0.0214679f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_330 N_A_215_47#_M1010_g N_A_549_47#_c_628_n 0.00636826f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_331 N_A_215_47#_M1012_g N_A_549_47#_c_628_n 0.00636826f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_332 N_A_215_47#_M1020_g N_A_549_47#_c_628_n 5.23702e-19 $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_333 N_A_215_47#_c_416_n N_A_549_47#_c_628_n 0.00518536f $X=2.04 $Y=0.4 $X2=0
+ $Y2=0
cc_334 N_A_215_47#_M1013_g N_A_549_47#_c_629_n 0.0102729f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_215_47#_M1014_g N_A_549_47#_c_629_n 0.0106215f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A_215_47#_M1019_g N_A_549_47#_c_629_n 7.66249e-19 $X=3.51 $Y=1.985
+ $X2=0 $Y2=0
cc_337 N_A_215_47#_c_419_n N_A_549_47#_c_629_n 0.00518536f $X=2.04 $Y=1.63 $X2=0
+ $Y2=0
cc_338 N_A_215_47#_M1012_g N_A_549_47#_c_596_n 0.00850187f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_339 N_A_215_47#_M1020_g N_A_549_47#_c_596_n 0.00850187f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_340 N_A_215_47#_c_377_n N_A_549_47#_c_596_n 0.0359512f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_341 N_A_215_47#_c_380_n N_A_549_47#_c_596_n 0.00205431f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_342 N_A_215_47#_M1010_g N_A_549_47#_c_597_n 0.00240257f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_343 N_A_215_47#_M1012_g N_A_549_47#_c_597_n 0.00109384f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_344 N_A_215_47#_c_377_n N_A_549_47#_c_597_n 0.0265235f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_345 N_A_215_47#_c_378_n N_A_549_47#_c_597_n 0.00795337f $X=2.46 $Y=0.82 $X2=0
+ $Y2=0
cc_346 N_A_215_47#_c_380_n N_A_549_47#_c_597_n 0.00213376f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_347 N_A_215_47#_M1014_g N_A_549_47#_c_622_n 0.0107189f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_A_215_47#_M1019_g N_A_549_47#_c_622_n 0.0107189f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_215_47#_c_377_n N_A_549_47#_c_622_n 0.0359514f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_350 N_A_215_47#_c_380_n N_A_549_47#_c_622_n 0.00198252f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_351 N_A_215_47#_M1013_g N_A_549_47#_c_623_n 0.00265135f $X=2.67 $Y=1.985
+ $X2=0 $Y2=0
cc_352 N_A_215_47#_M1014_g N_A_549_47#_c_623_n 0.00134262f $X=3.09 $Y=1.985
+ $X2=0 $Y2=0
cc_353 N_A_215_47#_c_377_n N_A_549_47#_c_623_n 0.026643f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_354 N_A_215_47#_c_391_n N_A_549_47#_c_623_n 0.0088897f $X=2.46 $Y=1.53 $X2=0
+ $Y2=0
cc_355 N_A_215_47#_c_380_n N_A_549_47#_c_623_n 0.00206439f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_356 N_A_215_47#_M1012_g N_A_549_47#_c_658_n 5.23702e-19 $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_357 N_A_215_47#_M1020_g N_A_549_47#_c_658_n 0.00636826f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_358 N_A_215_47#_M1021_g N_A_549_47#_c_658_n 0.00636826f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_359 N_A_215_47#_M1023_g N_A_549_47#_c_658_n 5.23702e-19 $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_360 N_A_215_47#_M1014_g N_A_549_47#_c_662_n 7.66249e-19 $X=3.09 $Y=1.985
+ $X2=0 $Y2=0
cc_361 N_A_215_47#_M1019_g N_A_549_47#_c_662_n 0.0106215f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_362 N_A_215_47#_M1024_g N_A_549_47#_c_662_n 0.0106215f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_363 N_A_215_47#_M1025_g N_A_549_47#_c_662_n 7.66249e-19 $X=4.35 $Y=1.985
+ $X2=0 $Y2=0
cc_364 N_A_215_47#_M1021_g N_A_549_47#_c_598_n 0.00850187f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_A_215_47#_M1023_g N_A_549_47#_c_598_n 0.00850187f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_366 N_A_215_47#_c_377_n N_A_549_47#_c_598_n 0.0568321f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_367 N_A_215_47#_c_380_n N_A_549_47#_c_598_n 0.00205431f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_368 N_A_215_47#_M1024_g N_A_549_47#_c_624_n 0.0107189f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_A_215_47#_M1025_g N_A_549_47#_c_624_n 0.0107189f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A_215_47#_c_377_n N_A_549_47#_c_624_n 0.0568326f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_371 N_A_215_47#_c_380_n N_A_549_47#_c_624_n 0.00198252f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_372 N_A_215_47#_M1021_g N_A_549_47#_c_674_n 5.24491e-19 $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_373 N_A_215_47#_M1023_g N_A_549_47#_c_674_n 0.00647394f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_374 N_A_215_47#_M1033_g N_A_549_47#_c_674_n 0.00647394f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_375 N_A_215_47#_M1024_g N_A_549_47#_c_677_n 7.67038e-19 $X=3.93 $Y=1.985
+ $X2=0 $Y2=0
cc_376 N_A_215_47#_M1025_g N_A_549_47#_c_677_n 0.0107272f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_377 N_A_215_47#_M1045_g N_A_549_47#_c_677_n 0.0107272f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_378 N_A_215_47#_M1033_g N_A_549_47#_c_599_n 0.00417409f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_379 N_A_215_47#_c_380_n N_A_549_47#_c_600_n 0.00412038f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_380 N_A_215_47#_M1020_g N_A_549_47#_c_602_n 0.00110541f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_381 N_A_215_47#_M1021_g N_A_549_47#_c_602_n 0.00110541f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_382 N_A_215_47#_c_377_n N_A_549_47#_c_602_n 0.0265235f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_383 N_A_215_47#_c_380_n N_A_549_47#_c_602_n 0.00213376f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_384 N_A_215_47#_M1019_g N_A_549_47#_c_626_n 0.00135419f $X=3.51 $Y=1.985
+ $X2=0 $Y2=0
cc_385 N_A_215_47#_M1024_g N_A_549_47#_c_626_n 0.00135419f $X=3.93 $Y=1.985
+ $X2=0 $Y2=0
cc_386 N_A_215_47#_c_377_n N_A_549_47#_c_626_n 0.026643f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_387 N_A_215_47#_c_380_n N_A_549_47#_c_626_n 0.00206439f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_388 N_A_215_47#_M1023_g N_A_549_47#_c_603_n 0.00123754f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_389 N_A_215_47#_M1033_g N_A_549_47#_c_603_n 0.0110598f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_390 N_A_215_47#_c_380_n N_A_549_47#_c_603_n 0.00205431f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_391 N_A_215_47#_M1025_g N_A_549_47#_c_627_n 0.00139111f $X=4.35 $Y=1.985
+ $X2=0 $Y2=0
cc_392 N_A_215_47#_M1045_g N_A_549_47#_c_627_n 0.0134729f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_393 N_A_215_47#_c_380_n N_A_549_47#_c_627_n 0.00198252f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_394 N_A_215_47#_c_377_n N_A_549_47#_c_604_n 0.015316f $X=4.5 $Y=1.16 $X2=0
+ $Y2=0
cc_395 N_A_215_47#_c_380_n N_A_549_47#_c_604_n 0.00217042f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_396 N_A_215_47#_c_380_n N_A_549_47#_c_605_n 0.0214679f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_397 N_A_215_47#_c_388_n N_VPWR_M1003_d 0.00165831f $X=1.875 $Y=1.53 $X2=0
+ $Y2=0
cc_398 N_A_215_47#_c_391_n N_VPWR_M1044_d 0.00187252f $X=2.46 $Y=1.53 $X2=0
+ $Y2=0
cc_399 N_A_215_47#_c_388_n N_VPWR_c_1031_n 0.0126919f $X=1.875 $Y=1.53 $X2=0
+ $Y2=0
cc_400 N_A_215_47#_M1013_g N_VPWR_c_1032_n 0.00154685f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_401 N_A_215_47#_c_391_n N_VPWR_c_1032_n 0.0126919f $X=2.46 $Y=1.53 $X2=0
+ $Y2=0
cc_402 N_A_215_47#_M1014_g N_VPWR_c_1033_n 0.00146448f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_403 N_A_215_47#_M1019_g N_VPWR_c_1033_n 0.00146448f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_404 N_A_215_47#_M1024_g N_VPWR_c_1034_n 0.00146448f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_405 N_A_215_47#_M1025_g N_VPWR_c_1034_n 0.00146448f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_406 N_A_215_47#_M1045_g N_VPWR_c_1035_n 0.00146448f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_407 N_A_215_47#_c_419_n N_VPWR_c_1047_n 0.0189039f $X=2.04 $Y=1.63 $X2=0
+ $Y2=0
cc_408 N_A_215_47#_M1013_g N_VPWR_c_1049_n 0.00541359f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A_215_47#_M1014_g N_VPWR_c_1049_n 0.00541359f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_410 N_A_215_47#_M1019_g N_VPWR_c_1051_n 0.00541359f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_411 N_A_215_47#_M1024_g N_VPWR_c_1051_n 0.00541359f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_412 N_A_215_47#_M1025_g N_VPWR_c_1053_n 0.00541359f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_413 N_A_215_47#_M1045_g N_VPWR_c_1053_n 0.00541359f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_414 N_A_215_47#_c_387_n N_VPWR_c_1065_n 0.0210382f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_415 N_A_215_47#_M1003_s N_VPWR_c_1028_n 0.00209319f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_416 N_A_215_47#_M1034_s N_VPWR_c_1028_n 0.00215201f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_417 N_A_215_47#_M1013_g N_VPWR_c_1028_n 0.00952874f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_A_215_47#_M1014_g N_VPWR_c_1028_n 0.00950154f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_419 N_A_215_47#_M1019_g N_VPWR_c_1028_n 0.00950154f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A_215_47#_M1024_g N_VPWR_c_1028_n 0.00950154f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_421 N_A_215_47#_M1025_g N_VPWR_c_1028_n 0.00950154f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_422 N_A_215_47#_M1045_g N_VPWR_c_1028_n 0.00952874f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_423 N_A_215_47#_c_387_n N_VPWR_c_1028_n 0.0124268f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_424 N_A_215_47#_c_419_n N_VPWR_c_1028_n 0.0122217f $X=2.04 $Y=1.63 $X2=0
+ $Y2=0
cc_425 N_A_215_47#_M1033_g N_X_c_1255_n 4.74777e-19 $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_426 N_A_215_47#_M1045_g N_X_c_1256_n 7.66249e-19 $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_427 N_A_215_47#_c_373_n N_VGND_M1006_s 0.00162006f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_428 N_A_215_47#_c_378_n N_VGND_M1011_s 0.00186748f $X=2.46 $Y=0.82 $X2=0
+ $Y2=0
cc_429 N_A_215_47#_c_373_n N_VGND_c_1559_n 0.0122414f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_430 N_A_215_47#_M1010_g N_VGND_c_1560_n 0.00146448f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_431 N_A_215_47#_c_378_n N_VGND_c_1560_n 0.0122414f $X=2.46 $Y=0.82 $X2=0
+ $Y2=0
cc_432 N_A_215_47#_M1012_g N_VGND_c_1561_n 0.00146448f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_433 N_A_215_47#_M1020_g N_VGND_c_1561_n 0.00146448f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_434 N_A_215_47#_M1021_g N_VGND_c_1562_n 0.00146448f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_435 N_A_215_47#_M1023_g N_VGND_c_1562_n 0.00146448f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_436 N_A_215_47#_M1033_g N_VGND_c_1563_n 0.00146448f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_437 N_A_215_47#_c_373_n N_VGND_c_1575_n 0.00390702f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_438 N_A_215_47#_c_416_n N_VGND_c_1575_n 0.0179571f $X=2.04 $Y=0.4 $X2=0 $Y2=0
cc_439 N_A_215_47#_M1010_g N_VGND_c_1577_n 0.00541562f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_440 N_A_215_47#_M1012_g N_VGND_c_1577_n 0.00424619f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_441 N_A_215_47#_M1020_g N_VGND_c_1579_n 0.00424619f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_442 N_A_215_47#_M1021_g N_VGND_c_1579_n 0.00424619f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_443 N_A_215_47#_M1023_g N_VGND_c_1581_n 0.00423644f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_444 N_A_215_47#_M1033_g N_VGND_c_1581_n 0.00423644f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_445 N_A_215_47#_c_372_n N_VGND_c_1593_n 0.020318f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_446 N_A_215_47#_c_373_n N_VGND_c_1593_n 0.00193763f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_447 N_A_215_47#_M1006_d N_VGND_c_1598_n 0.0020946f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_448 N_A_215_47#_M1007_d N_VGND_c_1598_n 0.00215347f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_449 N_A_215_47#_M1010_g N_VGND_c_1598_n 0.00952891f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_450 N_A_215_47#_M1012_g N_VGND_c_1598_n 0.00573624f $X=3.09 $Y=0.56 $X2=0
+ $Y2=0
cc_451 N_A_215_47#_M1020_g N_VGND_c_1598_n 0.00573624f $X=3.51 $Y=0.56 $X2=0
+ $Y2=0
cc_452 N_A_215_47#_M1021_g N_VGND_c_1598_n 0.00573624f $X=3.93 $Y=0.56 $X2=0
+ $Y2=0
cc_453 N_A_215_47#_M1023_g N_VGND_c_1598_n 0.00575105f $X=4.35 $Y=0.56 $X2=0
+ $Y2=0
cc_454 N_A_215_47#_M1033_g N_VGND_c_1598_n 0.00577825f $X=4.77 $Y=0.56 $X2=0
+ $Y2=0
cc_455 N_A_215_47#_c_372_n N_VGND_c_1598_n 0.0123792f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_456 N_A_215_47#_c_373_n N_VGND_c_1598_n 0.012122f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_457 N_A_215_47#_c_416_n N_VGND_c_1598_n 0.0120759f $X=2.04 $Y=0.4 $X2=0 $Y2=0
cc_458 N_A_215_47#_c_378_n N_VGND_c_1598_n 6.28727e-19 $X=2.46 $Y=0.82 $X2=0
+ $Y2=0
cc_459 N_A_549_47#_c_622_n N_VPWR_M1014_d 0.00185611f $X=3.555 $Y=1.53 $X2=0
+ $Y2=0
cc_460 N_A_549_47#_c_624_n N_VPWR_M1024_d 0.00185611f $X=4.395 $Y=1.53 $X2=0
+ $Y2=0
cc_461 N_A_549_47#_c_627_n N_VPWR_M1045_d 0.00207031f $X=4.977 $Y=1.53 $X2=0
+ $Y2=0
cc_462 N_A_549_47#_c_622_n N_VPWR_c_1033_n 0.0104788f $X=3.555 $Y=1.53 $X2=0
+ $Y2=0
cc_463 N_A_549_47#_c_624_n N_VPWR_c_1034_n 0.0104788f $X=4.395 $Y=1.53 $X2=0
+ $Y2=0
cc_464 N_A_549_47#_M1001_g N_VPWR_c_1035_n 0.00146448f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_465 N_A_549_47#_c_627_n N_VPWR_c_1035_n 0.0104788f $X=4.977 $Y=1.53 $X2=0
+ $Y2=0
cc_466 N_A_549_47#_M1001_g N_VPWR_c_1036_n 0.00541359f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_467 N_A_549_47#_M1002_g N_VPWR_c_1036_n 0.00541359f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_468 N_A_549_47#_M1002_g N_VPWR_c_1037_n 0.00146448f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_469 N_A_549_47#_M1004_g N_VPWR_c_1037_n 0.00146448f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_470 N_A_549_47#_M1005_g N_VPWR_c_1038_n 0.00146448f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_471 N_A_549_47#_M1008_g N_VPWR_c_1038_n 0.00146448f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_472 N_A_549_47#_M1015_g N_VPWR_c_1039_n 0.00146448f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_A_549_47#_M1016_g N_VPWR_c_1039_n 0.00146448f $X=7.71 $Y=1.985 $X2=0
+ $Y2=0
cc_474 N_A_549_47#_M1022_g N_VPWR_c_1040_n 0.00146448f $X=8.13 $Y=1.985 $X2=0
+ $Y2=0
cc_475 N_A_549_47#_M1030_g N_VPWR_c_1040_n 0.00146448f $X=8.55 $Y=1.985 $X2=0
+ $Y2=0
cc_476 N_A_549_47#_M1031_g N_VPWR_c_1041_n 0.00146448f $X=8.97 $Y=1.985 $X2=0
+ $Y2=0
cc_477 N_A_549_47#_M1036_g N_VPWR_c_1041_n 0.00146448f $X=9.39 $Y=1.985 $X2=0
+ $Y2=0
cc_478 N_A_549_47#_M1037_g N_VPWR_c_1042_n 0.00146448f $X=9.81 $Y=1.985 $X2=0
+ $Y2=0
cc_479 N_A_549_47#_M1039_g N_VPWR_c_1042_n 0.00146448f $X=10.23 $Y=1.985 $X2=0
+ $Y2=0
cc_480 N_A_549_47#_M1039_g N_VPWR_c_1043_n 0.00541359f $X=10.23 $Y=1.985 $X2=0
+ $Y2=0
cc_481 N_A_549_47#_M1047_g N_VPWR_c_1043_n 0.00541359f $X=10.65 $Y=1.985 $X2=0
+ $Y2=0
cc_482 N_A_549_47#_M1047_g N_VPWR_c_1044_n 0.00146448f $X=10.65 $Y=1.985 $X2=0
+ $Y2=0
cc_483 N_A_549_47#_M1048_g N_VPWR_c_1044_n 0.00146448f $X=11.07 $Y=1.985 $X2=0
+ $Y2=0
cc_484 N_A_549_47#_M1050_g N_VPWR_c_1046_n 0.00316354f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_A_549_47#_c_629_n N_VPWR_c_1049_n 0.0189039f $X=2.88 $Y=1.63 $X2=0
+ $Y2=0
cc_486 N_A_549_47#_c_662_n N_VPWR_c_1051_n 0.0189039f $X=3.72 $Y=1.63 $X2=0
+ $Y2=0
cc_487 N_A_549_47#_c_677_n N_VPWR_c_1053_n 0.0189039f $X=4.56 $Y=1.63 $X2=0
+ $Y2=0
cc_488 N_A_549_47#_M1004_g N_VPWR_c_1055_n 0.00541359f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_489 N_A_549_47#_M1005_g N_VPWR_c_1055_n 0.00541359f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_490 N_A_549_47#_M1008_g N_VPWR_c_1057_n 0.00541359f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_491 N_A_549_47#_M1015_g N_VPWR_c_1057_n 0.00541359f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_492 N_A_549_47#_M1016_g N_VPWR_c_1059_n 0.00541359f $X=7.71 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_A_549_47#_M1022_g N_VPWR_c_1059_n 0.00541359f $X=8.13 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_A_549_47#_M1030_g N_VPWR_c_1061_n 0.00541359f $X=8.55 $Y=1.985 $X2=0
+ $Y2=0
cc_495 N_A_549_47#_M1031_g N_VPWR_c_1061_n 0.00541359f $X=8.97 $Y=1.985 $X2=0
+ $Y2=0
cc_496 N_A_549_47#_M1036_g N_VPWR_c_1063_n 0.00541359f $X=9.39 $Y=1.985 $X2=0
+ $Y2=0
cc_497 N_A_549_47#_M1037_g N_VPWR_c_1063_n 0.00541359f $X=9.81 $Y=1.985 $X2=0
+ $Y2=0
cc_498 N_A_549_47#_M1048_g N_VPWR_c_1066_n 0.00541359f $X=11.07 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A_549_47#_M1050_g N_VPWR_c_1066_n 0.00541359f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_500 N_A_549_47#_M1013_s N_VPWR_c_1028_n 0.00215201f $X=2.745 $Y=1.485 $X2=0
+ $Y2=0
cc_501 N_A_549_47#_M1019_s N_VPWR_c_1028_n 0.00215201f $X=3.585 $Y=1.485 $X2=0
+ $Y2=0
cc_502 N_A_549_47#_M1025_s N_VPWR_c_1028_n 0.00215201f $X=4.425 $Y=1.485 $X2=0
+ $Y2=0
cc_503 N_A_549_47#_M1001_g N_VPWR_c_1028_n 0.00952874f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_504 N_A_549_47#_M1002_g N_VPWR_c_1028_n 0.00950154f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_505 N_A_549_47#_M1004_g N_VPWR_c_1028_n 0.00950154f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_506 N_A_549_47#_M1005_g N_VPWR_c_1028_n 0.00950154f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_507 N_A_549_47#_M1008_g N_VPWR_c_1028_n 0.00950154f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_508 N_A_549_47#_M1015_g N_VPWR_c_1028_n 0.00950154f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_509 N_A_549_47#_M1016_g N_VPWR_c_1028_n 0.00950154f $X=7.71 $Y=1.985 $X2=0
+ $Y2=0
cc_510 N_A_549_47#_M1022_g N_VPWR_c_1028_n 0.00950154f $X=8.13 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_A_549_47#_M1030_g N_VPWR_c_1028_n 0.00950154f $X=8.55 $Y=1.985 $X2=0
+ $Y2=0
cc_512 N_A_549_47#_M1031_g N_VPWR_c_1028_n 0.00950154f $X=8.97 $Y=1.985 $X2=0
+ $Y2=0
cc_513 N_A_549_47#_M1036_g N_VPWR_c_1028_n 0.00950154f $X=9.39 $Y=1.985 $X2=0
+ $Y2=0
cc_514 N_A_549_47#_M1037_g N_VPWR_c_1028_n 0.00950154f $X=9.81 $Y=1.985 $X2=0
+ $Y2=0
cc_515 N_A_549_47#_M1039_g N_VPWR_c_1028_n 0.00950154f $X=10.23 $Y=1.985 $X2=0
+ $Y2=0
cc_516 N_A_549_47#_M1047_g N_VPWR_c_1028_n 0.00950154f $X=10.65 $Y=1.985 $X2=0
+ $Y2=0
cc_517 N_A_549_47#_M1048_g N_VPWR_c_1028_n 0.00950154f $X=11.07 $Y=1.985 $X2=0
+ $Y2=0
cc_518 N_A_549_47#_M1050_g N_VPWR_c_1028_n 0.0104557f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_519 N_A_549_47#_c_629_n N_VPWR_c_1028_n 0.0122217f $X=2.88 $Y=1.63 $X2=0
+ $Y2=0
cc_520 N_A_549_47#_c_662_n N_VPWR_c_1028_n 0.0122217f $X=3.72 $Y=1.63 $X2=0
+ $Y2=0
cc_521 N_A_549_47#_c_677_n N_VPWR_c_1028_n 0.0122217f $X=4.56 $Y=1.63 $X2=0
+ $Y2=0
cc_522 N_A_549_47#_M1000_g N_X_c_1257_n 0.00202914f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_523 N_A_549_47#_M1009_g N_X_c_1257_n 0.00198339f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_524 N_A_549_47#_M1000_g N_X_c_1255_n 0.00439074f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_525 N_A_549_47#_M1009_g N_X_c_1255_n 0.00439074f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_526 N_A_549_47#_M1017_g N_X_c_1255_n 4.74777e-19 $X=6.03 $Y=0.56 $X2=0 $Y2=0
cc_527 N_A_549_47#_c_674_n N_X_c_1255_n 0.00518536f $X=4.56 $Y=0.4 $X2=0 $Y2=0
cc_528 N_A_549_47#_M1001_g N_X_c_1256_n 0.0106215f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_529 N_A_549_47#_M1002_g N_X_c_1256_n 0.0106215f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_530 N_A_549_47#_M1004_g N_X_c_1256_n 7.66249e-19 $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_531 N_A_549_47#_c_677_n N_X_c_1256_n 0.00671496f $X=4.56 $Y=1.63 $X2=0 $Y2=0
cc_532 N_A_549_47#_M1009_g N_X_c_1220_n 0.00850187f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_533 N_A_549_47#_M1017_g N_X_c_1220_n 0.00850187f $X=6.03 $Y=0.56 $X2=0 $Y2=0
cc_534 N_A_549_47#_c_601_n N_X_c_1220_n 0.0359512f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_535 N_A_549_47#_c_605_n N_X_c_1220_n 0.00205431f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_536 N_A_549_47#_M1000_g N_X_c_1221_n 0.00241717f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_537 N_A_549_47#_M1009_g N_X_c_1221_n 0.0011083f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_538 N_A_549_47#_c_601_n N_X_c_1221_n 0.0265361f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_539 N_A_549_47#_c_603_n N_X_c_1221_n 0.00795337f $X=4.977 $Y=0.82 $X2=0 $Y2=0
cc_540 N_A_549_47#_c_605_n N_X_c_1221_n 0.00213429f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_541 N_A_549_47#_M1002_g N_X_c_1237_n 0.0107189f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_542 N_A_549_47#_M1004_g N_X_c_1237_n 0.0107189f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_543 N_A_549_47#_c_601_n N_X_c_1237_n 0.0359514f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_544 N_A_549_47#_c_605_n N_X_c_1237_n 0.00198252f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_545 N_A_549_47#_M1001_g N_X_c_1238_n 0.00265135f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_546 N_A_549_47#_M1002_g N_X_c_1238_n 0.00134262f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_547 N_A_549_47#_c_601_n N_X_c_1238_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_548 N_A_549_47#_c_627_n N_X_c_1238_n 0.0088897f $X=4.977 $Y=1.53 $X2=0 $Y2=0
cc_549 N_A_549_47#_c_605_n N_X_c_1238_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_550 N_A_549_47#_M1017_g N_X_c_1285_n 0.00198339f $X=6.03 $Y=0.56 $X2=0 $Y2=0
cc_551 N_A_549_47#_M1018_g N_X_c_1285_n 0.00198339f $X=6.45 $Y=0.56 $X2=0 $Y2=0
cc_552 N_A_549_47#_M1009_g N_X_c_1287_n 4.74777e-19 $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_553 N_A_549_47#_M1017_g N_X_c_1287_n 0.00439074f $X=6.03 $Y=0.56 $X2=0 $Y2=0
cc_554 N_A_549_47#_M1018_g N_X_c_1287_n 0.00439074f $X=6.45 $Y=0.56 $X2=0 $Y2=0
cc_555 N_A_549_47#_M1026_g N_X_c_1287_n 4.74777e-19 $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_556 N_A_549_47#_M1002_g N_X_c_1291_n 7.66249e-19 $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_557 N_A_549_47#_M1004_g N_X_c_1291_n 0.0106215f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_558 N_A_549_47#_M1005_g N_X_c_1291_n 0.0106215f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_559 N_A_549_47#_M1008_g N_X_c_1291_n 7.66249e-19 $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_560 N_A_549_47#_M1018_g N_X_c_1222_n 0.00850187f $X=6.45 $Y=0.56 $X2=0 $Y2=0
cc_561 N_A_549_47#_M1026_g N_X_c_1222_n 0.00850187f $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_562 N_A_549_47#_c_601_n N_X_c_1222_n 0.0359512f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_563 N_A_549_47#_c_605_n N_X_c_1222_n 0.00205431f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_564 N_A_549_47#_M1005_g N_X_c_1239_n 0.0107189f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_565 N_A_549_47#_M1008_g N_X_c_1239_n 0.0107189f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_566 N_A_549_47#_c_601_n N_X_c_1239_n 0.0359514f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_567 N_A_549_47#_c_605_n N_X_c_1239_n 0.00198252f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_568 N_A_549_47#_M1026_g N_X_c_1303_n 0.00198339f $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_569 N_A_549_47#_M1027_g N_X_c_1303_n 0.00198339f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_570 N_A_549_47#_M1018_g N_X_c_1305_n 4.74777e-19 $X=6.45 $Y=0.56 $X2=0 $Y2=0
cc_571 N_A_549_47#_M1026_g N_X_c_1305_n 0.00439074f $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_572 N_A_549_47#_M1027_g N_X_c_1305_n 0.00439074f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_573 N_A_549_47#_M1028_g N_X_c_1305_n 4.74777e-19 $X=7.71 $Y=0.56 $X2=0 $Y2=0
cc_574 N_A_549_47#_M1005_g N_X_c_1309_n 7.66249e-19 $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_575 N_A_549_47#_M1008_g N_X_c_1309_n 0.0106215f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_576 N_A_549_47#_M1015_g N_X_c_1309_n 0.0106215f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_577 N_A_549_47#_M1016_g N_X_c_1309_n 7.66249e-19 $X=7.71 $Y=1.985 $X2=0 $Y2=0
cc_578 N_A_549_47#_M1027_g N_X_c_1223_n 0.00850187f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_579 N_A_549_47#_M1028_g N_X_c_1223_n 0.00850187f $X=7.71 $Y=0.56 $X2=0 $Y2=0
cc_580 N_A_549_47#_c_601_n N_X_c_1223_n 0.0359512f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_581 N_A_549_47#_c_605_n N_X_c_1223_n 0.00205431f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_582 N_A_549_47#_M1015_g N_X_c_1240_n 0.0107189f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_583 N_A_549_47#_M1016_g N_X_c_1240_n 0.0107189f $X=7.71 $Y=1.985 $X2=0 $Y2=0
cc_584 N_A_549_47#_c_601_n N_X_c_1240_n 0.0359514f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_585 N_A_549_47#_c_605_n N_X_c_1240_n 0.00198252f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_586 N_A_549_47#_M1027_g N_X_c_1321_n 5.23702e-19 $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_587 N_A_549_47#_M1028_g N_X_c_1321_n 0.00636826f $X=7.71 $Y=0.56 $X2=0 $Y2=0
cc_588 N_A_549_47#_M1029_g N_X_c_1321_n 0.00636826f $X=8.13 $Y=0.56 $X2=0 $Y2=0
cc_589 N_A_549_47#_M1035_g N_X_c_1321_n 5.23702e-19 $X=8.55 $Y=0.56 $X2=0 $Y2=0
cc_590 N_A_549_47#_M1015_g N_X_c_1325_n 7.66249e-19 $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_591 N_A_549_47#_M1016_g N_X_c_1325_n 0.0106215f $X=7.71 $Y=1.985 $X2=0 $Y2=0
cc_592 N_A_549_47#_M1022_g N_X_c_1325_n 0.0106215f $X=8.13 $Y=1.985 $X2=0 $Y2=0
cc_593 N_A_549_47#_M1030_g N_X_c_1325_n 7.66249e-19 $X=8.55 $Y=1.985 $X2=0 $Y2=0
cc_594 N_A_549_47#_M1029_g N_X_c_1224_n 0.00850187f $X=8.13 $Y=0.56 $X2=0 $Y2=0
cc_595 N_A_549_47#_M1035_g N_X_c_1224_n 0.00850187f $X=8.55 $Y=0.56 $X2=0 $Y2=0
cc_596 N_A_549_47#_c_601_n N_X_c_1224_n 0.0359512f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_597 N_A_549_47#_c_605_n N_X_c_1224_n 0.00205431f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_598 N_A_549_47#_M1022_g N_X_c_1241_n 0.0107189f $X=8.13 $Y=1.985 $X2=0 $Y2=0
cc_599 N_A_549_47#_M1030_g N_X_c_1241_n 0.0107189f $X=8.55 $Y=1.985 $X2=0 $Y2=0
cc_600 N_A_549_47#_c_601_n N_X_c_1241_n 0.0359514f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_601 N_A_549_47#_c_605_n N_X_c_1241_n 0.00198252f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_602 N_A_549_47#_M1029_g N_X_c_1337_n 5.23702e-19 $X=8.13 $Y=0.56 $X2=0 $Y2=0
cc_603 N_A_549_47#_M1035_g N_X_c_1337_n 0.00636826f $X=8.55 $Y=0.56 $X2=0 $Y2=0
cc_604 N_A_549_47#_M1038_g N_X_c_1337_n 0.00636826f $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_605 N_A_549_47#_M1040_g N_X_c_1337_n 5.23702e-19 $X=9.39 $Y=0.56 $X2=0 $Y2=0
cc_606 N_A_549_47#_M1022_g N_X_c_1341_n 7.66249e-19 $X=8.13 $Y=1.985 $X2=0 $Y2=0
cc_607 N_A_549_47#_M1030_g N_X_c_1341_n 0.0106215f $X=8.55 $Y=1.985 $X2=0 $Y2=0
cc_608 N_A_549_47#_M1031_g N_X_c_1341_n 0.0106215f $X=8.97 $Y=1.985 $X2=0 $Y2=0
cc_609 N_A_549_47#_M1036_g N_X_c_1341_n 7.66249e-19 $X=9.39 $Y=1.985 $X2=0 $Y2=0
cc_610 N_A_549_47#_M1038_g N_X_c_1225_n 0.00850187f $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_611 N_A_549_47#_M1040_g N_X_c_1225_n 0.00850187f $X=9.39 $Y=0.56 $X2=0 $Y2=0
cc_612 N_A_549_47#_c_601_n N_X_c_1225_n 0.0359512f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_613 N_A_549_47#_c_605_n N_X_c_1225_n 0.00205431f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_614 N_A_549_47#_M1031_g N_X_c_1242_n 0.0107189f $X=8.97 $Y=1.985 $X2=0 $Y2=0
cc_615 N_A_549_47#_M1036_g N_X_c_1242_n 0.0107189f $X=9.39 $Y=1.985 $X2=0 $Y2=0
cc_616 N_A_549_47#_c_601_n N_X_c_1242_n 0.0359514f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_617 N_A_549_47#_c_605_n N_X_c_1242_n 0.00198252f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_618 N_A_549_47#_M1038_g N_X_c_1353_n 5.23702e-19 $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_619 N_A_549_47#_M1040_g N_X_c_1353_n 0.00636826f $X=9.39 $Y=0.56 $X2=0 $Y2=0
cc_620 N_A_549_47#_M1041_g N_X_c_1353_n 0.00636826f $X=9.81 $Y=0.56 $X2=0 $Y2=0
cc_621 N_A_549_47#_M1042_g N_X_c_1353_n 5.23702e-19 $X=10.23 $Y=0.56 $X2=0 $Y2=0
cc_622 N_A_549_47#_M1031_g N_X_c_1357_n 7.66249e-19 $X=8.97 $Y=1.985 $X2=0 $Y2=0
cc_623 N_A_549_47#_M1036_g N_X_c_1357_n 0.0106215f $X=9.39 $Y=1.985 $X2=0 $Y2=0
cc_624 N_A_549_47#_M1037_g N_X_c_1357_n 0.0106215f $X=9.81 $Y=1.985 $X2=0 $Y2=0
cc_625 N_A_549_47#_M1039_g N_X_c_1357_n 7.66249e-19 $X=10.23 $Y=1.985 $X2=0
+ $Y2=0
cc_626 N_A_549_47#_M1041_g N_X_c_1226_n 0.00850187f $X=9.81 $Y=0.56 $X2=0 $Y2=0
cc_627 N_A_549_47#_M1042_g N_X_c_1226_n 0.00850187f $X=10.23 $Y=0.56 $X2=0 $Y2=0
cc_628 N_A_549_47#_c_601_n N_X_c_1226_n 0.0359512f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_629 N_A_549_47#_c_605_n N_X_c_1226_n 0.00205431f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_630 N_A_549_47#_M1037_g N_X_c_1243_n 0.0107189f $X=9.81 $Y=1.985 $X2=0 $Y2=0
cc_631 N_A_549_47#_M1039_g N_X_c_1243_n 0.0107189f $X=10.23 $Y=1.985 $X2=0 $Y2=0
cc_632 N_A_549_47#_c_601_n N_X_c_1243_n 0.0359514f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_633 N_A_549_47#_c_605_n N_X_c_1243_n 0.00198252f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_634 N_A_549_47#_M1041_g N_X_c_1369_n 5.23702e-19 $X=9.81 $Y=0.56 $X2=0 $Y2=0
cc_635 N_A_549_47#_M1042_g N_X_c_1369_n 0.00636826f $X=10.23 $Y=0.56 $X2=0 $Y2=0
cc_636 N_A_549_47#_M1043_g N_X_c_1369_n 0.00636826f $X=10.65 $Y=0.56 $X2=0 $Y2=0
cc_637 N_A_549_47#_M1046_g N_X_c_1369_n 5.23702e-19 $X=11.07 $Y=0.56 $X2=0 $Y2=0
cc_638 N_A_549_47#_M1037_g N_X_c_1373_n 7.66249e-19 $X=9.81 $Y=1.985 $X2=0 $Y2=0
cc_639 N_A_549_47#_M1039_g N_X_c_1373_n 0.0106215f $X=10.23 $Y=1.985 $X2=0 $Y2=0
cc_640 N_A_549_47#_M1047_g N_X_c_1373_n 0.0106215f $X=10.65 $Y=1.985 $X2=0 $Y2=0
cc_641 N_A_549_47#_M1048_g N_X_c_1373_n 7.66249e-19 $X=11.07 $Y=1.985 $X2=0
+ $Y2=0
cc_642 N_A_549_47#_M1043_g N_X_c_1227_n 0.00850187f $X=10.65 $Y=0.56 $X2=0 $Y2=0
cc_643 N_A_549_47#_M1046_g N_X_c_1227_n 0.00850187f $X=11.07 $Y=0.56 $X2=0 $Y2=0
cc_644 N_A_549_47#_c_601_n N_X_c_1227_n 0.0359512f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_645 N_A_549_47#_c_605_n N_X_c_1227_n 0.00205431f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_646 N_A_549_47#_M1047_g N_X_c_1244_n 0.0107189f $X=10.65 $Y=1.985 $X2=0 $Y2=0
cc_647 N_A_549_47#_M1048_g N_X_c_1244_n 0.0107189f $X=11.07 $Y=1.985 $X2=0 $Y2=0
cc_648 N_A_549_47#_c_601_n N_X_c_1244_n 0.0359514f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_649 N_A_549_47#_c_605_n N_X_c_1244_n 0.00198252f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_650 N_A_549_47#_M1043_g N_X_c_1385_n 5.23702e-19 $X=10.65 $Y=0.56 $X2=0 $Y2=0
cc_651 N_A_549_47#_M1046_g N_X_c_1385_n 0.00636826f $X=11.07 $Y=0.56 $X2=0 $Y2=0
cc_652 N_A_549_47#_M1051_g N_X_c_1385_n 0.0109928f $X=11.49 $Y=0.56 $X2=0 $Y2=0
cc_653 N_A_549_47#_M1047_g N_X_c_1388_n 7.66249e-19 $X=10.65 $Y=1.985 $X2=0
+ $Y2=0
cc_654 N_A_549_47#_M1048_g N_X_c_1388_n 0.0106215f $X=11.07 $Y=1.985 $X2=0 $Y2=0
cc_655 N_A_549_47#_M1050_g N_X_c_1388_n 0.0167471f $X=11.49 $Y=1.985 $X2=0 $Y2=0
cc_656 N_A_549_47#_M1051_g N_X_c_1228_n 0.011222f $X=11.49 $Y=0.56 $X2=0 $Y2=0
cc_657 N_A_549_47#_c_601_n N_X_c_1228_n 3.09302e-19 $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_658 N_A_549_47#_M1050_g N_X_c_1245_n 0.013439f $X=11.49 $Y=1.985 $X2=0 $Y2=0
cc_659 N_A_549_47#_c_601_n N_X_c_1245_n 3.09302e-19 $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_660 N_A_549_47#_M1017_g N_X_c_1229_n 0.00111988f $X=6.03 $Y=0.56 $X2=0 $Y2=0
cc_661 N_A_549_47#_M1018_g N_X_c_1229_n 0.00111988f $X=6.45 $Y=0.56 $X2=0 $Y2=0
cc_662 N_A_549_47#_c_601_n N_X_c_1229_n 0.0265319f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_663 N_A_549_47#_c_605_n N_X_c_1229_n 0.00213429f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_664 N_A_549_47#_M1004_g N_X_c_1246_n 0.00135419f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_665 N_A_549_47#_M1005_g N_X_c_1246_n 0.00135419f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_666 N_A_549_47#_c_601_n N_X_c_1246_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_667 N_A_549_47#_c_605_n N_X_c_1246_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_668 N_A_549_47#_M1026_g N_X_c_1230_n 0.00111988f $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_669 N_A_549_47#_M1027_g N_X_c_1230_n 0.00111988f $X=7.29 $Y=0.56 $X2=0 $Y2=0
cc_670 N_A_549_47#_c_601_n N_X_c_1230_n 0.0265319f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_671 N_A_549_47#_c_605_n N_X_c_1230_n 0.00213429f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_672 N_A_549_47#_M1008_g N_X_c_1247_n 0.00135419f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_673 N_A_549_47#_M1015_g N_X_c_1247_n 0.00135419f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_674 N_A_549_47#_c_601_n N_X_c_1247_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_675 N_A_549_47#_c_605_n N_X_c_1247_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_676 N_A_549_47#_M1028_g N_X_c_1231_n 0.00110541f $X=7.71 $Y=0.56 $X2=0 $Y2=0
cc_677 N_A_549_47#_M1029_g N_X_c_1231_n 0.00110541f $X=8.13 $Y=0.56 $X2=0 $Y2=0
cc_678 N_A_549_47#_c_601_n N_X_c_1231_n 0.0265235f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_679 N_A_549_47#_c_605_n N_X_c_1231_n 0.00213376f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_680 N_A_549_47#_M1016_g N_X_c_1248_n 0.00135419f $X=7.71 $Y=1.985 $X2=0 $Y2=0
cc_681 N_A_549_47#_M1022_g N_X_c_1248_n 0.00135419f $X=8.13 $Y=1.985 $X2=0 $Y2=0
cc_682 N_A_549_47#_c_601_n N_X_c_1248_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_683 N_A_549_47#_c_605_n N_X_c_1248_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_684 N_A_549_47#_M1035_g N_X_c_1232_n 0.00110541f $X=8.55 $Y=0.56 $X2=0 $Y2=0
cc_685 N_A_549_47#_M1038_g N_X_c_1232_n 0.00110541f $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_686 N_A_549_47#_c_601_n N_X_c_1232_n 0.0265235f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_687 N_A_549_47#_c_605_n N_X_c_1232_n 0.00213376f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_688 N_A_549_47#_M1030_g N_X_c_1249_n 0.00135419f $X=8.55 $Y=1.985 $X2=0 $Y2=0
cc_689 N_A_549_47#_M1031_g N_X_c_1249_n 0.00135419f $X=8.97 $Y=1.985 $X2=0 $Y2=0
cc_690 N_A_549_47#_c_601_n N_X_c_1249_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_691 N_A_549_47#_c_605_n N_X_c_1249_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_692 N_A_549_47#_M1040_g N_X_c_1233_n 0.00110541f $X=9.39 $Y=0.56 $X2=0 $Y2=0
cc_693 N_A_549_47#_M1041_g N_X_c_1233_n 0.00110541f $X=9.81 $Y=0.56 $X2=0 $Y2=0
cc_694 N_A_549_47#_c_601_n N_X_c_1233_n 0.0265235f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_695 N_A_549_47#_c_605_n N_X_c_1233_n 0.00213376f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_696 N_A_549_47#_M1036_g N_X_c_1250_n 0.00135419f $X=9.39 $Y=1.985 $X2=0 $Y2=0
cc_697 N_A_549_47#_M1037_g N_X_c_1250_n 0.00135419f $X=9.81 $Y=1.985 $X2=0 $Y2=0
cc_698 N_A_549_47#_c_601_n N_X_c_1250_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_699 N_A_549_47#_c_605_n N_X_c_1250_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_700 N_A_549_47#_M1042_g N_X_c_1234_n 0.00110541f $X=10.23 $Y=0.56 $X2=0 $Y2=0
cc_701 N_A_549_47#_M1043_g N_X_c_1234_n 0.00110541f $X=10.65 $Y=0.56 $X2=0 $Y2=0
cc_702 N_A_549_47#_c_601_n N_X_c_1234_n 0.0265235f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_703 N_A_549_47#_c_605_n N_X_c_1234_n 0.00213376f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_704 N_A_549_47#_M1039_g N_X_c_1251_n 0.00135419f $X=10.23 $Y=1.985 $X2=0
+ $Y2=0
cc_705 N_A_549_47#_M1047_g N_X_c_1251_n 0.00135419f $X=10.65 $Y=1.985 $X2=0
+ $Y2=0
cc_706 N_A_549_47#_c_601_n N_X_c_1251_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_707 N_A_549_47#_c_605_n N_X_c_1251_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_708 N_A_549_47#_M1046_g N_X_c_1235_n 0.00110541f $X=11.07 $Y=0.56 $X2=0 $Y2=0
cc_709 N_A_549_47#_M1051_g N_X_c_1235_n 0.00110541f $X=11.49 $Y=0.56 $X2=0 $Y2=0
cc_710 N_A_549_47#_c_601_n N_X_c_1235_n 0.0265235f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_711 N_A_549_47#_c_605_n N_X_c_1235_n 0.00213376f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_712 N_A_549_47#_M1048_g N_X_c_1252_n 0.00135419f $X=11.07 $Y=1.985 $X2=0
+ $Y2=0
cc_713 N_A_549_47#_M1050_g N_X_c_1252_n 0.00135419f $X=11.49 $Y=1.985 $X2=0
+ $Y2=0
cc_714 N_A_549_47#_c_601_n N_X_c_1252_n 0.026643f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_715 N_A_549_47#_c_605_n N_X_c_1252_n 0.00206439f $X=11.49 $Y=1.16 $X2=0 $Y2=0
cc_716 N_A_549_47#_M1051_g X 0.0204688f $X=11.49 $Y=0.56 $X2=0 $Y2=0
cc_717 N_A_549_47#_c_601_n X 0.0162963f $X=11.08 $Y=1.16 $X2=0 $Y2=0
cc_718 N_A_549_47#_c_596_n N_VGND_M1012_d 0.00162006f $X=3.555 $Y=0.82 $X2=0
+ $Y2=0
cc_719 N_A_549_47#_c_598_n N_VGND_M1021_d 0.00162006f $X=4.395 $Y=0.82 $X2=0
+ $Y2=0
cc_720 N_A_549_47#_c_603_n N_VGND_M1033_d 0.00186748f $X=4.977 $Y=0.82 $X2=0
+ $Y2=0
cc_721 N_A_549_47#_c_596_n N_VGND_c_1561_n 0.0122414f $X=3.555 $Y=0.82 $X2=0
+ $Y2=0
cc_722 N_A_549_47#_c_598_n N_VGND_c_1562_n 0.0122414f $X=4.395 $Y=0.82 $X2=0
+ $Y2=0
cc_723 N_A_549_47#_M1000_g N_VGND_c_1563_n 0.00146448f $X=5.19 $Y=0.56 $X2=0
+ $Y2=0
cc_724 N_A_549_47#_c_603_n N_VGND_c_1563_n 0.0122414f $X=4.977 $Y=0.82 $X2=0
+ $Y2=0
cc_725 N_A_549_47#_M1000_g N_VGND_c_1564_n 0.00539841f $X=5.19 $Y=0.56 $X2=0
+ $Y2=0
cc_726 N_A_549_47#_M1009_g N_VGND_c_1564_n 0.00423108f $X=5.61 $Y=0.56 $X2=0
+ $Y2=0
cc_727 N_A_549_47#_M1009_g N_VGND_c_1565_n 0.00146448f $X=5.61 $Y=0.56 $X2=0
+ $Y2=0
cc_728 N_A_549_47#_M1017_g N_VGND_c_1565_n 0.00146448f $X=6.03 $Y=0.56 $X2=0
+ $Y2=0
cc_729 N_A_549_47#_M1018_g N_VGND_c_1566_n 0.00146448f $X=6.45 $Y=0.56 $X2=0
+ $Y2=0
cc_730 N_A_549_47#_M1026_g N_VGND_c_1566_n 0.00146448f $X=6.87 $Y=0.56 $X2=0
+ $Y2=0
cc_731 N_A_549_47#_M1027_g N_VGND_c_1567_n 0.00146448f $X=7.29 $Y=0.56 $X2=0
+ $Y2=0
cc_732 N_A_549_47#_M1028_g N_VGND_c_1567_n 0.00146448f $X=7.71 $Y=0.56 $X2=0
+ $Y2=0
cc_733 N_A_549_47#_M1029_g N_VGND_c_1568_n 0.00146448f $X=8.13 $Y=0.56 $X2=0
+ $Y2=0
cc_734 N_A_549_47#_M1035_g N_VGND_c_1568_n 0.00146448f $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_735 N_A_549_47#_M1038_g N_VGND_c_1569_n 0.00146448f $X=8.97 $Y=0.56 $X2=0
+ $Y2=0
cc_736 N_A_549_47#_M1040_g N_VGND_c_1569_n 0.00146448f $X=9.39 $Y=0.56 $X2=0
+ $Y2=0
cc_737 N_A_549_47#_M1041_g N_VGND_c_1570_n 0.00146448f $X=9.81 $Y=0.56 $X2=0
+ $Y2=0
cc_738 N_A_549_47#_M1042_g N_VGND_c_1570_n 0.00146448f $X=10.23 $Y=0.56 $X2=0
+ $Y2=0
cc_739 N_A_549_47#_M1042_g N_VGND_c_1571_n 0.00424619f $X=10.23 $Y=0.56 $X2=0
+ $Y2=0
cc_740 N_A_549_47#_M1043_g N_VGND_c_1571_n 0.00424619f $X=10.65 $Y=0.56 $X2=0
+ $Y2=0
cc_741 N_A_549_47#_M1043_g N_VGND_c_1572_n 0.00146448f $X=10.65 $Y=0.56 $X2=0
+ $Y2=0
cc_742 N_A_549_47#_M1046_g N_VGND_c_1572_n 0.00146448f $X=11.07 $Y=0.56 $X2=0
+ $Y2=0
cc_743 N_A_549_47#_M1051_g N_VGND_c_1574_n 0.00316354f $X=11.49 $Y=0.56 $X2=0
+ $Y2=0
cc_744 N_A_549_47#_c_628_n N_VGND_c_1577_n 0.0182681f $X=2.88 $Y=0.4 $X2=0 $Y2=0
cc_745 N_A_549_47#_c_596_n N_VGND_c_1577_n 0.00193763f $X=3.555 $Y=0.82 $X2=0
+ $Y2=0
cc_746 N_A_549_47#_c_596_n N_VGND_c_1579_n 0.00193763f $X=3.555 $Y=0.82 $X2=0
+ $Y2=0
cc_747 N_A_549_47#_c_658_n N_VGND_c_1579_n 0.0182681f $X=3.72 $Y=0.4 $X2=0 $Y2=0
cc_748 N_A_549_47#_c_598_n N_VGND_c_1579_n 0.00193763f $X=4.395 $Y=0.82 $X2=0
+ $Y2=0
cc_749 N_A_549_47#_c_598_n N_VGND_c_1581_n 0.00390702f $X=4.395 $Y=0.82 $X2=0
+ $Y2=0
cc_750 N_A_549_47#_c_674_n N_VGND_c_1581_n 0.0179571f $X=4.56 $Y=0.4 $X2=0 $Y2=0
cc_751 N_A_549_47#_M1017_g N_VGND_c_1583_n 0.00423108f $X=6.03 $Y=0.56 $X2=0
+ $Y2=0
cc_752 N_A_549_47#_M1018_g N_VGND_c_1583_n 0.00423108f $X=6.45 $Y=0.56 $X2=0
+ $Y2=0
cc_753 N_A_549_47#_M1026_g N_VGND_c_1585_n 0.00423108f $X=6.87 $Y=0.56 $X2=0
+ $Y2=0
cc_754 N_A_549_47#_M1027_g N_VGND_c_1585_n 0.00423108f $X=7.29 $Y=0.56 $X2=0
+ $Y2=0
cc_755 N_A_549_47#_M1028_g N_VGND_c_1587_n 0.00424619f $X=7.71 $Y=0.56 $X2=0
+ $Y2=0
cc_756 N_A_549_47#_M1029_g N_VGND_c_1587_n 0.00424619f $X=8.13 $Y=0.56 $X2=0
+ $Y2=0
cc_757 N_A_549_47#_M1035_g N_VGND_c_1589_n 0.00424619f $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_758 N_A_549_47#_M1038_g N_VGND_c_1589_n 0.00424619f $X=8.97 $Y=0.56 $X2=0
+ $Y2=0
cc_759 N_A_549_47#_M1040_g N_VGND_c_1591_n 0.00424619f $X=9.39 $Y=0.56 $X2=0
+ $Y2=0
cc_760 N_A_549_47#_M1041_g N_VGND_c_1591_n 0.00424619f $X=9.81 $Y=0.56 $X2=0
+ $Y2=0
cc_761 N_A_549_47#_M1046_g N_VGND_c_1594_n 0.00424619f $X=11.07 $Y=0.56 $X2=0
+ $Y2=0
cc_762 N_A_549_47#_M1051_g N_VGND_c_1594_n 0.00424619f $X=11.49 $Y=0.56 $X2=0
+ $Y2=0
cc_763 N_A_549_47#_M1010_s N_VGND_c_1598_n 0.00215347f $X=2.745 $Y=0.235 $X2=0
+ $Y2=0
cc_764 N_A_549_47#_M1020_s N_VGND_c_1598_n 0.00215347f $X=3.585 $Y=0.235 $X2=0
+ $Y2=0
cc_765 N_A_549_47#_M1023_s N_VGND_c_1598_n 0.00215347f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_766 N_A_549_47#_M1000_g N_VGND_c_1598_n 0.00949176f $X=5.19 $Y=0.56 $X2=0
+ $Y2=0
cc_767 N_A_549_47#_M1009_g N_VGND_c_1598_n 0.00574532f $X=5.61 $Y=0.56 $X2=0
+ $Y2=0
cc_768 N_A_549_47#_M1017_g N_VGND_c_1598_n 0.00574532f $X=6.03 $Y=0.56 $X2=0
+ $Y2=0
cc_769 N_A_549_47#_M1018_g N_VGND_c_1598_n 0.00574532f $X=6.45 $Y=0.56 $X2=0
+ $Y2=0
cc_770 N_A_549_47#_M1026_g N_VGND_c_1598_n 0.00574532f $X=6.87 $Y=0.56 $X2=0
+ $Y2=0
cc_771 N_A_549_47#_M1027_g N_VGND_c_1598_n 0.00574532f $X=7.29 $Y=0.56 $X2=0
+ $Y2=0
cc_772 N_A_549_47#_M1028_g N_VGND_c_1598_n 0.00573624f $X=7.71 $Y=0.56 $X2=0
+ $Y2=0
cc_773 N_A_549_47#_M1029_g N_VGND_c_1598_n 0.00573624f $X=8.13 $Y=0.56 $X2=0
+ $Y2=0
cc_774 N_A_549_47#_M1035_g N_VGND_c_1598_n 0.00573624f $X=8.55 $Y=0.56 $X2=0
+ $Y2=0
cc_775 N_A_549_47#_M1038_g N_VGND_c_1598_n 0.00573624f $X=8.97 $Y=0.56 $X2=0
+ $Y2=0
cc_776 N_A_549_47#_M1040_g N_VGND_c_1598_n 0.00573624f $X=9.39 $Y=0.56 $X2=0
+ $Y2=0
cc_777 N_A_549_47#_M1041_g N_VGND_c_1598_n 0.00573624f $X=9.81 $Y=0.56 $X2=0
+ $Y2=0
cc_778 N_A_549_47#_M1042_g N_VGND_c_1598_n 0.00573624f $X=10.23 $Y=0.56 $X2=0
+ $Y2=0
cc_779 N_A_549_47#_M1043_g N_VGND_c_1598_n 0.00573624f $X=10.65 $Y=0.56 $X2=0
+ $Y2=0
cc_780 N_A_549_47#_M1046_g N_VGND_c_1598_n 0.00573624f $X=11.07 $Y=0.56 $X2=0
+ $Y2=0
cc_781 N_A_549_47#_M1051_g N_VGND_c_1598_n 0.00669045f $X=11.49 $Y=0.56 $X2=0
+ $Y2=0
cc_782 N_A_549_47#_c_628_n N_VGND_c_1598_n 0.0121741f $X=2.88 $Y=0.4 $X2=0 $Y2=0
cc_783 N_A_549_47#_c_596_n N_VGND_c_1598_n 0.00825759f $X=3.555 $Y=0.82 $X2=0
+ $Y2=0
cc_784 N_A_549_47#_c_658_n N_VGND_c_1598_n 0.0121741f $X=3.72 $Y=0.4 $X2=0 $Y2=0
cc_785 N_A_549_47#_c_598_n N_VGND_c_1598_n 0.012122f $X=4.395 $Y=0.82 $X2=0
+ $Y2=0
cc_786 N_A_549_47#_c_674_n N_VGND_c_1598_n 0.0120759f $X=4.56 $Y=0.4 $X2=0 $Y2=0
cc_787 N_A_549_47#_c_603_n N_VGND_c_1598_n 6.28727e-19 $X=4.977 $Y=0.82 $X2=0
+ $Y2=0
cc_788 N_VPWR_c_1028_n N_X_M1001_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_789 N_VPWR_c_1028_n N_X_M1004_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_790 N_VPWR_c_1028_n N_X_M1008_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_791 N_VPWR_c_1028_n N_X_M1016_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_792 N_VPWR_c_1028_n N_X_M1030_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_793 N_VPWR_c_1028_n N_X_M1036_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_794 N_VPWR_c_1028_n N_X_M1039_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_795 N_VPWR_c_1028_n N_X_M1048_d 0.00215201f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_796 N_VPWR_c_1036_n N_X_c_1256_n 0.0189039f $X=5.735 $Y=2.72 $X2=0 $Y2=0
cc_797 N_VPWR_c_1028_n N_X_c_1256_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_798 N_VPWR_M1002_s N_X_c_1237_n 0.00185611f $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_799 N_VPWR_c_1037_n N_X_c_1237_n 0.0104788f $X=5.82 $Y=2 $X2=0 $Y2=0
cc_800 N_VPWR_c_1055_n N_X_c_1291_n 0.0189039f $X=6.575 $Y=2.72 $X2=0 $Y2=0
cc_801 N_VPWR_c_1028_n N_X_c_1291_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_802 N_VPWR_M1005_s N_X_c_1239_n 0.00185611f $X=6.525 $Y=1.485 $X2=0 $Y2=0
cc_803 N_VPWR_c_1038_n N_X_c_1239_n 0.0104788f $X=6.66 $Y=2 $X2=0 $Y2=0
cc_804 N_VPWR_c_1057_n N_X_c_1309_n 0.0189039f $X=7.415 $Y=2.72 $X2=0 $Y2=0
cc_805 N_VPWR_c_1028_n N_X_c_1309_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_806 N_VPWR_M1015_s N_X_c_1240_n 0.00185611f $X=7.365 $Y=1.485 $X2=0 $Y2=0
cc_807 N_VPWR_c_1039_n N_X_c_1240_n 0.0104788f $X=7.5 $Y=2 $X2=0 $Y2=0
cc_808 N_VPWR_c_1059_n N_X_c_1325_n 0.0189039f $X=8.255 $Y=2.72 $X2=0 $Y2=0
cc_809 N_VPWR_c_1028_n N_X_c_1325_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_810 N_VPWR_M1022_s N_X_c_1241_n 0.00185611f $X=8.205 $Y=1.485 $X2=0 $Y2=0
cc_811 N_VPWR_c_1040_n N_X_c_1241_n 0.0104788f $X=8.34 $Y=2 $X2=0 $Y2=0
cc_812 N_VPWR_c_1061_n N_X_c_1341_n 0.0189039f $X=9.095 $Y=2.72 $X2=0 $Y2=0
cc_813 N_VPWR_c_1028_n N_X_c_1341_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_814 N_VPWR_M1031_s N_X_c_1242_n 0.00185611f $X=9.045 $Y=1.485 $X2=0 $Y2=0
cc_815 N_VPWR_c_1041_n N_X_c_1242_n 0.0104788f $X=9.18 $Y=2 $X2=0 $Y2=0
cc_816 N_VPWR_c_1063_n N_X_c_1357_n 0.0189039f $X=9.935 $Y=2.72 $X2=0 $Y2=0
cc_817 N_VPWR_c_1028_n N_X_c_1357_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_818 N_VPWR_M1037_s N_X_c_1243_n 0.00185611f $X=9.885 $Y=1.485 $X2=0 $Y2=0
cc_819 N_VPWR_c_1042_n N_X_c_1243_n 0.0104788f $X=10.02 $Y=2 $X2=0 $Y2=0
cc_820 N_VPWR_c_1043_n N_X_c_1373_n 0.0189039f $X=10.775 $Y=2.72 $X2=0 $Y2=0
cc_821 N_VPWR_c_1028_n N_X_c_1373_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_822 N_VPWR_M1047_s N_X_c_1244_n 0.00185611f $X=10.725 $Y=1.485 $X2=0 $Y2=0
cc_823 N_VPWR_c_1044_n N_X_c_1244_n 0.0104788f $X=10.86 $Y=2 $X2=0 $Y2=0
cc_824 N_VPWR_c_1066_n N_X_c_1388_n 0.0189039f $X=11.615 $Y=2.72 $X2=0 $Y2=0
cc_825 N_VPWR_c_1028_n N_X_c_1388_n 0.0122217f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_826 N_VPWR_M1050_s X 0.00443391f $X=11.565 $Y=1.485 $X2=0 $Y2=0
cc_827 N_VPWR_c_1046_n X 0.0120465f $X=11.7 $Y=2 $X2=0 $Y2=0
cc_828 N_X_c_1220_n N_VGND_M1009_d 0.00162006f $X=6.075 $Y=0.82 $X2=0 $Y2=0
cc_829 N_X_c_1222_n N_VGND_M1018_d 0.00162006f $X=6.915 $Y=0.82 $X2=0 $Y2=0
cc_830 N_X_c_1223_n N_VGND_M1027_d 0.00162006f $X=7.755 $Y=0.82 $X2=0 $Y2=0
cc_831 N_X_c_1224_n N_VGND_M1029_d 0.00162006f $X=8.595 $Y=0.82 $X2=0 $Y2=0
cc_832 N_X_c_1225_n N_VGND_M1038_d 0.00162006f $X=9.435 $Y=0.82 $X2=0 $Y2=0
cc_833 N_X_c_1226_n N_VGND_M1041_d 0.00162006f $X=10.275 $Y=0.82 $X2=0 $Y2=0
cc_834 N_X_c_1227_n N_VGND_M1043_d 0.00162006f $X=11.115 $Y=0.82 $X2=0 $Y2=0
cc_835 N_X_c_1228_n N_VGND_M1051_d 0.00322906f $X=11.62 $Y=0.82 $X2=0 $Y2=0
cc_836 N_X_c_1257_n N_VGND_c_1564_n 0.0188753f $X=5.4 $Y=0.425 $X2=0 $Y2=0
cc_837 N_X_c_1220_n N_VGND_c_1564_n 0.00193763f $X=6.075 $Y=0.82 $X2=0 $Y2=0
cc_838 N_X_c_1220_n N_VGND_c_1565_n 0.0122414f $X=6.075 $Y=0.82 $X2=0 $Y2=0
cc_839 N_X_c_1222_n N_VGND_c_1566_n 0.0122414f $X=6.915 $Y=0.82 $X2=0 $Y2=0
cc_840 N_X_c_1223_n N_VGND_c_1567_n 0.0122414f $X=7.755 $Y=0.82 $X2=0 $Y2=0
cc_841 N_X_c_1224_n N_VGND_c_1568_n 0.0122414f $X=8.595 $Y=0.82 $X2=0 $Y2=0
cc_842 N_X_c_1225_n N_VGND_c_1569_n 0.0122414f $X=9.435 $Y=0.82 $X2=0 $Y2=0
cc_843 N_X_c_1226_n N_VGND_c_1570_n 0.0122414f $X=10.275 $Y=0.82 $X2=0 $Y2=0
cc_844 N_X_c_1226_n N_VGND_c_1571_n 0.00193763f $X=10.275 $Y=0.82 $X2=0 $Y2=0
cc_845 N_X_c_1369_n N_VGND_c_1571_n 0.0182681f $X=10.44 $Y=0.4 $X2=0 $Y2=0
cc_846 N_X_c_1227_n N_VGND_c_1571_n 0.00193763f $X=11.115 $Y=0.82 $X2=0 $Y2=0
cc_847 N_X_c_1227_n N_VGND_c_1572_n 0.0122414f $X=11.115 $Y=0.82 $X2=0 $Y2=0
cc_848 N_X_c_1228_n N_VGND_c_1573_n 0.00146941f $X=11.62 $Y=0.82 $X2=0 $Y2=0
cc_849 N_X_c_1228_n N_VGND_c_1574_n 0.0140453f $X=11.62 $Y=0.82 $X2=0 $Y2=0
cc_850 N_X_c_1220_n N_VGND_c_1583_n 0.00193763f $X=6.075 $Y=0.82 $X2=0 $Y2=0
cc_851 N_X_c_1285_n N_VGND_c_1583_n 0.0187595f $X=6.24 $Y=0.425 $X2=0 $Y2=0
cc_852 N_X_c_1222_n N_VGND_c_1583_n 0.00193763f $X=6.915 $Y=0.82 $X2=0 $Y2=0
cc_853 N_X_c_1222_n N_VGND_c_1585_n 0.00193763f $X=6.915 $Y=0.82 $X2=0 $Y2=0
cc_854 N_X_c_1303_n N_VGND_c_1585_n 0.0187595f $X=7.08 $Y=0.425 $X2=0 $Y2=0
cc_855 N_X_c_1223_n N_VGND_c_1585_n 0.00193763f $X=7.755 $Y=0.82 $X2=0 $Y2=0
cc_856 N_X_c_1223_n N_VGND_c_1587_n 0.00193763f $X=7.755 $Y=0.82 $X2=0 $Y2=0
cc_857 N_X_c_1321_n N_VGND_c_1587_n 0.0182681f $X=7.92 $Y=0.4 $X2=0 $Y2=0
cc_858 N_X_c_1224_n N_VGND_c_1587_n 0.00193763f $X=8.595 $Y=0.82 $X2=0 $Y2=0
cc_859 N_X_c_1224_n N_VGND_c_1589_n 0.00193763f $X=8.595 $Y=0.82 $X2=0 $Y2=0
cc_860 N_X_c_1337_n N_VGND_c_1589_n 0.0182681f $X=8.76 $Y=0.4 $X2=0 $Y2=0
cc_861 N_X_c_1225_n N_VGND_c_1589_n 0.00193763f $X=9.435 $Y=0.82 $X2=0 $Y2=0
cc_862 N_X_c_1225_n N_VGND_c_1591_n 0.00193763f $X=9.435 $Y=0.82 $X2=0 $Y2=0
cc_863 N_X_c_1353_n N_VGND_c_1591_n 0.0182681f $X=9.6 $Y=0.4 $X2=0 $Y2=0
cc_864 N_X_c_1226_n N_VGND_c_1591_n 0.00193763f $X=10.275 $Y=0.82 $X2=0 $Y2=0
cc_865 N_X_c_1227_n N_VGND_c_1594_n 0.00193763f $X=11.115 $Y=0.82 $X2=0 $Y2=0
cc_866 N_X_c_1385_n N_VGND_c_1594_n 0.0182681f $X=11.28 $Y=0.4 $X2=0 $Y2=0
cc_867 N_X_c_1228_n N_VGND_c_1594_n 0.00193763f $X=11.62 $Y=0.82 $X2=0 $Y2=0
cc_868 N_X_M1000_s N_VGND_c_1598_n 0.00215228f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_869 N_X_M1017_s N_VGND_c_1598_n 0.00215254f $X=6.105 $Y=0.235 $X2=0 $Y2=0
cc_870 N_X_M1026_s N_VGND_c_1598_n 0.00215254f $X=6.945 $Y=0.235 $X2=0 $Y2=0
cc_871 N_X_M1028_s N_VGND_c_1598_n 0.00215347f $X=7.785 $Y=0.235 $X2=0 $Y2=0
cc_872 N_X_M1035_s N_VGND_c_1598_n 0.00215347f $X=8.625 $Y=0.235 $X2=0 $Y2=0
cc_873 N_X_M1040_s N_VGND_c_1598_n 0.00215347f $X=9.465 $Y=0.235 $X2=0 $Y2=0
cc_874 N_X_M1042_s N_VGND_c_1598_n 0.00215347f $X=10.305 $Y=0.235 $X2=0 $Y2=0
cc_875 N_X_M1046_s N_VGND_c_1598_n 0.00215347f $X=11.145 $Y=0.235 $X2=0 $Y2=0
cc_876 N_X_c_1257_n N_VGND_c_1598_n 0.0122666f $X=5.4 $Y=0.425 $X2=0 $Y2=0
cc_877 N_X_c_1220_n N_VGND_c_1598_n 0.00825759f $X=6.075 $Y=0.82 $X2=0 $Y2=0
cc_878 N_X_c_1285_n N_VGND_c_1598_n 0.0122584f $X=6.24 $Y=0.425 $X2=0 $Y2=0
cc_879 N_X_c_1222_n N_VGND_c_1598_n 0.00825759f $X=6.915 $Y=0.82 $X2=0 $Y2=0
cc_880 N_X_c_1303_n N_VGND_c_1598_n 0.0122584f $X=7.08 $Y=0.425 $X2=0 $Y2=0
cc_881 N_X_c_1223_n N_VGND_c_1598_n 0.00825759f $X=7.755 $Y=0.82 $X2=0 $Y2=0
cc_882 N_X_c_1321_n N_VGND_c_1598_n 0.0121741f $X=7.92 $Y=0.4 $X2=0 $Y2=0
cc_883 N_X_c_1224_n N_VGND_c_1598_n 0.00825759f $X=8.595 $Y=0.82 $X2=0 $Y2=0
cc_884 N_X_c_1337_n N_VGND_c_1598_n 0.0121741f $X=8.76 $Y=0.4 $X2=0 $Y2=0
cc_885 N_X_c_1225_n N_VGND_c_1598_n 0.00825759f $X=9.435 $Y=0.82 $X2=0 $Y2=0
cc_886 N_X_c_1353_n N_VGND_c_1598_n 0.0121741f $X=9.6 $Y=0.4 $X2=0 $Y2=0
cc_887 N_X_c_1226_n N_VGND_c_1598_n 0.00825759f $X=10.275 $Y=0.82 $X2=0 $Y2=0
cc_888 N_X_c_1369_n N_VGND_c_1598_n 0.0121741f $X=10.44 $Y=0.4 $X2=0 $Y2=0
cc_889 N_X_c_1227_n N_VGND_c_1598_n 0.00825759f $X=11.115 $Y=0.82 $X2=0 $Y2=0
cc_890 N_X_c_1385_n N_VGND_c_1598_n 0.0121741f $X=11.28 $Y=0.4 $X2=0 $Y2=0
cc_891 N_X_c_1228_n N_VGND_c_1598_n 0.00706467f $X=11.62 $Y=0.82 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o221ai_1.spice
* Created: Tue Sep  1 19:22:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o221ai_1.pex.spice"
.subckt sky130_fd_sc_hd__o221ai_1  VNB VPB C1 B1 B2 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1008 N_A_109_47#_M1008_d N_C1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1654 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_109_47#_M1006_d N_B1_M1006_g N_A_213_123#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.1652 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1000 N_A_213_123#_M1000_d N_B2_M1000_g N_A_109_47#_M1006_d VNB NSHORT L=0.15
+ W=0.65 AD=0.117 AS=0.08775 PD=1.01 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_213_123#_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.117 PD=0.92 PS=1.01 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_213_123#_M1004_d N_A1_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_C1_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.38
+ AS=0.28 PD=1.76 PS=2.56 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002.4
+ A=0.15 P=2.3 MULT=1
MM1003 A_295_297# N_B1_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1 AD=0.12
+ AS=0.38 PD=1.24 PS=1.76 NRD=12.7853 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g A_295_297# VPB PHIGHVT L=0.15 W=1 AD=0.225
+ AS=0.12 PD=1.45 PS=1.24 NRD=0 NRS=12.7853 M=1 R=6.66667 SA=75001.5 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1007 A_493_297# N_A2_M1007_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.225 PD=1.21 PS=1.45 NRD=9.8303 NRS=34.4553 M=1 R=6.66667 SA=75002.1
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_493_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__o221ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdfxtp_1.spice.SKY130_FD_SC_HD__SDFXTP_1.pxi
* Created: Thu Aug 27 14:47:17 2020
* 
x_PM_SKY130_FD_SC_HD__SDFXTP_1%CLK N_CLK_c_216_n N_CLK_c_220_n N_CLK_c_217_n
+ N_CLK_M1029_g N_CLK_c_221_n N_CLK_M1005_g N_CLK_c_222_n CLK
+ PM_SKY130_FD_SC_HD__SDFXTP_1%CLK
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_27_47# N_A_27_47#_M1029_s N_A_27_47#_M1005_s
+ N_A_27_47#_M1015_g N_A_27_47#_M1028_g N_A_27_47#_M1030_g N_A_27_47#_c_260_n
+ N_A_27_47#_c_261_n N_A_27_47#_M1006_g N_A_27_47#_M1026_g N_A_27_47#_c_262_n
+ N_A_27_47#_M1003_g N_A_27_47#_c_496_p N_A_27_47#_c_264_n N_A_27_47#_c_265_n
+ N_A_27_47#_c_277_n N_A_27_47#_c_266_n N_A_27_47#_c_386_p N_A_27_47#_c_278_n
+ N_A_27_47#_c_279_n N_A_27_47#_c_267_n N_A_27_47#_c_280_n N_A_27_47#_c_281_n
+ N_A_27_47#_c_282_n N_A_27_47#_c_283_n N_A_27_47#_c_284_n N_A_27_47#_c_285_n
+ N_A_27_47#_c_268_n N_A_27_47#_c_287_n N_A_27_47#_c_288_n N_A_27_47#_c_269_n
+ N_A_27_47#_c_270_n PM_SKY130_FD_SC_HD__SDFXTP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%SCE N_SCE_M1018_g N_SCE_M1031_g N_SCE_c_517_n
+ N_SCE_M1010_g N_SCE_M1025_g N_SCE_c_505_n N_SCE_c_506_n N_SCE_c_507_n
+ N_SCE_c_520_n N_SCE_c_508_n N_SCE_c_509_n N_SCE_c_510_n N_SCE_c_511_n
+ N_SCE_c_512_n N_SCE_c_513_n SCE N_SCE_c_514_n N_SCE_c_515_n
+ PM_SKY130_FD_SC_HD__SDFXTP_1%SCE
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_299_47# N_A_299_47#_M1031_s N_A_299_47#_M1018_s
+ N_A_299_47#_M1013_g N_A_299_47#_M1012_g N_A_299_47#_c_630_n
+ N_A_299_47#_c_639_n N_A_299_47#_c_647_n N_A_299_47#_c_631_n
+ N_A_299_47#_c_649_n N_A_299_47#_c_641_n N_A_299_47#_c_632_n
+ N_A_299_47#_c_642_n N_A_299_47#_c_633_n N_A_299_47#_c_634_n
+ N_A_299_47#_c_654_n N_A_299_47#_c_635_n N_A_299_47#_c_636_n
+ PM_SKY130_FD_SC_HD__SDFXTP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%D N_D_M1021_g N_D_M1014_g D N_D_c_771_n
+ N_D_c_772_n PM_SKY130_FD_SC_HD__SDFXTP_1%D
x_PM_SKY130_FD_SC_HD__SDFXTP_1%SCD N_SCD_M1011_g N_SCD_M1009_g N_SCD_c_820_n
+ N_SCD_c_823_n N_SCD_c_824_n N_SCD_c_825_n SCD N_SCD_c_822_n
+ PM_SKY130_FD_SC_HD__SDFXTP_1%SCD
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_193_47# N_A_193_47#_M1015_d N_A_193_47#_M1028_d
+ N_A_193_47#_M1023_g N_A_193_47#_M1027_g N_A_193_47#_c_875_n
+ N_A_193_47#_M1002_g N_A_193_47#_M1019_g N_A_193_47#_c_876_n
+ N_A_193_47#_c_893_n N_A_193_47#_c_877_n N_A_193_47#_c_878_n
+ N_A_193_47#_c_879_n N_A_193_47#_c_880_n N_A_193_47#_c_895_n
+ N_A_193_47#_c_896_n N_A_193_47#_c_881_n N_A_193_47#_c_882_n
+ N_A_193_47#_c_883_n N_A_193_47#_c_1017_p N_A_193_47#_c_884_n
+ N_A_193_47#_c_885_n N_A_193_47#_c_886_n N_A_193_47#_c_887_n
+ N_A_193_47#_c_888_n N_A_193_47#_c_889_n PM_SKY130_FD_SC_HD__SDFXTP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_1092_183# N_A_1092_183#_M1016_d
+ N_A_1092_183#_M1008_d N_A_1092_183#_M1022_g N_A_1092_183#_M1007_g
+ N_A_1092_183#_c_1093_n N_A_1092_183#_c_1119_n N_A_1092_183#_c_1139_p
+ N_A_1092_183#_c_1120_n N_A_1092_183#_c_1094_n N_A_1092_183#_c_1095_n
+ N_A_1092_183#_c_1107_n N_A_1092_183#_c_1096_n N_A_1092_183#_c_1097_n
+ PM_SKY130_FD_SC_HD__SDFXTP_1%A_1092_183#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_933_413# N_A_933_413#_M1030_d
+ N_A_933_413#_M1023_d N_A_933_413#_c_1186_n N_A_933_413#_M1008_g
+ N_A_933_413#_c_1187_n N_A_933_413#_M1016_g N_A_933_413#_c_1188_n
+ N_A_933_413#_c_1189_n N_A_933_413#_c_1190_n N_A_933_413#_c_1204_n
+ N_A_933_413#_c_1230_n N_A_933_413#_c_1191_n N_A_933_413#_c_1196_n
+ N_A_933_413#_c_1192_n PM_SKY130_FD_SC_HD__SDFXTP_1%A_933_413#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_1520_315# N_A_1520_315#_M1004_s
+ N_A_1520_315#_M1020_s N_A_1520_315#_M1001_g N_A_1520_315#_M1017_g
+ N_A_1520_315#_M1000_g N_A_1520_315#_M1024_g N_A_1520_315#_c_1305_n
+ N_A_1520_315#_c_1306_n N_A_1520_315#_c_1318_p N_A_1520_315#_c_1297_n
+ N_A_1520_315#_c_1307_n N_A_1520_315#_c_1298_n N_A_1520_315#_c_1299_n
+ N_A_1520_315#_c_1300_n N_A_1520_315#_c_1320_p N_A_1520_315#_c_1325_p
+ N_A_1520_315#_c_1301_n PM_SKY130_FD_SC_HD__SDFXTP_1%A_1520_315#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_1349_413# N_A_1349_413#_M1002_d
+ N_A_1349_413#_M1026_d N_A_1349_413#_c_1382_n N_A_1349_413#_M1004_g
+ N_A_1349_413#_M1020_g N_A_1349_413#_c_1383_n N_A_1349_413#_c_1384_n
+ N_A_1349_413#_c_1394_n N_A_1349_413#_c_1397_n N_A_1349_413#_c_1391_n
+ N_A_1349_413#_c_1385_n N_A_1349_413#_c_1386_n N_A_1349_413#_c_1387_n
+ PM_SKY130_FD_SC_HD__SDFXTP_1%A_1349_413#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%VPWR N_VPWR_M1005_d N_VPWR_M1018_d N_VPWR_M1009_d
+ N_VPWR_M1022_d N_VPWR_M1001_d N_VPWR_M1020_d N_VPWR_c_1471_n N_VPWR_c_1472_n
+ N_VPWR_c_1473_n N_VPWR_c_1474_n N_VPWR_c_1475_n N_VPWR_c_1476_n
+ N_VPWR_c_1477_n N_VPWR_c_1478_n N_VPWR_c_1479_n N_VPWR_c_1480_n
+ N_VPWR_c_1481_n N_VPWR_c_1482_n VPWR N_VPWR_c_1483_n N_VPWR_c_1484_n
+ N_VPWR_c_1485_n N_VPWR_c_1486_n N_VPWR_c_1470_n N_VPWR_c_1488_n
+ N_VPWR_c_1489_n N_VPWR_c_1490_n PM_SKY130_FD_SC_HD__SDFXTP_1%VPWR
x_PM_SKY130_FD_SC_HD__SDFXTP_1%A_556_369# N_A_556_369#_M1014_d
+ N_A_556_369#_M1030_s N_A_556_369#_M1021_d N_A_556_369#_M1023_s
+ N_A_556_369#_c_1637_n N_A_556_369#_c_1647_n N_A_556_369#_c_1660_n
+ N_A_556_369#_c_1628_n N_A_556_369#_c_1633_n N_A_556_369#_c_1634_n
+ N_A_556_369#_c_1629_n N_A_556_369#_c_1630_n N_A_556_369#_c_1631_n
+ N_A_556_369#_c_1632_n N_A_556_369#_c_1636_n
+ PM_SKY130_FD_SC_HD__SDFXTP_1%A_556_369#
x_PM_SKY130_FD_SC_HD__SDFXTP_1%Q N_Q_M1000_d N_Q_M1024_d N_Q_c_1746_n
+ N_Q_c_1744_n Q Q Q N_Q_c_1745_n PM_SKY130_FD_SC_HD__SDFXTP_1%Q
x_PM_SKY130_FD_SC_HD__SDFXTP_1%VGND N_VGND_M1029_d N_VGND_M1031_d N_VGND_M1011_d
+ N_VGND_M1007_d N_VGND_M1017_d N_VGND_M1004_d N_VGND_c_1771_n N_VGND_c_1772_n
+ N_VGND_c_1773_n N_VGND_c_1774_n N_VGND_c_1775_n N_VGND_c_1776_n
+ N_VGND_c_1777_n N_VGND_c_1778_n N_VGND_c_1779_n N_VGND_c_1780_n
+ N_VGND_c_1781_n VGND N_VGND_c_1782_n N_VGND_c_1783_n N_VGND_c_1784_n
+ N_VGND_c_1785_n N_VGND_c_1786_n N_VGND_c_1787_n N_VGND_c_1788_n
+ N_VGND_c_1789_n N_VGND_c_1790_n PM_SKY130_FD_SC_HD__SDFXTP_1%VGND
cc_1 VNB N_CLK_c_216_n 0.0573151f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_217_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0185843f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1015_g 0.0381832f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1030_g 0.0527519f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_6 VNB N_A_27_47#_c_260_n 0.0135588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_261_n 0.00284024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_262_n 0.0158261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1003_g 0.043789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_264_n 0.00318927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_265_n 0.00642096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_266_n 8.11193e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_267_n 0.00238348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_268_n 0.0228343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_269_n 0.00981039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_270_n 0.00148891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_SCE_c_505_n 0.0180512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_SCE_c_506_n 0.00617327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_SCE_c_507_n 0.00400614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_SCE_c_508_n 0.00238737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_509_n 0.0021066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_510_n 0.00268887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_511_n 0.0012149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_512_n 0.0268957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_SCE_c_513_n 0.00148358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_SCE_c_514_n 0.0277002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_SCE_c_515_n 0.0159686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_299_47#_M1013_g 0.0216077f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_29 VNB N_A_299_47#_c_630_n 0.0135235f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_30 VNB N_A_299_47#_c_631_n 0.00220603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_299_47#_c_632_n 0.00311043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_299_47#_c_633_n 0.00336447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_299_47#_c_634_n 0.0298258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_299_47#_c_635_n 0.00128446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_299_47#_c_636_n 0.00378082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_D_M1014_g 0.0462579f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_37 VNB N_SCD_M1011_g 0.0389108f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_38 VNB N_SCD_c_820_n 0.012101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB SCD 0.00442462f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_40 VNB N_SCD_c_822_n 0.0117071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_193_47#_c_875_n 0.0180432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_193_47#_c_876_n 0.00308215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_193_47#_c_877_n 0.00369255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_193_47#_c_878_n 0.00368817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_193_47#_c_879_n 0.0024951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_193_47#_c_880_n 0.00632811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_193_47#_c_881_n 0.0491774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_193_47#_c_882_n 0.00644541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_193_47#_c_883_n 0.0106143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_193_47#_c_884_n 0.0111044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_193_47#_c_885_n 4.77479e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_193_47#_c_886_n 0.0266741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_193_47#_c_887_n 0.00229326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_193_47#_c_888_n 0.0176132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_193_47#_c_889_n 0.0285203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1092_183#_M1022_g 0.0146965f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_57 VNB N_A_1092_183#_M1007_g 0.0210316f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_58 VNB N_A_1092_183#_c_1093_n 0.00354578f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_59 VNB N_A_1092_183#_c_1094_n 0.00364457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1092_183#_c_1095_n 0.00130744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1092_183#_c_1096_n 0.00302393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1092_183#_c_1097_n 0.0338642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_933_413#_c_1186_n 0.0118275f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_64 VNB N_A_933_413#_c_1187_n 0.0158415f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_65 VNB N_A_933_413#_c_1188_n 0.0152351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_933_413#_c_1189_n 0.00913873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_933_413#_c_1190_n 8.51874e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_933_413#_c_1191_n 0.0118116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_933_413#_c_1192_n 0.00180949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1520_315#_M1017_g 0.0482636f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_71 VNB N_A_1520_315#_c_1297_n 0.00161491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1520_315#_c_1298_n 0.00425124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1520_315#_c_1299_n 0.0267742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1520_315#_c_1300_n 0.00701384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1520_315#_c_1301_n 0.0198034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1349_413#_c_1382_n 0.0205013f $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=2.135
cc_77 VNB N_A_1349_413#_c_1383_n 0.0393229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1349_413#_c_1384_n 0.00807254f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_79 VNB N_A_1349_413#_c_1385_n 0.00998398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1349_413#_c_1386_n 0.00584041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1349_413#_c_1387_n 0.00344545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VPWR_c_1470_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_556_369#_c_1628_n 3.48728e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_556_369#_c_1629_n 0.0117265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_556_369#_c_1630_n 0.00196322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_556_369#_c_1631_n 0.0099948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_556_369#_c_1632_n 0.00880987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_Q_c_1744_n 0.0222649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_Q_c_1745_n 0.020756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1771_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1772_n 0.00278376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1773_n 0.00486519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1774_n 0.0457988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1775_n 0.0058544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1776_n 0.00237946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1777_n 0.00470745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1778_n 0.0430904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1779_n 0.00513917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1780_n 0.0220776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1781_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1782_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1783_n 0.0284383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1784_n 0.0345259f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1785_n 0.0187875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1786_n 0.46424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1787_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1788_n 0.00529791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1789_n 0.0038195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1790_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VPB N_CLK_c_216_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_111 VPB N_CLK_c_220_n 0.0162394f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_112 VPB N_CLK_c_221_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.74
cc_113 VPB N_CLK_c_222_n 0.0235707f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_114 VPB CLK 0.0178159f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_115 VPB N_A_27_47#_M1028_g 0.03676f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_116 VPB N_A_27_47#_c_260_n 0.0143056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_261_n 0.0057729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_M1006_g 0.0191311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_M1026_g 0.033754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_262_n 0.0211567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_277_n 0.00174908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_278_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_27_47#_c_279_n 0.00356676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_47#_c_280_n 0.0581087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_27_47#_c_281_n 0.00148899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_27_47#_c_282_n 7.65147e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_47#_c_283_n 0.00123715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_284_n 0.00853708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_285_n 0.00543917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_268_n 0.0115869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_287_n 0.0266783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_288_n 0.0106236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_269_n 0.0208929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_270_n 0.00437972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_SCE_M1018_g 0.0237177f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_136 VPB N_SCE_c_517_n 0.0172012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_SCE_M1010_g 0.019421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_SCE_c_507_n 0.0010385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_SCE_c_520_n 0.0256568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_SCE_c_514_n 0.00509844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_299_47#_M1012_g 0.0208907f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_142 VPB N_A_299_47#_c_630_n 0.0105295f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_143 VPB N_A_299_47#_c_639_n 0.00436811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_299_47#_c_631_n 0.00421481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_299_47#_c_641_n 0.00208743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_299_47#_c_642_n 0.00191659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_299_47#_c_635_n 5.84774e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_299_47#_c_636_n 0.0278256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_D_M1021_g 0.0189345f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_150 VPB N_D_M1014_g 0.00289755f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.135
cc_151 VPB N_D_c_771_n 0.0270664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_D_c_772_n 0.00443211f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_153 VPB N_SCD_c_823_n 0.0120745f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_154 VPB N_SCD_c_824_n 0.0223039f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_SCD_c_825_n 0.0133451f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_156 VPB SCD 0.0055368f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_157 VPB N_SCD_c_822_n 0.00546905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_193_47#_M1023_g 0.024991f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_159 VPB N_A_193_47#_M1019_g 0.0221869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_193_47#_c_876_n 0.00462988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_193_47#_c_893_n 0.032806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_193_47#_c_877_n 0.00311128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_193_47#_c_895_n 0.00568481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_193_47#_c_896_n 0.0266658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_193_47#_c_884_n 0.0122297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_1092_183#_M1022_g 0.049805f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_167 VPB N_A_1092_183#_c_1096_n 0.00255179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_933_413#_M1008_g 0.0226707f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_169 VPB N_A_933_413#_c_1189_n 0.0189969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_933_413#_c_1190_n 0.00681499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_933_413#_c_1196_n 0.00161138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_933_413#_c_1192_n 0.0087987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_1520_315#_M1001_g 0.0253795f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_174 VPB N_A_1520_315#_M1017_g 0.0179972f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_175 VPB N_A_1520_315#_M1024_g 0.0234525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1520_315#_c_1305_n 0.0128431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1520_315#_c_1306_n 0.0409149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1520_315#_c_1307_n 0.00235569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1520_315#_c_1298_n 0.00425124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1520_315#_c_1299_n 0.00728901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_1349_413#_M1020_g 0.0237342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1349_413#_c_1383_n 0.014657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1349_413#_c_1384_n 5.1131e-19 $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_184 VPB N_A_1349_413#_c_1391_n 0.0126839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1349_413#_c_1385_n 0.00386833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1349_413#_c_1386_n 0.0050339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1471_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1472_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1473_n 0.00484684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1474_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1475_n 0.00548992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1476_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1477_n 0.0515047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1478_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1479_n 0.0452789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1480_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1481_n 0.022285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1482_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1483_n 0.0156572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1484_n 0.0255057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1485_n 0.0371253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1486_n 0.0188998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1470_n 0.061048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1488_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1489_n 0.00436214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1490_n 0.00372368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_556_369#_c_1633_n 0.00847906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_556_369#_c_1634_n 0.00174955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_556_369#_c_1632_n 0.0110955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_556_369#_c_1636_n 0.00873933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_Q_c_1746_n 0.00678872f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_212 VPB N_Q_c_1744_n 0.00944121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB Q 0.028744f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 N_CLK_c_216_n N_A_27_47#_M1015_g 0.0049062f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_215 N_CLK_c_217_n N_A_27_47#_M1015_g 0.0187731f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_216 CLK N_A_27_47#_M1015_g 3.14819e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_217 N_CLK_c_220_n N_A_27_47#_M1028_g 0.00531917f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_218 N_CLK_c_222_n N_A_27_47#_M1028_g 0.0276478f $X=0.475 $Y=1.665 $X2=0 $Y2=0
cc_219 CLK N_A_27_47#_M1028_g 5.73308e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_220 N_CLK_c_216_n N_A_27_47#_c_264_n 0.00761961f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_221 N_CLK_c_217_n N_A_27_47#_c_264_n 0.00668648f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_222 CLK N_A_27_47#_c_264_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_223 N_CLK_c_216_n N_A_27_47#_c_265_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_224 CLK N_A_27_47#_c_265_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_225 N_CLK_c_221_n N_A_27_47#_c_277_n 0.0128144f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_226 N_CLK_c_222_n N_A_27_47#_c_277_n 0.0013816f $X=0.475 $Y=1.665 $X2=0 $Y2=0
cc_227 CLK N_A_27_47#_c_277_n 0.00728212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_228 N_CLK_c_216_n N_A_27_47#_c_266_n 3.98708e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_229 CLK N_A_27_47#_c_266_n 0.0516739f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_230 N_CLK_c_216_n N_A_27_47#_c_278_n 2.90926e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_231 N_CLK_c_220_n N_A_27_47#_c_278_n 7.09762e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_232 N_CLK_c_222_n N_A_27_47#_c_278_n 0.00440146f $X=0.475 $Y=1.665 $X2=0
+ $Y2=0
cc_233 N_CLK_c_216_n N_A_27_47#_c_279_n 2.26313e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_234 N_CLK_c_221_n N_A_27_47#_c_279_n 2.17882e-19 $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_235 N_CLK_c_222_n N_A_27_47#_c_279_n 0.00358837f $X=0.475 $Y=1.665 $X2=0
+ $Y2=0
cc_236 CLK N_A_27_47#_c_279_n 0.0153364f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_237 N_CLK_c_216_n N_A_27_47#_c_267_n 0.00381855f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_238 N_CLK_c_221_n N_A_27_47#_c_281_n 0.00101286f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_239 N_CLK_c_216_n N_A_27_47#_c_268_n 0.0169285f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_240 CLK N_A_27_47#_c_268_n 0.00161876f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_241 N_CLK_c_221_n N_VPWR_c_1471_n 0.00946555f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_221_n N_VPWR_c_1483_n 0.00332278f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_243 N_CLK_c_221_n N_VPWR_c_1470_n 0.00485269f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_244 N_CLK_c_217_n N_VGND_c_1771_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_245 N_CLK_c_216_n N_VGND_c_1782_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_246 N_CLK_c_217_n N_VGND_c_1782_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_247 N_CLK_c_217_n N_VGND_c_1786_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_280_n N_SCE_M1018_g 0.00256669f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_280_n N_SCE_M1010_g 0.00122494f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_280_n N_SCE_c_507_n 0.00406375f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_280_n N_SCE_c_520_n 0.0034961f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_280_n N_A_299_47#_M1012_g 3.67555e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_280_n N_A_299_47#_c_630_n 0.0120796f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_280_n N_A_299_47#_c_647_n 0.0162863f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_280_n N_A_299_47#_c_631_n 0.00918627f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_280_n N_A_299_47#_c_649_n 0.0355887f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_280_n N_A_299_47#_c_641_n 0.0116459f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1015_g N_A_299_47#_c_632_n 0.00126581f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_280_n N_A_299_47#_c_642_n 0.0138552f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_280_n N_A_299_47#_c_634_n 0.0024684f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_280_n N_A_299_47#_c_654_n 0.00478262f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_280_n N_A_299_47#_c_635_n 0.00152384f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_280_n N_A_299_47#_c_636_n 0.00124511f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_280_n N_D_M1021_g 0.00200411f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_280_n N_D_c_771_n 0.00308822f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_280_n N_D_c_772_n 0.00836282f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_267 N_A_27_47#_M1030_g N_SCD_c_820_n 0.00132967f $X=4.595 $Y=0.415 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_280_n N_SCD_c_824_n 0.00226525f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_280_n SCD 0.0116881f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_261_n N_SCD_c_822_n 0.00132967f $X=4.67 $Y=1.32 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_280_n N_A_193_47#_M1028_d 6.81311e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_280_n N_A_193_47#_M1023_g 0.00371812f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_284_n N_A_193_47#_M1023_g 9.60176e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_287_n N_A_193_47#_M1023_g 0.0144159f $X=5.115 $Y=1.74 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1003_g N_A_193_47#_c_875_n 0.0144677f $X=7.315 $Y=0.415 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1026_g N_A_193_47#_M1019_g 0.0175056f $X=6.67 $Y=2.275 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_285_n N_A_193_47#_M1019_g 0.00135837f $X=6.675 $Y=1.87 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_270_n N_A_193_47#_M1019_g 5.16255e-19 $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1030_g N_A_193_47#_c_876_n 0.00723459f $X=4.595 $Y=0.415
+ $X2=0 $Y2=0
cc_280 N_A_27_47#_c_260_n N_A_193_47#_c_876_n 0.00724741f $X=4.98 $Y=1.32 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_261_n N_A_193_47#_c_876_n 0.00418731f $X=4.67 $Y=1.32 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_280_n N_A_193_47#_c_876_n 0.0139192f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_283_n N_A_193_47#_c_876_n 2.04934e-19 $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_284_n N_A_193_47#_c_876_n 0.0169135f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_287_n N_A_193_47#_c_876_n 7.29366e-19 $X=5.115 $Y=1.74 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_288_n N_A_193_47#_c_876_n 0.00604391f $X=5.115 $Y=1.575
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_c_261_n N_A_193_47#_c_893_n 0.016259f $X=4.67 $Y=1.32 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_280_n N_A_193_47#_c_893_n 0.00545515f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_284_n N_A_193_47#_c_893_n 0.00118389f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_287_n N_A_193_47#_c_893_n 0.0174998f $X=5.115 $Y=1.74 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_262_n N_A_193_47#_c_877_n 0.0117161f $X=7.24 $Y=1.32 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_M1003_g N_A_193_47#_c_877_n 0.00430042f $X=7.315 $Y=0.415
+ $X2=0 $Y2=0
cc_293 N_A_27_47#_c_269_n N_A_193_47#_c_877_n 0.00402309f $X=6.665 $Y=1.32 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_270_n N_A_193_47#_c_877_n 0.0234373f $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1015_g N_A_193_47#_c_878_n 0.00136206f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_264_n N_A_193_47#_c_878_n 0.00440816f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_M1030_g N_A_193_47#_c_879_n 0.0112301f $X=4.595 $Y=0.415 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1003_g N_A_193_47#_c_880_n 0.0020279f $X=7.315 $Y=0.415 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_269_n N_A_193_47#_c_880_n 0.00222109f $X=6.665 $Y=1.32 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_270_n N_A_193_47#_c_880_n 0.0119224f $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1026_g N_A_193_47#_c_895_n 0.00117691f $X=6.67 $Y=2.275 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_262_n N_A_193_47#_c_895_n 0.00338756f $X=7.24 $Y=1.32 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_285_n N_A_193_47#_c_895_n 0.00508223f $X=6.675 $Y=1.87 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_270_n N_A_193_47#_c_895_n 0.0245744f $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_M1026_g N_A_193_47#_c_896_n 0.0130792f $X=6.67 $Y=2.275 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_262_n N_A_193_47#_c_896_n 0.0212127f $X=7.24 $Y=1.32 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_270_n N_A_193_47#_c_896_n 6.54911e-19 $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_M1030_g N_A_193_47#_c_881_n 0.00407284f $X=4.595 $Y=0.415
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_M1015_g N_A_193_47#_c_882_n 0.00666063f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_264_n N_A_193_47#_c_882_n 0.00223754f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_267_n N_A_193_47#_c_882_n 0.00522408f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_269_n N_A_193_47#_c_883_n 8.71689e-19 $X=6.665 $Y=1.32 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_M1015_g N_A_193_47#_c_884_n 0.0085043f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_264_n N_A_193_47#_c_884_n 0.00552566f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_266_n N_A_193_47#_c_884_n 0.0594418f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_386_p N_A_193_47#_c_884_n 0.00825932f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_267_n N_A_193_47#_c_884_n 0.00881475f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_280_n N_A_193_47#_c_884_n 0.0231935f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_281_n N_A_193_47#_c_884_n 0.00244175f $X=0.87 $Y=1.87 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_268_n N_A_193_47#_c_884_n 0.0174534f $X=0.895 $Y=1.235 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_269_n N_A_193_47#_c_885_n 2.55286e-19 $X=6.665 $Y=1.32 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_270_n N_A_193_47#_c_885_n 0.00125233f $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_M1030_g N_A_193_47#_c_886_n 0.0213113f $X=4.595 $Y=0.415 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_260_n N_A_193_47#_c_886_n 0.0174066f $X=4.98 $Y=1.32 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_284_n N_A_193_47#_c_886_n 4.76262e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_287_n N_A_193_47#_c_886_n 5.43883e-19 $X=5.115 $Y=1.74 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_260_n N_A_193_47#_c_887_n 0.00542986f $X=4.98 $Y=1.32 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_284_n N_A_193_47#_c_887_n 0.00398178f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_M1030_g N_A_193_47#_c_888_n 0.010243f $X=4.595 $Y=0.415 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_M1003_g N_A_193_47#_c_889_n 0.0193601f $X=7.315 $Y=0.415 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_269_n N_A_193_47#_c_889_n 0.020308f $X=6.665 $Y=1.32 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_282_n N_A_1092_183#_M1008_d 0.00523078f $X=6.53 $Y=1.87
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_260_n N_A_1092_183#_M1022_g 0.0113457f $X=4.98 $Y=1.32 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_M1006_g N_A_1092_183#_M1022_g 0.0276008f $X=5.055 $Y=2.275
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_282_n N_A_1092_183#_M1022_g 0.00281129f $X=6.53 $Y=1.87
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_283_n N_A_1092_183#_M1022_g 0.00151609f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_284_n N_A_1092_183#_M1022_g 0.0022f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_287_n N_A_1092_183#_M1022_g 0.0206011f $X=5.115 $Y=1.74
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_c_282_n N_A_1092_183#_c_1107_n 0.00261642f $X=6.53 $Y=1.87
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_M1026_g N_A_1092_183#_c_1096_n 0.00455971f $X=6.67 $Y=2.275
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_282_n N_A_1092_183#_c_1096_n 0.0193938f $X=6.53 $Y=1.87
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_c_285_n N_A_1092_183#_c_1096_n 0.00314501f $X=6.675 $Y=1.87
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_c_269_n N_A_1092_183#_c_1096_n 0.00225153f $X=6.665 $Y=1.32
+ $X2=0 $Y2=0
cc_344 N_A_27_47#_c_270_n N_A_1092_183#_c_1096_n 0.0517078f $X=6.665 $Y=1.41
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_269_n N_A_933_413#_c_1186_n 0.0158005f $X=6.665 $Y=1.32
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_c_270_n N_A_933_413#_c_1186_n 3.03019e-19 $X=6.665 $Y=1.41
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_M1026_g N_A_933_413#_M1008_g 0.0247799f $X=6.67 $Y=2.275 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_282_n N_A_933_413#_M1008_g 0.00700233f $X=6.53 $Y=1.87 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_270_n N_A_933_413#_M1008_g 8.29633e-19 $X=6.665 $Y=1.41
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_282_n N_A_933_413#_c_1189_n 0.00109659f $X=6.53 $Y=1.87
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_M1006_g N_A_933_413#_c_1204_n 0.00859956f $X=5.055 $Y=2.275
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_c_280_n N_A_933_413#_c_1204_n 0.00708547f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_282_n N_A_933_413#_c_1204_n 0.00299508f $X=6.53 $Y=1.87
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_283_n N_A_933_413#_c_1204_n 0.00236799f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_284_n N_A_933_413#_c_1204_n 0.0252894f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_287_n N_A_933_413#_c_1204_n 5.38487e-19 $X=5.115 $Y=1.74
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_M1030_g N_A_933_413#_c_1191_n 0.00106635f $X=4.595 $Y=0.415
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_c_260_n N_A_933_413#_c_1191_n 8.14452e-19 $X=4.98 $Y=1.32
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_M1006_g N_A_933_413#_c_1196_n 9.97608e-19 $X=5.055 $Y=2.275
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_c_282_n N_A_933_413#_c_1196_n 0.0183205f $X=6.53 $Y=1.87 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_283_n N_A_933_413#_c_1196_n 0.00266197f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_284_n N_A_933_413#_c_1196_n 0.0249845f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_287_n N_A_933_413#_c_1196_n 7.00613e-19 $X=5.115 $Y=1.74
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_260_n N_A_933_413#_c_1192_n 0.00225879f $X=4.98 $Y=1.32
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_282_n N_A_933_413#_c_1192_n 0.0162495f $X=6.53 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_283_n N_A_933_413#_c_1192_n 0.00303482f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_c_284_n N_A_933_413#_c_1192_n 0.00980238f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_c_288_n N_A_933_413#_c_1192_n 4.44848e-19 $X=5.115 $Y=1.575
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_M1003_g N_A_1520_315#_M1017_g 0.0463015f $X=7.315 $Y=0.415
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_M1026_g N_A_1349_413#_c_1394_n 0.00281529f $X=6.67 $Y=2.275
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_285_n N_A_1349_413#_c_1394_n 0.00210372f $X=6.675 $Y=1.87
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_270_n N_A_1349_413#_c_1394_n 0.0022468f $X=6.665 $Y=1.41
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_M1003_g N_A_1349_413#_c_1397_n 0.00800808f $X=7.315 $Y=0.415
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_285_n N_A_1349_413#_c_1391_n 0.00228172f $X=6.675 $Y=1.87
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_270_n N_A_1349_413#_c_1391_n 9.63849e-19 $X=6.665 $Y=1.41
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_M1003_g N_A_1349_413#_c_1385_n 3.1587e-19 $X=7.315 $Y=0.415
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_262_n N_A_1349_413#_c_1386_n 0.00558094f $X=7.24 $Y=1.32
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_M1003_g N_A_1349_413#_c_1386_n 0.0061466f $X=7.315 $Y=0.415
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_M1003_g N_A_1349_413#_c_1387_n 0.0110495f $X=7.315 $Y=0.415
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_386_p N_VPWR_M1005_d 6.91013e-19 $X=0.73 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_381 N_A_27_47#_c_281_n N_VPWR_M1005_d 0.00178771f $X=0.87 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_27_47#_c_282_n N_VPWR_M1022_d 0.00678497f $X=6.53 $Y=1.87 $X2=0 $Y2=0
cc_383 N_A_27_47#_M1028_g N_VPWR_c_1471_n 0.00937841f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_277_n N_VPWR_c_1471_n 0.0031092f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_386_p N_VPWR_c_1471_n 0.0133497f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_279_n N_VPWR_c_1471_n 0.012721f $X=0.265 $Y=1.96 $X2=0 $Y2=0
cc_387 N_A_27_47#_c_281_n N_VPWR_c_1471_n 0.00330948f $X=0.87 $Y=1.87 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_280_n N_VPWR_c_1472_n 0.00124401f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_280_n N_VPWR_c_1473_n 9.19647e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_282_n N_VPWR_c_1474_n 0.00950843f $X=6.53 $Y=1.87 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_M1006_g N_VPWR_c_1477_n 0.0037886f $X=5.055 $Y=2.275 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_M1026_g N_VPWR_c_1479_n 0.00430107f $X=6.67 $Y=2.275 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_270_n N_VPWR_c_1479_n 0.00157744f $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_277_n N_VPWR_c_1483_n 0.0018545f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_279_n N_VPWR_c_1483_n 0.0120313f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1028_g N_VPWR_c_1484_n 0.00442511f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_M1028_g N_VPWR_c_1470_n 0.00534571f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_M1006_g N_VPWR_c_1470_n 0.00557714f $X=5.055 $Y=2.275 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_M1026_g N_VPWR_c_1470_n 0.0057371f $X=6.67 $Y=2.275 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_277_n N_VPWR_c_1470_n 0.00403677f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_279_n N_VPWR_c_1470_n 0.00646745f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_280_n N_VPWR_c_1470_n 0.199094f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_403 N_A_27_47#_c_281_n N_VPWR_c_1470_n 0.0145601f $X=0.87 $Y=1.87 $X2=0 $Y2=0
cc_404 N_A_27_47#_c_282_n N_VPWR_c_1470_n 0.0517485f $X=6.53 $Y=1.87 $X2=0 $Y2=0
cc_405 N_A_27_47#_c_283_n N_VPWR_c_1470_n 0.0148452f $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_285_n N_VPWR_c_1470_n 0.0159329f $X=6.675 $Y=1.87 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_270_n N_VPWR_c_1470_n 0.00100625f $X=6.665 $Y=1.41 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_c_280_n N_A_556_369#_c_1637_n 0.00544764f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_280_n N_A_556_369#_c_1633_n 0.0227214f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_280_n N_A_556_369#_c_1634_n 0.0106068f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_M1030_g N_A_556_369#_c_1631_n 0.0100896f $X=4.595 $Y=0.415
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_M1030_g N_A_556_369#_c_1632_n 0.00550322f $X=4.595 $Y=0.415
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_280_n N_A_556_369#_c_1632_n 0.0104876f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_280_n N_A_556_369#_c_1636_n 0.0111926f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_415 N_A_27_47#_c_284_n N_A_556_369#_c_1636_n 0.00314032f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_280_n A_640_369# 0.00134881f $X=5.145 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_417 N_A_27_47#_c_264_n N_VGND_M1029_d 0.00166329f $X=0.615 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_418 N_A_27_47#_M1015_g N_VGND_c_1771_n 0.00965468f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_264_n N_VGND_c_1771_n 0.0150403f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_266_n N_VGND_c_1771_n 0.00108069f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_268_n N_VGND_c_1771_n 5.70216e-19 $X=0.895 $Y=1.235 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1030_g N_VGND_c_1773_n 0.00293607f $X=4.595 $Y=0.415 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_M1030_g N_VGND_c_1774_n 0.00545274f $X=4.595 $Y=0.415 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_M1003_g N_VGND_c_1776_n 0.00230753f $X=7.315 $Y=0.415 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_M1003_g N_VGND_c_1778_n 0.00379696f $X=7.315 $Y=0.415 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_c_496_p N_VGND_c_1782_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_264_n N_VGND_c_1782_n 0.00243651f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_M1015_g N_VGND_c_1783_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_M1029_s N_VGND_c_1786_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_M1015_g N_VGND_c_1786_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_M1030_g N_VGND_c_1786_n 0.00731459f $X=4.595 $Y=0.415 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_M1003_g N_VGND_c_1786_n 0.00575728f $X=7.315 $Y=0.415 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_496_p N_VGND_c_1786_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_264_n N_VGND_c_1786_n 0.00564532f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_435 N_SCE_c_505_n N_A_299_47#_M1013_g 0.0186561f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_436 N_SCE_c_507_n N_A_299_47#_M1013_g 9.16072e-19 $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_437 N_SCE_c_508_n N_A_299_47#_M1013_g 0.0105179f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_438 N_SCE_c_509_n N_A_299_47#_M1013_g 7.13575e-19 $X=1.99 $Y=0.7 $X2=0 $Y2=0
cc_439 SCE N_A_299_47#_M1013_g 0.00483914f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_440 N_SCE_c_514_n N_A_299_47#_M1013_g 0.00330265f $X=1.855 $Y=1.385 $X2=0
+ $Y2=0
cc_441 N_SCE_M1018_g N_A_299_47#_c_630_n 0.00425611f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_442 N_SCE_c_505_n N_A_299_47#_c_630_n 0.00426868f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_443 N_SCE_c_506_n N_A_299_47#_c_630_n 0.012036f $X=1.84 $Y=0.815 $X2=0 $Y2=0
cc_444 N_SCE_c_507_n N_A_299_47#_c_630_n 0.0602583f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_445 N_SCE_c_520_n N_A_299_47#_c_630_n 0.00698249f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_446 N_SCE_c_509_n N_A_299_47#_c_630_n 0.0157003f $X=1.99 $Y=0.7 $X2=0 $Y2=0
cc_447 N_SCE_M1018_g N_A_299_47#_c_647_n 0.0122756f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_448 N_SCE_c_507_n N_A_299_47#_c_647_n 0.0105401f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_449 N_SCE_c_520_n N_A_299_47#_c_647_n 0.00408496f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_450 N_SCE_M1018_g N_A_299_47#_c_631_n 0.00147664f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_451 N_SCE_c_517_n N_A_299_47#_c_631_n 0.00774359f $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_452 N_SCE_M1010_g N_A_299_47#_c_631_n 0.00579344f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_453 N_SCE_c_507_n N_A_299_47#_c_631_n 0.0376646f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_454 N_SCE_c_520_n N_A_299_47#_c_631_n 0.00129015f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_455 N_SCE_c_514_n N_A_299_47#_c_631_n 0.00132872f $X=1.855 $Y=1.385 $X2=0
+ $Y2=0
cc_456 N_SCE_M1010_g N_A_299_47#_c_649_n 0.0054673f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_457 N_SCE_c_505_n N_A_299_47#_c_632_n 0.00242797f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_458 N_SCE_c_509_n N_A_299_47#_c_632_n 9.9503e-19 $X=1.99 $Y=0.7 $X2=0 $Y2=0
cc_459 N_SCE_c_520_n N_A_299_47#_c_642_n 2.83838e-19 $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_460 N_SCE_c_517_n N_A_299_47#_c_633_n 3.99992e-19 $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_461 N_SCE_c_507_n N_A_299_47#_c_633_n 0.0119415f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_462 N_SCE_c_508_n N_A_299_47#_c_633_n 0.0201957f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_463 N_SCE_c_511_n N_A_299_47#_c_633_n 0.00390849f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_464 N_SCE_c_514_n N_A_299_47#_c_633_n 2.03234e-19 $X=1.855 $Y=1.385 $X2=0
+ $Y2=0
cc_465 N_SCE_c_517_n N_A_299_47#_c_634_n 0.00856869f $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_466 N_SCE_c_507_n N_A_299_47#_c_634_n 0.00176299f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_467 N_SCE_c_508_n N_A_299_47#_c_634_n 0.00317862f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_468 N_SCE_c_514_n N_A_299_47#_c_634_n 0.0172737f $X=1.855 $Y=1.385 $X2=0
+ $Y2=0
cc_469 N_SCE_M1010_g N_A_299_47#_c_654_n 0.00682561f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_470 N_SCE_c_510_n N_A_299_47#_c_635_n 2.16874e-19 $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_471 N_SCE_c_511_n N_A_299_47#_c_635_n 0.0115929f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_472 N_SCE_c_512_n N_A_299_47#_c_635_n 4.48662e-19 $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_473 N_SCE_c_511_n N_A_299_47#_c_636_n 2.28784e-19 $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_474 N_SCE_c_512_n N_A_299_47#_c_636_n 0.015542f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_475 N_SCE_M1010_g N_D_M1021_g 0.0406154f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_476 N_SCE_c_510_n N_D_M1014_g 0.0124861f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_477 N_SCE_c_511_n N_D_M1014_g 0.0019752f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_478 N_SCE_c_512_n N_D_M1014_g 0.0214615f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_479 N_SCE_c_515_n N_D_M1014_g 0.0129735f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_480 N_SCE_c_517_n N_D_c_771_n 0.00996826f $X=2.185 $Y=1.58 $X2=0 $Y2=0
cc_481 N_SCE_c_520_n N_D_c_771_n 0.00174797f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_482 N_SCE_c_510_n N_D_c_771_n 7.89925e-19 $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_483 N_SCE_c_513_n N_D_c_771_n 0.00128987f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_484 N_SCE_c_514_n N_D_c_771_n 3.28065e-19 $X=1.855 $Y=1.385 $X2=0 $Y2=0
cc_485 N_SCE_c_517_n N_D_c_772_n 0.0012389f $X=2.185 $Y=1.58 $X2=0 $Y2=0
cc_486 N_SCE_c_508_n N_D_c_772_n 2.69368e-19 $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_487 N_SCE_c_510_n N_D_c_772_n 0.00184567f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_488 N_SCE_c_513_n N_D_c_772_n 0.00314298f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_489 N_SCE_c_511_n N_SCD_M1011_g 0.00141715f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_490 N_SCE_c_515_n N_SCD_M1011_g 0.0560917f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_491 N_SCE_c_511_n SCD 0.00198147f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_492 N_SCE_c_517_n N_A_193_47#_c_881_n 0.00184114f $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_493 N_SCE_c_506_n N_A_193_47#_c_881_n 5.97087e-19 $X=1.84 $Y=0.815 $X2=0
+ $Y2=0
cc_494 N_SCE_c_507_n N_A_193_47#_c_881_n 0.0135865f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_495 N_SCE_c_520_n N_A_193_47#_c_881_n 0.00293807f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_496 N_SCE_c_508_n N_A_193_47#_c_881_n 0.0148275f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_497 N_SCE_c_509_n N_A_193_47#_c_881_n 0.00951232f $X=1.99 $Y=0.7 $X2=0 $Y2=0
cc_498 N_SCE_c_510_n N_A_193_47#_c_881_n 0.0196688f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_499 N_SCE_c_511_n N_A_193_47#_c_881_n 0.0108237f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_500 N_SCE_c_512_n N_A_193_47#_c_881_n 0.00367465f $X=3.15 $Y=0.93 $X2=0 $Y2=0
cc_501 N_SCE_c_513_n N_A_193_47#_c_881_n 0.00735012f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_502 N_SCE_c_514_n N_A_193_47#_c_881_n 0.00192272f $X=1.855 $Y=1.385 $X2=0
+ $Y2=0
cc_503 N_SCE_M1018_g N_A_193_47#_c_884_n 0.00154779f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_504 N_SCE_M1018_g N_VPWR_c_1472_n 0.00870017f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_505 N_SCE_M1010_g N_VPWR_c_1472_n 0.0092033f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_506 N_SCE_M1018_g N_VPWR_c_1484_n 0.00340533f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_507 N_SCE_M1010_g N_VPWR_c_1485_n 0.00354675f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_508 N_SCE_M1018_g N_VPWR_c_1470_n 0.00515557f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_509 N_SCE_M1010_g N_VPWR_c_1470_n 0.00400283f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_510 N_SCE_c_510_n N_A_556_369#_M1014_d 0.00218877f $X=3.065 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_511 N_SCE_M1010_g N_A_556_369#_c_1637_n 5.52806e-19 $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_512 N_SCE_c_510_n N_A_556_369#_c_1647_n 0.0214191f $X=3.065 $Y=0.7 $X2=0
+ $Y2=0
cc_513 N_SCE_c_512_n N_A_556_369#_c_1647_n 5.06463e-19 $X=3.15 $Y=0.93 $X2=0
+ $Y2=0
cc_514 N_SCE_c_515_n N_A_556_369#_c_1647_n 0.00756611f $X=3.15 $Y=0.765 $X2=0
+ $Y2=0
cc_515 N_SCE_c_510_n N_A_556_369#_c_1628_n 0.0079009f $X=3.065 $Y=0.7 $X2=0
+ $Y2=0
cc_516 N_SCE_c_515_n N_A_556_369#_c_1628_n 0.0040848f $X=3.15 $Y=0.765 $X2=0
+ $Y2=0
cc_517 N_SCE_c_510_n N_A_556_369#_c_1630_n 0.00610516f $X=3.065 $Y=0.7 $X2=0
+ $Y2=0
cc_518 N_SCE_c_511_n N_A_556_369#_c_1630_n 0.00694211f $X=3.15 $Y=0.93 $X2=0
+ $Y2=0
cc_519 N_SCE_c_515_n N_A_556_369#_c_1630_n 9.24156e-19 $X=3.15 $Y=0.765 $X2=0
+ $Y2=0
cc_520 N_SCE_c_508_n N_VGND_M1031_d 0.00221059f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_521 N_SCE_c_505_n N_VGND_c_1772_n 0.00416942f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_522 N_SCE_c_508_n N_VGND_c_1772_n 0.0178763f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_523 N_SCE_c_509_n N_VGND_c_1772_n 5.78103e-19 $X=1.99 $Y=0.7 $X2=0 $Y2=0
cc_524 SCE N_VGND_c_1772_n 0.0103951f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_525 N_SCE_c_505_n N_VGND_c_1783_n 0.00417177f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_526 N_SCE_c_509_n N_VGND_c_1783_n 0.00282365f $X=1.99 $Y=0.7 $X2=0 $Y2=0
cc_527 N_SCE_c_508_n N_VGND_c_1784_n 0.0024952f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_528 N_SCE_c_510_n N_VGND_c_1784_n 0.00277894f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_529 SCE N_VGND_c_1784_n 0.00772962f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_530 N_SCE_c_515_n N_VGND_c_1784_n 0.00362032f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_531 N_SCE_c_505_n N_VGND_c_1786_n 0.00687852f $X=1.84 $Y=0.73 $X2=0 $Y2=0
cc_532 N_SCE_c_508_n N_VGND_c_1786_n 0.0027377f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_533 N_SCE_c_509_n N_VGND_c_1786_n 0.00220581f $X=1.99 $Y=0.7 $X2=0 $Y2=0
cc_534 N_SCE_c_510_n N_VGND_c_1786_n 0.00226167f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_535 SCE N_VGND_c_1786_n 0.00302552f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_536 N_SCE_c_515_n N_VGND_c_1786_n 0.00526606f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_537 SCE A_483_47# 0.00514624f $X=2.475 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_538 N_A_299_47#_M1012_g N_D_M1021_g 0.0283246f $X=3.125 $Y=2.165 $X2=0 $Y2=0
cc_539 N_A_299_47#_c_631_n N_D_M1021_g 0.00115294f $X=2.202 $Y=1.86 $X2=0 $Y2=0
cc_540 N_A_299_47#_c_649_n N_D_M1021_g 0.0118022f $X=3.05 $Y=1.967 $X2=0 $Y2=0
cc_541 N_A_299_47#_c_641_n N_D_M1021_g 0.00129689f $X=3.135 $Y=1.86 $X2=0 $Y2=0
cc_542 N_A_299_47#_M1013_g N_D_M1014_g 0.0415208f $X=2.34 $Y=0.445 $X2=0 $Y2=0
cc_543 N_A_299_47#_c_631_n N_D_M1014_g 0.00511189f $X=2.202 $Y=1.86 $X2=0 $Y2=0
cc_544 N_A_299_47#_c_633_n N_D_M1014_g 0.0020825f $X=2.28 $Y=1.045 $X2=0 $Y2=0
cc_545 N_A_299_47#_c_634_n N_D_M1014_g 0.0168022f $X=2.28 $Y=1.045 $X2=0 $Y2=0
cc_546 N_A_299_47#_c_635_n N_D_M1014_g 3.21995e-19 $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_547 N_A_299_47#_c_636_n N_D_M1014_g 0.00266404f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_548 N_A_299_47#_c_631_n N_D_c_771_n 6.16226e-19 $X=2.202 $Y=1.86 $X2=0 $Y2=0
cc_549 N_A_299_47#_c_649_n N_D_c_771_n 0.00294687f $X=3.05 $Y=1.967 $X2=0 $Y2=0
cc_550 N_A_299_47#_c_635_n N_D_c_771_n 0.00116042f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_551 N_A_299_47#_c_636_n N_D_c_771_n 0.0195382f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_552 N_A_299_47#_c_631_n N_D_c_772_n 0.0254671f $X=2.202 $Y=1.86 $X2=0 $Y2=0
cc_553 N_A_299_47#_c_649_n N_D_c_772_n 0.0194959f $X=3.05 $Y=1.967 $X2=0 $Y2=0
cc_554 N_A_299_47#_c_635_n N_D_c_772_n 0.0169894f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_555 N_A_299_47#_c_636_n N_D_c_772_n 0.00100629f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_556 N_A_299_47#_M1012_g N_SCD_c_823_n 0.00264946f $X=3.125 $Y=2.165 $X2=0
+ $Y2=0
cc_557 N_A_299_47#_c_641_n N_SCD_c_823_n 0.00118569f $X=3.135 $Y=1.86 $X2=0
+ $Y2=0
cc_558 N_A_299_47#_M1012_g N_SCD_c_824_n 0.0341472f $X=3.125 $Y=2.165 $X2=0
+ $Y2=0
cc_559 N_A_299_47#_c_649_n N_SCD_c_824_n 2.09833e-19 $X=3.05 $Y=1.967 $X2=0
+ $Y2=0
cc_560 N_A_299_47#_c_641_n N_SCD_c_824_n 0.00185718f $X=3.135 $Y=1.86 $X2=0
+ $Y2=0
cc_561 N_A_299_47#_c_641_n SCD 9.59643e-19 $X=3.135 $Y=1.86 $X2=0 $Y2=0
cc_562 N_A_299_47#_c_635_n SCD 0.017508f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_563 N_A_299_47#_c_636_n SCD 0.00114843f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_564 N_A_299_47#_c_635_n N_SCD_c_822_n 9.90326e-19 $X=3.185 $Y=1.47 $X2=0
+ $Y2=0
cc_565 N_A_299_47#_c_636_n N_SCD_c_822_n 0.0193339f $X=3.185 $Y=1.47 $X2=0 $Y2=0
cc_566 N_A_299_47#_c_630_n N_A_193_47#_c_878_n 0.0959385f $X=1.505 $Y=1.86 $X2=0
+ $Y2=0
cc_567 N_A_299_47#_c_632_n N_A_193_47#_c_878_n 0.00899224f $X=1.625 $Y=0.38
+ $X2=0 $Y2=0
cc_568 N_A_299_47#_M1013_g N_A_193_47#_c_881_n 0.00179873f $X=2.34 $Y=0.445
+ $X2=0 $Y2=0
cc_569 N_A_299_47#_c_630_n N_A_193_47#_c_881_n 0.0179969f $X=1.505 $Y=1.86 $X2=0
+ $Y2=0
cc_570 N_A_299_47#_c_632_n N_A_193_47#_c_881_n 0.00483511f $X=1.625 $Y=0.38
+ $X2=0 $Y2=0
cc_571 N_A_299_47#_c_633_n N_A_193_47#_c_881_n 0.00870823f $X=2.28 $Y=1.045
+ $X2=0 $Y2=0
cc_572 N_A_299_47#_c_634_n N_A_193_47#_c_881_n 0.00446499f $X=2.28 $Y=1.045
+ $X2=0 $Y2=0
cc_573 N_A_299_47#_c_635_n N_A_193_47#_c_881_n 0.00194601f $X=3.185 $Y=1.47
+ $X2=0 $Y2=0
cc_574 N_A_299_47#_c_636_n N_A_193_47#_c_881_n 8.21137e-19 $X=3.185 $Y=1.47
+ $X2=0 $Y2=0
cc_575 N_A_299_47#_c_630_n N_A_193_47#_c_882_n 0.00266292f $X=1.505 $Y=1.86
+ $X2=0 $Y2=0
cc_576 N_A_299_47#_c_639_n N_A_193_47#_c_884_n 0.0267023f $X=1.625 $Y=2.175
+ $X2=0 $Y2=0
cc_577 N_A_299_47#_c_642_n N_A_193_47#_c_884_n 0.0154783f $X=1.565 $Y=1.967
+ $X2=0 $Y2=0
cc_578 N_A_299_47#_c_647_n N_VPWR_M1018_d 0.00402367f $X=2.115 $Y=1.967 $X2=0
+ $Y2=0
cc_579 N_A_299_47#_c_647_n N_VPWR_c_1472_n 0.0125181f $X=2.115 $Y=1.967 $X2=0
+ $Y2=0
cc_580 N_A_299_47#_c_654_n N_VPWR_c_1472_n 0.00272071f $X=2.202 $Y=1.967 $X2=0
+ $Y2=0
cc_581 N_A_299_47#_c_639_n N_VPWR_c_1484_n 0.0177913f $X=1.625 $Y=2.175 $X2=0
+ $Y2=0
cc_582 N_A_299_47#_c_647_n N_VPWR_c_1484_n 0.00240758f $X=2.115 $Y=1.967 $X2=0
+ $Y2=0
cc_583 N_A_299_47#_M1012_g N_VPWR_c_1485_n 0.00368123f $X=3.125 $Y=2.165 $X2=0
+ $Y2=0
cc_584 N_A_299_47#_c_649_n N_VPWR_c_1485_n 0.00593225f $X=3.05 $Y=1.967 $X2=0
+ $Y2=0
cc_585 N_A_299_47#_c_654_n N_VPWR_c_1485_n 0.00138725f $X=2.202 $Y=1.967 $X2=0
+ $Y2=0
cc_586 N_A_299_47#_M1018_s N_VPWR_c_1470_n 0.00184114f $X=1.5 $Y=1.845 $X2=0
+ $Y2=0
cc_587 N_A_299_47#_M1012_g N_VPWR_c_1470_n 0.00536624f $X=3.125 $Y=2.165 $X2=0
+ $Y2=0
cc_588 N_A_299_47#_c_639_n N_VPWR_c_1470_n 0.00521387f $X=1.625 $Y=2.175 $X2=0
+ $Y2=0
cc_589 N_A_299_47#_c_647_n N_VPWR_c_1470_n 0.00246602f $X=2.115 $Y=1.967 $X2=0
+ $Y2=0
cc_590 N_A_299_47#_c_649_n N_VPWR_c_1470_n 0.00540738f $X=3.05 $Y=1.967 $X2=0
+ $Y2=0
cc_591 N_A_299_47#_c_654_n N_VPWR_c_1470_n 0.00123093f $X=2.202 $Y=1.967 $X2=0
+ $Y2=0
cc_592 N_A_299_47#_c_649_n A_467_369# 0.00491631f $X=3.05 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_593 N_A_299_47#_c_649_n N_A_556_369#_M1021_d 0.00422263f $X=3.05 $Y=1.967
+ $X2=0 $Y2=0
cc_594 N_A_299_47#_M1012_g N_A_556_369#_c_1637_n 0.00815124f $X=3.125 $Y=2.165
+ $X2=0 $Y2=0
cc_595 N_A_299_47#_c_649_n N_A_556_369#_c_1637_n 0.0257062f $X=3.05 $Y=1.967
+ $X2=0 $Y2=0
cc_596 N_A_299_47#_c_635_n N_A_556_369#_c_1637_n 3.10199e-19 $X=3.185 $Y=1.47
+ $X2=0 $Y2=0
cc_597 N_A_299_47#_c_636_n N_A_556_369#_c_1637_n 0.00134649f $X=3.185 $Y=1.47
+ $X2=0 $Y2=0
cc_598 N_A_299_47#_M1012_g N_A_556_369#_c_1660_n 0.00372978f $X=3.125 $Y=2.165
+ $X2=0 $Y2=0
cc_599 N_A_299_47#_M1012_g N_A_556_369#_c_1634_n 5.59945e-19 $X=3.125 $Y=2.165
+ $X2=0 $Y2=0
cc_600 N_A_299_47#_c_649_n N_A_556_369#_c_1634_n 0.00683182f $X=3.05 $Y=1.967
+ $X2=0 $Y2=0
cc_601 N_A_299_47#_c_641_n N_A_556_369#_c_1634_n 0.00221463f $X=3.135 $Y=1.86
+ $X2=0 $Y2=0
cc_602 N_A_299_47#_c_632_n N_VGND_c_1771_n 0.00268339f $X=1.625 $Y=0.38 $X2=0
+ $Y2=0
cc_603 N_A_299_47#_M1013_g N_VGND_c_1772_n 0.00857304f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_604 N_A_299_47#_c_632_n N_VGND_c_1783_n 0.0214549f $X=1.625 $Y=0.38 $X2=0
+ $Y2=0
cc_605 N_A_299_47#_M1013_g N_VGND_c_1784_n 0.0030886f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_606 N_A_299_47#_M1031_s N_VGND_c_1786_n 0.00186095f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_607 N_A_299_47#_M1013_g N_VGND_c_1786_n 0.00342951f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_608 N_A_299_47#_c_632_n N_VGND_c_1786_n 0.00629155f $X=1.625 $Y=0.38 $X2=0
+ $Y2=0
cc_609 N_D_M1014_g N_SCD_M1011_g 0.00211944f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_610 N_D_M1014_g N_A_193_47#_c_881_n 0.00392332f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_611 N_D_c_771_n N_A_193_47#_c_881_n 0.00255857f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_612 N_D_c_772_n N_A_193_47#_c_881_n 0.00699833f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_613 N_D_M1021_g N_VPWR_c_1472_n 0.00183225f $X=2.705 $Y=2.165 $X2=0 $Y2=0
cc_614 N_D_M1021_g N_VPWR_c_1485_n 0.00391499f $X=2.705 $Y=2.165 $X2=0 $Y2=0
cc_615 N_D_M1021_g N_VPWR_c_1470_n 0.00546297f $X=2.705 $Y=2.165 $X2=0 $Y2=0
cc_616 N_D_M1021_g N_A_556_369#_c_1637_n 0.00569061f $X=2.705 $Y=2.165 $X2=0
+ $Y2=0
cc_617 N_D_M1014_g N_VGND_c_1772_n 0.00144868f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_618 N_D_M1014_g N_VGND_c_1784_n 0.00422112f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_619 N_D_M1014_g N_VGND_c_1786_n 0.0056538f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_620 N_SCD_M1011_g N_A_193_47#_c_881_n 0.00245396f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_621 SCD N_A_193_47#_c_881_n 0.011855f $X=3.745 $Y=1.105 $X2=0 $Y2=0
cc_622 N_SCD_c_824_n N_VPWR_c_1473_n 0.00641619f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_623 N_SCD_c_824_n N_VPWR_c_1485_n 0.00419204f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_624 N_SCD_c_824_n N_VPWR_c_1470_n 0.00692748f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_625 N_SCD_c_824_n N_A_556_369#_c_1637_n 0.00465107f $X=3.6 $Y=1.77 $X2=0
+ $Y2=0
cc_626 N_SCD_M1011_g N_A_556_369#_c_1647_n 0.00475738f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_627 N_SCD_c_824_n N_A_556_369#_c_1660_n 0.00666112f $X=3.6 $Y=1.77 $X2=0
+ $Y2=0
cc_628 N_SCD_M1011_g N_A_556_369#_c_1628_n 0.00675657f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_629 N_SCD_c_824_n N_A_556_369#_c_1633_n 0.00958108f $X=3.6 $Y=1.77 $X2=0
+ $Y2=0
cc_630 N_SCD_c_825_n N_A_556_369#_c_1633_n 5.4464e-19 $X=3.665 $Y=1.52 $X2=0
+ $Y2=0
cc_631 SCD N_A_556_369#_c_1633_n 0.0302269f $X=3.745 $Y=1.105 $X2=0 $Y2=0
cc_632 N_SCD_c_824_n N_A_556_369#_c_1634_n 0.00237391f $X=3.6 $Y=1.77 $X2=0
+ $Y2=0
cc_633 SCD N_A_556_369#_c_1634_n 0.00193305f $X=3.745 $Y=1.105 $X2=0 $Y2=0
cc_634 N_SCD_M1011_g N_A_556_369#_c_1629_n 0.00756932f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_635 N_SCD_c_820_n N_A_556_369#_c_1629_n 7.71914e-19 $X=3.657 $Y=1.19 $X2=0
+ $Y2=0
cc_636 SCD N_A_556_369#_c_1629_n 0.0282592f $X=3.745 $Y=1.105 $X2=0 $Y2=0
cc_637 N_SCD_M1011_g N_A_556_369#_c_1630_n 0.00276697f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_638 SCD N_A_556_369#_c_1630_n 0.00392519f $X=3.745 $Y=1.105 $X2=0 $Y2=0
cc_639 N_SCD_M1011_g N_A_556_369#_c_1631_n 0.00271689f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_640 N_SCD_M1011_g N_A_556_369#_c_1632_n 0.00388747f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_641 N_SCD_c_820_n N_A_556_369#_c_1632_n 0.00135976f $X=3.657 $Y=1.19 $X2=0
+ $Y2=0
cc_642 N_SCD_c_823_n N_A_556_369#_c_1632_n 0.00327354f $X=3.6 $Y=1.715 $X2=0
+ $Y2=0
cc_643 N_SCD_c_824_n N_A_556_369#_c_1632_n 0.00107219f $X=3.6 $Y=1.77 $X2=0
+ $Y2=0
cc_644 SCD N_A_556_369#_c_1632_n 0.0451792f $X=3.745 $Y=1.105 $X2=0 $Y2=0
cc_645 N_SCD_c_824_n N_A_556_369#_c_1636_n 0.00283443f $X=3.6 $Y=1.77 $X2=0
+ $Y2=0
cc_646 N_SCD_M1011_g N_VGND_c_1773_n 0.00553893f $X=3.59 $Y=0.445 $X2=0 $Y2=0
cc_647 N_SCD_M1011_g N_VGND_c_1784_n 0.00399156f $X=3.59 $Y=0.445 $X2=0 $Y2=0
cc_648 N_SCD_M1011_g N_VGND_c_1786_n 0.00665835f $X=3.59 $Y=0.445 $X2=0 $Y2=0
cc_649 N_A_193_47#_c_880_n N_A_1092_183#_M1016_d 0.00133652f $X=6.94 $Y=0.87
+ $X2=-0.19 $Y2=-0.24
cc_650 N_A_193_47#_c_883_n N_A_1092_183#_M1016_d 0.00119173f $X=6.57 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_651 N_A_193_47#_c_885_n N_A_1092_183#_M1016_d 4.46878e-19 $X=6.715 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_652 N_A_193_47#_c_883_n N_A_1092_183#_M1007_g 0.00208483f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_653 N_A_193_47#_c_888_n N_A_1092_183#_M1007_g 0.013781f $X=5.015 $Y=0.705
+ $X2=0 $Y2=0
cc_654 N_A_193_47#_c_883_n N_A_1092_183#_c_1093_n 0.0221014f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_655 N_A_193_47#_c_885_n N_A_1092_183#_c_1119_n 8.64715e-19 $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_656 N_A_193_47#_c_880_n N_A_1092_183#_c_1120_n 0.00716698f $X=6.94 $Y=0.87
+ $X2=0 $Y2=0
cc_657 N_A_193_47#_c_883_n N_A_1092_183#_c_1120_n 0.00447852f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_658 N_A_193_47#_c_885_n N_A_1092_183#_c_1120_n 7.91937e-19 $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_659 N_A_193_47#_c_883_n N_A_1092_183#_c_1094_n 0.00899288f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_660 N_A_193_47#_c_877_n N_A_1092_183#_c_1095_n 0.00114045f $X=7.035 $Y=1.575
+ $X2=0 $Y2=0
cc_661 N_A_193_47#_c_880_n N_A_1092_183#_c_1095_n 0.0187533f $X=6.94 $Y=0.87
+ $X2=0 $Y2=0
cc_662 N_A_193_47#_c_883_n N_A_1092_183#_c_1095_n 0.0176435f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_663 N_A_193_47#_c_885_n N_A_1092_183#_c_1095_n 0.00179169f $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_664 N_A_193_47#_c_889_n N_A_1092_183#_c_1095_n 5.82389e-19 $X=6.895 $Y=0.87
+ $X2=0 $Y2=0
cc_665 N_A_193_47#_c_877_n N_A_1092_183#_c_1096_n 0.00620052f $X=7.035 $Y=1.575
+ $X2=0 $Y2=0
cc_666 N_A_193_47#_c_883_n N_A_1092_183#_c_1097_n 0.00299829f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_667 N_A_193_47#_c_886_n N_A_1092_183#_c_1097_n 0.0179412f $X=5.015 $Y=0.87
+ $X2=0 $Y2=0
cc_668 N_A_193_47#_c_877_n N_A_933_413#_c_1186_n 6.31337e-19 $X=7.035 $Y=1.575
+ $X2=0 $Y2=0
cc_669 N_A_193_47#_c_875_n N_A_933_413#_c_1187_n 0.00957285f $X=6.8 $Y=0.705
+ $X2=0 $Y2=0
cc_670 N_A_193_47#_c_880_n N_A_933_413#_c_1187_n 0.00100831f $X=6.94 $Y=0.87
+ $X2=0 $Y2=0
cc_671 N_A_193_47#_c_877_n N_A_933_413#_c_1188_n 3.37852e-19 $X=7.035 $Y=1.575
+ $X2=0 $Y2=0
cc_672 N_A_193_47#_c_889_n N_A_933_413#_c_1188_n 0.00957285f $X=6.895 $Y=0.87
+ $X2=0 $Y2=0
cc_673 N_A_193_47#_M1023_g N_A_933_413#_c_1204_n 0.00186646f $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_674 N_A_193_47#_c_876_n N_A_933_413#_c_1204_n 0.00286257f $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_675 N_A_193_47#_c_893_n N_A_933_413#_c_1204_n 6.94615e-19 $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_676 N_A_193_47#_c_879_n N_A_933_413#_c_1230_n 0.00356905f $X=4.76 $Y=0.87
+ $X2=0 $Y2=0
cc_677 N_A_193_47#_c_883_n N_A_933_413#_c_1230_n 0.00495571f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_678 N_A_193_47#_c_1017_p N_A_933_413#_c_1230_n 0.0011267f $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_679 N_A_193_47#_c_886_n N_A_933_413#_c_1230_n 0.00256542f $X=5.015 $Y=0.87
+ $X2=0 $Y2=0
cc_680 N_A_193_47#_c_887_n N_A_933_413#_c_1230_n 0.0204344f $X=5.015 $Y=0.87
+ $X2=0 $Y2=0
cc_681 N_A_193_47#_c_888_n N_A_933_413#_c_1230_n 0.00840911f $X=5.015 $Y=0.705
+ $X2=0 $Y2=0
cc_682 N_A_193_47#_c_876_n N_A_933_413#_c_1191_n 0.00979504f $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_683 N_A_193_47#_c_883_n N_A_933_413#_c_1191_n 0.0188221f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_684 N_A_193_47#_c_1017_p N_A_933_413#_c_1191_n 4.96697e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_685 N_A_193_47#_c_887_n N_A_933_413#_c_1191_n 0.0238568f $X=5.015 $Y=0.87
+ $X2=0 $Y2=0
cc_686 N_A_193_47#_c_888_n N_A_933_413#_c_1191_n 0.00604394f $X=5.015 $Y=0.705
+ $X2=0 $Y2=0
cc_687 N_A_193_47#_c_876_n N_A_933_413#_c_1192_n 0.00649323f $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_688 N_A_193_47#_c_883_n N_A_933_413#_c_1192_n 0.00803733f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_689 N_A_193_47#_M1019_g N_A_1520_315#_c_1306_n 0.0180347f $X=7.09 $Y=2.275
+ $X2=0 $Y2=0
cc_690 N_A_193_47#_c_896_n N_A_1520_315#_c_1306_n 0.0119764f $X=7.175 $Y=1.74
+ $X2=0 $Y2=0
cc_691 N_A_193_47#_M1019_g N_A_1349_413#_c_1394_n 0.00974744f $X=7.09 $Y=2.275
+ $X2=0 $Y2=0
cc_692 N_A_193_47#_c_895_n N_A_1349_413#_c_1394_n 0.012999f $X=7.175 $Y=1.74
+ $X2=0 $Y2=0
cc_693 N_A_193_47#_c_896_n N_A_1349_413#_c_1394_n 0.00300896f $X=7.175 $Y=1.74
+ $X2=0 $Y2=0
cc_694 N_A_193_47#_c_880_n N_A_1349_413#_c_1397_n 0.0153172f $X=6.94 $Y=0.87
+ $X2=0 $Y2=0
cc_695 N_A_193_47#_c_889_n N_A_1349_413#_c_1397_n 8.54271e-19 $X=6.895 $Y=0.87
+ $X2=0 $Y2=0
cc_696 N_A_193_47#_M1019_g N_A_1349_413#_c_1391_n 0.0046302f $X=7.09 $Y=2.275
+ $X2=0 $Y2=0
cc_697 N_A_193_47#_c_877_n N_A_1349_413#_c_1391_n 0.00868218f $X=7.035 $Y=1.575
+ $X2=0 $Y2=0
cc_698 N_A_193_47#_c_895_n N_A_1349_413#_c_1391_n 0.0246912f $X=7.175 $Y=1.74
+ $X2=0 $Y2=0
cc_699 N_A_193_47#_c_896_n N_A_1349_413#_c_1391_n 0.00187857f $X=7.175 $Y=1.74
+ $X2=0 $Y2=0
cc_700 N_A_193_47#_c_877_n N_A_1349_413#_c_1386_n 0.0272384f $X=7.035 $Y=1.575
+ $X2=0 $Y2=0
cc_701 N_A_193_47#_c_896_n N_A_1349_413#_c_1386_n 0.00102186f $X=7.175 $Y=1.74
+ $X2=0 $Y2=0
cc_702 N_A_193_47#_c_875_n N_A_1349_413#_c_1387_n 8.96907e-19 $X=6.8 $Y=0.705
+ $X2=0 $Y2=0
cc_703 N_A_193_47#_c_880_n N_A_1349_413#_c_1387_n 0.0255572f $X=6.94 $Y=0.87
+ $X2=0 $Y2=0
cc_704 N_A_193_47#_c_885_n N_A_1349_413#_c_1387_n 8.61155e-19 $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_705 N_A_193_47#_c_889_n N_A_1349_413#_c_1387_n 3.08898e-19 $X=6.895 $Y=0.87
+ $X2=0 $Y2=0
cc_706 N_A_193_47#_c_884_n N_VPWR_c_1471_n 0.012732f $X=1.125 $Y=0.85 $X2=0
+ $Y2=0
cc_707 N_A_193_47#_c_884_n N_VPWR_c_1472_n 5.34357e-19 $X=1.125 $Y=0.85 $X2=0
+ $Y2=0
cc_708 N_A_193_47#_M1023_g N_VPWR_c_1473_n 0.00275573f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_709 N_A_193_47#_M1023_g N_VPWR_c_1477_n 0.005785f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_710 N_A_193_47#_M1019_g N_VPWR_c_1479_n 0.00383564f $X=7.09 $Y=2.275 $X2=0
+ $Y2=0
cc_711 N_A_193_47#_c_884_n N_VPWR_c_1484_n 0.0149126f $X=1.125 $Y=0.85 $X2=0
+ $Y2=0
cc_712 N_A_193_47#_M1023_g N_VPWR_c_1470_n 0.00734982f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_713 N_A_193_47#_M1019_g N_VPWR_c_1470_n 0.00579176f $X=7.09 $Y=2.275 $X2=0
+ $Y2=0
cc_714 N_A_193_47#_c_876_n N_VPWR_c_1470_n 0.00189161f $X=4.605 $Y=1.74 $X2=0
+ $Y2=0
cc_715 N_A_193_47#_c_893_n N_VPWR_c_1470_n 4.15345e-19 $X=4.605 $Y=1.74 $X2=0
+ $Y2=0
cc_716 N_A_193_47#_c_884_n N_VPWR_c_1470_n 0.00381577f $X=1.125 $Y=0.85 $X2=0
+ $Y2=0
cc_717 N_A_193_47#_c_881_n N_A_556_369#_c_1647_n 0.00542704f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_718 N_A_193_47#_c_881_n N_A_556_369#_c_1629_n 0.0215404f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_719 N_A_193_47#_c_881_n N_A_556_369#_c_1630_n 0.00999898f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_720 N_A_193_47#_c_879_n N_A_556_369#_c_1631_n 0.0114096f $X=4.76 $Y=0.87
+ $X2=0 $Y2=0
cc_721 N_A_193_47#_c_881_n N_A_556_369#_c_1631_n 0.0115743f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_722 N_A_193_47#_c_1017_p N_A_556_369#_c_1631_n 3.33018e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_723 N_A_193_47#_c_876_n N_A_556_369#_c_1632_n 0.0585452f $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_724 N_A_193_47#_c_893_n N_A_556_369#_c_1632_n 0.0052844f $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_725 N_A_193_47#_c_879_n N_A_556_369#_c_1632_n 0.0112291f $X=4.76 $Y=0.87
+ $X2=0 $Y2=0
cc_726 N_A_193_47#_c_881_n N_A_556_369#_c_1632_n 0.011116f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_727 N_A_193_47#_c_1017_p N_A_556_369#_c_1632_n 2.28604e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_728 N_A_193_47#_M1023_g N_A_556_369#_c_1636_n 0.00999238f $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_729 N_A_193_47#_c_876_n N_A_556_369#_c_1636_n 0.00558861f $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_730 N_A_193_47#_c_893_n N_A_556_369#_c_1636_n 9.82843e-19 $X=4.605 $Y=1.74
+ $X2=0 $Y2=0
cc_731 N_A_193_47#_c_881_n N_VGND_c_1772_n 0.00122509f $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_732 N_A_193_47#_c_881_n N_VGND_c_1773_n 9.19202e-19 $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_733 N_A_193_47#_c_879_n N_VGND_c_1774_n 0.00114596f $X=4.76 $Y=0.87 $X2=0
+ $Y2=0
cc_734 N_A_193_47#_c_888_n N_VGND_c_1774_n 0.0037981f $X=5.015 $Y=0.705 $X2=0
+ $Y2=0
cc_735 N_A_193_47#_c_883_n N_VGND_c_1775_n 0.00197288f $X=6.57 $Y=0.85 $X2=0
+ $Y2=0
cc_736 N_A_193_47#_c_875_n N_VGND_c_1778_n 0.00435108f $X=6.8 $Y=0.705 $X2=0
+ $Y2=0
cc_737 N_A_193_47#_c_880_n N_VGND_c_1778_n 0.00341023f $X=6.94 $Y=0.87 $X2=0
+ $Y2=0
cc_738 N_A_193_47#_c_889_n N_VGND_c_1778_n 8.04624e-19 $X=6.895 $Y=0.87 $X2=0
+ $Y2=0
cc_739 N_A_193_47#_c_878_n N_VGND_c_1783_n 0.00933042f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_740 N_A_193_47#_M1015_d N_VGND_c_1786_n 0.0025245f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_741 N_A_193_47#_c_875_n N_VGND_c_1786_n 0.00615106f $X=6.8 $Y=0.705 $X2=0
+ $Y2=0
cc_742 N_A_193_47#_c_878_n N_VGND_c_1786_n 0.00355905f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_743 N_A_193_47#_c_879_n N_VGND_c_1786_n 0.00249883f $X=4.76 $Y=0.87 $X2=0
+ $Y2=0
cc_744 N_A_193_47#_c_880_n N_VGND_c_1786_n 0.00363841f $X=6.94 $Y=0.87 $X2=0
+ $Y2=0
cc_745 N_A_193_47#_c_881_n N_VGND_c_1786_n 0.157258f $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_746 N_A_193_47#_c_882_n N_VGND_c_1786_n 0.0152176f $X=1.27 $Y=0.85 $X2=0
+ $Y2=0
cc_747 N_A_193_47#_c_883_n N_VGND_c_1786_n 0.0733748f $X=6.57 $Y=0.85 $X2=0
+ $Y2=0
cc_748 N_A_193_47#_c_1017_p N_VGND_c_1786_n 0.0146f $X=4.975 $Y=0.85 $X2=0 $Y2=0
cc_749 N_A_193_47#_c_885_n N_VGND_c_1786_n 0.0146166f $X=6.715 $Y=0.85 $X2=0
+ $Y2=0
cc_750 N_A_193_47#_c_888_n N_VGND_c_1786_n 0.00563926f $X=5.015 $Y=0.705 $X2=0
+ $Y2=0
cc_751 N_A_193_47#_c_889_n N_VGND_c_1786_n 0.00134095f $X=6.895 $Y=0.87 $X2=0
+ $Y2=0
cc_752 N_A_1092_183#_c_1096_n N_A_933_413#_c_1186_n 0.00595764f $X=6.365
+ $Y=2.135 $X2=0 $Y2=0
cc_753 N_A_1092_183#_M1022_g N_A_933_413#_M1008_g 0.0139082f $X=5.535 $Y=2.275
+ $X2=0 $Y2=0
cc_754 N_A_1092_183#_c_1107_n N_A_933_413#_M1008_g 0.00378805f $X=6.405 $Y=2.3
+ $X2=0 $Y2=0
cc_755 N_A_1092_183#_c_1096_n N_A_933_413#_M1008_g 0.0122998f $X=6.365 $Y=2.135
+ $X2=0 $Y2=0
cc_756 N_A_1092_183#_M1007_g N_A_933_413#_c_1187_n 0.0109128f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_757 N_A_1092_183#_c_1093_n N_A_933_413#_c_1187_n 0.00351053f $X=6.24 $Y=0.915
+ $X2=0 $Y2=0
cc_758 N_A_1092_183#_c_1119_n N_A_933_413#_c_1187_n 0.00675936f $X=6.325
+ $Y=0.765 $X2=0 $Y2=0
cc_759 N_A_1092_183#_c_1139_p N_A_933_413#_c_1187_n 0.004701f $X=6.41 $Y=0.45
+ $X2=0 $Y2=0
cc_760 N_A_1092_183#_c_1095_n N_A_933_413#_c_1187_n 0.00333126f $X=6.325
+ $Y=0.915 $X2=0 $Y2=0
cc_761 N_A_1092_183#_c_1097_n N_A_933_413#_c_1187_n 0.00500517f $X=5.565 $Y=0.93
+ $X2=0 $Y2=0
cc_762 N_A_1092_183#_M1022_g N_A_933_413#_c_1188_n 0.00398999f $X=5.535 $Y=2.275
+ $X2=0 $Y2=0
cc_763 N_A_1092_183#_c_1093_n N_A_933_413#_c_1188_n 0.00996228f $X=6.24 $Y=0.915
+ $X2=0 $Y2=0
cc_764 N_A_1092_183#_c_1094_n N_A_933_413#_c_1188_n 2.46578e-19 $X=5.78 $Y=0.93
+ $X2=0 $Y2=0
cc_765 N_A_1092_183#_c_1095_n N_A_933_413#_c_1188_n 0.00234347f $X=6.325
+ $Y=0.915 $X2=0 $Y2=0
cc_766 N_A_1092_183#_c_1096_n N_A_933_413#_c_1188_n 0.00394884f $X=6.365
+ $Y=2.135 $X2=0 $Y2=0
cc_767 N_A_1092_183#_c_1097_n N_A_933_413#_c_1188_n 0.00573363f $X=5.565 $Y=0.93
+ $X2=0 $Y2=0
cc_768 N_A_1092_183#_M1022_g N_A_933_413#_c_1189_n 0.0173592f $X=5.535 $Y=2.275
+ $X2=0 $Y2=0
cc_769 N_A_1092_183#_c_1093_n N_A_933_413#_c_1189_n 0.00400764f $X=6.24 $Y=0.915
+ $X2=0 $Y2=0
cc_770 N_A_1092_183#_c_1097_n N_A_933_413#_c_1189_n 0.00238133f $X=5.565 $Y=0.93
+ $X2=0 $Y2=0
cc_771 N_A_1092_183#_c_1096_n N_A_933_413#_c_1190_n 0.00611615f $X=6.365
+ $Y=2.135 $X2=0 $Y2=0
cc_772 N_A_1092_183#_M1022_g N_A_933_413#_c_1204_n 0.0101048f $X=5.535 $Y=2.275
+ $X2=0 $Y2=0
cc_773 N_A_1092_183#_M1007_g N_A_933_413#_c_1191_n 0.00441151f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_774 N_A_1092_183#_c_1094_n N_A_933_413#_c_1191_n 0.0243525f $X=5.78 $Y=0.93
+ $X2=0 $Y2=0
cc_775 N_A_1092_183#_c_1097_n N_A_933_413#_c_1191_n 0.0095167f $X=5.565 $Y=0.93
+ $X2=0 $Y2=0
cc_776 N_A_1092_183#_M1022_g N_A_933_413#_c_1196_n 0.0153761f $X=5.535 $Y=2.275
+ $X2=0 $Y2=0
cc_777 N_A_1092_183#_c_1096_n N_A_933_413#_c_1196_n 0.00754007f $X=6.365
+ $Y=2.135 $X2=0 $Y2=0
cc_778 N_A_1092_183#_M1022_g N_A_933_413#_c_1192_n 0.0138593f $X=5.535 $Y=2.275
+ $X2=0 $Y2=0
cc_779 N_A_1092_183#_c_1093_n N_A_933_413#_c_1192_n 0.0186614f $X=6.24 $Y=0.915
+ $X2=0 $Y2=0
cc_780 N_A_1092_183#_c_1094_n N_A_933_413#_c_1192_n 0.0112018f $X=5.78 $Y=0.93
+ $X2=0 $Y2=0
cc_781 N_A_1092_183#_c_1096_n N_A_933_413#_c_1192_n 0.0245884f $X=6.365 $Y=2.135
+ $X2=0 $Y2=0
cc_782 N_A_1092_183#_c_1097_n N_A_933_413#_c_1192_n 0.00213749f $X=5.565 $Y=0.93
+ $X2=0 $Y2=0
cc_783 N_A_1092_183#_c_1107_n N_A_1349_413#_c_1394_n 0.0109209f $X=6.405 $Y=2.3
+ $X2=0 $Y2=0
cc_784 N_A_1092_183#_M1022_g N_VPWR_c_1474_n 0.0057281f $X=5.535 $Y=2.275 $X2=0
+ $Y2=0
cc_785 N_A_1092_183#_c_1096_n N_VPWR_c_1474_n 0.0237f $X=6.365 $Y=2.135 $X2=0
+ $Y2=0
cc_786 N_A_1092_183#_M1022_g N_VPWR_c_1477_n 0.00378797f $X=5.535 $Y=2.275 $X2=0
+ $Y2=0
cc_787 N_A_1092_183#_c_1107_n N_VPWR_c_1479_n 0.015079f $X=6.405 $Y=2.3 $X2=0
+ $Y2=0
cc_788 N_A_1092_183#_M1008_d N_VPWR_c_1470_n 0.00285154f $X=6.27 $Y=1.735 $X2=0
+ $Y2=0
cc_789 N_A_1092_183#_M1022_g N_VPWR_c_1470_n 0.00596544f $X=5.535 $Y=2.275 $X2=0
+ $Y2=0
cc_790 N_A_1092_183#_c_1107_n N_VPWR_c_1470_n 0.00439826f $X=6.405 $Y=2.3 $X2=0
+ $Y2=0
cc_791 N_A_1092_183#_c_1093_n N_VGND_M1007_d 0.00306998f $X=6.24 $Y=0.915 $X2=0
+ $Y2=0
cc_792 N_A_1092_183#_M1007_g N_VGND_c_1774_n 0.00585385f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_793 N_A_1092_183#_M1007_g N_VGND_c_1775_n 0.00603751f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_794 N_A_1092_183#_c_1119_n N_VGND_c_1775_n 0.00354103f $X=6.325 $Y=0.765
+ $X2=0 $Y2=0
cc_795 N_A_1092_183#_c_1139_p N_VGND_c_1775_n 0.013122f $X=6.41 $Y=0.45 $X2=0
+ $Y2=0
cc_796 N_A_1092_183#_c_1094_n N_VGND_c_1775_n 0.0258565f $X=5.78 $Y=0.93 $X2=0
+ $Y2=0
cc_797 N_A_1092_183#_c_1097_n N_VGND_c_1775_n 0.00122075f $X=5.565 $Y=0.93 $X2=0
+ $Y2=0
cc_798 N_A_1092_183#_c_1139_p N_VGND_c_1778_n 0.00594819f $X=6.41 $Y=0.45 $X2=0
+ $Y2=0
cc_799 N_A_1092_183#_c_1120_n N_VGND_c_1778_n 0.0100275f $X=6.535 $Y=0.45 $X2=0
+ $Y2=0
cc_800 N_A_1092_183#_M1016_d N_VGND_c_1786_n 0.0024731f $X=6.37 $Y=0.235 $X2=0
+ $Y2=0
cc_801 N_A_1092_183#_M1007_g N_VGND_c_1786_n 0.0070154f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_802 N_A_1092_183#_c_1093_n N_VGND_c_1786_n 0.0042145f $X=6.24 $Y=0.915 $X2=0
+ $Y2=0
cc_803 N_A_1092_183#_c_1139_p N_VGND_c_1786_n 0.00261981f $X=6.41 $Y=0.45 $X2=0
+ $Y2=0
cc_804 N_A_1092_183#_c_1120_n N_VGND_c_1786_n 0.00443994f $X=6.535 $Y=0.45 $X2=0
+ $Y2=0
cc_805 N_A_1092_183#_c_1094_n N_VGND_c_1786_n 0.00269026f $X=5.78 $Y=0.93 $X2=0
+ $Y2=0
cc_806 N_A_933_413#_c_1204_n N_VPWR_M1022_d 0.00236303f $X=5.56 $Y=2.275 $X2=0
+ $Y2=0
cc_807 N_A_933_413#_c_1196_n N_VPWR_M1022_d 0.00412006f $X=5.645 $Y=2.19 $X2=0
+ $Y2=0
cc_808 N_A_933_413#_M1008_g N_VPWR_c_1474_n 0.00314007f $X=6.195 $Y=2.11 $X2=0
+ $Y2=0
cc_809 N_A_933_413#_c_1189_n N_VPWR_c_1474_n 9.53331e-19 $X=6.12 $Y=1.41 $X2=0
+ $Y2=0
cc_810 N_A_933_413#_c_1204_n N_VPWR_c_1474_n 0.0138309f $X=5.56 $Y=2.275 $X2=0
+ $Y2=0
cc_811 N_A_933_413#_c_1196_n N_VPWR_c_1474_n 0.025225f $X=5.645 $Y=2.19 $X2=0
+ $Y2=0
cc_812 N_A_933_413#_c_1192_n N_VPWR_c_1474_n 0.00741701f $X=5.645 $Y=1.41 $X2=0
+ $Y2=0
cc_813 N_A_933_413#_c_1204_n N_VPWR_c_1477_n 0.0359536f $X=5.56 $Y=2.275 $X2=0
+ $Y2=0
cc_814 N_A_933_413#_M1008_g N_VPWR_c_1479_n 0.00541359f $X=6.195 $Y=2.11 $X2=0
+ $Y2=0
cc_815 N_A_933_413#_M1023_d N_VPWR_c_1470_n 0.00217001f $X=4.665 $Y=2.065 $X2=0
+ $Y2=0
cc_816 N_A_933_413#_M1008_g N_VPWR_c_1470_n 0.00665748f $X=6.195 $Y=2.11 $X2=0
+ $Y2=0
cc_817 N_A_933_413#_c_1204_n N_VPWR_c_1470_n 0.0161651f $X=5.56 $Y=2.275 $X2=0
+ $Y2=0
cc_818 N_A_933_413#_c_1204_n N_A_556_369#_c_1636_n 0.0104003f $X=5.56 $Y=2.275
+ $X2=0 $Y2=0
cc_819 N_A_933_413#_c_1204_n A_1026_413# 0.0045944f $X=5.56 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_820 N_A_933_413#_c_1230_n N_VGND_c_1774_n 0.0255873f $X=5.27 $Y=0.45 $X2=0
+ $Y2=0
cc_821 N_A_933_413#_c_1187_n N_VGND_c_1775_n 0.00816054f $X=6.295 $Y=0.95 $X2=0
+ $Y2=0
cc_822 N_A_933_413#_c_1187_n N_VGND_c_1778_n 0.00407056f $X=6.295 $Y=0.95 $X2=0
+ $Y2=0
cc_823 N_A_933_413#_M1030_d N_VGND_c_1786_n 0.00228029f $X=4.67 $Y=0.235 $X2=0
+ $Y2=0
cc_824 N_A_933_413#_c_1187_n N_VGND_c_1786_n 0.00620172f $X=6.295 $Y=0.95 $X2=0
+ $Y2=0
cc_825 N_A_933_413#_c_1230_n N_VGND_c_1786_n 0.0113042f $X=5.27 $Y=0.45 $X2=0
+ $Y2=0
cc_826 N_A_933_413#_c_1230_n A_1030_47# 0.00455507f $X=5.27 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_827 N_A_933_413#_c_1191_n A_1030_47# 0.00200718f $X=5.355 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_828 N_A_1520_315#_c_1297_n N_A_1349_413#_c_1382_n 0.00505396f $X=8.62
+ $Y=0.995 $X2=0 $Y2=0
cc_829 N_A_1520_315#_c_1300_n N_A_1349_413#_c_1382_n 0.00768498f $X=8.52
+ $Y=0.385 $X2=0 $Y2=0
cc_830 N_A_1520_315#_c_1301_n N_A_1349_413#_c_1382_n 0.0193264f $X=9.175
+ $Y=0.995 $X2=0 $Y2=0
cc_831 N_A_1520_315#_M1024_g N_A_1349_413#_M1020_g 0.0196432f $X=9.185 $Y=1.985
+ $X2=0 $Y2=0
cc_832 N_A_1520_315#_c_1306_n N_A_1349_413#_M1020_g 0.00198604f $X=7.855 $Y=1.74
+ $X2=0 $Y2=0
cc_833 N_A_1520_315#_c_1318_p N_A_1349_413#_M1020_g 0.0104955f $X=8.52 $Y=2.29
+ $X2=0 $Y2=0
cc_834 N_A_1520_315#_c_1307_n N_A_1349_413#_M1020_g 0.00742753f $X=8.62 $Y=1.575
+ $X2=0 $Y2=0
cc_835 N_A_1520_315#_c_1320_p N_A_1349_413#_M1020_g 0.00489897f $X=8.52 $Y=1.68
+ $X2=0 $Y2=0
cc_836 N_A_1520_315#_M1017_g N_A_1349_413#_c_1383_n 0.0149936f $X=7.79 $Y=0.445
+ $X2=0 $Y2=0
cc_837 N_A_1520_315#_c_1305_n N_A_1349_413#_c_1383_n 0.00734699f $X=8.435
+ $Y=1.74 $X2=0 $Y2=0
cc_838 N_A_1520_315#_c_1300_n N_A_1349_413#_c_1383_n 0.00747686f $X=8.52
+ $Y=0.385 $X2=0 $Y2=0
cc_839 N_A_1520_315#_c_1320_p N_A_1349_413#_c_1383_n 0.00407845f $X=8.52 $Y=1.68
+ $X2=0 $Y2=0
cc_840 N_A_1520_315#_c_1325_p N_A_1349_413#_c_1383_n 0.01406f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_841 N_A_1520_315#_c_1298_n N_A_1349_413#_c_1384_n 0.0155195f $X=9.15 $Y=1.16
+ $X2=0 $Y2=0
cc_842 N_A_1520_315#_c_1299_n N_A_1349_413#_c_1384_n 0.0215061f $X=9.15 $Y=1.16
+ $X2=0 $Y2=0
cc_843 N_A_1520_315#_c_1325_p N_A_1349_413#_c_1384_n 0.00155371f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_844 N_A_1520_315#_M1001_g N_A_1349_413#_c_1394_n 0.0019846f $X=7.675 $Y=2.275
+ $X2=0 $Y2=0
cc_845 N_A_1520_315#_M1017_g N_A_1349_413#_c_1397_n 0.00114979f $X=7.79 $Y=0.445
+ $X2=0 $Y2=0
cc_846 N_A_1520_315#_c_1305_n N_A_1349_413#_c_1391_n 0.0262086f $X=8.435 $Y=1.74
+ $X2=0 $Y2=0
cc_847 N_A_1520_315#_c_1306_n N_A_1349_413#_c_1391_n 0.00865902f $X=7.855
+ $Y=1.74 $X2=0 $Y2=0
cc_848 N_A_1520_315#_M1017_g N_A_1349_413#_c_1385_n 0.018366f $X=7.79 $Y=0.445
+ $X2=0 $Y2=0
cc_849 N_A_1520_315#_c_1305_n N_A_1349_413#_c_1385_n 0.0355898f $X=8.435 $Y=1.74
+ $X2=0 $Y2=0
cc_850 N_A_1520_315#_c_1306_n N_A_1349_413#_c_1385_n 0.00739167f $X=7.855
+ $Y=1.74 $X2=0 $Y2=0
cc_851 N_A_1520_315#_c_1300_n N_A_1349_413#_c_1385_n 7.42989e-19 $X=8.52
+ $Y=0.385 $X2=0 $Y2=0
cc_852 N_A_1520_315#_c_1325_p N_A_1349_413#_c_1385_n 0.0278269f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_853 N_A_1520_315#_M1017_g N_A_1349_413#_c_1386_n 0.00880678f $X=7.79 $Y=0.445
+ $X2=0 $Y2=0
cc_854 N_A_1520_315#_M1017_g N_A_1349_413#_c_1387_n 0.00779225f $X=7.79 $Y=0.445
+ $X2=0 $Y2=0
cc_855 N_A_1520_315#_M1001_g N_VPWR_c_1475_n 0.0114377f $X=7.675 $Y=2.275 $X2=0
+ $Y2=0
cc_856 N_A_1520_315#_c_1305_n N_VPWR_c_1475_n 0.0186057f $X=8.435 $Y=1.74 $X2=0
+ $Y2=0
cc_857 N_A_1520_315#_c_1306_n N_VPWR_c_1475_n 0.00469579f $X=7.855 $Y=1.74 $X2=0
+ $Y2=0
cc_858 N_A_1520_315#_c_1318_p N_VPWR_c_1475_n 0.0151041f $X=8.52 $Y=2.29 $X2=0
+ $Y2=0
cc_859 N_A_1520_315#_M1024_g N_VPWR_c_1476_n 0.00711113f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_860 N_A_1520_315#_c_1318_p N_VPWR_c_1476_n 0.0399488f $X=8.52 $Y=2.29 $X2=0
+ $Y2=0
cc_861 N_A_1520_315#_c_1298_n N_VPWR_c_1476_n 0.00956157f $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_862 N_A_1520_315#_c_1299_n N_VPWR_c_1476_n 6.26814e-19 $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_863 N_A_1520_315#_c_1320_p N_VPWR_c_1476_n 0.0220075f $X=8.52 $Y=1.68 $X2=0
+ $Y2=0
cc_864 N_A_1520_315#_M1001_g N_VPWR_c_1479_n 0.00585385f $X=7.675 $Y=2.275 $X2=0
+ $Y2=0
cc_865 N_A_1520_315#_c_1318_p N_VPWR_c_1481_n 0.0157187f $X=8.52 $Y=2.29 $X2=0
+ $Y2=0
cc_866 N_A_1520_315#_M1024_g N_VPWR_c_1486_n 0.0054411f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_867 N_A_1520_315#_M1020_s N_VPWR_c_1470_n 0.00234057f $X=8.395 $Y=1.485 $X2=0
+ $Y2=0
cc_868 N_A_1520_315#_M1001_g N_VPWR_c_1470_n 0.012435f $X=7.675 $Y=2.275 $X2=0
+ $Y2=0
cc_869 N_A_1520_315#_M1024_g N_VPWR_c_1470_n 0.0106959f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_870 N_A_1520_315#_c_1305_n N_VPWR_c_1470_n 0.0145003f $X=8.435 $Y=1.74 $X2=0
+ $Y2=0
cc_871 N_A_1520_315#_c_1306_n N_VPWR_c_1470_n 0.00103388f $X=7.855 $Y=1.74 $X2=0
+ $Y2=0
cc_872 N_A_1520_315#_c_1318_p N_VPWR_c_1470_n 0.00997475f $X=8.52 $Y=2.29 $X2=0
+ $Y2=0
cc_873 N_A_1520_315#_M1024_g N_Q_c_1746_n 0.00415546f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_874 N_A_1520_315#_c_1307_n N_Q_c_1746_n 0.00198007f $X=8.62 $Y=1.575 $X2=0
+ $Y2=0
cc_875 N_A_1520_315#_c_1299_n N_Q_c_1746_n 0.00193312f $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_876 N_A_1520_315#_c_1320_p N_Q_c_1746_n 0.00158627f $X=8.52 $Y=1.68 $X2=0
+ $Y2=0
cc_877 N_A_1520_315#_M1024_g N_Q_c_1744_n 0.00455553f $X=9.185 $Y=1.985 $X2=0
+ $Y2=0
cc_878 N_A_1520_315#_c_1298_n N_Q_c_1744_n 0.0262705f $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_879 N_A_1520_315#_c_1299_n N_Q_c_1744_n 0.00830784f $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_880 N_A_1520_315#_c_1301_n N_Q_c_1744_n 0.00411924f $X=9.175 $Y=0.995 $X2=0
+ $Y2=0
cc_881 N_A_1520_315#_M1024_g Q 0.00809632f $X=9.185 $Y=1.985 $X2=0 $Y2=0
cc_882 N_A_1520_315#_c_1299_n N_Q_c_1745_n 0.00191171f $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_883 N_A_1520_315#_c_1300_n N_Q_c_1745_n 0.00375716f $X=8.52 $Y=0.385 $X2=0
+ $Y2=0
cc_884 N_A_1520_315#_c_1301_n N_Q_c_1745_n 0.00816502f $X=9.175 $Y=0.995 $X2=0
+ $Y2=0
cc_885 N_A_1520_315#_M1017_g N_VGND_c_1776_n 0.0215676f $X=7.79 $Y=0.445 $X2=0
+ $Y2=0
cc_886 N_A_1520_315#_c_1300_n N_VGND_c_1776_n 0.0187345f $X=8.52 $Y=0.385 $X2=0
+ $Y2=0
cc_887 N_A_1520_315#_c_1298_n N_VGND_c_1777_n 0.00956157f $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_888 N_A_1520_315#_c_1299_n N_VGND_c_1777_n 6.26814e-19 $X=9.15 $Y=1.16 $X2=0
+ $Y2=0
cc_889 N_A_1520_315#_c_1300_n N_VGND_c_1777_n 0.0292994f $X=8.52 $Y=0.385 $X2=0
+ $Y2=0
cc_890 N_A_1520_315#_c_1301_n N_VGND_c_1777_n 0.00556109f $X=9.175 $Y=0.995
+ $X2=0 $Y2=0
cc_891 N_A_1520_315#_c_1300_n N_VGND_c_1780_n 0.0172098f $X=8.52 $Y=0.385 $X2=0
+ $Y2=0
cc_892 N_A_1520_315#_c_1301_n N_VGND_c_1785_n 0.00543342f $X=9.175 $Y=0.995
+ $X2=0 $Y2=0
cc_893 N_A_1520_315#_M1004_s N_VGND_c_1786_n 0.00212021f $X=8.395 $Y=0.235 $X2=0
+ $Y2=0
cc_894 N_A_1520_315#_M1017_g N_VGND_c_1786_n 9.61436e-19 $X=7.79 $Y=0.445 $X2=0
+ $Y2=0
cc_895 N_A_1520_315#_c_1300_n N_VGND_c_1786_n 0.0127495f $X=8.52 $Y=0.385 $X2=0
+ $Y2=0
cc_896 N_A_1520_315#_c_1301_n N_VGND_c_1786_n 0.010693f $X=9.175 $Y=0.995 $X2=0
+ $Y2=0
cc_897 N_A_1349_413#_M1020_g N_VPWR_c_1475_n 0.00220635f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_898 N_A_1349_413#_M1020_g N_VPWR_c_1476_n 0.00587825f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_899 N_A_1349_413#_c_1394_n N_VPWR_c_1479_n 0.0273845f $X=7.43 $Y=2.25 $X2=0
+ $Y2=0
cc_900 N_A_1349_413#_M1020_g N_VPWR_c_1481_n 0.00511679f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_901 N_A_1349_413#_M1026_d N_VPWR_c_1470_n 0.00219484f $X=6.745 $Y=2.065 $X2=0
+ $Y2=0
cc_902 N_A_1349_413#_M1020_g N_VPWR_c_1470_n 0.0103298f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_903 N_A_1349_413#_c_1394_n N_VPWR_c_1470_n 0.0276628f $X=7.43 $Y=2.25 $X2=0
+ $Y2=0
cc_904 N_A_1349_413#_c_1394_n A_1433_413# 0.0105858f $X=7.43 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_905 N_A_1349_413#_c_1391_n A_1433_413# 0.00184879f $X=7.515 $Y=2.165
+ $X2=-0.19 $Y2=-0.24
cc_906 N_A_1349_413#_M1020_g N_Q_c_1746_n 5.14267e-19 $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_907 N_A_1349_413#_c_1382_n N_Q_c_1745_n 4.19418e-19 $X=8.73 $Y=0.995 $X2=0
+ $Y2=0
cc_908 N_A_1349_413#_c_1382_n N_VGND_c_1776_n 0.00268732f $X=8.73 $Y=0.995 $X2=0
+ $Y2=0
cc_909 N_A_1349_413#_c_1397_n N_VGND_c_1776_n 0.0104892f $X=7.3 $Y=0.45 $X2=0
+ $Y2=0
cc_910 N_A_1349_413#_c_1385_n N_VGND_c_1776_n 0.0154767f $X=8.28 $Y=1.16 $X2=0
+ $Y2=0
cc_911 N_A_1349_413#_c_1387_n N_VGND_c_1776_n 0.00447237f $X=7.45 $Y=0.995 $X2=0
+ $Y2=0
cc_912 N_A_1349_413#_c_1382_n N_VGND_c_1777_n 0.00534404f $X=8.73 $Y=0.995 $X2=0
+ $Y2=0
cc_913 N_A_1349_413#_c_1397_n N_VGND_c_1778_n 0.0184388f $X=7.3 $Y=0.45 $X2=0
+ $Y2=0
cc_914 N_A_1349_413#_c_1382_n N_VGND_c_1780_n 0.00514019f $X=8.73 $Y=0.995 $X2=0
+ $Y2=0
cc_915 N_A_1349_413#_M1002_d N_VGND_c_1786_n 0.00333348f $X=6.875 $Y=0.235 $X2=0
+ $Y2=0
cc_916 N_A_1349_413#_c_1382_n N_VGND_c_1786_n 0.0103347f $X=8.73 $Y=0.995 $X2=0
+ $Y2=0
cc_917 N_A_1349_413#_c_1397_n N_VGND_c_1786_n 0.0182474f $X=7.3 $Y=0.45 $X2=0
+ $Y2=0
cc_918 N_A_1349_413#_c_1397_n A_1478_47# 0.00201232f $X=7.3 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_919 N_A_1349_413#_c_1387_n A_1478_47# 0.00127737f $X=7.45 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_920 N_VPWR_c_1470_n A_467_369# 0.00261295f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_921 N_VPWR_c_1470_n N_A_556_369#_M1021_d 0.00179277f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1470_n N_A_556_369#_M1023_s 0.00262146f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1472_n N_A_556_369#_c_1637_n 0.00574717f $X=2.045 $Y=2.33 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1473_n N_A_556_369#_c_1637_n 0.0134906f $X=3.815 $Y=2.33 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1485_n N_A_556_369#_c_1637_n 0.0371081f $X=3.73 $Y=2.72 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1470_n N_A_556_369#_c_1637_n 0.013847f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1473_n N_A_556_369#_c_1660_n 0.00564282f $X=3.815 $Y=2.33 $X2=0
+ $Y2=0
cc_928 N_VPWR_M1009_d N_A_556_369#_c_1633_n 0.00303203f $X=3.67 $Y=1.845 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1473_n N_A_556_369#_c_1633_n 0.0136785f $X=3.815 $Y=2.33 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1477_n N_A_556_369#_c_1633_n 0.00385977f $X=5.9 $Y=2.72 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1485_n N_A_556_369#_c_1633_n 0.00194486f $X=3.73 $Y=2.72 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1470_n N_A_556_369#_c_1633_n 0.00501574f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1473_n N_A_556_369#_c_1636_n 0.0158431f $X=3.815 $Y=2.33 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1477_n N_A_556_369#_c_1636_n 0.0143719f $X=5.9 $Y=2.72 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1470_n N_A_556_369#_c_1636_n 0.004301f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_936 N_VPWR_c_1470_n A_640_369# 0.00214028f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_937 N_VPWR_c_1470_n A_1026_413# 0.00220276f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_938 N_VPWR_c_1470_n A_1433_413# 0.00377587f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_939 N_VPWR_c_1470_n N_Q_M1024_d 0.00214872f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_940 N_VPWR_c_1476_n N_Q_c_1746_n 0.0534068f $X=8.96 $Y=1.79 $X2=0 $Y2=0
cc_941 N_VPWR_c_1486_n Q 0.0152684f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_942 N_VPWR_c_1470_n Q 0.0125286f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_943 N_A_556_369#_c_1637_n A_640_369# 0.00372468f $X=3.39 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_944 N_A_556_369#_c_1660_n A_640_369# 0.0026432f $X=3.475 $Y=2.245 $X2=-0.19
+ $Y2=-0.24
cc_945 N_A_556_369#_c_1634_n A_640_369# 9.23695e-19 $X=3.56 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_946 N_A_556_369#_c_1647_n N_VGND_c_1773_n 0.0135147f $X=3.42 $Y=0.36 $X2=0
+ $Y2=0
cc_947 N_A_556_369#_c_1628_n N_VGND_c_1773_n 0.00707612f $X=3.505 $Y=0.715 $X2=0
+ $Y2=0
cc_948 N_A_556_369#_c_1629_n N_VGND_c_1773_n 0.0142754f $X=4.18 $Y=0.8 $X2=0
+ $Y2=0
cc_949 N_A_556_369#_c_1631_n N_VGND_c_1773_n 0.0168771f $X=4.265 $Y=0.885 $X2=0
+ $Y2=0
cc_950 N_A_556_369#_c_1629_n N_VGND_c_1774_n 0.00340284f $X=4.18 $Y=0.8 $X2=0
+ $Y2=0
cc_951 N_A_556_369#_c_1631_n N_VGND_c_1774_n 0.0162661f $X=4.265 $Y=0.885 $X2=0
+ $Y2=0
cc_952 N_A_556_369#_c_1647_n N_VGND_c_1784_n 0.0382345f $X=3.42 $Y=0.36 $X2=0
+ $Y2=0
cc_953 N_A_556_369#_c_1629_n N_VGND_c_1784_n 0.00248845f $X=4.18 $Y=0.8 $X2=0
+ $Y2=0
cc_954 N_A_556_369#_M1014_d N_VGND_c_1786_n 0.00220178f $X=2.805 $Y=0.235 $X2=0
+ $Y2=0
cc_955 N_A_556_369#_M1030_s N_VGND_c_1786_n 0.00230714f $X=4.245 $Y=0.235 $X2=0
+ $Y2=0
cc_956 N_A_556_369#_c_1647_n N_VGND_c_1786_n 0.0126483f $X=3.42 $Y=0.36 $X2=0
+ $Y2=0
cc_957 N_A_556_369#_c_1629_n N_VGND_c_1786_n 0.00475725f $X=4.18 $Y=0.8 $X2=0
+ $Y2=0
cc_958 N_A_556_369#_c_1631_n N_VGND_c_1786_n 0.00497919f $X=4.265 $Y=0.885 $X2=0
+ $Y2=0
cc_959 N_A_556_369#_c_1647_n A_657_47# 0.00233635f $X=3.42 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_960 N_A_556_369#_c_1628_n A_657_47# 0.00224071f $X=3.505 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_961 N_Q_c_1745_n N_VGND_c_1777_n 0.0270681f $X=9.395 $Y=0.395 $X2=0 $Y2=0
cc_962 N_Q_c_1745_n N_VGND_c_1785_n 0.0166398f $X=9.395 $Y=0.395 $X2=0 $Y2=0
cc_963 N_Q_M1000_d N_VGND_c_1786_n 0.00212516f $X=9.26 $Y=0.235 $X2=0 $Y2=0
cc_964 N_Q_c_1745_n N_VGND_c_1786_n 0.0126182f $X=9.395 $Y=0.395 $X2=0 $Y2=0
cc_965 N_VGND_c_1786_n A_483_47# 0.00171756f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_966 N_VGND_c_1786_n A_657_47# 0.00152416f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_967 N_VGND_c_1786_n A_1030_47# 0.00272292f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24
cc_968 N_VGND_c_1786_n A_1478_47# 0.0111093f $X=9.43 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__dlymetal6s6s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s6s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.575000 1.700000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.080000 0.255000 4.515000 0.825000 ;
        RECT 4.080000 1.495000 4.515000 2.465000 ;
        RECT 4.155000 0.825000 4.515000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.525000 0.655000 ;
      RECT 0.085000  0.655000 1.080000 0.825000 ;
      RECT 0.085000  1.870000 1.080000 2.040000 ;
      RECT 0.085000  2.040000 0.525000 2.465000 ;
      RECT 0.695000  0.085000 1.080000 0.485000 ;
      RECT 0.695000  2.210000 1.080000 2.635000 ;
      RECT 0.745000  0.825000 1.080000 0.995000 ;
      RECT 0.745000  0.995000 1.155000 1.325000 ;
      RECT 0.745000  1.325000 1.080000 1.870000 ;
      RECT 1.250000  0.255000 1.520000 0.825000 ;
      RECT 1.250000  1.495000 1.975000 1.675000 ;
      RECT 1.250000  1.675000 1.520000 2.465000 ;
      RECT 1.325000  0.825000 1.520000 0.995000 ;
      RECT 1.325000  0.995000 1.975000 1.495000 ;
      RECT 1.690000  0.255000 1.940000 0.655000 ;
      RECT 1.690000  0.655000 2.495000 0.825000 ;
      RECT 1.690000  1.845000 2.495000 2.040000 ;
      RECT 1.690000  2.040000 1.940000 2.465000 ;
      RECT 2.110000  0.085000 2.495000 0.485000 ;
      RECT 2.110000  2.210000 2.495000 2.635000 ;
      RECT 2.145000  0.825000 2.495000 0.995000 ;
      RECT 2.145000  0.995000 2.570000 1.325000 ;
      RECT 2.145000  1.325000 2.495000 1.845000 ;
      RECT 2.665000  0.255000 2.915000 0.825000 ;
      RECT 2.665000  1.495000 3.390000 1.675000 ;
      RECT 2.665000  1.675000 2.915000 2.465000 ;
      RECT 2.740000  0.825000 2.915000 0.995000 ;
      RECT 2.740000  0.995000 3.390000 1.495000 ;
      RECT 3.085000  0.255000 3.355000 0.655000 ;
      RECT 3.085000  0.655000 3.910000 0.825000 ;
      RECT 3.085000  1.845000 3.910000 2.040000 ;
      RECT 3.085000  2.040000 3.355000 2.465000 ;
      RECT 3.525000  0.085000 3.910000 0.485000 ;
      RECT 3.525000  2.210000 3.910000 2.635000 ;
      RECT 3.560000  0.825000 3.910000 0.995000 ;
      RECT 3.560000  0.995000 3.985000 1.325000 ;
      RECT 3.560000  1.325000 3.910000 1.845000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__dlymetal6s6s_1
END LIBRARY

* File: sky130_fd_sc_hd__conb_1.spice
* Created: Thu Aug 27 14:13:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__conb_1.pex.spice"
.subckt sky130_fd_sc_hd__conb_1  VNB VPB HI VPWR VGND LO
* 
* LO	LO
* VGND	VGND
* VPWR	VPWR
* HI	HI
* VPB	VPB
* VNB	VNB
DX0_noxref VNB VPB NWDIODE A=2.8248 P=6.73
R1 N_HI_R1_pos N_VPWR_R1_neg SHORT 0.01 M=1
R0 N_VGND_R0_pos N_LO_R0_neg SHORT 0.01 M=1
*
.include "sky130_fd_sc_hd__conb_1.pxi.spice"
*
.ends
*
*

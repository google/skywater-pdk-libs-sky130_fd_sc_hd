* File: sky130_fd_sc_hd__inv_2.spice
* Created: Tue Sep  1 19:10:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__inv_2.pex.spice"
.subckt sky130_fd_sc_hd__inv_2  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1001_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX4_noxref VNB VPB NWDIODE A=2.8248 P=6.73
*
.include "sky130_fd_sc_hd__inv_2.pxi.spice"
*
.ends
*
*

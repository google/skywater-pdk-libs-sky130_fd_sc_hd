* File: sky130_fd_sc_hd__a2bb2o_2.spice
* Created: Thu Aug 27 14:03:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2bb2o_2.pex.spice"
.subckt sky130_fd_sc_hd__a2bb2o_2  VNB VPB A1_N A2_N B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_82_21#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.08775 PD=1.83 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_82_21#_M1008_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.145916 AS=0.08775 PD=1.31822 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1011 N_A_313_47#_M1011_d N_A1_N_M1011_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0942841 PD=0.69 PS=0.851776 NRD=0 NRS=45.708 M=1 R=2.8
+ SA=75001.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_N_M1000_g N_A_313_47#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.14175 AS=0.0567 PD=1.095 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_82_21#_M1001_d N_A_313_47#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.14175 PD=0.69 PS=1.095 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_646_47# N_B2_M1004_g N_A_82_21#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=22.848 NRS=0 M=1 R=2.8 SA=75002.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g A_646_47# VNB NSHORT L=0.15 W=0.42 AD=0.1092
+ AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=22.848 M=1 R=2.8 SA=75003.3 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_82_21#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.265 PD=1.27 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1012 N_X_M1002_d N_A_82_21#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.226829 PD=1.27 PS=1.75 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 A_313_297# N_A1_N_M1005_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.145171 PD=0.85 PS=1.12 NRD=15.3857 NRS=52.8748 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_313_47#_M1006_d N_A2_N_M1006_g A_313_297# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_574_369#_M1009_d N_A_313_47#_M1009_g N_A_82_21#_M1009_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0976 AS=0.1664 PD=0.945 PS=1.8 NRD=9.2196 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1013 N_VPWR_M1013_d N_B2_M1013_g N_A_574_369#_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.0976 PD=0.91 PS=0.945 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_574_369#_M1010_d N_B1_M1010_g N_VPWR_M1013_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_75 VPB 0 1.32536e-19 $X=0.125 $Y=2.635
*
.include "sky130_fd_sc_hd__a2bb2o_2.pxi.spice"
*
.ends
*
*

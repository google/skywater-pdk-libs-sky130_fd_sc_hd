* File: sky130_fd_sc_hd__mux2i_4.pxi.spice
* Created: Tue Sep  1 19:14:54 2020
* 
x_PM_SKY130_FD_SC_HD__MUX2I_4%A0 N_A0_c_113_n N_A0_M1015_g N_A0_M1004_g
+ N_A0_c_114_n N_A0_M1018_g N_A0_M1006_g N_A0_c_115_n N_A0_M1023_g N_A0_M1024_g
+ N_A0_c_116_n N_A0_M1033_g N_A0_M1030_g A0 A0 N_A0_c_117_n N_A0_c_133_p
+ PM_SKY130_FD_SC_HD__MUX2I_4%A0
x_PM_SKY130_FD_SC_HD__MUX2I_4%A1 N_A1_c_177_n N_A1_M1019_g N_A1_M1000_g
+ N_A1_c_178_n N_A1_M1025_g N_A1_M1007_g N_A1_c_179_n N_A1_M1028_g N_A1_M1027_g
+ N_A1_c_180_n N_A1_M1029_g N_A1_M1031_g A1 A1 A1 A1 N_A1_c_182_n
+ PM_SKY130_FD_SC_HD__MUX2I_4%A1
x_PM_SKY130_FD_SC_HD__MUX2I_4%S N_S_c_248_n N_S_M1012_g N_S_M1001_g N_S_c_249_n
+ N_S_M1016_g N_S_M1011_g N_S_c_250_n N_S_M1020_g N_S_M1014_g N_S_c_251_n
+ N_S_M1026_g N_S_M1032_g N_S_M1010_g N_S_M1017_g N_S_c_262_n N_S_c_252_n
+ N_S_c_253_n S S S S S N_S_c_254_n N_S_c_255_n N_S_c_256_n
+ PM_SKY130_FD_SC_HD__MUX2I_4%S
x_PM_SKY130_FD_SC_HD__MUX2I_4%A_1191_21# N_A_1191_21#_M1010_d
+ N_A_1191_21#_M1017_d N_A_1191_21#_c_382_n N_A_1191_21#_M1003_g
+ N_A_1191_21#_M1002_g N_A_1191_21#_c_383_n N_A_1191_21#_M1009_g
+ N_A_1191_21#_M1005_g N_A_1191_21#_c_384_n N_A_1191_21#_M1013_g
+ N_A_1191_21#_M1008_g N_A_1191_21#_c_385_n N_A_1191_21#_M1021_g
+ N_A_1191_21#_M1022_g N_A_1191_21#_c_386_n N_A_1191_21#_c_387_n
+ N_A_1191_21#_c_416_n N_A_1191_21#_c_459_p N_A_1191_21#_c_388_n
+ N_A_1191_21#_c_396_n N_A_1191_21#_c_397_n N_A_1191_21#_c_389_n
+ N_A_1191_21#_c_390_n N_A_1191_21#_c_391_n
+ PM_SKY130_FD_SC_HD__MUX2I_4%A_1191_21#
x_PM_SKY130_FD_SC_HD__MUX2I_4%Y N_Y_M1015_d N_Y_M1018_d N_Y_M1033_d N_Y_M1025_s
+ N_Y_M1029_s N_Y_M1004_s N_Y_M1006_s N_Y_M1030_s N_Y_M1007_s N_Y_M1031_s
+ N_Y_c_493_n N_Y_c_494_n Y Y Y Y Y N_Y_c_497_n Y N_Y_c_498_n
+ PM_SKY130_FD_SC_HD__MUX2I_4%Y
x_PM_SKY130_FD_SC_HD__MUX2I_4%A_109_297# N_A_109_297#_M1004_d
+ N_A_109_297#_M1024_d N_A_109_297#_M1001_d N_A_109_297#_M1014_d
+ N_A_109_297#_c_564_n PM_SKY130_FD_SC_HD__MUX2I_4%A_109_297#
x_PM_SKY130_FD_SC_HD__MUX2I_4%A_445_297# N_A_445_297#_M1000_d
+ N_A_445_297#_M1027_d N_A_445_297#_M1002_d N_A_445_297#_M1008_d
+ N_A_445_297#_c_606_n N_A_445_297#_c_648_p N_A_445_297#_c_620_n
+ N_A_445_297#_c_621_n N_A_445_297#_c_651_p N_A_445_297#_c_622_n
+ PM_SKY130_FD_SC_HD__MUX2I_4%A_445_297#
x_PM_SKY130_FD_SC_HD__MUX2I_4%VPWR N_VPWR_M1001_s N_VPWR_M1011_s N_VPWR_M1032_s
+ N_VPWR_M1005_s N_VPWR_M1022_s N_VPWR_c_661_n N_VPWR_c_662_n N_VPWR_c_663_n
+ N_VPWR_c_664_n N_VPWR_c_665_n N_VPWR_c_666_n N_VPWR_c_667_n N_VPWR_c_668_n
+ VPWR N_VPWR_c_669_n N_VPWR_c_670_n N_VPWR_c_671_n N_VPWR_c_672_n
+ N_VPWR_c_660_n N_VPWR_c_674_n N_VPWR_c_675_n N_VPWR_c_676_n N_VPWR_c_677_n
+ PM_SKY130_FD_SC_HD__MUX2I_4%VPWR
x_PM_SKY130_FD_SC_HD__MUX2I_4%A_109_47# N_A_109_47#_M1015_s N_A_109_47#_M1023_s
+ N_A_109_47#_M1003_s N_A_109_47#_M1013_s N_A_109_47#_c_856_p
+ N_A_109_47#_c_776_n N_A_109_47#_c_777_n N_A_109_47#_c_778_n
+ N_A_109_47#_c_779_n N_A_109_47#_c_780_n N_A_109_47#_c_781_n
+ N_A_109_47#_c_791_n N_A_109_47#_c_782_n PM_SKY130_FD_SC_HD__MUX2I_4%A_109_47#
x_PM_SKY130_FD_SC_HD__MUX2I_4%A_445_47# N_A_445_47#_M1019_d N_A_445_47#_M1028_d
+ N_A_445_47#_M1012_d N_A_445_47#_M1020_d N_A_445_47#_c_871_n
+ N_A_445_47#_c_906_p N_A_445_47#_c_882_n N_A_445_47#_c_911_p
+ N_A_445_47#_c_887_n PM_SKY130_FD_SC_HD__MUX2I_4%A_445_47#
x_PM_SKY130_FD_SC_HD__MUX2I_4%VGND N_VGND_M1012_s N_VGND_M1016_s N_VGND_M1026_s
+ N_VGND_M1009_d N_VGND_M1021_d N_VGND_c_920_n N_VGND_c_921_n N_VGND_c_922_n
+ N_VGND_c_923_n N_VGND_c_924_n N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n
+ VGND N_VGND_c_928_n N_VGND_c_929_n N_VGND_c_930_n N_VGND_c_931_n
+ N_VGND_c_932_n N_VGND_c_933_n N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n
+ PM_SKY130_FD_SC_HD__MUX2I_4%VGND
cc_1 VNB N_A0_c_113_n 0.0191796f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A0_c_114_n 0.0159976f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A0_c_115_n 0.0157837f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A0_c_116_n 0.0157133f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A0_c_117_n 0.0666495f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_6 VNB N_A1_c_177_n 0.0159188f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_7 VNB N_A1_c_178_n 0.0157218f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_8 VNB N_A1_c_179_n 0.0157218f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_9 VNB N_A1_c_180_n 0.0213742f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_10 VNB A1 0.00843821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_182_n 0.0631588f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.16
cc_12 VNB N_S_c_248_n 0.0204799f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_S_c_249_n 0.0154946f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_14 VNB N_S_c_250_n 0.0154946f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_15 VNB N_S_c_251_n 0.0156473f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_16 VNB N_S_c_252_n 5.06002e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_17 VNB N_S_c_253_n 0.02429f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_S_c_254_n 0.0807893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_S_c_255_n 0.0195927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_S_c_256_n 0.0119128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_1191_21#_c_382_n 0.0154937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_1191_21#_c_383_n 0.0155532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_1191_21#_c_384_n 0.0162883f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_1191_21#_c_385_n 0.0165157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_1191_21#_c_386_n 0.00188285f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_26 VNB N_A_1191_21#_c_387_n 0.00134493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_1191_21#_c_388_n 0.0155218f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_28 VNB N_A_1191_21#_c_389_n 0.00723806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_1191_21#_c_390_n 0.0216914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_1191_21#_c_391_n 0.0657303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_493_n 0.00229201f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_32 VNB N_Y_c_494_n 0.00749881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB Y 0.0362141f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_660_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_109_47#_c_776_n 0.00358387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_109_47#_c_777_n 0.00128994f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_37 VNB N_A_109_47#_c_778_n 0.032359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_109_47#_c_779_n 0.00270558f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_39 VNB N_A_109_47#_c_780_n 0.00277693f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_40 VNB N_A_109_47#_c_781_n 0.00309796f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_41 VNB N_A_109_47#_c_782_n 0.00245739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_445_47#_c_871_n 0.0069465f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_43 VNB N_VGND_c_920_n 0.00556396f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_44 VNB N_VGND_c_921_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_45 VNB N_VGND_c_922_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_46 VNB N_VGND_c_923_n 3.11529e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_924_n 0.00395754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_925_n 0.00224165f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_49 VNB N_VGND_c_926_n 0.0970139f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_50 VNB N_VGND_c_927_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_51 VNB N_VGND_c_928_n 0.0117571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_929_n 0.0143953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_930_n 0.0181756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_931_n 0.0143233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_932_n 0.392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_933_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_934_n 0.00430185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_935_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_936_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VPB N_A0_M1004_g 0.0218974f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_A0_M1006_g 0.0185007f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_A0_M1024_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_63 VPB N_A0_M1030_g 0.0188371f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_64 VPB A0 9.56887e-19 $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_65 VPB N_A0_c_117_n 0.011016f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_66 VPB N_A1_M1000_g 0.0188371f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_A1_M1007_g 0.0185065f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_A1_M1027_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_69 VPB N_A1_M1031_g 0.0259842f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_70 VPB A1 0.00246857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A1_c_182_n 0.0104929f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.16
cc_72 VPB N_S_M1001_g 0.02509f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_73 VPB N_S_M1011_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_74 VPB N_S_M1014_g 0.0182735f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_75 VPB N_S_M1032_g 0.0185151f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_76 VPB N_S_M1017_g 0.021582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_S_c_262_n 0.0124079f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.16
cc_78 VPB N_S_c_252_n 0.00101908f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_79 VPB N_S_c_253_n 0.00484543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_S_c_254_n 0.0186308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_S_c_256_n 0.00284529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_1191_21#_M1002_g 0.0178983f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_83 VPB N_A_1191_21#_M1005_g 0.0177381f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_84 VPB N_A_1191_21#_M1008_g 0.0183807f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_85 VPB N_A_1191_21#_M1022_g 0.0192986f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_86 VPB N_A_1191_21#_c_396_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_1191_21#_c_397_n 0.0208429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_1191_21#_c_390_n 0.01957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_1191_21#_c_391_n 0.011431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB Y 0.0379757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_Y_c_497_n 0.00747992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_Y_c_498_n 0.00218948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_109_297#_c_564_n 0.00939914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_445_297#_c_606_n 0.00721458f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_95 VPB N_VPWR_c_661_n 0.00551074f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_96 VPB N_VPWR_c_662_n 0.011815f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_97 VPB N_VPWR_c_663_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_98 VPB N_VPWR_c_664_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_665_n 3.18775e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_666_n 0.00220674f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.16
cc_101 VPB N_VPWR_c_667_n 0.0957431f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.16
cc_102 VPB N_VPWR_c_668_n 0.00507168f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_103 VPB N_VPWR_c_669_n 0.011815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_670_n 0.0109642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_671_n 0.0159568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_672_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_660_n 0.0470842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_674_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_675_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_676_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_677_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 N_A0_c_116_n N_A1_c_177_n 0.0300515f $X=1.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_113 N_A0_M1030_g N_A1_M1000_g 0.0300515f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A0_c_117_n A1 0.00968937f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A0_c_117_n N_A1_c_182_n 0.0300515f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A0_c_113_n N_Y_c_493_n 0.0116557f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A0_c_114_n N_Y_c_493_n 0.00802124f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A0_c_115_n N_Y_c_493_n 0.00796648f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A0_c_116_n N_Y_c_493_n 0.00838304f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A0_c_113_n Y 0.0566596f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A0_c_133_p Y 0.0204711f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A0_M1004_g N_Y_c_498_n 0.0118662f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A0_M1006_g N_Y_c_498_n 0.00958166f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A0_M1024_g N_Y_c_498_n 0.00958166f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A0_M1030_g N_Y_c_498_n 0.00958166f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A0_M1004_g N_A_109_297#_c_564_n 0.00397177f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A0_M1006_g N_A_109_297#_c_564_n 0.0105345f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A0_M1024_g N_A_109_297#_c_564_n 0.0140195f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A0_M1030_g N_A_109_297#_c_564_n 0.0126559f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_130 A0 N_A_109_297#_c_564_n 0.0148933f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_131 N_A0_c_117_n N_A_109_297#_c_564_n 0.00470231f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A0_c_133_p N_A_109_297#_c_564_n 0.0159649f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A0_M1030_g N_A_445_297#_c_606_n 8.22884e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A0_M1004_g N_VPWR_c_667_n 0.00366111f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A0_M1006_g N_VPWR_c_667_n 0.00366111f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A0_M1024_g N_VPWR_c_667_n 0.00366111f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A0_M1030_g N_VPWR_c_667_n 0.00366111f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A0_M1004_g N_VPWR_c_660_n 0.00619429f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A0_M1006_g N_VPWR_c_660_n 0.00524008f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A0_M1024_g N_VPWR_c_660_n 0.00524008f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A0_M1030_g N_VPWR_c_660_n 0.00526729f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A0_c_116_n N_A_109_47#_c_778_n 0.00314568f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A0_c_115_n N_A_109_47#_c_779_n 4.99997e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A0_c_116_n N_A_109_47#_c_779_n 0.00354096f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A0_c_117_n N_A_109_47#_c_779_n 0.00252992f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A0_c_114_n N_A_109_47#_c_781_n 5.39464e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A0_c_115_n N_A_109_47#_c_781_n 0.00432443f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A0_c_116_n N_A_109_47#_c_781_n 0.00724554f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A0_c_117_n N_A_109_47#_c_781_n 0.00273752f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A0_c_113_n N_A_109_47#_c_791_n 0.00363882f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A0_c_114_n N_A_109_47#_c_791_n 0.00835735f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A0_c_115_n N_A_109_47#_c_791_n 0.0105707f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_153 A0 N_A_109_47#_c_791_n 0.0168981f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A0_c_117_n N_A_109_47#_c_791_n 0.00389845f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A0_c_133_p N_A_109_47#_c_791_n 0.0215892f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A0_c_116_n N_A_445_47#_c_871_n 5.0821e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A0_c_113_n N_VGND_c_926_n 0.00370116f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A0_c_114_n N_VGND_c_926_n 0.00370116f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A0_c_115_n N_VGND_c_926_n 0.00370116f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A0_c_116_n N_VGND_c_926_n 0.00370116f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A0_c_113_n N_VGND_c_932_n 0.00620778f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A0_c_114_n N_VGND_c_932_n 0.00525357f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A0_c_115_n N_VGND_c_932_n 0.00525357f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A0_c_116_n N_VGND_c_932_n 0.00518598f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_165 A1 N_S_c_254_n 0.0034512f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A1_c_182_n N_S_c_254_n 0.00656311f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_167 A1 N_S_c_256_n 0.0135622f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A1_c_182_n N_S_c_256_n 9.26194e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A1_c_177_n N_Y_c_493_n 0.00918142f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_c_178_n N_Y_c_493_n 0.00797825f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A1_c_179_n N_Y_c_493_n 0.00797825f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A1_c_180_n N_Y_c_493_n 0.00797825f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_173 A1 N_Y_c_493_n 0.00295891f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A1_M1000_g N_Y_c_498_n 0.00924135f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A1_M1007_g N_Y_c_498_n 0.00789149f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A1_M1027_g N_Y_c_498_n 0.00789149f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A1_M1031_g N_Y_c_498_n 0.00789149f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A1_M1000_g N_A_109_297#_c_564_n 0.0121541f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A1_M1007_g N_A_109_297#_c_564_n 0.0108371f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A1_M1027_g N_A_109_297#_c_564_n 0.0108371f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A1_M1031_g N_A_109_297#_c_564_n 0.0129401f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_182 A1 N_A_109_297#_c_564_n 0.0744382f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_183 N_A1_c_182_n N_A_109_297#_c_564_n 0.00573337f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A1_M1000_g N_A_445_297#_c_606_n 0.00414626f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A1_M1007_g N_A_445_297#_c_606_n 0.00835694f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A1_M1027_g N_A_445_297#_c_606_n 0.00835694f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A1_M1031_g N_A_445_297#_c_606_n 0.0104599f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A1_M1031_g N_VPWR_c_661_n 0.00294182f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A1_M1000_g N_VPWR_c_667_n 0.00366111f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A1_M1007_g N_VPWR_c_667_n 0.00366111f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A1_M1027_g N_VPWR_c_667_n 0.00366111f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A1_M1031_g N_VPWR_c_667_n 0.00366111f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A1_M1000_g N_VPWR_c_660_n 0.00526729f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A1_M1007_g N_VPWR_c_660_n 0.00524008f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A1_M1027_g N_VPWR_c_660_n 0.00524008f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A1_M1031_g N_VPWR_c_660_n 0.00656615f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A1_c_177_n N_A_109_47#_c_778_n 0.00365431f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A1_c_178_n N_A_109_47#_c_778_n 0.00200334f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_179_n N_A_109_47#_c_778_n 0.00200334f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_180_n N_A_109_47#_c_778_n 0.00296219f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_201 A1 N_A_109_47#_c_778_n 0.0440177f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A1_c_182_n N_A_109_47#_c_778_n 0.00689377f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A1_c_177_n N_A_109_47#_c_779_n 4.48188e-19 $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A1_c_177_n N_A_109_47#_c_781_n 0.00148704f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A1_c_177_n N_A_445_47#_c_871_n 0.00328646f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A1_c_178_n N_A_445_47#_c_871_n 0.00744623f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_c_179_n N_A_445_47#_c_871_n 0.00744623f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A1_c_180_n N_A_445_47#_c_871_n 0.00954923f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_209 A1 N_A_445_47#_c_871_n 0.0790641f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_210 N_A1_c_182_n N_A_445_47#_c_871_n 0.00592732f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A1_c_180_n N_VGND_c_920_n 0.00323055f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A1_c_177_n N_VGND_c_926_n 0.00370116f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A1_c_178_n N_VGND_c_926_n 0.00370116f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A1_c_179_n N_VGND_c_926_n 0.00370116f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A1_c_180_n N_VGND_c_926_n 0.00370116f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A1_c_177_n N_VGND_c_932_n 0.00522046f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A1_c_178_n N_VGND_c_932_n 0.00519326f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A1_c_179_n N_VGND_c_932_n 0.00519326f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A1_c_180_n N_VGND_c_932_n 0.00651933f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_220 N_S_c_251_n N_A_1191_21#_c_382_n 0.0281996f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_221 N_S_M1032_g N_A_1191_21#_M1002_g 0.0281996f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_222 N_S_c_262_n N_A_1191_21#_M1002_g 0.0111161f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_223 N_S_c_256_n N_A_1191_21#_M1002_g 4.73289e-19 $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_224 N_S_c_262_n N_A_1191_21#_M1005_g 0.0128436f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_225 N_S_c_262_n N_A_1191_21#_M1008_g 0.0115952f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_226 N_S_c_255_n N_A_1191_21#_c_385_n 0.0208288f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_227 N_S_M1017_g N_A_1191_21#_M1022_g 0.0367345f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_228 N_S_c_262_n N_A_1191_21#_M1022_g 0.0155447f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_229 N_S_c_252_n N_A_1191_21#_M1022_g 0.00186804f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_230 N_S_c_262_n N_A_1191_21#_c_386_n 0.0538621f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_231 N_S_c_252_n N_A_1191_21#_c_386_n 0.0137152f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_232 N_S_c_253_n N_A_1191_21#_c_386_n 0.00112698f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_233 N_S_c_252_n N_A_1191_21#_c_387_n 0.00568392f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_234 N_S_c_253_n N_A_1191_21#_c_387_n 4.51858e-19 $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_235 N_S_c_255_n N_A_1191_21#_c_387_n 0.00144115f $X=7.765 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_S_c_262_n N_A_1191_21#_c_416_n 0.00499447f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_237 N_S_c_252_n N_A_1191_21#_c_416_n 0.0108252f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_238 N_S_c_253_n N_A_1191_21#_c_416_n 0.00134547f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_239 N_S_c_255_n N_A_1191_21#_c_416_n 0.0143161f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_240 N_S_M1017_g N_A_1191_21#_c_390_n 0.0119502f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_241 N_S_c_262_n N_A_1191_21#_c_390_n 0.0134681f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_242 N_S_c_252_n N_A_1191_21#_c_390_n 0.0307572f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_243 N_S_c_253_n N_A_1191_21#_c_390_n 0.00753785f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_244 N_S_c_255_n N_A_1191_21#_c_390_n 0.00401066f $X=7.765 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_S_c_262_n N_A_1191_21#_c_391_n 0.00865217f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_246 N_S_c_252_n N_A_1191_21#_c_391_n 7.94023e-19 $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_247 N_S_c_253_n N_A_1191_21#_c_391_n 0.0210442f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_248 N_S_c_254_n N_A_1191_21#_c_391_n 0.0281996f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_249 N_S_c_256_n N_A_1191_21#_c_391_n 0.00911724f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_250 N_S_M1001_g N_A_109_297#_c_564_n 0.0111391f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_251 N_S_M1011_g N_A_109_297#_c_564_n 0.00903607f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_252 N_S_M1014_g N_A_109_297#_c_564_n 0.00903607f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_253 N_S_M1032_g N_A_109_297#_c_564_n 0.00475469f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_254 N_S_c_254_n N_A_109_297#_c_564_n 0.0117992f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_255 N_S_c_256_n N_A_109_297#_c_564_n 0.0744898f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_256 N_S_c_262_n N_A_445_297#_M1002_d 0.00177804f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_257 N_S_c_262_n N_A_445_297#_M1008_d 0.00368929f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_258 N_S_M1001_g N_A_445_297#_c_606_n 0.0135546f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_259 N_S_M1011_g N_A_445_297#_c_606_n 0.0114516f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_260 N_S_M1014_g N_A_445_297#_c_606_n 0.0114516f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_261 N_S_M1032_g N_A_445_297#_c_606_n 0.0128972f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_262 N_S_c_262_n N_A_445_297#_c_606_n 0.00610735f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_263 N_S_c_256_n N_A_445_297#_c_606_n 0.0107246f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_264 N_S_c_262_n N_A_445_297#_c_620_n 0.0193328f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_265 N_S_c_262_n N_A_445_297#_c_621_n 0.0117344f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_266 N_S_c_262_n N_A_445_297#_c_622_n 0.0112304f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_267 N_S_c_256_n N_VPWR_M1032_s 0.00327615f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_268 N_S_c_262_n N_VPWR_M1005_s 0.00222979f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_269 N_S_c_262_n N_VPWR_M1022_s 0.0042052f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_270 N_S_M1001_g N_VPWR_c_661_n 0.00921014f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_271 N_S_M1011_g N_VPWR_c_661_n 0.00110281f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_272 N_S_M1001_g N_VPWR_c_662_n 0.00339367f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_273 N_S_M1011_g N_VPWR_c_662_n 0.00339367f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_274 N_S_M1001_g N_VPWR_c_663_n 0.00110281f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_275 N_S_M1011_g N_VPWR_c_663_n 0.00810864f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_276 N_S_M1014_g N_VPWR_c_663_n 0.00810864f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_277 N_S_M1032_g N_VPWR_c_663_n 0.00110281f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_278 N_S_M1014_g N_VPWR_c_664_n 0.00110281f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_279 N_S_M1032_g N_VPWR_c_664_n 0.00807474f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_280 N_S_M1017_g N_VPWR_c_666_n 0.00874183f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_281 N_S_c_262_n N_VPWR_c_666_n 0.00652775f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_282 N_S_M1014_g N_VPWR_c_669_n 0.00339367f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_283 N_S_M1032_g N_VPWR_c_669_n 0.00339367f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_284 N_S_M1017_g N_VPWR_c_672_n 0.0046653f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_285 N_S_M1001_g N_VPWR_c_660_n 0.00398704f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_286 N_S_M1011_g N_VPWR_c_660_n 0.00398704f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_287 N_S_M1014_g N_VPWR_c_660_n 0.00398704f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_288 N_S_M1032_g N_VPWR_c_660_n 0.00398704f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_289 N_S_M1017_g N_VPWR_c_660_n 0.008846f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_290 N_S_c_262_n N_A_109_47#_c_776_n 0.0091871f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_291 N_S_c_248_n N_A_109_47#_c_778_n 0.00339216f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_292 N_S_c_249_n N_A_109_47#_c_778_n 0.00243331f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_293 N_S_c_250_n N_A_109_47#_c_778_n 0.00243331f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_294 N_S_c_251_n N_A_109_47#_c_778_n 0.00590253f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_295 N_S_c_262_n N_A_109_47#_c_778_n 0.00433579f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_296 N_S_c_254_n N_A_109_47#_c_778_n 0.0141705f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_297 N_S_c_256_n N_A_109_47#_c_778_n 0.0571674f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_298 N_S_c_251_n N_A_109_47#_c_780_n 4.04423e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_299 N_S_c_262_n N_A_109_47#_c_780_n 0.00735336f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_300 N_S_c_262_n N_A_109_47#_c_782_n 0.00709898f $X=7.68 $Y=1.51 $X2=0 $Y2=0
cc_301 N_S_c_248_n N_A_445_47#_c_871_n 0.0132343f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_302 N_S_c_254_n N_A_445_47#_c_871_n 0.00639383f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_303 N_S_c_256_n N_A_445_47#_c_871_n 0.0245762f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_304 N_S_c_249_n N_A_445_47#_c_882_n 0.0110872f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_305 N_S_c_250_n N_A_445_47#_c_882_n 0.0106549f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_306 N_S_c_251_n N_A_445_47#_c_882_n 8.79528e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_307 N_S_c_254_n N_A_445_47#_c_882_n 0.00411986f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_308 N_S_c_256_n N_A_445_47#_c_882_n 0.0309697f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_309 N_S_c_254_n N_A_445_47#_c_887_n 0.00207868f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_310 N_S_c_256_n N_A_445_47#_c_887_n 0.00684798f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_311 N_S_c_248_n N_VGND_c_920_n 0.00776101f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_312 N_S_c_249_n N_VGND_c_920_n 5.08801e-19 $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_313 N_S_c_248_n N_VGND_c_921_n 0.00341689f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_314 N_S_c_249_n N_VGND_c_921_n 0.00341689f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_315 N_S_c_248_n N_VGND_c_922_n 5.08801e-19 $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_316 N_S_c_249_n N_VGND_c_922_n 0.00665951f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_317 N_S_c_250_n N_VGND_c_922_n 0.00665951f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_318 N_S_c_251_n N_VGND_c_922_n 5.08801e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_319 N_S_c_250_n N_VGND_c_923_n 5.45345e-19 $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_320 N_S_c_251_n N_VGND_c_923_n 0.00817595f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_321 N_S_c_256_n N_VGND_c_923_n 0.00409219f $X=5.76 $Y=1.182 $X2=0 $Y2=0
cc_322 N_S_c_255_n N_VGND_c_925_n 0.00832147f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_323 N_S_c_250_n N_VGND_c_928_n 0.00341689f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_324 N_S_c_251_n N_VGND_c_928_n 0.0046653f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_325 N_S_c_255_n N_VGND_c_931_n 0.00341689f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_326 N_S_c_248_n N_VGND_c_932_n 0.00374793f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_327 N_S_c_249_n N_VGND_c_932_n 0.00374793f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_328 N_S_c_250_n N_VGND_c_932_n 0.00374793f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_329 N_S_c_251_n N_VGND_c_932_n 0.00439268f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_330 N_S_c_255_n N_VGND_c_932_n 0.00493711f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_1191_21#_M1002_g N_A_109_297#_c_564_n 7.53608e-19 $X=6.03 $Y=1.985
+ $X2=0 $Y2=0
cc_332 N_A_1191_21#_M1002_g N_A_445_297#_c_606_n 0.0102478f $X=6.03 $Y=1.985
+ $X2=0 $Y2=0
cc_333 N_A_1191_21#_M1005_g N_A_445_297#_c_620_n 0.0102478f $X=6.45 $Y=1.985
+ $X2=0 $Y2=0
cc_334 N_A_1191_21#_M1008_g N_A_445_297#_c_620_n 0.010292f $X=6.87 $Y=1.985
+ $X2=0 $Y2=0
cc_335 N_A_1191_21#_M1002_g N_VPWR_c_664_n 0.00661031f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A_1191_21#_M1005_g N_VPWR_c_664_n 5.08801e-19 $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A_1191_21#_M1002_g N_VPWR_c_665_n 5.08801e-19 $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A_1191_21#_M1005_g N_VPWR_c_665_n 0.00664421f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A_1191_21#_M1008_g N_VPWR_c_665_n 0.00689755f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_1191_21#_M1022_g N_VPWR_c_665_n 5.10067e-19 $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_1191_21#_M1022_g N_VPWR_c_666_n 0.00169441f $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_1191_21#_M1002_g N_VPWR_c_670_n 0.00339367f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_1191_21#_M1005_g N_VPWR_c_670_n 0.00339367f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_1191_21#_M1008_g N_VPWR_c_671_n 0.00339367f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_345 N_A_1191_21#_M1022_g N_VPWR_c_671_n 0.00585385f $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_A_1191_21#_c_397_n N_VPWR_c_672_n 0.0179951f $X=8.02 $Y=1.96 $X2=0
+ $Y2=0
cc_347 N_A_1191_21#_M1017_d N_VPWR_c_660_n 0.00382897f $X=7.885 $Y=1.485 $X2=0
+ $Y2=0
cc_348 N_A_1191_21#_M1002_g N_VPWR_c_660_n 0.00394406f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_1191_21#_M1005_g N_VPWR_c_660_n 0.00394406f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_350 N_A_1191_21#_M1008_g N_VPWR_c_660_n 0.00408307f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_351 N_A_1191_21#_M1022_g N_VPWR_c_660_n 0.0107224f $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A_1191_21#_c_397_n N_VPWR_c_660_n 0.00993477f $X=8.02 $Y=1.96 $X2=0
+ $Y2=0
cc_353 N_A_1191_21#_c_383_n N_A_109_47#_c_776_n 0.00717432f $X=6.45 $Y=0.995
+ $X2=0 $Y2=0
cc_354 N_A_1191_21#_c_384_n N_A_109_47#_c_776_n 0.0107582f $X=6.87 $Y=0.995
+ $X2=0 $Y2=0
cc_355 N_A_1191_21#_c_386_n N_A_109_47#_c_776_n 0.0185558f $X=7.34 $Y=1.16 $X2=0
+ $Y2=0
cc_356 N_A_1191_21#_c_391_n N_A_109_47#_c_776_n 0.00261365f $X=7.345 $Y=1.16
+ $X2=0 $Y2=0
cc_357 N_A_1191_21#_c_385_n N_A_109_47#_c_777_n 0.00349008f $X=7.345 $Y=0.995
+ $X2=0 $Y2=0
cc_358 N_A_1191_21#_c_386_n N_A_109_47#_c_777_n 0.0129401f $X=7.34 $Y=1.16 $X2=0
+ $Y2=0
cc_359 N_A_1191_21#_c_387_n N_A_109_47#_c_777_n 0.00548541f $X=7.425 $Y=1.075
+ $X2=0 $Y2=0
cc_360 N_A_1191_21#_c_459_p N_A_109_47#_c_777_n 0.0130629f $X=7.51 $Y=0.74 $X2=0
+ $Y2=0
cc_361 N_A_1191_21#_c_391_n N_A_109_47#_c_777_n 0.00325298f $X=7.345 $Y=1.16
+ $X2=0 $Y2=0
cc_362 N_A_1191_21#_c_382_n N_A_109_47#_c_778_n 0.00528324f $X=6.03 $Y=0.995
+ $X2=0 $Y2=0
cc_363 N_A_1191_21#_c_382_n N_A_109_47#_c_780_n 0.00320288f $X=6.03 $Y=0.995
+ $X2=0 $Y2=0
cc_364 N_A_1191_21#_c_383_n N_A_109_47#_c_780_n 7.95234e-19 $X=6.45 $Y=0.995
+ $X2=0 $Y2=0
cc_365 N_A_1191_21#_c_391_n N_A_109_47#_c_780_n 0.00252992f $X=7.345 $Y=1.16
+ $X2=0 $Y2=0
cc_366 N_A_1191_21#_c_382_n N_A_109_47#_c_782_n 0.00274919f $X=6.03 $Y=0.995
+ $X2=0 $Y2=0
cc_367 N_A_1191_21#_c_383_n N_A_109_47#_c_782_n 0.00759988f $X=6.45 $Y=0.995
+ $X2=0 $Y2=0
cc_368 N_A_1191_21#_c_391_n N_A_109_47#_c_782_n 0.00259382f $X=7.345 $Y=1.16
+ $X2=0 $Y2=0
cc_369 N_A_1191_21#_c_387_n N_VGND_M1021_d 7.39312e-19 $X=7.425 $Y=1.075 $X2=0
+ $Y2=0
cc_370 N_A_1191_21#_c_416_n N_VGND_M1021_d 0.00484187f $X=7.935 $Y=0.74 $X2=0
+ $Y2=0
cc_371 N_A_1191_21#_c_459_p N_VGND_M1021_d 3.67444e-19 $X=7.51 $Y=0.74 $X2=0
+ $Y2=0
cc_372 N_A_1191_21#_c_382_n N_VGND_c_923_n 0.00781141f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_373 N_A_1191_21#_c_383_n N_VGND_c_923_n 5.60997e-19 $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_A_1191_21#_c_383_n N_VGND_c_924_n 0.00150347f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A_1191_21#_c_384_n N_VGND_c_924_n 0.00167094f $X=6.87 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A_1191_21#_c_385_n N_VGND_c_925_n 0.00173437f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A_1191_21#_c_416_n N_VGND_c_925_n 0.0134931f $X=7.935 $Y=0.74 $X2=0
+ $Y2=0
cc_378 N_A_1191_21#_c_459_p N_VGND_c_925_n 0.00250582f $X=7.51 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_1191_21#_c_382_n N_VGND_c_929_n 0.00486043f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_380 N_A_1191_21#_c_383_n N_VGND_c_929_n 0.00436487f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_381 N_A_1191_21#_c_384_n N_VGND_c_930_n 0.00435702f $X=6.87 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A_1191_21#_c_385_n N_VGND_c_930_n 0.0050138f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_383 N_A_1191_21#_c_459_p N_VGND_c_930_n 0.00149044f $X=7.51 $Y=0.74 $X2=0
+ $Y2=0
cc_384 N_A_1191_21#_c_416_n N_VGND_c_931_n 0.0023303f $X=7.935 $Y=0.74 $X2=0
+ $Y2=0
cc_385 N_A_1191_21#_c_388_n N_VGND_c_931_n 0.0179308f $X=8.02 $Y=0.42 $X2=0
+ $Y2=0
cc_386 N_A_1191_21#_M1010_d N_VGND_c_932_n 0.00227813f $X=7.885 $Y=0.235 $X2=0
+ $Y2=0
cc_387 N_A_1191_21#_c_382_n N_VGND_c_932_n 0.00454278f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_388 N_A_1191_21#_c_383_n N_VGND_c_932_n 0.00572899f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_389 N_A_1191_21#_c_384_n N_VGND_c_932_n 0.00591942f $X=6.87 $Y=0.995 $X2=0
+ $Y2=0
cc_390 N_A_1191_21#_c_385_n N_VGND_c_932_n 0.00822896f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_391 N_A_1191_21#_c_416_n N_VGND_c_932_n 0.00525664f $X=7.935 $Y=0.74 $X2=0
+ $Y2=0
cc_392 N_A_1191_21#_c_459_p N_VGND_c_932_n 0.00272271f $X=7.51 $Y=0.74 $X2=0
+ $Y2=0
cc_393 N_A_1191_21#_c_388_n N_VGND_c_932_n 0.00992122f $X=8.02 $Y=0.42 $X2=0
+ $Y2=0
cc_394 N_Y_c_498_n N_A_109_297#_M1004_d 0.00444362f $X=3.62 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_395 N_Y_c_498_n N_A_109_297#_M1024_d 0.00444362f $X=3.62 $Y=2.34 $X2=0 $Y2=0
cc_396 N_Y_M1006_s N_A_109_297#_c_564_n 0.00458555f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_397 N_Y_M1030_s N_A_109_297#_c_564_n 0.00719351f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_398 N_Y_M1007_s N_A_109_297#_c_564_n 0.00340334f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_399 N_Y_M1031_s N_A_109_297#_c_564_n 0.0104487f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_400 Y N_A_109_297#_c_564_n 0.0121051f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_401 N_Y_c_498_n N_A_109_297#_c_564_n 0.0365499f $X=3.62 $Y=2.34 $X2=0 $Y2=0
cc_402 N_Y_c_498_n N_A_445_297#_M1000_d 0.00325828f $X=3.62 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_403 N_Y_c_498_n N_A_445_297#_M1027_d 0.00325828f $X=3.62 $Y=2.34 $X2=0 $Y2=0
cc_404 N_Y_M1007_s N_A_445_297#_c_606_n 0.0031771f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_405 N_Y_M1031_s N_A_445_297#_c_606_n 0.00498799f $X=3.485 $Y=1.485 $X2=0
+ $Y2=0
cc_406 N_Y_c_498_n N_A_445_297#_c_606_n 0.0797617f $X=3.62 $Y=2.34 $X2=0 $Y2=0
cc_407 N_Y_c_498_n N_VPWR_c_661_n 0.0137364f $X=3.62 $Y=2.34 $X2=0 $Y2=0
cc_408 N_Y_c_497_n N_VPWR_c_667_n 0.0125737f $X=0.207 $Y=2.255 $X2=0 $Y2=0
cc_409 N_Y_c_498_n N_VPWR_c_667_n 0.152999f $X=3.62 $Y=2.34 $X2=0 $Y2=0
cc_410 N_Y_M1004_s N_VPWR_c_660_n 0.00211589f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_411 N_Y_M1006_s N_VPWR_c_660_n 0.00217615f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_412 N_Y_M1030_s N_VPWR_c_660_n 0.00217615f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_413 N_Y_M1007_s N_VPWR_c_660_n 0.00217615f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_414 N_Y_M1031_s N_VPWR_c_660_n 0.00211652f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_415 N_Y_c_497_n N_VPWR_c_660_n 0.00848224f $X=0.207 $Y=2.255 $X2=0 $Y2=0
cc_416 N_Y_c_498_n N_VPWR_c_660_n 0.119789f $X=3.62 $Y=2.34 $X2=0 $Y2=0
cc_417 N_Y_c_493_n N_A_109_47#_M1015_s 0.00321971f $X=3.62 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_418 N_Y_c_493_n N_A_109_47#_M1023_s 0.00313041f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_419 N_Y_M1033_d N_A_109_47#_c_778_n 0.00213469f $X=1.805 $Y=0.235 $X2=0 $Y2=0
cc_420 N_Y_c_493_n N_A_109_47#_c_778_n 0.0127962f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_421 N_Y_c_493_n N_A_109_47#_c_779_n 0.00221805f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_422 N_Y_M1018_d N_A_109_47#_c_791_n 0.00328781f $X=0.965 $Y=0.235 $X2=0 $Y2=0
cc_423 N_Y_c_493_n N_A_109_47#_c_791_n 0.0559591f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_424 Y N_A_109_47#_c_791_n 0.0121051f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_425 N_Y_c_493_n N_A_445_47#_M1019_d 0.00312714f $X=3.62 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_426 N_Y_c_493_n N_A_445_47#_M1028_d 0.00312714f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_427 N_Y_M1025_s N_A_445_47#_c_871_n 0.00234448f $X=2.645 $Y=0.235 $X2=0 $Y2=0
cc_428 N_Y_M1029_s N_A_445_47#_c_871_n 0.00619269f $X=3.485 $Y=0.235 $X2=0 $Y2=0
cc_429 N_Y_c_493_n N_A_445_47#_c_871_n 0.0741865f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_430 N_Y_c_493_n N_VGND_c_920_n 0.0121829f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_431 N_Y_c_493_n N_VGND_c_926_n 0.138967f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_432 N_Y_c_494_n N_VGND_c_926_n 0.0114485f $X=0.207 $Y=0.485 $X2=0 $Y2=0
cc_433 N_Y_M1015_d N_VGND_c_932_n 0.00213654f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_434 N_Y_M1018_d N_VGND_c_932_n 0.00219774f $X=0.965 $Y=0.235 $X2=0 $Y2=0
cc_435 N_Y_M1033_d N_VGND_c_932_n 0.00180037f $X=1.805 $Y=0.235 $X2=0 $Y2=0
cc_436 N_Y_M1025_s N_VGND_c_932_n 0.00180037f $X=2.645 $Y=0.235 $X2=0 $Y2=0
cc_437 N_Y_M1029_s N_VGND_c_932_n 0.00175336f $X=3.485 $Y=0.235 $X2=0 $Y2=0
cc_438 N_Y_c_493_n N_VGND_c_932_n 0.0746967f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_439 N_Y_c_494_n N_VGND_c_932_n 0.00840192f $X=0.207 $Y=0.485 $X2=0 $Y2=0
cc_440 N_A_109_297#_c_564_n N_A_445_297#_M1000_d 0.00340334f $X=5.4 $Y=1.66
+ $X2=-0.19 $Y2=1.305
cc_441 N_A_109_297#_c_564_n N_A_445_297#_M1027_d 0.00340334f $X=5.4 $Y=1.66
+ $X2=0 $Y2=0
cc_442 N_A_109_297#_M1001_d N_A_445_297#_c_606_n 0.00429879f $X=4.425 $Y=1.485
+ $X2=0 $Y2=0
cc_443 N_A_109_297#_M1014_d N_A_445_297#_c_606_n 0.00429879f $X=5.265 $Y=1.485
+ $X2=0 $Y2=0
cc_444 N_A_109_297#_c_564_n N_A_445_297#_c_606_n 0.18362f $X=5.4 $Y=1.66 $X2=0
+ $Y2=0
cc_445 N_A_109_297#_c_564_n N_VPWR_M1001_s 0.00506752f $X=5.4 $Y=1.66 $X2=-0.19
+ $Y2=1.305
cc_446 N_A_109_297#_c_564_n N_VPWR_M1011_s 0.00351036f $X=5.4 $Y=1.66 $X2=0
+ $Y2=0
cc_447 N_A_109_297#_M1004_d N_VPWR_c_660_n 0.00219239f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_A_109_297#_M1024_d N_VPWR_c_660_n 0.00219239f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_449 N_A_109_297#_M1001_d N_VPWR_c_660_n 0.00315309f $X=4.425 $Y=1.485 $X2=0
+ $Y2=0
cc_450 N_A_109_297#_M1014_d N_VPWR_c_660_n 0.00315309f $X=5.265 $Y=1.485 $X2=0
+ $Y2=0
cc_451 N_A_109_297#_c_564_n N_A_109_47#_c_779_n 0.00605413f $X=5.4 $Y=1.66 $X2=0
+ $Y2=0
cc_452 N_A_109_297#_c_564_n N_A_109_47#_c_781_n 0.0053371f $X=5.4 $Y=1.66 $X2=0
+ $Y2=0
cc_453 N_A_445_297#_c_606_n N_VPWR_M1001_s 0.00479287f $X=6.155 $Y=2 $X2=-0.19
+ $Y2=1.305
cc_454 N_A_445_297#_c_606_n N_VPWR_M1011_s 0.00317338f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_455 N_A_445_297#_c_606_n N_VPWR_M1032_s 0.00391669f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_456 N_A_445_297#_c_620_n N_VPWR_M1005_s 0.00368869f $X=6.995 $Y=2 $X2=0 $Y2=0
cc_457 N_A_445_297#_c_606_n N_VPWR_c_661_n 0.0206068f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_458 N_A_445_297#_c_606_n N_VPWR_c_662_n 0.0077537f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_459 N_A_445_297#_c_606_n N_VPWR_c_663_n 0.0159625f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_460 N_A_445_297#_c_606_n N_VPWR_c_664_n 0.0159625f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_461 N_A_445_297#_c_620_n N_VPWR_c_665_n 0.0159625f $X=6.995 $Y=2 $X2=0 $Y2=0
cc_462 N_A_445_297#_c_606_n N_VPWR_c_667_n 0.00346265f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_463 N_A_445_297#_c_606_n N_VPWR_c_669_n 0.0077537f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_464 N_A_445_297#_c_606_n N_VPWR_c_670_n 0.00243651f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_465 N_A_445_297#_c_648_p N_VPWR_c_670_n 0.0113839f $X=6.24 $Y=2.3 $X2=0 $Y2=0
cc_466 N_A_445_297#_c_620_n N_VPWR_c_670_n 0.00243651f $X=6.995 $Y=2 $X2=0 $Y2=0
cc_467 N_A_445_297#_c_620_n N_VPWR_c_671_n 0.00243651f $X=6.995 $Y=2 $X2=0 $Y2=0
cc_468 N_A_445_297#_c_651_p N_VPWR_c_671_n 0.0115924f $X=7.08 $Y=2.3 $X2=0 $Y2=0
cc_469 N_A_445_297#_M1000_d N_VPWR_c_660_n 0.00219239f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_470 N_A_445_297#_M1027_d N_VPWR_c_660_n 0.00219239f $X=3.065 $Y=1.485 $X2=0
+ $Y2=0
cc_471 N_A_445_297#_M1002_d N_VPWR_c_660_n 0.00249348f $X=6.105 $Y=1.485 $X2=0
+ $Y2=0
cc_472 N_A_445_297#_M1008_d N_VPWR_c_660_n 0.00640954f $X=6.945 $Y=1.485 $X2=0
+ $Y2=0
cc_473 N_A_445_297#_c_606_n N_VPWR_c_660_n 0.0434736f $X=6.155 $Y=2 $X2=0 $Y2=0
cc_474 N_A_445_297#_c_648_p N_VPWR_c_660_n 0.00646745f $X=6.24 $Y=2.3 $X2=0
+ $Y2=0
cc_475 N_A_445_297#_c_620_n N_VPWR_c_660_n 0.00998922f $X=6.995 $Y=2 $X2=0 $Y2=0
cc_476 N_A_445_297#_c_651_p N_VPWR_c_660_n 0.00646745f $X=7.08 $Y=2.3 $X2=0
+ $Y2=0
cc_477 N_A_109_47#_c_778_n N_A_445_47#_M1020_d 6.95505e-19 $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_478 N_A_109_47#_c_778_n N_A_445_47#_c_871_n 0.0687817f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_479 N_A_109_47#_c_779_n N_A_445_47#_c_871_n 9.61573e-19 $X=1.76 $Y=0.85 $X2=0
+ $Y2=0
cc_480 N_A_109_47#_c_781_n N_A_445_47#_c_871_n 0.00429899f $X=1.52 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A_109_47#_c_778_n N_A_445_47#_c_882_n 0.0279268f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_482 N_A_109_47#_c_780_n N_A_445_47#_c_882_n 8.86792e-19 $X=6.235 $Y=0.85
+ $X2=0 $Y2=0
cc_483 N_A_109_47#_c_782_n N_A_445_47#_c_882_n 5.15816e-19 $X=6.45 $Y=0.825
+ $X2=0 $Y2=0
cc_484 N_A_109_47#_c_778_n N_A_445_47#_c_887_n 0.00672952f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_485 N_A_109_47#_c_778_n N_VGND_M1026_s 0.0019359f $X=6.09 $Y=0.85 $X2=0 $Y2=0
cc_486 N_A_109_47#_c_776_n N_VGND_M1009_d 0.00162148f $X=6.995 $Y=0.81 $X2=0
+ $Y2=0
cc_487 N_A_109_47#_c_778_n N_VGND_c_920_n 0.00133167f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_488 N_A_109_47#_c_778_n N_VGND_c_922_n 0.0013116f $X=6.09 $Y=0.85 $X2=0 $Y2=0
cc_489 N_A_109_47#_c_778_n N_VGND_c_923_n 0.00617756f $X=6.09 $Y=0.85 $X2=0
+ $Y2=0
cc_490 N_A_109_47#_c_776_n N_VGND_c_924_n 0.0122675f $X=6.995 $Y=0.81 $X2=0
+ $Y2=0
cc_491 N_A_109_47#_c_856_p N_VGND_c_929_n 0.0112671f $X=6.24 $Y=0.42 $X2=0 $Y2=0
cc_492 N_A_109_47#_c_782_n N_VGND_c_929_n 0.0026358f $X=6.45 $Y=0.825 $X2=0
+ $Y2=0
cc_493 N_A_109_47#_c_776_n N_VGND_c_930_n 0.00245083f $X=6.995 $Y=0.81 $X2=0
+ $Y2=0
cc_494 N_A_109_47#_c_777_n N_VGND_c_930_n 0.00413931f $X=7.08 $Y=0.675 $X2=0
+ $Y2=0
cc_495 N_A_109_47#_M1015_s N_VGND_c_932_n 0.00221414f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_496 N_A_109_47#_M1023_s N_VGND_c_932_n 0.00189607f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_497 N_A_109_47#_M1003_s N_VGND_c_932_n 0.00215893f $X=6.105 $Y=0.235 $X2=0
+ $Y2=0
cc_498 N_A_109_47#_M1013_s N_VGND_c_932_n 0.00684785f $X=6.945 $Y=0.235 $X2=0
+ $Y2=0
cc_499 N_A_109_47#_c_856_p N_VGND_c_932_n 0.00295874f $X=6.24 $Y=0.42 $X2=0
+ $Y2=0
cc_500 N_A_109_47#_c_776_n N_VGND_c_932_n 0.00555922f $X=6.995 $Y=0.81 $X2=0
+ $Y2=0
cc_501 N_A_109_47#_c_777_n N_VGND_c_932_n 0.00540999f $X=7.08 $Y=0.675 $X2=0
+ $Y2=0
cc_502 N_A_109_47#_c_778_n N_VGND_c_932_n 0.196992f $X=6.09 $Y=0.85 $X2=0 $Y2=0
cc_503 N_A_109_47#_c_779_n N_VGND_c_932_n 0.0147197f $X=1.76 $Y=0.85 $X2=0 $Y2=0
cc_504 N_A_109_47#_c_780_n N_VGND_c_932_n 0.0147888f $X=6.235 $Y=0.85 $X2=0
+ $Y2=0
cc_505 N_A_109_47#_c_782_n N_VGND_c_932_n 0.00427567f $X=6.45 $Y=0.825 $X2=0
+ $Y2=0
cc_506 N_A_445_47#_c_871_n N_VGND_M1012_s 0.00430513f $X=4.475 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_507 N_A_445_47#_c_882_n N_VGND_M1016_s 0.00273671f $X=5.315 $Y=0.74 $X2=0
+ $Y2=0
cc_508 N_A_445_47#_c_871_n N_VGND_c_920_n 0.0170446f $X=4.475 $Y=0.74 $X2=0
+ $Y2=0
cc_509 N_A_445_47#_c_871_n N_VGND_c_921_n 0.0023303f $X=4.475 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_445_47#_c_906_p N_VGND_c_921_n 0.0112554f $X=4.56 $Y=0.42 $X2=0 $Y2=0
cc_511 N_A_445_47#_c_882_n N_VGND_c_921_n 0.0023303f $X=5.315 $Y=0.74 $X2=0
+ $Y2=0
cc_512 N_A_445_47#_c_882_n N_VGND_c_922_n 0.0131836f $X=5.315 $Y=0.74 $X2=0
+ $Y2=0
cc_513 N_A_445_47#_c_871_n N_VGND_c_926_n 0.00332039f $X=4.475 $Y=0.74 $X2=0
+ $Y2=0
cc_514 N_A_445_47#_c_882_n N_VGND_c_928_n 0.0023303f $X=5.315 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_445_47#_c_911_p N_VGND_c_928_n 0.0112554f $X=5.4 $Y=0.42 $X2=0 $Y2=0
cc_516 N_A_445_47#_M1019_d N_VGND_c_932_n 0.00181381f $X=2.225 $Y=0.235 $X2=0
+ $Y2=0
cc_517 N_A_445_47#_M1028_d N_VGND_c_932_n 0.00181381f $X=3.065 $Y=0.235 $X2=0
+ $Y2=0
cc_518 N_A_445_47#_M1012_d N_VGND_c_932_n 0.00198522f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_519 N_A_445_47#_M1020_d N_VGND_c_932_n 0.00226669f $X=5.265 $Y=0.235 $X2=0
+ $Y2=0
cc_520 N_A_445_47#_c_871_n N_VGND_c_932_n 0.00779802f $X=4.475 $Y=0.74 $X2=0
+ $Y2=0
cc_521 N_A_445_47#_c_906_p N_VGND_c_932_n 0.00305234f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_522 N_A_445_47#_c_882_n N_VGND_c_932_n 0.00445205f $X=5.315 $Y=0.74 $X2=0
+ $Y2=0
cc_523 N_A_445_47#_c_911_p N_VGND_c_932_n 0.00305234f $X=5.4 $Y=0.42 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s18_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
M1000 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=6.814e+11p pd=5.94e+06u as=1.134e+11p ps=1.38e+06u
M1001 VGND a_334_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1002 VPWR a_334_47# X VPB phighvt w=1e+06u l=150000u
+  ad=1.1825e+12p pd=8.5e+06u as=2.8e+11p ps=2.56e+06u
M1003 a_227_47# a_27_47# VGND VNB nshort w=650000u l=180000u
+  ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1004 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 VGND a_227_47# a_334_47# VNB nshort w=650000u l=180000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1006 X a_334_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_227_47# a_334_47# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=2.173e+11p ps=2.17e+06u
M1008 X a_334_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_227_47# a_27_47# VPWR VPB phighvt w=820000u l=180000u
+  ad=2.173e+11p pd=2.17e+06u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__a2111o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 0.955000 3.775000 1.740000 ;
        RECT 3.505000 0.290000 3.995000 0.825000 ;
        RECT 3.505000 0.825000 3.775000 0.955000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945000 0.995000 4.515000 1.740000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.995000 3.195000 1.740000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 0.995000 2.735000 2.355000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.995000 2.255000 1.325000 ;
        RECT 1.960000 1.325000 2.255000 2.355000 ;
    END
  END D1
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.255000 0.895000 2.390000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.085000 0.435000 0.885000 ;
      RECT 0.085000  1.635000 0.435000 2.635000 ;
      RECT 1.065000  0.085000 2.010000 0.445000 ;
      RECT 1.065000  0.445000 1.325000 0.865000 ;
      RECT 1.065000  1.075000 1.705000 1.325000 ;
      RECT 1.065000  1.495000 1.315000 2.635000 ;
      RECT 1.495000  0.615000 3.335000 0.785000 ;
      RECT 1.495000  0.785000 1.705000 1.075000 ;
      RECT 1.495000  1.325000 1.705000 1.495000 ;
      RECT 1.495000  1.495000 1.785000 2.465000 ;
      RECT 2.180000  0.255000 2.420000 0.615000 ;
      RECT 2.590000  0.085000 2.920000 0.445000 ;
      RECT 3.070000  1.915000 4.515000 2.085000 ;
      RECT 3.070000  2.085000 3.400000 2.465000 ;
      RECT 3.090000  0.255000 3.335000 0.615000 ;
      RECT 3.590000  2.255000 3.920000 2.635000 ;
      RECT 4.090000  2.085000 4.515000 2.465000 ;
      RECT 4.165000  0.085000 4.515000 0.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111o_2
END LIBRARY

* NGSPICE file created from sky130_fd_sc_hd__o311ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 VGND A2 a_138_47# VNB nshort w=650000u l=150000u
+  ad=3.575e+11p pd=3.7e+06u as=5.72e+11p ps=4.36e+06u
M1001 Y A3 a_222_297# VPB phighvt w=1e+06u l=150000u
+  ad=7.6e+11p pd=5.52e+06u as=2.7e+11p ps=2.54e+06u
M1002 a_222_297# A2 a_138_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 a_138_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1005 Y C1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_138_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C1 a_458_47# VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=1.365e+11p ps=1.72e+06u
M1008 a_458_47# B1 a_138_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_138_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


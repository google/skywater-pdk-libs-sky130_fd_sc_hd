* File: sky130_fd_sc_hd__inv_6.pxi.spice
* Created: Thu Aug 27 14:22:53 2020
* 
x_PM_SKY130_FD_SC_HD__INV_6%A N_A_c_52_n N_A_M1004_g N_A_M1000_g N_A_c_53_n
+ N_A_M1005_g N_A_M1001_g N_A_c_54_n N_A_M1007_g N_A_M1002_g N_A_c_55_n
+ N_A_M1008_g N_A_M1003_g N_A_c_56_n N_A_M1010_g N_A_M1006_g N_A_c_57_n
+ N_A_M1011_g N_A_M1009_g A A A A N_A_c_59_n N_A_c_60_n
+ PM_SKY130_FD_SC_HD__INV_6%A
x_PM_SKY130_FD_SC_HD__INV_6%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_M1009_d N_VPWR_c_162_n N_VPWR_c_163_n N_VPWR_c_164_n N_VPWR_c_165_n
+ N_VPWR_c_166_n N_VPWR_c_167_n N_VPWR_c_168_n N_VPWR_c_169_n N_VPWR_c_170_n
+ VPWR N_VPWR_c_171_n N_VPWR_c_172_n N_VPWR_c_161_n
+ PM_SKY130_FD_SC_HD__INV_6%VPWR
x_PM_SKY130_FD_SC_HD__INV_6%Y N_Y_M1004_d N_Y_M1007_d N_Y_M1010_d N_Y_M1000_s
+ N_Y_M1002_s N_Y_M1006_s N_Y_c_220_n N_Y_c_224_n N_Y_c_298_p N_Y_c_212_n
+ N_Y_c_213_n N_Y_c_234_n N_Y_c_238_n N_Y_c_293_p N_Y_c_214_n N_Y_c_246_n
+ N_Y_c_301_p N_Y_c_249_n N_Y_c_215_n Y Y Y N_Y_c_217_n N_Y_c_219_n N_Y_c_266_n
+ PM_SKY130_FD_SC_HD__INV_6%Y
x_PM_SKY130_FD_SC_HD__INV_6%VGND N_VGND_M1004_s N_VGND_M1005_s N_VGND_M1008_s
+ N_VGND_M1011_s N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n
+ N_VGND_c_315_n N_VGND_c_316_n N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n
+ VGND N_VGND_c_320_n N_VGND_c_321_n N_VGND_c_322_n
+ PM_SKY130_FD_SC_HD__INV_6%VGND
cc_1 VNB N_A_c_52_n 0.0219754f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=0.995
cc_2 VNB N_A_c_53_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=1.06 $Y2=0.995
cc_3 VNB N_A_c_54_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_4 VNB N_A_c_55_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_5 VNB N_A_c_56_n 0.0157808f $X=-0.19 $Y=-0.24 $X2=2.32 $Y2=0.995
cc_6 VNB N_A_c_57_n 0.0189107f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=0.995
cc_7 VNB A 0.00932659f $X=-0.19 $Y=-0.24 $X2=2.405 $Y2=1.105
cc_8 VNB N_A_c_59_n 0.0438762f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.16
cc_9 VNB N_A_c_60_n 0.0933498f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=1.16
cc_10 VNB N_VPWR_c_161_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_11 VNB N_Y_c_212_n 0.00308196f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.985
cc_12 VNB N_Y_c_213_n 0.00148844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_Y_c_214_n 0.00308196f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=1.325
cc_14 VNB N_Y_c_215_n 0.00126815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB Y 0.0179825f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.16
cc_16 VNB N_Y_c_217_n 0.0112303f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=1.16
cc_17 VNB N_VGND_c_311_n 0.011417f $X=-0.19 $Y=-0.24 $X2=1.06 $Y2=1.985
cc_18 VNB N_VGND_c_312_n 0.0176196f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_19 VNB N_VGND_c_313_n 0.00419608f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=1.985
cc_20 VNB N_VGND_c_314_n 0.0178019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_315_n 0.00358448f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.325
cc_22 VNB N_VGND_c_316_n 0.0112684f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.985
cc_23 VNB N_VGND_c_317_n 0.00229341f $X=-0.19 $Y=-0.24 $X2=2.32 $Y2=0.995
cc_24 VNB N_VGND_c_318_n 0.0225579f $X=-0.19 $Y=-0.24 $X2=2.32 $Y2=0.56
cc_25 VNB N_VGND_c_319_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=2.32 $Y2=1.325
cc_26 VNB N_VGND_c_320_n 0.0145246f $X=-0.19 $Y=-0.24 $X2=2.74 $Y2=1.325
cc_27 VNB N_VGND_c_321_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_322_n 0.181603f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_29 VPB N_A_M1000_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.985
cc_30 VPB N_A_M1001_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.985
cc_31 VPB N_A_M1002_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.985
cc_32 VPB N_A_M1003_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.985
cc_33 VPB N_A_M1006_g 0.0184947f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=1.985
cc_34 VPB N_A_M1009_g 0.0230192f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=1.985
cc_35 VPB A 7.73822e-19 $X=-0.19 $Y=1.305 $X2=2.405 $Y2=1.105
cc_36 VPB N_A_c_59_n 0.0170655f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_37 VPB N_A_c_60_n 0.0162192f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=1.16
cc_38 VPB N_VPWR_c_162_n 0.0119961f $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.985
cc_39 VPB N_VPWR_c_163_n 0.0418654f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_40 VPB N_VPWR_c_164_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_165_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_42 VPB N_VPWR_c_166_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.985
cc_43 VPB N_VPWR_c_167_n 0.0113416f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=0.995
cc_44 VPB N_VPWR_c_168_n 0.00416524f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=0.56
cc_45 VPB N_VPWR_c_169_n 0.0208097f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=1.985
cc_46 VPB N_VPWR_c_170_n 0.00323736f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=1.985
cc_47 VPB N_VPWR_c_171_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.74 $Y2=1.985
cc_48 VPB N_VPWR_c_172_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_161_n 0.046138f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_50 VPB Y 0.00821566f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.16
cc_51 VPB N_Y_c_219_n 0.00985087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_A_M1000_g N_VPWR_c_163_n 0.0252634f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_53 A N_VPWR_c_163_n 0.023743f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A_c_59_n N_VPWR_c_163_n 0.00682563f $X=0.565 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_M1001_g N_VPWR_c_164_n 0.00268723f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_56 N_A_M1002_g N_VPWR_c_164_n 0.00146448f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A_M1002_g N_VPWR_c_165_n 0.00541359f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_58 N_A_M1003_g N_VPWR_c_165_n 0.00541359f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_VPWR_c_166_n 0.00146448f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_60 N_A_M1006_g N_VPWR_c_166_n 0.00146448f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_M1009_g N_VPWR_c_168_n 0.00316354f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VPWR_c_169_n 0.00541359f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_M1001_g N_VPWR_c_169_n 0.00541359f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_64 N_A_M1006_g N_VPWR_c_171_n 0.00541359f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_65 N_A_M1009_g N_VPWR_c_171_n 0.00541359f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1000_g N_VPWR_c_161_n 0.0108239f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_VPWR_c_161_n 0.00950154f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_M1002_g N_VPWR_c_161_n 0.00950154f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A_M1003_g N_VPWR_c_161_n 0.00950154f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A_M1006_g N_VPWR_c_161_n 0.00950154f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_M1009_g N_VPWR_c_161_n 0.0104652f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_Y_c_220_n 0.00269551f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A_M1001_g N_Y_c_220_n 8.84614e-19 $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_74 A N_Y_c_220_n 0.0213676f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_60_n N_Y_c_220_n 0.00209661f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_Y_c_224_n 0.0108991f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_M1001_g N_Y_c_224_n 0.00975139f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1002_g N_Y_c_224_n 6.1949e-19 $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_c_53_n N_Y_c_212_n 0.0119895f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_c_54_n N_Y_c_212_n 0.0124475f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_81 A N_Y_c_212_n 0.0483239f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A_c_60_n N_Y_c_212_n 0.00222133f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_c_52_n N_Y_c_213_n 0.00126679f $X=0.64 $Y=0.995 $X2=0 $Y2=0
cc_84 A N_Y_c_213_n 0.0140175f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_85 N_A_c_60_n N_Y_c_213_n 0.00230339f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_M1001_g N_Y_c_234_n 0.0107189f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_Y_c_234_n 0.0107189f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_88 A N_Y_c_234_n 0.0320704f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A_c_60_n N_Y_c_234_n 0.00201785f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_Y_c_238_n 6.1949e-19 $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_Y_c_238_n 0.00975139f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_M1003_g N_Y_c_238_n 0.00973632f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_M1006_g N_Y_c_238_n 6.21474e-19 $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_c_55_n N_Y_c_214_n 0.0124942f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_c_56_n N_Y_c_214_n 0.0124942f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_96 A N_Y_c_214_n 0.0608913f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_97 N_A_c_60_n N_Y_c_214_n 0.00222133f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_M1003_g N_Y_c_246_n 5.61575e-19 $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_M1006_g N_Y_c_246_n 0.00950901f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_M1009_g N_Y_c_246_n 0.0249522f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_M1002_g N_Y_c_249_n 8.84614e-19 $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_M1003_g N_Y_c_249_n 8.84614e-19 $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_103 A N_Y_c_249_n 0.0213676f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A_c_60_n N_Y_c_249_n 0.00209661f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_105 A N_Y_c_215_n 0.0140175f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_106 N_A_c_60_n N_Y_c_215_n 0.00230339f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_c_56_n Y 4.3959e-19 $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_M1006_g Y 8.13266e-19 $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_c_57_n Y 0.00357285f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_M1009_g Y 0.00670223f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_111 A Y 0.0198811f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_112 N_A_c_60_n Y 0.0150247f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_c_57_n N_Y_c_217_n 0.0149435f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_c_60_n N_Y_c_217_n 0.00222133f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_M1006_g N_Y_c_219_n 0.00128027f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_M1009_g N_Y_c_219_n 0.0152528f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_c_60_n N_Y_c_219_n 0.00202298f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_M1003_g N_Y_c_266_n 0.0107189f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_M1006_g N_Y_c_266_n 0.0107189f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_120 A N_Y_c_266_n 0.0478206f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A_c_60_n N_Y_c_266_n 0.00201785f $X=2.74 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_c_52_n N_VGND_c_312_n 0.0106174f $X=0.64 $Y=0.995 $X2=0 $Y2=0
cc_123 A N_VGND_c_312_n 0.00883493f $X=2.405 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_c_59_n N_VGND_c_312_n 0.00524994f $X=0.565 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_53_n N_VGND_c_313_n 0.00268723f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_54_n N_VGND_c_313_n 0.00146448f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_54_n N_VGND_c_314_n 0.00437852f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_55_n N_VGND_c_314_n 0.00437852f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_55_n N_VGND_c_315_n 0.00146448f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_56_n N_VGND_c_315_n 0.00137415f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_56_n N_VGND_c_317_n 5.60631e-19 $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_57_n N_VGND_c_317_n 0.00865f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_52_n N_VGND_c_318_n 0.00585385f $X=0.64 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_53_n N_VGND_c_318_n 0.00437852f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_56_n N_VGND_c_320_n 0.00437852f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_57_n N_VGND_c_320_n 0.00349488f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_52_n N_VGND_c_322_n 0.0118594f $X=0.64 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_c_53_n N_VGND_c_322_n 0.00588671f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_c_54_n N_VGND_c_322_n 0.00588671f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_55_n N_VGND_c_322_n 0.00588671f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_c_56_n N_VGND_c_322_n 0.00588671f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_57_n N_VGND_c_322_n 0.00412119f $X=2.74 $Y=0.995 $X2=0 $Y2=0
cc_143 N_VPWR_c_161_n N_Y_M1000_s 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_144 N_VPWR_c_161_n N_Y_M1002_s 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_145 N_VPWR_c_161_n N_Y_M1006_s 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_146 N_VPWR_c_163_n N_Y_c_220_n 0.0100071f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_147 N_VPWR_c_163_n N_Y_c_224_n 0.0444181f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_148 N_VPWR_c_169_n N_Y_c_224_n 0.0189039f $X=1.185 $Y=2.72 $X2=0 $Y2=0
cc_149 N_VPWR_c_161_n N_Y_c_224_n 0.0122217f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_150 N_VPWR_M1001_d N_Y_c_234_n 0.00311483f $X=1.135 $Y=1.485 $X2=0 $Y2=0
cc_151 N_VPWR_c_164_n N_Y_c_234_n 0.0126919f $X=1.27 $Y=2 $X2=0 $Y2=0
cc_152 N_VPWR_c_165_n N_Y_c_238_n 0.0189039f $X=2.025 $Y=2.72 $X2=0 $Y2=0
cc_153 N_VPWR_c_161_n N_Y_c_238_n 0.0122217f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_c_171_n N_Y_c_246_n 0.0189039f $X=2.865 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_161_n N_Y_c_246_n 0.0122217f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_M1009_d Y 6.79636e-19 $X=2.815 $Y=1.485 $X2=0 $Y2=0
cc_157 N_VPWR_M1009_d N_Y_c_219_n 0.00644124f $X=2.815 $Y=1.485 $X2=0 $Y2=0
cc_158 N_VPWR_c_168_n N_Y_c_219_n 0.00601237f $X=2.95 $Y=2.34 $X2=0 $Y2=0
cc_159 N_VPWR_M1003_d N_Y_c_266_n 0.00311483f $X=1.975 $Y=1.485 $X2=0 $Y2=0
cc_160 N_VPWR_c_166_n N_Y_c_266_n 0.0126919f $X=2.11 $Y=2 $X2=0 $Y2=0
cc_161 N_Y_c_212_n N_VGND_M1005_s 0.001659f $X=1.605 $Y=0.815 $X2=0 $Y2=0
cc_162 N_Y_c_214_n N_VGND_M1008_s 0.001659f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_163 N_Y_c_217_n N_VGND_M1011_s 0.00345636f $X=2.96 $Y=0.905 $X2=0 $Y2=0
cc_164 N_Y_c_212_n N_VGND_c_313_n 0.0116647f $X=1.605 $Y=0.815 $X2=0 $Y2=0
cc_165 N_Y_c_212_n N_VGND_c_314_n 0.00278354f $X=1.605 $Y=0.815 $X2=0 $Y2=0
cc_166 N_Y_c_293_p N_VGND_c_314_n 0.0113595f $X=1.69 $Y=0.42 $X2=0 $Y2=0
cc_167 N_Y_c_214_n N_VGND_c_314_n 0.00278354f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_168 N_Y_c_214_n N_VGND_c_315_n 0.0116647f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_169 N_Y_c_217_n N_VGND_c_316_n 0.00149611f $X=2.96 $Y=0.905 $X2=0 $Y2=0
cc_170 N_Y_c_217_n N_VGND_c_317_n 0.0144491f $X=2.96 $Y=0.905 $X2=0 $Y2=0
cc_171 N_Y_c_298_p N_VGND_c_318_n 0.0113595f $X=0.85 $Y=0.42 $X2=0 $Y2=0
cc_172 N_Y_c_212_n N_VGND_c_318_n 0.00278354f $X=1.605 $Y=0.815 $X2=0 $Y2=0
cc_173 N_Y_c_214_n N_VGND_c_320_n 0.00479168f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_174 N_Y_c_301_p N_VGND_c_320_n 0.0111061f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_175 N_Y_M1004_d N_VGND_c_322_n 0.00412336f $X=0.715 $Y=0.235 $X2=0 $Y2=0
cc_176 N_Y_M1007_d N_VGND_c_322_n 0.00262315f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_177 N_Y_M1010_d N_VGND_c_322_n 0.00264915f $X=2.395 $Y=0.235 $X2=0 $Y2=0
cc_178 N_Y_c_298_p N_VGND_c_322_n 0.0064623f $X=0.85 $Y=0.42 $X2=0 $Y2=0
cc_179 N_Y_c_212_n N_VGND_c_322_n 0.0122342f $X=1.605 $Y=0.815 $X2=0 $Y2=0
cc_180 N_Y_c_293_p N_VGND_c_322_n 0.0064623f $X=1.69 $Y=0.42 $X2=0 $Y2=0
cc_181 N_Y_c_214_n N_VGND_c_322_n 0.016186f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_182 N_Y_c_301_p N_VGND_c_322_n 0.00640911f $X=2.53 $Y=0.42 $X2=0 $Y2=0
cc_183 N_Y_c_217_n N_VGND_c_322_n 0.00363552f $X=2.96 $Y=0.905 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a32o_1.spice.pex
* Created: Thu Aug 27 14:05:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A32O_1%A_93_21# 1 2 9 12 17 18 19 20 21 23 24 26 30
+ 33 34 35 38
r95 34 39 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.627 $Y=1.16
+ $X2=0.627 $Y2=1.325
r96 34 38 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.627 $Y=1.16
+ $X2=0.627 $Y2=0.995
r97 33 36 8.47458 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.722 $Y=1.16
+ $X2=0.722 $Y2=1.325
r98 33 35 8.47458 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.722 $Y=1.16
+ $X2=0.722 $Y2=0.995
r99 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.655
+ $Y=1.16 $X2=0.655 $Y2=1.16
r100 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=1.665
+ $X2=2.99 $Y2=1.96
r101 24 26 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=1.265 $Y=0.4
+ $X2=2.545 $Y2=0.4
r102 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=0.485
+ $X2=1.265 $Y2=0.4
r103 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.18 $Y=0.485
+ $X2=1.18 $Y2=0.655
r104 20 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=1.58
+ $X2=2.99 $Y2=1.665
r105 20 21 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=2.905 $Y=1.58
+ $X2=0.875 $Y2=1.58
r106 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.095 $Y=0.74
+ $X2=1.18 $Y2=0.655
r107 18 19 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.095 $Y=0.74
+ $X2=0.875 $Y2=0.74
r108 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.79 $Y=1.495
+ $X2=0.875 $Y2=1.58
r109 17 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.79 $Y=1.495
+ $X2=0.79 $Y2=1.325
r110 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.79 $Y=0.825
+ $X2=0.875 $Y2=0.74
r111 14 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.79 $Y=0.825
+ $X2=0.79 $Y2=0.995
r112 12 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.54 $Y=1.985
+ $X2=0.54 $Y2=1.325
r113 9 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.56
+ $X2=0.54 $Y2=0.995
r114 2 30 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.485 $X2=2.99 $Y2=1.96
r115 1 26 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.235 $X2=2.545 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%A3 3 7 8 11 13
r37 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.235 $Y=1.16
+ $X2=1.235 $Y2=1.325
r38 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.235 $Y=1.16
+ $X2=1.235 $Y2=0.995
r39 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.235
+ $Y=1.16 $X2=1.235 $Y2=1.16
r40 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.205 $Y=0.56
+ $X2=1.205 $Y2=0.995
r41 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.175 $Y=1.985
+ $X2=1.175 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%A2 3 6 8 9 13 15
r37 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.16
+ $X2=1.715 $Y2=1.325
r38 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.16
+ $X2=1.715 $Y2=0.995
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.715
+ $Y=1.16 $X2=1.715 $Y2=1.16
r40 9 14 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=1.665 $Y=1.19 $X2=1.665
+ $Y2=1.16
r41 8 14 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.665 $Y=0.85
+ $X2=1.665 $Y2=1.16
r42 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.655 $Y=1.985
+ $X2=1.655 $Y2=1.325
r43 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.655 $Y=0.56
+ $X2=1.655 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%A1 3 6 8 9 13 15
r34 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.16
+ $X2=2.195 $Y2=1.325
r35 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.16
+ $X2=2.195 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.195
+ $Y=1.16 $X2=2.195 $Y2=1.16
r37 9 14 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=2.135 $Y=1.19 $X2=2.135
+ $Y2=1.16
r38 8 14 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.135 $Y=0.85
+ $X2=2.135 $Y2=1.16
r39 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.255 $Y=1.985
+ $X2=2.255 $Y2=1.325
r40 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.255 $Y=0.56
+ $X2=2.255 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%B1 3 7 8 9 13 15
r35 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.16
+ $X2=2.785 $Y2=1.325
r36 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.16
+ $X2=2.785 $Y2=0.995
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=1.16 $X2=2.785 $Y2=1.16
r38 9 14 0.823174 $w=4.18e-07 $l=3e-08 $layer=LI1_cond $X=2.66 $Y=1.19 $X2=2.66
+ $Y2=1.16
r39 8 14 8.50613 $w=4.18e-07 $l=3.1e-07 $layer=LI1_cond $X=2.66 $Y=0.85 $X2=2.66
+ $Y2=1.16
r40 7 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.845 $Y=0.56
+ $X2=2.845 $Y2=0.995
r41 3 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.775 $Y=1.985
+ $X2=2.775 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%B2 3 6 8 9 13 15
r24 17 23 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=3.427 $Y=1.325
+ $X2=3.427 $Y2=1.16
r25 14 23 5.65745 $w=3.28e-07 $l=1.62e-07 $layer=LI1_cond $X=3.265 $Y=1.16
+ $X2=3.427 $Y2=1.16
r26 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.265 $Y=1.16
+ $X2=3.265 $Y2=1.325
r27 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.265 $Y=1.16
+ $X2=3.265 $Y2=0.995
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.265
+ $Y=1.16 $X2=3.265 $Y2=1.16
r29 9 17 11.0909 $w=2.03e-07 $l=2.05e-07 $layer=LI1_cond $X=3.427 $Y=1.53
+ $X2=3.427 $Y2=1.325
r30 8 23 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=3.445 $Y=1.16
+ $X2=3.427 $Y2=1.16
r31 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.205 $Y=1.985
+ $X2=3.205 $Y2=1.325
r32 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.205 $Y=0.56
+ $X2=3.205 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%X 1 2 7 8 9 10 11 12 36 42 46
r18 46 47 2.40535 $w=3.33e-07 $l=5e-08 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.56
r19 36 49 2.03372 $w=2.53e-07 $l=4.5e-08 $layer=LI1_cond $X=0.217 $Y=1.87
+ $X2=0.217 $Y2=1.915
r20 12 37 4.40336 $w=3.33e-07 $l=1.28e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.082
r21 11 37 5.05699 $w=3.33e-07 $l=1.47e-07 $layer=LI1_cond $X=0.257 $Y=1.935
+ $X2=0.257 $Y2=2.082
r22 11 49 1.37331 $w=3.33e-07 $l=2e-08 $layer=LI1_cond $X=0.257 $Y=1.935
+ $X2=0.257 $Y2=1.915
r23 11 36 0.903877 $w=2.53e-07 $l=2e-08 $layer=LI1_cond $X=0.217 $Y=1.85
+ $X2=0.217 $Y2=1.87
r24 11 33 8.58683 $w=2.53e-07 $l=1.9e-07 $layer=LI1_cond $X=0.217 $Y=1.85
+ $X2=0.217 $Y2=1.66
r25 10 33 5.8752 $w=2.53e-07 $l=1.3e-07 $layer=LI1_cond $X=0.217 $Y=1.53
+ $X2=0.217 $Y2=1.66
r26 9 10 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.217 $Y=1.19
+ $X2=0.217 $Y2=1.53
r27 8 9 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.217 $Y2=1.19
r28 8 25 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.217 $Y2=0.725
r29 7 46 0.619223 $w=3.33e-07 $l=1.8e-08 $layer=LI1_cond $X=0.257 $Y=0.492
+ $X2=0.257 $Y2=0.51
r30 7 42 3.68094 $w=3.33e-07 $l=1.07e-07 $layer=LI1_cond $X=0.257 $Y=0.492
+ $X2=0.257 $Y2=0.385
r31 7 25 6.68869 $w=2.53e-07 $l=1.48e-07 $layer=LI1_cond $X=0.217 $Y=0.577
+ $X2=0.217 $Y2=0.725
r32 7 47 0.768295 $w=2.53e-07 $l=1.7e-08 $layer=LI1_cond $X=0.217 $Y=0.577
+ $X2=0.217 $Y2=0.56
r33 2 11 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
r34 2 33 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r35 1 42 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.385
r36 1 25 182 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%VPWR 1 2 11 15 17 19 26 27 30 33
r53 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 27 34 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=2.72
+ $X2=1.955 $Y2=2.72
r58 24 26 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=2.12 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 23 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 20 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=0.84 $Y2=2.72
r63 20 22 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=2.72
+ $X2=1.955 $Y2=2.72
r65 19 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.79 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 17 31 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=2.635
+ $X2=1.955 $Y2=2.72
r68 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.955 $Y=2.635
+ $X2=1.955 $Y2=2.34
r69 9 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=2.635 $X2=0.84
+ $Y2=2.72
r70 9 11 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.84 $Y=2.635
+ $X2=0.84 $Y2=2
r71 2 15 600 $w=1.7e-07 $l=9.60937e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=1.485 $X2=1.955 $Y2=2.34
r72 1 11 300 $w=1.7e-07 $l=6.17333e-07 $layer=licon1_PDIFF $count=2 $X=0.615
+ $Y=1.485 $X2=0.84 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%A_250_297# 1 2 3 10 12 14 16 18 19 22
r31 20 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.42 $Y=2.295
+ $X2=3.42 $Y2=1.96
r32 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=2.38
+ $X2=3.42 $Y2=2.295
r33 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.335 $Y=2.38
+ $X2=2.675 $Y2=2.38
r34 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.51 $Y=2.295
+ $X2=2.675 $Y2=2.38
r35 16 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=2.045 $X2=2.51
+ $Y2=1.96
r36 16 17 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.51 $Y=2.045
+ $X2=2.51 $Y2=2.295
r37 15 25 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.535 $Y=1.96
+ $X2=1.392 $Y2=1.96
r38 14 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=1.96
+ $X2=2.51 $Y2=1.96
r39 14 15 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.345 $Y=1.96
+ $X2=1.535 $Y2=1.96
r40 10 25 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.392 $Y=2.045
+ $X2=1.392 $Y2=1.96
r41 10 12 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=1.392 $Y=2.045
+ $X2=1.392 $Y2=2.3
r42 3 22 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=1.485 $X2=3.42 $Y2=1.96
r43 2 27 300 $w=1.7e-07 $l=5.98268e-07 $layer=licon1_PDIFF $count=2 $X=2.33
+ $Y=1.485 $X2=2.51 $Y2=2
r44 1 25 600 $w=1.7e-07 $l=5.51362e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.485 $X2=1.415 $Y2=1.96
r45 1 12 600 $w=1.7e-07 $l=8.937e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.485 $X2=1.415 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_1%VGND 1 2 9 11 13 15 17 22 31 35
r50 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r51 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r53 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r54 26 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r55 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r56 25 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r57 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.76
+ $Y2=0
r59 23 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.15
+ $Y2=0
r60 22 34 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.467
+ $Y2=0
r61 22 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r62 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.76
+ $Y2=0
r63 17 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r64 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r65 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 11 34 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.467 $Y2=0
r67 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.38
r68 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0
r69 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.4
r70 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.28
+ $Y=0.235 $X2=3.42 $Y2=0.38
r71 1 9 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.76 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__a21oi_1.pxi.spice
* Created: Thu Aug 27 14:01:16 2020
* 
x_PM_SKY130_FD_SC_HD__A21OI_1%B1 N_B1_c_38_n N_B1_M1003_g N_B1_M1002_g B1 B1
+ N_B1_c_40_n PM_SKY130_FD_SC_HD__A21OI_1%B1
x_PM_SKY130_FD_SC_HD__A21OI_1%A1 N_A1_M1005_g N_A1_M1004_g A1 A1 A1 N_A1_c_69_n
+ N_A1_c_70_n PM_SKY130_FD_SC_HD__A21OI_1%A1
x_PM_SKY130_FD_SC_HD__A21OI_1%A2 N_A2_c_106_n N_A2_M1001_g N_A2_M1000_g A2
+ N_A2_c_108_n PM_SKY130_FD_SC_HD__A21OI_1%A2
x_PM_SKY130_FD_SC_HD__A21OI_1%Y N_Y_M1003_d N_Y_M1002_s N_Y_c_133_n N_Y_c_135_n
+ N_Y_c_157_p N_Y_c_143_n Y Y PM_SKY130_FD_SC_HD__A21OI_1%Y
x_PM_SKY130_FD_SC_HD__A21OI_1%A_113_297# N_A_113_297#_M1002_d
+ N_A_113_297#_M1000_d N_A_113_297#_c_165_n N_A_113_297#_c_164_n
+ N_A_113_297#_c_162_n N_A_113_297#_c_163_n
+ PM_SKY130_FD_SC_HD__A21OI_1%A_113_297#
x_PM_SKY130_FD_SC_HD__A21OI_1%VPWR N_VPWR_M1004_d N_VPWR_c_192_n VPWR
+ N_VPWR_c_193_n N_VPWR_c_194_n N_VPWR_c_191_n N_VPWR_c_196_n
+ PM_SKY130_FD_SC_HD__A21OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A21OI_1%VGND N_VGND_M1003_s N_VGND_M1001_d N_VGND_c_219_n
+ N_VGND_c_220_n N_VGND_c_221_n N_VGND_c_222_n VGND N_VGND_c_223_n
+ N_VGND_c_224_n PM_SKY130_FD_SC_HD__A21OI_1%VGND
cc_1 VNB N_B1_c_38_n 0.0180023f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB B1 0.0240495f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B1_c_40_n 0.0366992f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_4 VNB A1 0.00237744f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_5 VNB A1 0.00241688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A1_c_69_n 0.0220581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A1_c_70_n 0.0167491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A2_c_106_n 0.0224156f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_9 VNB A2 0.011652f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_10 VNB N_A2_c_108_n 0.0345054f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_11 VNB N_Y_c_133_n 0.00267358f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_12 VNB N_VPWR_c_191_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=0.85
cc_13 VNB N_VGND_c_219_n 0.010754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_220_n 0.0123169f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_15 VNB N_VGND_c_221_n 0.0110018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_222_n 0.0278608f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_17 VNB N_VGND_c_223_n 0.0265996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_224_n 0.12296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VPB N_B1_M1002_g 0.0254851f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_20 VPB B1 0.00295004f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_21 VPB N_B1_c_40_n 0.0102765f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_22 VPB N_A1_M1004_g 0.0195193f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_23 VPB A1 0.0019321f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_A1_c_69_n 0.00430826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_A2_M1000_g 0.026592f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_26 VPB A2 9.93507e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_27 VPB N_A2_c_108_n 0.00839f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_28 VPB N_Y_c_133_n 0.00164814f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_29 VPB N_Y_c_135_n 0.00838917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB Y 0.0301226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_113_297#_c_162_n 0.0216381f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_A_113_297#_c_163_n 0.0168665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_192_n 0.00480811f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_34 VPB N_VPWR_c_193_n 0.0290088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_194_n 0.0176368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_191_n 0.0441211f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=0.85
cc_37 VPB N_VPWR_c_196_n 0.00372273f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.16
cc_38 N_B1_M1002_g N_A1_M1004_g 0.0239045f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_39 N_B1_c_40_n A1 3.13443e-19 $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_40 N_B1_c_40_n N_A1_c_69_n 0.0166148f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_41 N_B1_c_38_n N_A1_c_70_n 0.0211138f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_42 N_B1_c_38_n N_Y_c_133_n 0.00329281f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_43 N_B1_M1002_g N_Y_c_133_n 0.00860803f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_44 N_B1_c_40_n N_Y_c_133_n 0.00820724f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_45 N_B1_M1002_g N_Y_c_135_n 0.0164668f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_46 B1 N_Y_c_135_n 0.0188975f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_47 N_B1_c_40_n N_Y_c_135_n 0.00369264f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_48 N_B1_c_38_n N_Y_c_143_n 0.00547826f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_49 B1 N_Y_c_143_n 0.0467653f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_50 N_B1_M1002_g N_A_113_297#_c_164_n 0.00750868f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_51 N_B1_M1002_g N_VPWR_c_193_n 0.0054778f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_52 N_B1_M1002_g N_VPWR_c_191_n 0.0109105f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_53 B1 N_VGND_M1003_s 0.0052051f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_54 B1 N_VGND_c_219_n 2.61981e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_55 N_B1_c_38_n N_VGND_c_220_n 0.0096955f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_56 B1 N_VGND_c_220_n 0.0165104f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_B1_c_40_n N_VGND_c_220_n 0.00239977f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_58 N_B1_c_38_n N_VGND_c_223_n 0.00423516f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_59 N_B1_c_38_n N_VGND_c_224_n 0.0063961f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_60 B1 N_VGND_c_224_n 0.00158303f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_61 A1 N_A2_c_106_n 0.00527738f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_62 N_A1_c_70_n N_A2_c_106_n 0.0317591f $X=0.945 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_63 N_A1_M1004_g N_A2_M1000_g 0.0414946f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_64 A1 A2 0.0253572f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A1_c_69_n A2 2.34825e-19 $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_66 A1 N_A2_c_108_n 0.00268901f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A1_c_69_n N_A2_c_108_n 0.0206996f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A1_M1004_g N_Y_c_133_n 0.00355357f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_69 A1 N_Y_c_133_n 0.00631556f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_70 A1 N_Y_c_133_n 0.0252656f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A1_c_69_n N_Y_c_133_n 0.00202728f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A1_c_70_n N_Y_c_133_n 0.00129914f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A1_M1004_g N_Y_c_135_n 0.00177221f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A1_M1004_g N_A_113_297#_c_165_n 0.0168659f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_75 A1 N_A_113_297#_c_165_n 0.0249903f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A1_c_69_n N_A_113_297#_c_165_n 0.00175071f $X=0.945 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A1_M1004_g N_A_113_297#_c_164_n 0.0097318f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_78 A1 N_A_113_297#_c_164_n 0.00140072f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A1_M1004_g N_A_113_297#_c_163_n 5.13631e-19 $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A1_M1004_g N_VPWR_c_192_n 0.00278983f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A1_M1004_g N_VPWR_c_193_n 0.0042139f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A1_M1004_g N_VPWR_c_191_n 0.00581876f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A1_c_70_n N_VGND_c_220_n 0.00122243f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_84 A1 N_VGND_c_223_n 0.00807754f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_85 N_A1_c_70_n N_VGND_c_223_n 0.00585385f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_86 A1 N_VGND_c_224_n 0.00818989f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_87 N_A1_c_70_n N_VGND_c_224_n 0.0109563f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_88 A1 A_199_47# 0.00666314f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_89 N_A2_M1000_g N_A_113_297#_c_165_n 0.021141f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A2_M1000_g N_A_113_297#_c_164_n 5.11169e-19 $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_91 N_A2_M1000_g N_A_113_297#_c_162_n 0.00237594f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_92 A2 N_A_113_297#_c_162_n 0.0196095f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A2_c_108_n N_A_113_297#_c_162_n 0.00600404f $X=1.575 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A2_M1000_g N_A_113_297#_c_163_n 0.00590193f $X=1.365 $Y=1.985 $X2=0
+ $Y2=0
cc_95 N_A2_M1000_g N_VPWR_c_192_n 0.00273631f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A2_M1000_g N_VPWR_c_194_n 0.00422894f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A2_M1000_g N_VPWR_c_191_n 0.00674203f $X=1.365 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A2_c_106_n N_VGND_c_222_n 0.00875894f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_99 A2 N_VGND_c_222_n 0.021221f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A2_c_108_n N_VGND_c_222_n 0.0059591f $X=1.575 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A2_c_106_n N_VGND_c_223_n 0.00585385f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A2_c_106_n N_VGND_c_224_n 0.0116626f $X=1.365 $Y=0.995 $X2=0 $Y2=0
cc_103 N_Y_c_133_n N_A_113_297#_M1002_d 2.84554e-19 $X=0.592 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_104 N_Y_c_135_n N_A_113_297#_M1002_d 0.00253042f $X=0.592 $Y=1.59 $X2=-0.19
+ $Y2=-0.24
cc_105 N_Y_c_135_n N_A_113_297#_c_164_n 0.0202664f $X=0.592 $Y=1.59 $X2=0 $Y2=0
cc_106 Y N_VPWR_c_193_n 0.0177547f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_107 N_Y_M1002_s N_VPWR_c_191_n 0.00374186f $X=0.15 $Y=1.485 $X2=0 $Y2=0
cc_108 Y N_VPWR_c_191_n 0.010464f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_109 N_Y_c_157_p N_VGND_c_223_n 0.0127788f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_110 N_Y_c_143_n N_VGND_c_223_n 0.00145809f $X=0.67 $Y=0.825 $X2=0 $Y2=0
cc_111 N_Y_M1003_d N_VGND_c_224_n 0.00279501f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_112 N_Y_c_157_p N_VGND_c_224_n 0.00851675f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_113 N_Y_c_143_n N_VGND_c_224_n 0.00279001f $X=0.67 $Y=0.825 $X2=0 $Y2=0
cc_114 N_A_113_297#_c_165_n N_VPWR_M1004_d 0.00400065f $X=1.415 $Y=1.775
+ $X2=-0.19 $Y2=1.305
cc_115 N_A_113_297#_c_165_n N_VPWR_c_192_n 0.0151154f $X=1.415 $Y=1.775 $X2=0
+ $Y2=0
cc_116 N_A_113_297#_c_165_n N_VPWR_c_193_n 0.00228062f $X=1.415 $Y=1.775 $X2=0
+ $Y2=0
cc_117 N_A_113_297#_c_164_n N_VPWR_c_193_n 0.0178106f $X=0.87 $Y=1.775 $X2=0
+ $Y2=0
cc_118 N_A_113_297#_c_165_n N_VPWR_c_194_n 0.00236435f $X=1.415 $Y=1.775 $X2=0
+ $Y2=0
cc_119 N_A_113_297#_c_163_n N_VPWR_c_194_n 0.0197891f $X=1.58 $Y=2.33 $X2=0
+ $Y2=0
cc_120 N_A_113_297#_M1002_d N_VPWR_c_191_n 0.00223577f $X=0.565 $Y=1.485 $X2=0
+ $Y2=0
cc_121 N_A_113_297#_M1000_d N_VPWR_c_191_n 0.00213747f $X=1.44 $Y=1.485 $X2=0
+ $Y2=0
cc_122 N_A_113_297#_c_165_n N_VPWR_c_191_n 0.00940406f $X=1.415 $Y=1.775 $X2=0
+ $Y2=0
cc_123 N_A_113_297#_c_164_n N_VPWR_c_191_n 0.0122349f $X=0.87 $Y=1.775 $X2=0
+ $Y2=0
cc_124 N_A_113_297#_c_163_n N_VPWR_c_191_n 0.0123896f $X=1.58 $Y=2.33 $X2=0
+ $Y2=0
cc_125 N_VGND_c_224_n A_199_47# 0.00481717f $X=1.61 $Y=0 $X2=-0.19 $Y2=-0.24

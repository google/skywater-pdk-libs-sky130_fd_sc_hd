* File: sky130_fd_sc_hd__mux2i_2.pex.spice
* Created: Thu Aug 27 14:28:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX2I_2%S 1 3 6 8 10 13 15 17 20 22 23 32
r67 31 32 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r68 29 31 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.89 $Y2=1.16
r69 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r70 26 29 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.515 $Y2=1.16
r71 23 30 1.29787 $w=2.82e-07 $l=3e-08 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.16
r72 22 30 13.4113 $w=2.82e-07 $l=3.1e-07 $layer=LI1_cond $X=0.605 $Y=0.85
+ $X2=0.605 $Y2=1.16
r73 18 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r74 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r75 15 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r76 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r77 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r78 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r79 8 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r80 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r81 4 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r82 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r83 1 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r84 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%A_27_47# 1 2 9 13 17 21 24 27 30 32 34 37 39
+ 40 43 45 50
c95 32 0 1.34758e-19 $X=1.395 $Y=1.24
c96 21 0 1.47556e-19 $X=2.15 $Y=1.985
r97 44 50 65.9856 $w=3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.82 $Y=1.175 $X2=2.15
+ $Y2=1.175
r98 44 47 17.9961 $w=3e-07 $l=9e-08 $layer=POLY_cond $X=1.82 $Y=1.175 $X2=1.73
+ $Y2=1.175
r99 43 45 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=1.2
+ $X2=1.655 $Y2=1.2
r100 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.16 $X2=1.82 $Y2=1.16
r101 39 40 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=2.3
+ $X2=0.215 $Y2=2.135
r102 34 36 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=0.51
+ $X2=0.215 $Y2=0.675
r103 32 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.395 $Y=1.24
+ $X2=1.655 $Y2=1.24
r104 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.31 $Y=1.325
+ $X2=1.395 $Y2=1.24
r105 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.495
r106 28 37 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.26 $Y=1.58
+ $X2=0.172 $Y2=1.58
r107 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.225 $Y=1.58
+ $X2=1.31 $Y2=1.495
r108 27 28 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.225 $Y=1.58
+ $X2=0.26 $Y2=1.58
r109 25 37 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.172 $Y=1.665
+ $X2=0.172 $Y2=1.58
r110 25 40 29.787 $w=1.73e-07 $l=4.7e-07 $layer=LI1_cond $X=0.172 $Y=1.665
+ $X2=0.172 $Y2=2.135
r111 24 37 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.172 $Y=1.495
+ $X2=0.172 $Y2=1.58
r112 24 36 51.9688 $w=1.73e-07 $l=8.2e-07 $layer=LI1_cond $X=0.172 $Y=1.495
+ $X2=0.172 $Y2=0.675
r113 19 50 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.175
r114 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r115 15 50 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.175
r116 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r117 11 47 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.175
r118 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r119 7 47 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.175
r120 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r121 2 39 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.3
r122 1 34 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%A0 1 3 6 8 10 13 15 16 17 27 31
r55 29 31 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.315 $Y=1.16
+ $X2=3.51 $Y2=1.16
r56 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.315
+ $Y=1.16 $X2=3.315 $Y2=1.16
r57 26 29 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.09 $Y=1.16
+ $X2=3.315 $Y2=1.16
r58 26 27 13.7064 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.09 $Y=1.16
+ $X2=3.015 $Y2=1.16
r59 23 27 75.9834 $w=3e-07 $l=3.8e-07 $layer=POLY_cond $X=2.635 $Y=1.145
+ $X2=3.015 $Y2=1.145
r60 17 30 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.315 $Y2=1.175
r61 16 30 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.315 $Y2=1.175
r62 15 16 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=3.015 $Y2=1.175
r63 15 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.635
+ $Y=1.16 $X2=2.635 $Y2=1.16
r64 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=1.325
+ $X2=3.51 $Y2=1.16
r65 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.51 $Y=1.325
+ $X2=3.51 $Y2=1.985
r66 8 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.16
r67 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
r68 4 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.325
+ $X2=3.09 $Y2=1.16
r69 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.09 $Y=1.325 $X2=3.09
+ $Y2=1.985
r70 1 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=1.16
r71 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.09 $Y=0.995 $X2=3.09
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%A1 1 3 6 8 10 13 15 16 23 24
r45 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.55
+ $Y=1.16 $X2=4.55 $Y2=1.16
r46 21 23 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=4.395 $Y=1.16
+ $X2=4.55 $Y2=1.16
r47 19 21 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=3.97 $Y=1.16
+ $X2=4.395 $Y2=1.16
r48 15 16 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=4.472 $Y=1.19
+ $X2=4.472 $Y2=1.53
r49 15 24 1.06379 $w=3.23e-07 $l=3e-08 $layer=LI1_cond $X=4.472 $Y=1.19
+ $X2=4.472 $Y2=1.16
r50 11 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.325
+ $X2=4.395 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.395 $Y=1.325
+ $X2=4.395 $Y2=1.985
r52 8 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=0.995
+ $X2=4.395 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.395 $Y=0.995
+ $X2=4.395 $Y2=0.56
r54 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.97 $Y=1.325
+ $X2=3.97 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.97 $Y=1.325 $X2=3.97
+ $Y2=1.985
r56 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.97 $Y=0.995
+ $X2=3.97 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.97 $Y=0.995 $X2=3.97
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r71 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 46 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r73 44 47 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r74 43 46 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r75 43 44 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r76 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r78 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r79 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r81 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r82 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r84 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 28 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r87 26 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.4 $Y2=2.72
r89 25 43 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.53 $Y2=2.72
r90 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.4 $Y2=2.72
r91 23 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.15 $Y2=2.72
r92 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.52 $Y2=2.72
r93 22 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=2.07 $Y2=2.72
r94 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.52 $Y2=2.72
r95 18 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.635
+ $X2=2.4 $Y2=2.72
r96 18 20 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.4 $Y=2.635
+ $X2=2.4 $Y2=2.34
r97 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r98 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.34
r99 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r100 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r101 3 20 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.34
r102 2 16 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r103 1 12 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%A_193_297# 1 2 7 12 14 16 17
c48 7 0 1.47556e-19 $X=1.565 $Y=1.92
r49 16 17 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=1.605
+ $X2=3.135 $Y2=1.605
r50 14 17 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.735 $Y=1.58
+ $X2=3.135 $Y2=1.58
r51 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.735 $Y2=1.58
r52 11 12 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.835
r53 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.565 $Y=1.92
+ $X2=1.65 $Y2=1.835
r54 7 9 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.565 $Y=1.92 $X2=1.1
+ $Y2=1.92
r55 2 16 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=1.63
r56 1 9 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%A_361_297# 1 2 11 13 16 17
r36 16 17 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.715 $Y=1.96
+ $X2=2.885 $Y2=1.96
r37 13 15 23.4141 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=1.967 $Y=1.92
+ $X2=1.967 $Y2=2.3
r38 11 17 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=4.185 $Y=2 $X2=2.885
+ $Y2=2
r39 8 13 1.63057 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=2.08 $Y=1.92
+ $X2=1.967 $Y2=1.92
r40 8 16 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.08 $Y=1.92
+ $X2=2.715 $Y2=1.92
r41 2 11 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.485 $X2=4.185 $Y2=2
r42 1 15 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%Y 1 2 3 4 5 6 19 28 29 37 41 56
r55 47 49 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.74 $Y=2.34
+ $X2=4.61 $Y2=2.34
r56 44 47 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.88 $Y=2.34 $X2=3.74
+ $Y2=2.34
r57 37 41 2.30489 $w=2.23e-07 $l=4.5e-08 $layer=LI1_cond $X=4.862 $Y=2.255
+ $X2=4.862 $Y2=2.21
r58 36 56 1.38293 $w=2.23e-07 $l=2.7e-08 $layer=LI1_cond $X=4.862 $Y=1.897
+ $X2=4.862 $Y2=1.87
r59 29 37 3.0159 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.862 $Y=2.34
+ $X2=4.862 $Y2=2.255
r60 29 49 7.82882 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=4.75 $Y=2.34
+ $X2=4.61 $Y2=2.34
r61 29 41 1.02439 $w=2.23e-07 $l=2e-08 $layer=LI1_cond $X=4.862 $Y=2.19
+ $X2=4.862 $Y2=2.21
r62 28 56 1.48537 $w=2.23e-07 $l=2.9e-08 $layer=LI1_cond $X=4.862 $Y=1.841
+ $X2=4.862 $Y2=1.87
r63 28 29 13.522 $w=2.23e-07 $l=2.64e-07 $layer=LI1_cond $X=4.862 $Y=1.926
+ $X2=4.862 $Y2=2.19
r64 28 36 1.48537 $w=2.23e-07 $l=2.9e-08 $layer=LI1_cond $X=4.862 $Y=1.926
+ $X2=4.862 $Y2=1.897
r65 27 28 54.6137 $w=2.83e-07 $l=1.32e-06 $layer=LI1_cond $X=4.89 $Y=0.465
+ $X2=4.89 $Y2=1.785
r66 24 26 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=3.72 $Y=0.38
+ $X2=4.8 $Y2=0.38
r67 21 24 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.88 $Y=0.38
+ $X2=3.72 $Y2=0.38
r68 19 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.805 $Y=0.38
+ $X2=4.89 $Y2=0.465
r69 19 26 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.805 $Y=0.38 $X2=4.8
+ $Y2=0.38
r70 6 49 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.485 $X2=4.61 $Y2=2.34
r71 5 47 600 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.74 $Y2=2.34
r72 4 44 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.485 $X2=2.88 $Y2=2.34
r73 3 26 182 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_NDIFF $count=1 $X=4.47
+ $Y=0.235 $X2=4.8 $Y2=0.38
r74 2 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.38
r75 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.235 $X2=2.88 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r75 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r76 46 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r77 44 47 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r78 43 46 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r79 43 44 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r80 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r81 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r82 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r83 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r84 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r85 35 50 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.835 $Y=0 $X2=0.675
+ $Y2=0
r86 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.835 $Y=0 $X2=1.15
+ $Y2=0
r87 30 50 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.675
+ $Y2=0
r88 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r89 28 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r90 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r91 26 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.07
+ $Y2=0
r92 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.36
+ $Y2=0
r93 25 43 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.53
+ $Y2=0
r94 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.36
+ $Y2=0
r95 23 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.15
+ $Y2=0
r96 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.56
+ $Y2=0
r97 22 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=2.07
+ $Y2=0
r98 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.56
+ $Y2=0
r99 18 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0
r100 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.38
r101 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=0.085
+ $X2=1.56 $Y2=0
r102 14 16 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.56 $Y=0.085
+ $X2=1.56 $Y2=0.38
r103 10 50 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0
r104 10 12 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0.38
r105 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.38
r106 2 16 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r107 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%A_193_47# 1 2 7 8 14 15 18
r66 15 23 13.2257 $w=2.26e-07 $l=2.45e-07 $layer=LI1_cond $X=3.935 $Y=0.795
+ $X2=4.18 $Y2=0.795
r67 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.935 $Y=0.85
+ $X2=3.935 $Y2=0.85
r68 10 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=0.85
+ $X2=1.155 $Y2=0.85
r69 8 10 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=0.85
+ $X2=1.155 $Y2=0.85
r70 7 14 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.79 $Y=0.85
+ $X2=3.935 $Y2=0.85
r71 7 8 3.08168 $w=1.4e-07 $l=2.49e-06 $layer=MET1_cond $X=3.79 $Y=0.85 $X2=1.3
+ $Y2=0.85
r72 2 23 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.045
+ $Y=0.235 $X2=4.18 $Y2=0.74
r73 1 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2I_2%A_361_47# 1 2 9 12 14 15
r37 14 15 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=0.78
+ $X2=3.135 $Y2=0.78
r38 12 15 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.025 $Y=0.82
+ $X2=3.135 $Y2=0.82
r39 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=2.025 $Y2=0.82
r40 7 9 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.46
r41 2 14 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.74
r42 1 9 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.46
.ends


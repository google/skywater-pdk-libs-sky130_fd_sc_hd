* File: sky130_fd_sc_hd__buf_16.spice.pex
* Created: Thu Aug 27 14:09:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUF_16%A 3 7 11 15 19 23 27 31 35 39 43 47 49 50 64
+ 65
c125 64 0 1.39258e-19 $X=2.3 $Y=1.16
c126 47 0 1.25206e-19 $X=2.57 $Y=1.985
c127 43 0 1.25206e-19 $X=2.57 $Y=0.56
r128 63 65 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=2.3 $Y=1.16
+ $X2=2.57 $Y2=1.16
r129 63 64 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.3
+ $Y=1.16 $X2=2.3 $Y2=1.16
r130 61 63 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.3 $Y2=1.16
r131 60 61 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=2.15 $Y2=1.16
r132 59 60 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r133 58 59 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r134 56 58 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=0.6 $Y=1.16
+ $X2=0.89 $Y2=1.16
r135 56 57 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r136 53 56 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.6 $Y2=1.16
r137 50 64 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=2.3 $Y2=1.175
r138 49 50 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=2.075 $Y2=1.175
r139 49 57 56.2864 $w=1.98e-07 $l=1.015e-06 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=0.6 $Y2=1.175
r140 45 65 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r141 45 47 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r142 41 65 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r143 41 43 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r144 37 61 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r145 37 39 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r146 33 61 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r147 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r148 29 60 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r149 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r150 25 60 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r151 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r152 21 59 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r153 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r154 17 59 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r155 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r156 13 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r157 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r158 9 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.16
r159 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r160 5 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r161 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.985
r162 1 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r163 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_16%A_109_47# 1 2 3 4 5 6 21 25 29 33 37 41 45 49
+ 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 153 157 158 159 160 163 167 171 173 177 181 186 188 194 197 198
+ 200 203 205 224
c463 224 0 1.39258e-19 $X=9.29 $Y=1.16
r464 221 222 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.45 $Y=1.16
+ $X2=8.87 $Y2=1.16
r465 220 221 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.03 $Y=1.16
+ $X2=8.45 $Y2=1.16
r466 219 220 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.61 $Y=1.16
+ $X2=8.03 $Y2=1.16
r467 218 219 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.19 $Y=1.16
+ $X2=7.61 $Y2=1.16
r468 217 218 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.77 $Y=1.16
+ $X2=7.19 $Y2=1.16
r469 216 217 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.35 $Y=1.16
+ $X2=6.77 $Y2=1.16
r470 215 216 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.93 $Y=1.16
+ $X2=6.35 $Y2=1.16
r471 214 215 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.51 $Y=1.16
+ $X2=5.93 $Y2=1.16
r472 213 214 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.09 $Y=1.16
+ $X2=5.51 $Y2=1.16
r473 212 213 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.67 $Y=1.16
+ $X2=5.09 $Y2=1.16
r474 211 212 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.25 $Y=1.16
+ $X2=4.67 $Y2=1.16
r475 210 211 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.83 $Y=1.16
+ $X2=4.25 $Y2=1.16
r476 209 210 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.41 $Y=1.16
+ $X2=3.83 $Y2=1.16
r477 195 224 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=9.22 $Y=1.16
+ $X2=9.29 $Y2=1.16
r478 195 222 77.7608 $w=2.7e-07 $l=3.5e-07 $layer=POLY_cond $X=9.22 $Y=1.16
+ $X2=8.87 $Y2=1.16
r479 194 195 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=9.22
+ $Y=1.16 $X2=9.22 $Y2=1.16
r480 192 209 68.8738 $w=2.7e-07 $l=3.1e-07 $layer=POLY_cond $X=3.1 $Y=1.16
+ $X2=3.41 $Y2=1.16
r481 192 206 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=3.1 $Y=1.16
+ $X2=2.99 $Y2=1.16
r482 191 194 339.382 $w=1.98e-07 $l=6.12e-06 $layer=LI1_cond $X=3.1 $Y=1.175
+ $X2=9.22 $Y2=1.175
r483 191 192 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=3.1
+ $Y=1.16 $X2=3.1 $Y2=1.16
r484 189 205 0.866423 $w=2e-07 $l=8.8e-08 $layer=LI1_cond $X=2.865 $Y=1.175
+ $X2=2.777 $Y2=1.175
r485 189 191 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=2.865 $Y=1.175
+ $X2=3.1 $Y2=1.175
r486 188 203 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.777 $Y=1.445
+ $X2=2.777 $Y2=1.53
r487 187 205 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=2.777 $Y=1.275
+ $X2=2.777 $Y2=1.175
r488 187 188 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=2.777 $Y=1.275
+ $X2=2.777 $Y2=1.445
r489 186 205 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=2.777 $Y=1.075
+ $X2=2.777 $Y2=1.175
r490 185 200 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.777 $Y=0.905
+ $X2=2.777 $Y2=0.82
r491 185 186 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=2.777 $Y=0.905
+ $X2=2.777 $Y2=1.075
r492 181 183 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.36 $Y=1.63
+ $X2=2.36 $Y2=2.31
r493 179 203 27.2053 $w=1.68e-07 $l=4.17e-07 $layer=LI1_cond $X=2.36 $Y=1.53
+ $X2=2.777 $Y2=1.53
r494 179 181 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.36 $Y=1.615
+ $X2=2.36 $Y2=1.63
r495 175 200 27.2053 $w=1.68e-07 $l=4.17e-07 $layer=LI1_cond $X=2.36 $Y=0.82
+ $X2=2.777 $Y2=0.82
r496 175 177 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.36 $Y=0.735
+ $X2=2.36 $Y2=0.4
r497 174 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.53
+ $X2=1.52 $Y2=1.53
r498 173 179 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=1.53
+ $X2=2.36 $Y2=1.53
r499 173 174 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.195 $Y=1.53
+ $X2=1.685 $Y2=1.53
r500 172 197 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0.82
+ $X2=1.52 $Y2=0.82
r501 171 175 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=2.36 $Y2=0.82
r502 171 172 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=1.685 $Y2=0.82
r503 167 169 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.52 $Y=1.63
+ $X2=1.52 $Y2=2.31
r504 165 198 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.615
+ $X2=1.52 $Y2=1.53
r505 165 167 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.52 $Y=1.615
+ $X2=1.52 $Y2=1.63
r506 161 197 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.735
+ $X2=1.52 $Y2=0.82
r507 161 163 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=0.735
+ $X2=1.52 $Y2=0.4
r508 159 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.53
+ $X2=1.52 $Y2=1.53
r509 159 160 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.53
+ $X2=0.845 $Y2=1.53
r510 157 197 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0.82
+ $X2=1.52 $Y2=0.82
r511 157 158 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=0.82
+ $X2=0.845 $Y2=0.82
r512 153 155 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.68 $Y=1.63
+ $X2=0.68 $Y2=2.31
r513 151 160 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.68 $Y=1.615
+ $X2=0.845 $Y2=1.53
r514 151 153 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.68 $Y=1.615
+ $X2=0.68 $Y2=1.63
r515 147 158 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.68 $Y=0.735
+ $X2=0.845 $Y2=0.82
r516 147 149 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.735
+ $X2=0.68 $Y2=0.4
r517 143 224 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.29 $Y=1.295
+ $X2=9.29 $Y2=1.16
r518 143 145 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.29 $Y=1.295
+ $X2=9.29 $Y2=1.985
r519 139 224 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.29 $Y=1.025
+ $X2=9.29 $Y2=1.16
r520 139 141 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.29 $Y=1.025
+ $X2=9.29 $Y2=0.56
r521 135 222 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.87 $Y=1.295
+ $X2=8.87 $Y2=1.16
r522 135 137 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.87 $Y=1.295
+ $X2=8.87 $Y2=1.985
r523 131 222 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.87 $Y=1.025
+ $X2=8.87 $Y2=1.16
r524 131 133 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.87 $Y=1.025
+ $X2=8.87 $Y2=0.56
r525 127 221 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.45 $Y=1.295
+ $X2=8.45 $Y2=1.16
r526 127 129 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.45 $Y=1.295
+ $X2=8.45 $Y2=1.985
r527 123 221 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.45 $Y=1.025
+ $X2=8.45 $Y2=1.16
r528 123 125 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.45 $Y=1.025
+ $X2=8.45 $Y2=0.56
r529 119 220 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.03 $Y=1.295
+ $X2=8.03 $Y2=1.16
r530 119 121 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.03 $Y=1.295
+ $X2=8.03 $Y2=1.985
r531 115 220 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.03 $Y=1.025
+ $X2=8.03 $Y2=1.16
r532 115 117 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.03 $Y=1.025
+ $X2=8.03 $Y2=0.56
r533 111 219 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.61 $Y=1.295
+ $X2=7.61 $Y2=1.16
r534 111 113 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.61 $Y=1.295
+ $X2=7.61 $Y2=1.985
r535 107 219 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.61 $Y=1.025
+ $X2=7.61 $Y2=1.16
r536 107 109 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.61 $Y=1.025
+ $X2=7.61 $Y2=0.56
r537 103 218 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.19 $Y=1.295
+ $X2=7.19 $Y2=1.16
r538 103 105 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.19 $Y=1.295
+ $X2=7.19 $Y2=1.985
r539 99 218 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.19 $Y=1.025
+ $X2=7.19 $Y2=1.16
r540 99 101 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.19 $Y=1.025
+ $X2=7.19 $Y2=0.56
r541 95 217 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.16
r542 95 97 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.985
r543 91 217 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=1.16
r544 91 93 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=0.56
r545 87 216 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.16
r546 87 89 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.985
r547 83 216 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=1.16
r548 83 85 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=0.56
r549 79 215 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.16
r550 79 81 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.985
r551 75 215 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=1.16
r552 75 77 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=0.56
r553 71 214 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.16
r554 71 73 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.985
r555 67 214 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=1.16
r556 67 69 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=0.56
r557 63 213 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.16
r558 63 65 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.985
r559 59 213 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=1.16
r560 59 61 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=0.56
r561 55 212 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.16
r562 55 57 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.985
r563 51 212 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=1.16
r564 51 53 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=0.56
r565 47 211 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.16
r566 47 49 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.985
r567 43 211 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=1.16
r568 43 45 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=0.56
r569 39 210 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.16
r570 39 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.985
r571 35 210 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=1.16
r572 35 37 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=0.56
r573 31 209 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r574 31 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r575 27 209 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r576 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r577 23 206 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r578 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r579 19 206 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r580 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r581 6 183 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.31
r582 6 181 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.63
r583 5 169 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.31
r584 5 167 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.63
r585 4 155 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.31
r586 4 153 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.63
r587 3 177 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.4
r588 2 163 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r589 1 149 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37 39 45 49
+ 53 57 61 63 67 71 75 79 83 85 89 92 93 95 96 98 99 101 102 103 104 106 107 109
+ 110 112 113 114 115 116 149 150 156 159
r164 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r165 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r166 150 160 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r167 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r168 147 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.585 $Y=2.72
+ $X2=9.5 $Y2=2.72
r169 147 149 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.585 $Y=2.72
+ $X2=9.89 $Y2=2.72
r170 146 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r171 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r172 143 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r173 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r174 140 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r175 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r176 137 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r177 137 157 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r178 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r179 134 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.3 $Y2=2.72
r180 134 136 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.75 $Y2=2.72
r181 133 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r182 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r183 130 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r184 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r185 127 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r186 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r187 124 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r188 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r189 121 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r190 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r191 118 153 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r192 118 120 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r193 116 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r194 116 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r195 114 145 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.575 $Y=2.72
+ $X2=8.51 $Y2=2.72
r196 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=2.72
+ $X2=8.66 $Y2=2.72
r197 112 142 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.735 $Y=2.72
+ $X2=7.59 $Y2=2.72
r198 112 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.735 $Y=2.72
+ $X2=7.82 $Y2=2.72
r199 111 145 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.905 $Y=2.72
+ $X2=8.51 $Y2=2.72
r200 111 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=2.72
+ $X2=7.82 $Y2=2.72
r201 109 139 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.895 $Y=2.72
+ $X2=6.67 $Y2=2.72
r202 109 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.895 $Y=2.72
+ $X2=6.98 $Y2=2.72
r203 108 142 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.065 $Y=2.72
+ $X2=7.59 $Y2=2.72
r204 108 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=2.72
+ $X2=6.98 $Y2=2.72
r205 106 136 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=5.75 $Y2=2.72
r206 106 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=6.14 $Y2=2.72
r207 105 139 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.225 $Y=2.72
+ $X2=6.67 $Y2=2.72
r208 105 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=2.72
+ $X2=6.14 $Y2=2.72
r209 103 132 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.37 $Y2=2.72
r210 103 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=2.72
+ $X2=4.46 $Y2=2.72
r211 101 129 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.45 $Y2=2.72
r212 101 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.62 $Y2=2.72
r213 100 132 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.705 $Y=2.72
+ $X2=4.37 $Y2=2.72
r214 100 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=2.72
+ $X2=3.62 $Y2=2.72
r215 98 126 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.53 $Y2=2.72
r216 98 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.78 $Y2=2.72
r217 97 129 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.45 $Y2=2.72
r218 97 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.78 $Y2=2.72
r219 95 123 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r220 95 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.94 $Y2=2.72
r221 94 126 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.53 $Y2=2.72
r222 94 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.94 $Y2=2.72
r223 92 120 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r224 92 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r225 91 123 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r226 91 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r227 87 159 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.5 $Y=2.635
+ $X2=9.5 $Y2=2.72
r228 87 89 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.5 $Y=2.635
+ $X2=9.5 $Y2=2
r229 86 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=2.72
+ $X2=8.66 $Y2=2.72
r230 85 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.415 $Y=2.72
+ $X2=9.5 $Y2=2.72
r231 85 86 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.415 $Y=2.72
+ $X2=8.745 $Y2=2.72
r232 81 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.66 $Y=2.635
+ $X2=8.66 $Y2=2.72
r233 81 83 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.66 $Y=2.635
+ $X2=8.66 $Y2=2
r234 77 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.82 $Y=2.635
+ $X2=7.82 $Y2=2.72
r235 77 79 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.82 $Y=2.635
+ $X2=7.82 $Y2=2
r236 73 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=2.635
+ $X2=6.98 $Y2=2.72
r237 73 75 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.98 $Y=2.635
+ $X2=6.98 $Y2=2
r238 69 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=2.635
+ $X2=6.14 $Y2=2.72
r239 69 71 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.14 $Y=2.635
+ $X2=6.14 $Y2=2
r240 65 156 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.72
r241 65 67 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2
r242 64 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.46 $Y2=2.72
r243 63 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=2.72
+ $X2=5.3 $Y2=2.72
r244 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.215 $Y=2.72
+ $X2=4.545 $Y2=2.72
r245 59 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2.72
r246 59 61 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2
r247 55 102 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r248 55 57 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2
r249 51 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r250 51 53 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r251 47 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r252 47 49 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r253 43 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r254 43 45 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r255 39 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r256 37 153 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r257 37 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r258 12 89 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.365
+ $Y=1.485 $X2=9.5 $Y2=2
r259 11 83 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.525
+ $Y=1.485 $X2=8.66 $Y2=2
r260 10 79 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.685
+ $Y=1.485 $X2=7.82 $Y2=2
r261 9 75 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.845
+ $Y=1.485 $X2=6.98 $Y2=2
r262 8 71 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.005
+ $Y=1.485 $X2=6.14 $Y2=2
r263 7 67 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=2
r264 6 61 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=2
r265 5 57 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2
r266 4 53 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r267 3 49 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r268 2 45 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r269 1 42 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r270 1 39 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 49
+ 50 53 57 58 59 60 61 62 65 69 71 73 74 77 81 83 87 91 95 97 101 105 109 111
+ 115 119 123 125 129 133 137 139 143 147 151 153 161 162 165 166 167 168 169
+ 170 171 172 173 174 175 176 178 179 180 192
c348 60 0 1.25206e-19 $X=3.365 $Y=1.53
c349 58 0 1.25206e-19 $X=3.365 $Y=0.82
r350 180 192 2.90768 $w=3.27e-07 $l=1.07912e-07 $layer=LI1_cond $X=9.845 $Y=1.53
+ $X2=9.897 $Y2=1.615
r351 180 192 0.112383 $w=7.43e-07 $l=7e-09 $layer=LI1_cond $X=9.89 $Y=1.987
+ $X2=9.897 $Y2=1.987
r352 179 180 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=9.845 $Y=1.19
+ $X2=9.845 $Y2=1.445
r353 177 179 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=9.845 $Y=0.905
+ $X2=9.845 $Y2=1.19
r354 177 178 2.90768 $w=3.27e-07 $l=8.5e-08 $layer=LI1_cond $X=9.845 $Y=0.905
+ $X2=9.845 $Y2=0.82
r355 154 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.245 $Y=1.53
+ $X2=9.08 $Y2=1.53
r356 153 180 3.78066 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.655 $Y=1.53
+ $X2=9.845 $Y2=1.53
r357 153 154 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.655 $Y=1.53
+ $X2=9.245 $Y2=1.53
r358 152 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.245 $Y=0.82
+ $X2=9.08 $Y2=0.82
r359 151 178 3.78066 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.655 $Y=0.82
+ $X2=9.845 $Y2=0.82
r360 151 152 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.655 $Y=0.82
+ $X2=9.245 $Y2=0.82
r361 147 149 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.08 $Y=1.63
+ $X2=9.08 $Y2=2.31
r362 145 176 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.08 $Y=1.615
+ $X2=9.08 $Y2=1.53
r363 145 147 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=9.08 $Y=1.615
+ $X2=9.08 $Y2=1.63
r364 141 175 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.08 $Y=0.735
+ $X2=9.08 $Y2=0.82
r365 141 143 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.08 $Y=0.735
+ $X2=9.08 $Y2=0.4
r366 140 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=1.53
+ $X2=8.24 $Y2=1.53
r367 139 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.915 $Y=1.53
+ $X2=9.08 $Y2=1.53
r368 139 140 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.915 $Y=1.53
+ $X2=8.405 $Y2=1.53
r369 138 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=0.82
+ $X2=8.24 $Y2=0.82
r370 137 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.915 $Y=0.82
+ $X2=9.08 $Y2=0.82
r371 137 138 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.915 $Y=0.82
+ $X2=8.405 $Y2=0.82
r372 133 135 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.24 $Y=1.63
+ $X2=8.24 $Y2=2.31
r373 131 174 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=1.615
+ $X2=8.24 $Y2=1.53
r374 131 133 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.24 $Y=1.615
+ $X2=8.24 $Y2=1.63
r375 127 173 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=0.735
+ $X2=8.24 $Y2=0.82
r376 127 129 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.24 $Y=0.735
+ $X2=8.24 $Y2=0.4
r377 126 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.565 $Y=1.53
+ $X2=7.4 $Y2=1.53
r378 125 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=1.53
+ $X2=8.24 $Y2=1.53
r379 125 126 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.075 $Y=1.53
+ $X2=7.565 $Y2=1.53
r380 124 171 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.565 $Y=0.82
+ $X2=7.4 $Y2=0.82
r381 123 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0.82
+ $X2=8.24 $Y2=0.82
r382 123 124 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.075 $Y=0.82
+ $X2=7.565 $Y2=0.82
r383 119 121 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.4 $Y=1.63
+ $X2=7.4 $Y2=2.31
r384 117 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=1.615
+ $X2=7.4 $Y2=1.53
r385 117 119 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.4 $Y=1.615
+ $X2=7.4 $Y2=1.63
r386 113 171 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0.735
+ $X2=7.4 $Y2=0.82
r387 113 115 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.4 $Y=0.735
+ $X2=7.4 $Y2=0.4
r388 112 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=1.53
+ $X2=6.56 $Y2=1.53
r389 111 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=1.53
+ $X2=7.4 $Y2=1.53
r390 111 112 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.235 $Y=1.53
+ $X2=6.725 $Y2=1.53
r391 110 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=0.82
+ $X2=6.56 $Y2=0.82
r392 109 171 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=0.82
+ $X2=7.4 $Y2=0.82
r393 109 110 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.235 $Y=0.82
+ $X2=6.725 $Y2=0.82
r394 105 107 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.56 $Y=1.63
+ $X2=6.56 $Y2=2.31
r395 103 170 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=1.615
+ $X2=6.56 $Y2=1.53
r396 103 105 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.56 $Y=1.615
+ $X2=6.56 $Y2=1.63
r397 99 169 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=0.735
+ $X2=6.56 $Y2=0.82
r398 99 101 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.56 $Y=0.735
+ $X2=6.56 $Y2=0.4
r399 98 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.885 $Y=1.53
+ $X2=5.72 $Y2=1.53
r400 97 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=1.53
+ $X2=6.56 $Y2=1.53
r401 97 98 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.395 $Y=1.53
+ $X2=5.885 $Y2=1.53
r402 96 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.885 $Y=0.82
+ $X2=5.72 $Y2=0.82
r403 95 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=0.82
+ $X2=6.56 $Y2=0.82
r404 95 96 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.395 $Y=0.82
+ $X2=5.885 $Y2=0.82
r405 91 93 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.72 $Y=1.63
+ $X2=5.72 $Y2=2.31
r406 89 168 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=1.615
+ $X2=5.72 $Y2=1.53
r407 89 91 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.72 $Y=1.615
+ $X2=5.72 $Y2=1.63
r408 85 167 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=0.735
+ $X2=5.72 $Y2=0.82
r409 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.72 $Y=0.735
+ $X2=5.72 $Y2=0.4
r410 84 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=1.53
+ $X2=4.88 $Y2=1.53
r411 83 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.555 $Y=1.53
+ $X2=5.72 $Y2=1.53
r412 83 84 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.555 $Y=1.53
+ $X2=5.045 $Y2=1.53
r413 82 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=0.82
+ $X2=4.88 $Y2=0.82
r414 81 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.555 $Y=0.82
+ $X2=5.72 $Y2=0.82
r415 81 82 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.555 $Y=0.82
+ $X2=5.045 $Y2=0.82
r416 77 79 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.88 $Y=1.63
+ $X2=4.88 $Y2=2.31
r417 75 166 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=1.615
+ $X2=4.88 $Y2=1.53
r418 75 77 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.88 $Y=1.615
+ $X2=4.88 $Y2=1.63
r419 74 165 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.735
+ $X2=4.88 $Y2=0.82
r420 73 164 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=4.88 $Y=0.425
+ $X2=4.88 $Y2=0.4
r421 73 74 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=4.88 $Y=0.425
+ $X2=4.88 $Y2=0.735
r422 72 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=1.53
+ $X2=4.04 $Y2=1.53
r423 71 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=1.53
+ $X2=4.88 $Y2=1.53
r424 71 72 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.715 $Y=1.53
+ $X2=4.205 $Y2=1.53
r425 70 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0.82
+ $X2=4.04 $Y2=0.82
r426 69 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0.82
+ $X2=4.88 $Y2=0.82
r427 69 70 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.715 $Y=0.82
+ $X2=4.205 $Y2=0.82
r428 65 67 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.04 $Y=1.63
+ $X2=4.04 $Y2=2.31
r429 63 162 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.615
+ $X2=4.04 $Y2=1.53
r430 63 65 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.04 $Y=1.615
+ $X2=4.04 $Y2=1.63
r431 62 161 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.735
+ $X2=4.04 $Y2=0.82
r432 61 160 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=4.04 $Y=0.425
+ $X2=4.04 $Y2=0.4
r433 61 62 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=4.04 $Y=0.425
+ $X2=4.04 $Y2=0.735
r434 59 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=1.53
+ $X2=4.04 $Y2=1.53
r435 59 60 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.875 $Y=1.53
+ $X2=3.365 $Y2=1.53
r436 57 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=0.82
+ $X2=4.04 $Y2=0.82
r437 57 58 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.875 $Y=0.82
+ $X2=3.365 $Y2=0.82
r438 53 55 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.2 $Y=1.63 $X2=3.2
+ $Y2=2.31
r439 51 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.2 $Y=1.615
+ $X2=3.365 $Y2=1.53
r440 51 53 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.2 $Y=1.615
+ $X2=3.2 $Y2=1.63
r441 50 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.2 $Y=0.735
+ $X2=3.365 $Y2=0.82
r442 49 158 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=3.2 $Y=0.425
+ $X2=3.2 $Y2=0.4
r443 49 50 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.2 $Y=0.425 $X2=3.2
+ $Y2=0.735
r444 16 149 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=1.485 $X2=9.08 $Y2=2.31
r445 16 147 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.945
+ $Y=1.485 $X2=9.08 $Y2=1.63
r446 15 135 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.24 $Y2=2.31
r447 15 133 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.24 $Y2=1.63
r448 14 121 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.485 $X2=7.4 $Y2=2.31
r449 14 119 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.485 $X2=7.4 $Y2=1.63
r450 13 107 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.485 $X2=6.56 $Y2=2.31
r451 13 105 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.485 $X2=6.56 $Y2=1.63
r452 12 93 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=2.31
r453 12 91 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=1.63
r454 11 79 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=2.31
r455 11 77 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=1.63
r456 10 67 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=2.31
r457 10 65 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=1.63
r458 9 55 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.31
r459 9 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.63
r460 8 143 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.945
+ $Y=0.235 $X2=9.08 $Y2=0.4
r461 7 129 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.105
+ $Y=0.235 $X2=8.24 $Y2=0.4
r462 6 115 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=7.265
+ $Y=0.235 $X2=7.4 $Y2=0.4
r463 5 101 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=6.425
+ $Y=0.235 $X2=6.56 $Y2=0.4
r464 4 87 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.4
r465 3 164 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.4
r466 2 160 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.4
r467 1 158 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 37 39 43 47
+ 51 55 59 61 65 69 73 77 81 83 87 90 91 93 94 96 97 99 100 101 102 104 105 107
+ 108 110 111 112 113 114 147 148 154 157
r194 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r195 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r196 148 158 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=9.43 $Y2=0
r197 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r198 145 157 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.585 $Y=0 $X2=9.5
+ $Y2=0
r199 145 147 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.585 $Y=0
+ $X2=9.89 $Y2=0
r200 144 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r201 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r202 141 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r203 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r204 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r205 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r206 135 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r207 135 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r208 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r209 132 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.3
+ $Y2=0
r210 132 134 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.385 $Y=0
+ $X2=5.75 $Y2=0
r211 131 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r212 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r213 128 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r214 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r215 125 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r216 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r217 122 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r218 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r219 119 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r220 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r221 116 151 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r222 116 118 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.69 $Y2=0
r223 114 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r224 114 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r225 112 143 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.575 $Y=0
+ $X2=8.51 $Y2=0
r226 112 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=0
+ $X2=8.66 $Y2=0
r227 110 140 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.735 $Y=0
+ $X2=7.59 $Y2=0
r228 110 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.735 $Y=0
+ $X2=7.82 $Y2=0
r229 109 143 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.905 $Y=0
+ $X2=8.51 $Y2=0
r230 109 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=0
+ $X2=7.82 $Y2=0
r231 107 137 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.895 $Y=0
+ $X2=6.67 $Y2=0
r232 107 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.895 $Y=0
+ $X2=6.98 $Y2=0
r233 106 140 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.065 $Y=0
+ $X2=7.59 $Y2=0
r234 106 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=0
+ $X2=6.98 $Y2=0
r235 104 134 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.055 $Y=0
+ $X2=5.75 $Y2=0
r236 104 105 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=0
+ $X2=6.14 $Y2=0
r237 103 137 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.225 $Y=0
+ $X2=6.67 $Y2=0
r238 103 105 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=0
+ $X2=6.14 $Y2=0
r239 101 130 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=0
+ $X2=4.37 $Y2=0
r240 101 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=0
+ $X2=4.46 $Y2=0
r241 99 127 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0
+ $X2=3.45 $Y2=0
r242 99 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.62
+ $Y2=0
r243 98 130 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.705 $Y=0
+ $X2=4.37 $Y2=0
r244 98 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.62
+ $Y2=0
r245 96 124 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=2.53 $Y2=0
r246 96 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.78
+ $Y2=0
r247 95 127 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=3.45 $Y2=0
r248 95 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.78
+ $Y2=0
r249 93 121 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.61 $Y2=0
r250 93 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.94
+ $Y2=0
r251 92 124 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.53 $Y2=0
r252 92 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.94
+ $Y2=0
r253 90 118 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r254 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r255 89 121 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r256 89 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r257 85 157 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.5 $Y=0.085
+ $X2=9.5 $Y2=0
r258 85 87 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.5 $Y=0.085
+ $X2=9.5 $Y2=0.4
r259 84 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=0 $X2=8.66
+ $Y2=0
r260 83 157 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.415 $Y=0 $X2=9.5
+ $Y2=0
r261 83 84 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.415 $Y=0
+ $X2=8.745 $Y2=0
r262 79 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.66 $Y=0.085
+ $X2=8.66 $Y2=0
r263 79 81 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.66 $Y=0.085
+ $X2=8.66 $Y2=0.4
r264 75 111 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.82 $Y=0.085
+ $X2=7.82 $Y2=0
r265 75 77 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.82 $Y=0.085
+ $X2=7.82 $Y2=0.4
r266 71 108 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=0.085
+ $X2=6.98 $Y2=0
r267 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.98 $Y=0.085
+ $X2=6.98 $Y2=0.4
r268 67 105 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=0.085
+ $X2=6.14 $Y2=0
r269 67 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.14 $Y=0.085
+ $X2=6.14 $Y2=0.4
r270 63 154 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0
r271 63 65 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0.4
r272 62 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=0 $X2=4.46
+ $Y2=0
r273 61 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.3
+ $Y2=0
r274 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.215 $Y=0
+ $X2=4.545 $Y2=0
r275 57 102 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r276 57 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.4
r277 53 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0
r278 53 55 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0.4
r279 49 97 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r280 49 51 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.4
r281 45 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r282 45 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.4
r283 41 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r284 41 43 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.4
r285 37 151 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r286 37 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r287 12 87 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=9.365
+ $Y=0.235 $X2=9.5 $Y2=0.4
r288 11 81 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.525
+ $Y=0.235 $X2=8.66 $Y2=0.4
r289 10 77 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.235 $X2=7.82 $Y2=0.4
r290 9 73 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.845
+ $Y=0.235 $X2=6.98 $Y2=0.4
r291 8 69 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.005
+ $Y=0.235 $X2=6.14 $Y2=0.4
r292 7 65 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.165
+ $Y=0.235 $X2=5.3 $Y2=0.4
r293 6 59 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.4
r294 5 55 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.4
r295 4 51 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.4
r296 3 47 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.4
r297 2 43 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r298 1 39 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__sdfbbn_2.spice.SKY130_FD_SC_HD__SDFBBN_2.pxi
* Created: Thu Aug 27 14:45:25 2020
* 
x_PM_SKY130_FD_SC_HD__SDFBBN_2%CLK_N N_CLK_N_c_313_n N_CLK_N_c_308_n
+ N_CLK_N_M1048_g N_CLK_N_c_314_n N_CLK_N_M1027_g N_CLK_N_c_309_n
+ N_CLK_N_c_315_n CLK_N CLK_N N_CLK_N_c_311_n N_CLK_N_c_312_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%CLK_N
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_27_47# N_A_27_47#_M1048_s N_A_27_47#_M1027_s
+ N_A_27_47#_M1028_g N_A_27_47#_M1000_g N_A_27_47#_M1040_g N_A_27_47#_c_354_n
+ N_A_27_47#_c_355_n N_A_27_47#_M1020_g N_A_27_47#_c_357_n N_A_27_47#_c_358_n
+ N_A_27_47#_M1008_g N_A_27_47#_M1021_g N_A_27_47#_c_617_p N_A_27_47#_c_359_n
+ N_A_27_47#_c_360_n N_A_27_47#_c_380_n N_A_27_47#_c_361_n N_A_27_47#_c_362_n
+ N_A_27_47#_c_363_n N_A_27_47#_c_381_n N_A_27_47#_c_382_n N_A_27_47#_c_383_n
+ N_A_27_47#_c_364_n N_A_27_47#_c_365_n N_A_27_47#_c_366_n N_A_27_47#_c_367_n
+ N_A_27_47#_c_368_n N_A_27_47#_c_369_n N_A_27_47#_c_370_n N_A_27_47#_c_371_n
+ N_A_27_47#_c_372_n N_A_27_47#_c_373_n N_A_27_47#_c_374_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%SCD N_SCD_M1006_g N_SCD_M1034_g SCD SCD
+ N_SCD_c_636_n PM_SKY130_FD_SC_HD__SDFBBN_2%SCD
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_423_315# N_A_423_315#_M1013_s
+ N_A_423_315#_M1035_s N_A_423_315#_c_676_n N_A_423_315#_M1039_g
+ N_A_423_315#_c_677_n N_A_423_315#_c_678_n N_A_423_315#_M1023_g
+ N_A_423_315#_c_679_n N_A_423_315#_c_732_p N_A_423_315#_c_680_n
+ N_A_423_315#_c_669_n N_A_423_315#_c_670_n N_A_423_315#_c_671_n
+ N_A_423_315#_c_672_n N_A_423_315#_c_673_n N_A_423_315#_c_682_n
+ N_A_423_315#_c_674_n N_A_423_315#_c_675_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_423_315#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%SCE N_SCE_c_772_n N_SCE_M1012_g N_SCE_c_773_n
+ N_SCE_c_774_n N_SCE_M1013_g N_SCE_c_775_n N_SCE_c_782_n N_SCE_M1035_g
+ N_SCE_c_783_n N_SCE_c_784_n N_SCE_M1022_g N_SCE_c_776_n N_SCE_c_785_n
+ N_SCE_c_777_n SCE SCE SCE N_SCE_c_780_n PM_SKY130_FD_SC_HD__SDFBBN_2%SCE
x_PM_SKY130_FD_SC_HD__SDFBBN_2%D N_D_M1024_g N_D_M1019_g D D N_D_c_874_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%D
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_193_47# N_A_193_47#_M1028_d N_A_193_47#_M1000_d
+ N_A_193_47#_c_912_n N_A_193_47#_M1045_g N_A_193_47#_M1010_g
+ N_A_193_47#_M1032_g N_A_193_47#_c_913_n N_A_193_47#_c_914_n
+ N_A_193_47#_M1003_g N_A_193_47#_c_916_n N_A_193_47#_c_917_n
+ N_A_193_47#_c_924_n N_A_193_47#_c_925_n N_A_193_47#_c_926_n
+ N_A_193_47#_c_927_n N_A_193_47#_c_928_n N_A_193_47#_c_929_n
+ N_A_193_47#_c_930_n N_A_193_47#_c_931_n N_A_193_47#_c_932_n
+ N_A_193_47#_c_933_n N_A_193_47#_c_918_n PM_SKY130_FD_SC_HD__SDFBBN_2%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_1107_21# N_A_1107_21#_M1016_d
+ N_A_1107_21#_M1011_d N_A_1107_21#_M1038_g N_A_1107_21#_M1036_g
+ N_A_1107_21#_M1050_g N_A_1107_21#_c_1127_n N_A_1107_21#_M1041_g
+ N_A_1107_21#_c_1136_n N_A_1107_21#_c_1185_p N_A_1107_21#_c_1150_n
+ N_A_1107_21#_c_1128_n N_A_1107_21#_c_1129_n N_A_1107_21#_c_1130_n
+ N_A_1107_21#_c_1138_n N_A_1107_21#_c_1139_n N_A_1107_21#_c_1155_n
+ N_A_1107_21#_c_1131_n N_A_1107_21#_c_1132_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_1107_21#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%SET_B N_SET_B_c_1272_n N_SET_B_M1011_g
+ N_SET_B_M1047_g N_SET_B_M1004_g N_SET_B_M1007_g SET_B N_SET_B_c_1278_n
+ N_SET_B_c_1279_n N_SET_B_c_1280_n N_SET_B_c_1281_n N_SET_B_c_1282_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%SET_B
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_931_47# N_A_931_47#_M1045_d N_A_931_47#_M1040_d
+ N_A_931_47#_M1016_g N_A_931_47#_M1037_g N_A_931_47#_c_1414_n
+ N_A_931_47#_c_1415_n N_A_931_47#_c_1409_n N_A_931_47#_c_1404_n
+ N_A_931_47#_c_1405_n N_A_931_47#_c_1406_n N_A_931_47#_c_1407_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_931_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_1401_21# N_A_1401_21#_M1009_s
+ N_A_1401_21#_M1030_s N_A_1401_21#_c_1509_n N_A_1401_21#_M1014_g
+ N_A_1401_21#_c_1510_n N_A_1401_21#_M1031_g N_A_1401_21#_M1029_g
+ N_A_1401_21#_M1017_g N_A_1401_21#_c_1512_n N_A_1401_21#_c_1513_n
+ N_A_1401_21#_c_1521_n N_A_1401_21#_c_1522_n N_A_1401_21#_c_1514_n
+ N_A_1401_21#_c_1515_n N_A_1401_21#_c_1524_n N_A_1401_21#_c_1525_n
+ N_A_1401_21#_c_1526_n N_A_1401_21#_c_1527_n N_A_1401_21#_c_1516_n
+ N_A_1401_21#_c_1517_n PM_SKY130_FD_SC_HD__SDFBBN_2%A_1401_21#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_1888_21# N_A_1888_21#_M1001_d
+ N_A_1888_21#_M1007_d N_A_1888_21#_M1042_g N_A_1888_21#_M1043_g
+ N_A_1888_21#_c_1666_n N_A_1888_21#_M1049_g N_A_1888_21#_M1002_g
+ N_A_1888_21#_M1051_g N_A_1888_21#_M1046_g N_A_1888_21#_c_1669_n
+ N_A_1888_21#_c_1670_n N_A_1888_21#_c_1671_n N_A_1888_21#_c_1672_n
+ N_A_1888_21#_c_1673_n N_A_1888_21#_M1044_g N_A_1888_21#_c_1684_n
+ N_A_1888_21#_M1033_g N_A_1888_21#_c_1674_n N_A_1888_21#_c_1675_n
+ N_A_1888_21#_c_1685_n N_A_1888_21#_c_1686_n N_A_1888_21#_c_1687_n
+ N_A_1888_21#_c_1688_n N_A_1888_21#_c_1742_p N_A_1888_21#_c_1796_p
+ N_A_1888_21#_c_1714_n N_A_1888_21#_c_1676_n N_A_1888_21#_c_1690_n
+ N_A_1888_21#_c_1691_n N_A_1888_21#_c_1731_n N_A_1888_21#_c_1707_n
+ N_A_1888_21#_c_1733_n N_A_1888_21#_c_1677_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_1888_21#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_1714_47# N_A_1714_47#_M1008_d
+ N_A_1714_47#_M1032_d N_A_1714_47#_M1001_g N_A_1714_47#_M1025_g
+ N_A_1714_47#_c_1872_n N_A_1714_47#_c_1875_n N_A_1714_47#_c_1861_n
+ N_A_1714_47#_c_1867_n N_A_1714_47#_c_1862_n N_A_1714_47#_c_1863_n
+ N_A_1714_47#_c_1864_n N_A_1714_47#_c_1865_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_1714_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%RESET_B N_RESET_B_M1009_g N_RESET_B_M1030_g
+ RESET_B N_RESET_B_c_1961_n PM_SKY130_FD_SC_HD__SDFBBN_2%RESET_B
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_2696_47# N_A_2696_47#_M1044_s
+ N_A_2696_47#_M1033_s N_A_2696_47#_c_1995_n N_A_2696_47#_M1015_g
+ N_A_2696_47#_M1005_g N_A_2696_47#_c_1996_n N_A_2696_47#_M1026_g
+ N_A_2696_47#_M1018_g N_A_2696_47#_c_1997_n N_A_2696_47#_c_2003_n
+ N_A_2696_47#_c_1998_n N_A_2696_47#_c_1999_n N_A_2696_47#_c_2000_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_2696_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%VPWR N_VPWR_M1027_d N_VPWR_M1034_s N_VPWR_M1035_d
+ N_VPWR_M1036_d N_VPWR_M1031_d N_VPWR_M1043_d N_VPWR_M1029_d N_VPWR_M1030_d
+ N_VPWR_M1046_s N_VPWR_M1033_d N_VPWR_M1018_d N_VPWR_c_2071_n N_VPWR_c_2072_n
+ N_VPWR_c_2073_n N_VPWR_c_2074_n N_VPWR_c_2075_n N_VPWR_c_2076_n
+ N_VPWR_c_2077_n N_VPWR_c_2078_n N_VPWR_c_2079_n N_VPWR_c_2080_n
+ N_VPWR_c_2081_n N_VPWR_c_2082_n N_VPWR_c_2083_n N_VPWR_c_2084_n VPWR VPWR
+ N_VPWR_c_2085_n N_VPWR_c_2086_n N_VPWR_c_2087_n N_VPWR_c_2088_n
+ N_VPWR_c_2089_n N_VPWR_c_2090_n N_VPWR_c_2091_n N_VPWR_c_2092_n
+ N_VPWR_c_2093_n N_VPWR_c_2094_n N_VPWR_c_2095_n N_VPWR_c_2096_n
+ N_VPWR_c_2097_n N_VPWR_c_2098_n N_VPWR_c_2099_n N_VPWR_c_2100_n
+ N_VPWR_c_2070_n PM_SKY130_FD_SC_HD__SDFBBN_2%VPWR
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_453_47# N_A_453_47#_M1012_d N_A_453_47#_M1024_d
+ N_A_453_47#_M1039_d N_A_453_47#_M1019_d N_A_453_47#_c_2297_n
+ N_A_453_47#_c_2298_n N_A_453_47#_c_2306_n N_A_453_47#_c_2307_n
+ N_A_453_47#_c_2299_n N_A_453_47#_c_2300_n N_A_453_47#_c_2301_n
+ N_A_453_47#_c_2302_n N_A_453_47#_c_2303_n N_A_453_47#_c_2304_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%A_453_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%Q_N N_Q_N_M1049_s N_Q_N_M1002_d N_Q_N_c_2432_n
+ N_Q_N_c_2430_n Q_N Q_N Q_N N_Q_N_c_2443_n Q_N PM_SKY130_FD_SC_HD__SDFBBN_2%Q_N
x_PM_SKY130_FD_SC_HD__SDFBBN_2%Q N_Q_M1015_d N_Q_M1005_s N_Q_c_2457_n
+ N_Q_c_2455_n N_Q_c_2454_n Q Q Q PM_SKY130_FD_SC_HD__SDFBBN_2%Q
x_PM_SKY130_FD_SC_HD__SDFBBN_2%VGND N_VGND_M1048_d N_VGND_M1006_s N_VGND_M1013_d
+ N_VGND_M1038_d N_VGND_M1041_s N_VGND_M1042_d N_VGND_M1009_d N_VGND_M1051_d
+ N_VGND_M1044_d N_VGND_M1026_s N_VGND_c_2475_n N_VGND_c_2476_n N_VGND_c_2477_n
+ N_VGND_c_2478_n N_VGND_c_2479_n N_VGND_c_2480_n N_VGND_c_2481_n
+ N_VGND_c_2482_n N_VGND_c_2483_n N_VGND_c_2484_n N_VGND_c_2485_n
+ N_VGND_c_2486_n N_VGND_c_2487_n N_VGND_c_2488_n N_VGND_c_2489_n
+ N_VGND_c_2490_n N_VGND_c_2491_n N_VGND_c_2492_n VGND VGND N_VGND_c_2493_n
+ N_VGND_c_2494_n N_VGND_c_2495_n N_VGND_c_2496_n N_VGND_c_2497_n
+ N_VGND_c_2498_n N_VGND_c_2499_n N_VGND_c_2500_n N_VGND_c_2501_n
+ N_VGND_c_2502_n N_VGND_c_2503_n N_VGND_c_2504_n N_VGND_c_2505_n
+ PM_SKY130_FD_SC_HD__SDFBBN_2%VGND
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_1251_47# N_A_1251_47#_M1047_d
+ N_A_1251_47#_M1014_d N_A_1251_47#_c_2713_n N_A_1251_47#_c_2716_n
+ N_A_1251_47#_c_2723_n PM_SKY130_FD_SC_HD__SDFBBN_2%A_1251_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_2%A_2004_47# N_A_2004_47#_M1004_d
+ N_A_2004_47#_M1017_d N_A_2004_47#_c_2748_n N_A_2004_47#_c_2744_n
+ N_A_2004_47#_c_2749_n PM_SKY130_FD_SC_HD__SDFBBN_2%A_2004_47#
cc_1 VNB N_CLK_N_c_308_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_N_c_309_n 0.022961f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK_N 0.0187448f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_N_c_311_n 0.0195341f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_CLK_N_c_312_n 0.0141401f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1028_g 0.0382831f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_354_n 0.0133397f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_27_47#_c_355_n 0.00420241f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_9 VNB N_A_27_47#_M1020_g 0.0199586f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_10 VNB N_A_27_47#_c_357_n 0.00878847f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_11 VNB N_A_27_47#_c_358_n 0.018063f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_12 VNB N_A_27_47#_c_359_n 7.55444e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_360_n 0.00643757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_361_n 0.00302353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_362_n 0.0315468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_363_n 0.00458399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_364_n 0.0327022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_365_n 0.00310819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_366_n 0.0012554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_367_n 0.0212068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_368_n 0.00235584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_369_n 0.00292248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_370_n 0.00200585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_371_n 0.00147534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_372_n 0.0229605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_373_n 0.0249277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_374_n 0.00497848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_SCD_M1006_g 0.0513804f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_29 VNB SCD 0.00784766f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_30 VNB N_A_423_315#_c_669_n 0.00299978f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_31 VNB N_A_423_315#_c_670_n 6.97905e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_32 VNB N_A_423_315#_c_671_n 0.00186605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_423_315#_c_672_n 0.0282104f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_34 VNB N_A_423_315#_c_673_n 0.00348698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_423_315#_c_674_n 0.00275863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_423_315#_c_675_n 0.0162167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_SCE_c_772_n 0.0169394f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_38 VNB N_SCE_c_773_n 0.0467783f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.59
cc_39 VNB N_SCE_c_774_n 0.0183888f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_40 VNB N_SCE_c_775_n 0.0275048f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_41 VNB N_SCE_c_776_n 0.00477854f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_42 VNB N_SCE_c_777_n 0.00444822f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_43 VNB SCE 0.00142423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB SCE 0.00462988f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_45 VNB N_SCE_c_780_n 0.0296743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_D_M1024_g 0.0472628f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_47 VNB N_A_193_47#_c_912_n 0.0180417f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_48 VNB N_A_193_47#_c_913_n 0.0124337f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_49 VNB N_A_193_47#_c_914_n 0.00338665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_193_47#_M1003_g 0.0470935f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_51 VNB N_A_193_47#_c_916_n 0.0042958f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_52 VNB N_A_193_47#_c_917_n 0.0326251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_193_47#_c_918_n 0.0182675f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1107_21#_M1038_g 0.0422736f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_55 VNB N_A_1107_21#_c_1127_n 0.0192786f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_56 VNB N_A_1107_21#_c_1128_n 0.00190301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1107_21#_c_1129_n 0.00419998f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_58 VNB N_A_1107_21#_c_1130_n 0.0114386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1107_21#_c_1131_n 0.00587713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1107_21#_c_1132_n 0.0321305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_SET_B_c_1272_n 0.0324673f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_62 VNB N_SET_B_M1011_g 0.00696335f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_63 VNB N_SET_B_M1047_g 0.0204057f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_64 VNB N_SET_B_M1004_g 0.0200444f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_65 VNB N_SET_B_M1007_g 0.00793898f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_66 VNB SET_B 0.00764108f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_67 VNB N_SET_B_c_1278_n 0.0153139f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_68 VNB N_SET_B_c_1279_n 0.00193382f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_69 VNB N_SET_B_c_1280_n 0.00209085f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_70 VNB N_SET_B_c_1281_n 0.00538514f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_71 VNB N_SET_B_c_1282_n 0.0316983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_931_47#_M1016_g 0.025882f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_73 VNB N_A_931_47#_c_1404_n 0.00430594f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_74 VNB N_A_931_47#_c_1405_n 0.00748589f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_75 VNB N_A_931_47#_c_1406_n 0.00392752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_931_47#_c_1407_n 0.0142922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1401_21#_c_1509_n 0.0176574f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_78 VNB N_A_1401_21#_c_1510_n 0.0338404f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_79 VNB N_A_1401_21#_M1017_g 0.0281252f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_80 VNB N_A_1401_21#_c_1512_n 0.0133934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1401_21#_c_1513_n 0.00176366f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_82 VNB N_A_1401_21#_c_1514_n 0.00736663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1401_21#_c_1515_n 9.08783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1401_21#_c_1516_n 0.0197178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1401_21#_c_1517_n 0.00543093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1888_21#_M1042_g 0.0441996f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_87 VNB N_A_1888_21#_c_1666_n 0.0165362f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_88 VNB N_A_1888_21#_M1051_g 0.0213222f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_89 VNB N_A_1888_21#_M1046_g 5.23365e-19 $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_90 VNB N_A_1888_21#_c_1669_n 0.0538654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1888_21#_c_1670_n 0.0331492f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_92 VNB N_A_1888_21#_c_1671_n 0.00806382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_1888_21#_c_1672_n 4.83176e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_1888_21#_c_1673_n 0.01839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_1888_21#_c_1674_n 0.0183891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_1888_21#_c_1675_n 0.00820903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_1888_21#_c_1676_n 0.00321658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_1888_21#_c_1677_n 0.00365923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_1714_47#_M1001_g 0.0224258f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_100 VNB N_A_1714_47#_c_1861_n 0.0117849f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_101 VNB N_A_1714_47#_c_1862_n 0.0114143f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_102 VNB N_A_1714_47#_c_1863_n 4.91252e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_A_1714_47#_c_1864_n 0.00186712f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_104 VNB N_A_1714_47#_c_1865_n 0.017672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_RESET_B_M1009_g 0.0351078f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_106 VNB RESET_B 0.0040306f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_107 VNB N_RESET_B_c_1961_n 0.0302879f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_108 VNB N_A_2696_47#_c_1995_n 0.0168966f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_109 VNB N_A_2696_47#_c_1996_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_A_2696_47#_c_1997_n 0.00821385f $X=-0.19 $Y=-0.24 $X2=0.24
+ $Y2=1.235
cc_111 VNB N_A_2696_47#_c_1998_n 0.0051319f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_112 VNB N_A_2696_47#_c_1999_n 4.85991e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_A_2696_47#_c_2000_n 0.0519216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VPWR_c_2070_n 0.6303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_A_453_47#_c_2297_n 0.00547438f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_116 VNB N_A_453_47#_c_2298_n 0.00628769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_A_453_47#_c_2299_n 0.00688335f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_118 VNB N_A_453_47#_c_2300_n 0.00860491f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_119 VNB N_A_453_47#_c_2301_n 0.00217312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_A_453_47#_c_2302_n 0.00690765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_A_453_47#_c_2303_n 0.00279367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_A_453_47#_c_2304_n 0.0142904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_Q_N_c_2430_n 0.00127056f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_124 VNB N_Q_c_2454_n 0.00103626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2475_n 4.08532e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2476_n 0.00948744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2477_n 0.00280508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2478_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2479_n 0.00562135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2480_n 0.0024154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2481_n 0.00549276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2482_n 0.0125743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2483_n 0.019615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2484_n 0.00254394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2485_n 0.0101633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2486_n 0.0321728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2487_n 0.0568827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2488_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2489_n 0.0387378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2490_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2491_n 0.0404697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2492_n 0.00372951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2493_n 0.0153564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2494_n 0.0157857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2495_n 0.0448896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2496_n 0.0562803f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2497_n 0.0152053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2498_n 0.0152053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2499_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2500_n 0.00526527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2501_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2502_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2503_n 0.00451684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2504_n 0.00440331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2505_n 0.700949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_156 VPB N_CLK_N_c_313_n 0.0118979f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_157 VPB N_CLK_N_c_314_n 0.0186097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_158 VPB N_CLK_N_c_315_n 0.0238007f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_159 VPB CLK_N 0.0178201f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_160 VPB N_CLK_N_c_311_n 0.0100928f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_161 VPB N_A_27_47#_M1000_g 0.0375468f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_162 VPB N_A_27_47#_M1040_g 0.0466077f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_163 VPB N_A_27_47#_c_354_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_164 VPB N_A_27_47#_c_355_n 0.00338145f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_165 VPB N_A_27_47#_M1021_g 0.0222026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_27_47#_c_380_n 0.0018848f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_27_47#_c_381_n 0.00384216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_27_47#_c_382_n 0.0287783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_27_47#_c_383_n 0.00362242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_27_47#_c_369_n 0.00321856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_27_47#_c_371_n 2.53141e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_27_47#_c_372_n 0.0119012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_SCD_M1006_g 0.00110964f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_174 VPB N_SCD_M1034_g 0.0216746f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_175 VPB SCD 0.00529215f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_176 VPB N_SCD_c_636_n 0.0453337f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_177 VPB N_A_423_315#_c_676_n 0.0180115f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_178 VPB N_A_423_315#_c_677_n 0.0626142f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_179 VPB N_A_423_315#_c_678_n 0.0078776f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_180 VPB N_A_423_315#_c_679_n 0.00298811f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_181 VPB N_A_423_315#_c_680_n 0.0084158f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_182 VPB N_A_423_315#_c_673_n 0.00550351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_423_315#_c_682_n 0.00640598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_SCE_c_775_n 0.0317461f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_185 VPB N_SCE_c_782_n 0.0172669f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_186 VPB N_SCE_c_783_n 0.0252061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_SCE_c_784_n 0.0144423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_SCE_c_785_n 0.00545787f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_189 VPB SCE 0.0083231f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_190 VPB N_D_M1024_g 0.00324838f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_191 VPB N_D_M1019_g 0.036057f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_192 VPB D 0.0116166f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_193 VPB N_D_c_874_n 0.0385655f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_194 VPB N_A_193_47#_M1010_g 0.0215869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_193_47#_M1032_g 0.020906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_193_47#_c_913_n 0.0178865f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_197 VPB N_A_193_47#_c_914_n 0.00403646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_193_47#_c_916_n 0.00245106f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_199 VPB N_A_193_47#_c_924_n 0.0273903f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_200 VPB N_A_193_47#_c_925_n 0.00491076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_193_47#_c_926_n 0.00875464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_193_47#_c_927_n 0.00165292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_193_47#_c_928_n 0.00361706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_193_47#_c_929_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_193_47#_c_930_n 0.00575159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_193_47#_c_931_n 0.0282388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_193_47#_c_932_n 0.00514398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_193_47#_c_933_n 0.0125285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_193_47#_c_918_n 0.0180193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_1107_21#_M1038_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_211 VPB N_A_1107_21#_M1036_g 0.0210587f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_212 VPB N_A_1107_21#_M1050_g 0.0317411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_213 VPB N_A_1107_21#_c_1136_n 0.0055347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_1107_21#_c_1129_n 0.00619371f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_215 VPB N_A_1107_21#_c_1138_n 0.00575673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_1107_21#_c_1139_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_1107_21#_c_1132_n 0.00659461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_SET_B_M1011_g 0.0508831f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_219 VPB N_SET_B_M1007_g 0.0496547f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_220 VPB N_A_931_47#_M1037_g 0.0203673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_221 VPB N_A_931_47#_c_1409_n 0.0121994f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_222 VPB N_A_931_47#_c_1405_n 0.00789134f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_223 VPB N_A_931_47#_c_1406_n 0.00271559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_931_47#_c_1407_n 0.0166796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1401_21#_c_1510_n 0.0218089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_226 VPB N_A_1401_21#_M1031_g 0.0205161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1401_21#_M1029_g 0.0210664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1401_21#_c_1521_n 0.00188964f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_229 VPB N_A_1401_21#_c_1522_n 0.00746077f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_230 VPB N_A_1401_21#_c_1515_n 0.00162652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_1401_21#_c_1524_n 0.0329117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_1401_21#_c_1525_n 0.00261931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_1401_21#_c_1526_n 0.00737873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_1401_21#_c_1527_n 0.00339519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_1401_21#_c_1516_n 0.0263136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_1401_21#_c_1517_n 0.00369973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_A_1888_21#_M1042_g 0.0159543f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_238 VPB N_A_1888_21#_M1043_g 0.021027f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_239 VPB N_A_1888_21#_M1002_g 0.0200318f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_240 VPB N_A_1888_21#_M1046_g 0.0237065f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_241 VPB N_A_1888_21#_c_1670_n 0.00453783f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_242 VPB N_A_1888_21#_c_1672_n 0.0132086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_A_1888_21#_c_1684_n 0.018641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_A_1888_21#_c_1685_n 0.0184285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_A_1888_21#_c_1686_n 0.00421617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_A_1888_21#_c_1687_n 0.0324865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_A_1888_21#_c_1688_n 0.00304218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_A_1888_21#_c_1676_n 0.00331499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_A_1888_21#_c_1690_n 0.00915661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_A_1888_21#_c_1691_n 0.0015533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_A_1714_47#_M1025_g 0.021833f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_252 VPB N_A_1714_47#_c_1867_n 0.0118251f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_253 VPB N_A_1714_47#_c_1862_n 0.00584496f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_254 VPB N_A_1714_47#_c_1863_n 7.62954e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_A_1714_47#_c_1864_n 0.00126723f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_256 VPB N_A_1714_47#_c_1865_n 0.00899175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_RESET_B_M1030_g 0.0251875f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_258 VPB RESET_B 9.6982e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_259 VPB N_RESET_B_c_1961_n 0.0100579f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_260 VPB N_A_2696_47#_M1005_g 0.02086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_A_2696_47#_M1018_g 0.025289f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_262 VPB N_A_2696_47#_c_2003_n 0.0146779f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_263 VPB N_A_2696_47#_c_1998_n 0.00518989f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_264 VPB N_A_2696_47#_c_1999_n 2.42996e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_A_2696_47#_c_2000_n 0.00966347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_2071_n 0.00105358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_2072_n 0.00871789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_2073_n 4.89322e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_2074_n 0.00313724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_2075_n 0.00562862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_2076_n 0.0136158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_2077_n 0.0200059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_2078_n 0.00353766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_2079_n 0.0101374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_2080_n 0.0413727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_2081_n 0.0292737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_2082_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_2083_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_2084_n 0.022998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_2085_n 0.0154511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_2086_n 0.0156521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_2087_n 0.0416309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_2088_n 0.0534515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_2089_n 0.0591311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_2090_n 0.0341009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_2091_n 0.0151994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_2092_n 0.0152053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_2093_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_2094_n 0.00579271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_2095_n 0.00456344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_2096_n 0.00609488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_2097_n 0.00928062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_2098_n 0.00456443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_2099_n 0.00449095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_2100_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_2070_n 0.077822f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_297 VPB N_A_453_47#_c_2297_n 0.00263158f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_298 VPB N_A_453_47#_c_2306_n 0.00579707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_299 VPB N_A_453_47#_c_2307_n 0.00536501f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_300 VPB N_A_453_47#_c_2301_n 3.39779e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_301 VPB N_A_453_47#_c_2302_n 0.00407396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_302 VPB N_A_453_47#_c_2303_n 8.04394e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_303 VPB N_A_453_47#_c_2304_n 0.0146808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_304 VPB N_Q_N_c_2430_n 0.00118478f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_305 VPB N_Q_c_2455_n 9.73602e-19 $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_306 VPB N_Q_c_2454_n 0.00112104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_307 N_CLK_N_c_308_n N_A_27_47#_M1028_g 0.0205277f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_308 CLK_N N_A_27_47#_M1028_g 3.07529e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_309 N_CLK_N_c_312_n N_A_27_47#_M1028_g 0.00498861f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_310 N_CLK_N_c_315_n N_A_27_47#_M1000_g 0.0275641f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_311 CLK_N N_A_27_47#_M1000_g 5.68848e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_312 N_CLK_N_c_311_n N_A_27_47#_M1000_g 0.00521293f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_313 N_CLK_N_c_308_n N_A_27_47#_c_359_n 0.00685438f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_314 N_CLK_N_c_309_n N_A_27_47#_c_359_n 0.00799602f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_315 CLK_N N_A_27_47#_c_359_n 0.00698378f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_316 N_CLK_N_c_309_n N_A_27_47#_c_360_n 0.00621081f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_317 CLK_N N_A_27_47#_c_360_n 0.0148236f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_318 N_CLK_N_c_311_n N_A_27_47#_c_360_n 3.2891e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_319 N_CLK_N_c_314_n N_A_27_47#_c_380_n 0.0129431f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_320 N_CLK_N_c_315_n N_A_27_47#_c_380_n 0.0013404f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_321 CLK_N N_A_27_47#_c_380_n 0.00690269f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_322 N_CLK_N_c_314_n N_A_27_47#_c_383_n 2.18052e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_323 N_CLK_N_c_315_n N_A_27_47#_c_383_n 0.00374438f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_324 CLK_N N_A_27_47#_c_383_n 0.0157801f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_325 N_CLK_N_c_311_n N_A_27_47#_c_383_n 2.59784e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_326 N_CLK_N_c_309_n N_A_27_47#_c_365_n 0.0017166f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_327 N_CLK_N_c_312_n N_A_27_47#_c_365_n 0.00154887f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_328 N_CLK_N_c_309_n N_A_27_47#_c_369_n 0.00155723f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_329 N_CLK_N_c_315_n N_A_27_47#_c_369_n 0.0045823f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_330 CLK_N N_A_27_47#_c_369_n 0.0517134f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_331 N_CLK_N_c_311_n N_A_27_47#_c_369_n 0.00100166f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_332 N_CLK_N_c_312_n N_A_27_47#_c_369_n 0.00207651f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_333 CLK_N N_A_27_47#_c_372_n 0.00162145f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_334 N_CLK_N_c_311_n N_A_27_47#_c_372_n 0.0169859f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_335 N_CLK_N_c_314_n N_VPWR_c_2071_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_336 N_CLK_N_c_314_n N_VPWR_c_2085_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_337 N_CLK_N_c_314_n N_VPWR_c_2070_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_338 N_CLK_N_c_308_n N_VGND_c_2475_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_339 N_CLK_N_c_308_n N_VGND_c_2493_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_340 N_CLK_N_c_309_n N_VGND_c_2493_n 4.87495e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_341 N_CLK_N_c_308_n N_VGND_c_2505_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_342 N_A_27_47#_c_364_n N_SCD_M1006_g 0.0120872f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_343 N_A_27_47#_c_364_n SCD 0.00948568f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_344 N_A_27_47#_c_364_n N_SCD_c_636_n 0.00128241f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_345 N_A_27_47#_c_372_n N_SCD_c_636_n 0.00542368f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_364_n N_A_423_315#_c_669_n 0.0197158f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_364_n N_A_423_315#_c_670_n 0.00685013f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_364_n N_A_423_315#_c_671_n 0.014943f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_364_n N_A_423_315#_c_672_n 0.00180177f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_364_n N_SCE_c_773_n 0.00565864f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_351 N_A_27_47#_c_364_n N_SCE_c_775_n 0.00239268f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_352 N_A_27_47#_c_364_n N_SCE_c_776_n 4.50186e-19 $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_353 N_A_27_47#_c_364_n N_SCE_c_777_n 0.0291484f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_364_n SCE 0.00178707f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_364_n SCE 0.00106129f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_356 N_A_27_47#_c_364_n N_SCE_c_780_n 0.00371035f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_355_n N_D_M1024_g 0.0186046f $X=4.665 $Y=1.32 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_364_n N_D_M1024_g 0.00630058f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_359 N_A_27_47#_M1040_g N_D_c_874_n 0.0186046f $X=4.59 $Y=2.275 $X2=0 $Y2=0
cc_360 N_A_27_47#_M1020_g N_A_193_47#_c_912_n 0.0127842f $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_374_n N_A_193_47#_c_912_n 4.90539e-19 $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_M1040_g N_A_193_47#_M1010_g 0.0190155f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_363_n N_A_193_47#_c_913_n 0.0110561f $X=8.937 $Y=1.305 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_381_n N_A_193_47#_c_913_n 0.00853911f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_382_n N_A_193_47#_c_913_n 0.0216716f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_371_n N_A_193_47#_c_913_n 3.23054e-19 $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_361_n N_A_193_47#_c_914_n 2.62384e-19 $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_362_n N_A_193_47#_c_914_n 0.0209335f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_363_n N_A_193_47#_c_914_n 0.00356667f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_371_n N_A_193_47#_c_914_n 9.01357e-19 $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_358_n N_A_193_47#_M1003_g 0.0129153f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_361_n N_A_193_47#_M1003_g 0.00307377f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_362_n N_A_193_47#_M1003_g 0.021369f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_363_n N_A_193_47#_M1003_g 0.00622479f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_M1040_g N_A_193_47#_c_916_n 0.00534395f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_354_n N_A_193_47#_c_916_n 0.010154f $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_355_n N_A_193_47#_c_916_n 0.00203307f $X=4.665 $Y=1.32 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_M1020_g N_A_193_47#_c_916_n 4.45841e-19 $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_364_n N_A_193_47#_c_916_n 0.0155618f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_366_n N_A_193_47#_c_916_n 0.00934078f $X=5.327 $Y=1.12 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_370_n N_A_193_47#_c_916_n 4.74166e-19 $X=5.29 $Y=0.85 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_373_n N_A_193_47#_c_916_n 0.00674133f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_374_n N_A_193_47#_c_916_n 0.0210004f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_355_n N_A_193_47#_c_917_n 0.0232669f $X=4.665 $Y=1.32 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_M1020_g N_A_193_47#_c_917_n 0.0214266f $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_364_n N_A_193_47#_c_917_n 0.00553622f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_374_n N_A_193_47#_c_917_n 0.00154674f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_M1040_g N_A_193_47#_c_924_n 0.00696374f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1000_g N_A_193_47#_c_925_n 0.00459685f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_380_n N_A_193_47#_c_925_n 0.00561276f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_369_n N_A_193_47#_c_925_n 0.00113557f $X=0.69 $Y=0.85 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_354_n N_A_193_47#_c_926_n 3.83457e-19 $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_368_n N_A_193_47#_c_926_n 0.111295f $X=5.435 $Y=1.19 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_M1040_g N_A_193_47#_c_927_n 5.24592e-19 $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_M1021_g N_A_193_47#_c_928_n 0.00133927f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_c_381_n N_A_193_47#_c_928_n 0.00483121f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_382_n N_A_193_47#_c_928_n 0.00219663f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_M1040_g N_A_193_47#_c_929_n 0.0174486f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_354_n N_A_193_47#_c_929_n 0.0212221f $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_374_n N_A_193_47#_c_929_n 3.18577e-19 $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_M1040_g N_A_193_47#_c_930_n 0.00867228f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_354_n N_A_193_47#_c_930_n 0.00654686f $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_374_n N_A_193_47#_c_930_n 0.00339609f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_M1021_g N_A_193_47#_c_931_n 0.0192968f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_c_381_n N_A_193_47#_c_931_n 5.88448e-19 $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_382_n N_A_193_47#_c_931_n 0.0169266f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_367_n N_A_193_47#_c_931_n 2.37019e-19 $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_M1021_g N_A_193_47#_c_932_n 6.52047e-19 $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_363_n N_A_193_47#_c_932_n 0.00682571f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_381_n N_A_193_47#_c_932_n 0.0168759f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_c_382_n N_A_193_47#_c_932_n 0.00153059f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_c_371_n N_A_193_47#_c_932_n 0.00149027f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_381_n N_A_193_47#_c_933_n 0.00347329f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_M1028_g N_A_193_47#_c_918_n 0.023031f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_359_n N_A_193_47#_c_918_n 0.0113579f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_380_n N_A_193_47#_c_918_n 0.00860312f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_364_n N_A_193_47#_c_918_n 0.0271407f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_365_n N_A_193_47#_c_918_n 0.00145827f $X=0.835 $Y=0.85 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_369_n N_A_193_47#_c_918_n 0.0688642f $X=0.69 $Y=0.85 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_M1020_g N_A_1107_21#_M1038_g 0.0245694f $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_357_n N_A_1107_21#_M1038_g 0.0105189f $X=5.13 $Y=1.245 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_367_n N_A_1107_21#_M1038_g 7.74803e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_370_n N_A_1107_21#_M1038_g 0.00642269f $X=5.29 $Y=0.85 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_373_n N_A_1107_21#_M1038_g 0.0200662f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_374_n N_A_1107_21#_M1038_g 0.00189958f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_c_358_n N_A_1107_21#_c_1127_n 0.0187265f $X=8.495 $Y=0.705
+ $X2=0 $Y2=0
cc_427 N_A_27_47#_c_361_n N_A_1107_21#_c_1127_n 0.001702f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_367_n N_A_1107_21#_c_1136_n 0.00196084f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_367_n N_A_1107_21#_c_1150_n 0.00348372f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_367_n N_A_1107_21#_c_1128_n 0.0016677f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_367_n N_A_1107_21#_c_1129_n 0.016449f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_c_367_n N_A_1107_21#_c_1130_n 0.00904925f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_367_n N_A_1107_21#_c_1138_n 8.24776e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_c_367_n N_A_1107_21#_c_1155_n 6.83984e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_361_n N_A_1107_21#_c_1131_n 0.0111636f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_362_n N_A_1107_21#_c_1131_n 9.14426e-19 $X=8.62 $Y=0.87
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_363_n N_A_1107_21#_c_1131_n 0.00462764f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_367_n N_A_1107_21#_c_1131_n 0.0153364f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_371_n N_A_1107_21#_c_1131_n 0.00129536f $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_361_n N_A_1107_21#_c_1132_n 5.13187e-19 $X=8.62 $Y=0.87
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_362_n N_A_1107_21#_c_1132_n 0.0187265f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_363_n N_A_1107_21#_c_1132_n 0.00174717f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_367_n N_A_1107_21#_c_1132_n 0.00365485f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_371_n N_A_1107_21#_c_1132_n 6.8647e-19 $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_367_n N_SET_B_c_1272_n 0.00392015f $X=8.365 $Y=1.19
+ $X2=-0.19 $Y2=-0.24
cc_446 N_A_27_47#_c_367_n N_SET_B_M1011_g 0.0011704f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_367_n SET_B 0.00593372f $X=8.365 $Y=1.19 $X2=0 $Y2=0
cc_448 N_A_27_47#_c_361_n N_SET_B_c_1278_n 0.0194369f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_362_n N_SET_B_c_1278_n 0.0023282f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_363_n N_SET_B_c_1278_n 0.0053562f $X=8.937 $Y=1.305 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_367_n N_SET_B_c_1278_n 0.158116f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_371_n N_SET_B_c_1278_n 0.0254944f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_c_367_n N_SET_B_c_1279_n 0.0265123f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_367_n N_A_931_47#_M1016_g 0.00190146f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_M1040_g N_A_931_47#_c_1414_n 0.00264322f $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_456 N_A_27_47#_M1020_g N_A_931_47#_c_1415_n 0.00883573f $X=5.13 $Y=0.415
+ $X2=0 $Y2=0
cc_457 N_A_27_47#_c_364_n N_A_931_47#_c_1415_n 0.00579266f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_458 N_A_27_47#_c_370_n N_A_931_47#_c_1415_n 0.00257401f $X=5.29 $Y=0.85 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_373_n N_A_931_47#_c_1415_n 5.24878e-19 $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_374_n N_A_931_47#_c_1415_n 0.0194937f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_M1040_g N_A_931_47#_c_1409_n 8.73767e-19 $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_462 N_A_27_47#_c_368_n N_A_931_47#_c_1409_n 3.03433e-19 $X=5.435 $Y=1.19
+ $X2=0 $Y2=0
cc_463 N_A_27_47#_M1020_g N_A_931_47#_c_1404_n 0.00119254f $X=5.13 $Y=0.415
+ $X2=0 $Y2=0
cc_464 N_A_27_47#_c_357_n N_A_931_47#_c_1404_n 8.54957e-19 $X=5.13 $Y=1.245
+ $X2=0 $Y2=0
cc_465 N_A_27_47#_c_367_n N_A_931_47#_c_1404_n 0.0145635f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_370_n N_A_931_47#_c_1404_n 0.0138897f $X=5.29 $Y=0.85 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_373_n N_A_931_47#_c_1404_n 7.78235e-19 $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_374_n N_A_931_47#_c_1404_n 0.0244377f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_c_367_n N_A_931_47#_c_1405_n 0.0375702f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_357_n N_A_931_47#_c_1406_n 0.00268952f $X=5.13 $Y=1.245
+ $X2=0 $Y2=0
cc_471 N_A_27_47#_c_367_n N_A_931_47#_c_1406_n 0.0109965f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_368_n N_A_931_47#_c_1406_n 0.00666557f $X=5.435 $Y=1.19
+ $X2=0 $Y2=0
cc_473 N_A_27_47#_c_373_n N_A_931_47#_c_1406_n 5.70846e-19 $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_374_n N_A_931_47#_c_1406_n 0.0053097f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_367_n N_A_931_47#_c_1407_n 0.00390921f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_476 N_A_27_47#_c_367_n N_A_1401_21#_c_1510_n 0.0075896f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_477 N_A_27_47#_c_367_n N_A_1401_21#_c_1515_n 0.0122882f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_478 N_A_27_47#_c_363_n N_A_1401_21#_c_1524_n 0.00715591f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_479 N_A_27_47#_c_381_n N_A_1401_21#_c_1524_n 0.0157692f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_480 N_A_27_47#_c_382_n N_A_1401_21#_c_1524_n 0.00184742f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_481 N_A_27_47#_c_367_n N_A_1401_21#_c_1524_n 0.014133f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_371_n N_A_1401_21#_c_1524_n 0.027417f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_367_n N_A_1401_21#_c_1525_n 0.0276968f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_484 N_A_27_47#_c_381_n N_A_1401_21#_c_1526_n 0.00264766f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_485 N_A_27_47#_c_367_n N_A_1401_21#_c_1526_n 0.00618009f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_486 N_A_27_47#_c_381_n N_A_1888_21#_M1042_g 3.51933e-19 $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_487 N_A_27_47#_M1021_g N_A_1888_21#_c_1687_n 0.0162278f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_488 N_A_27_47#_c_382_n N_A_1888_21#_c_1687_n 0.00879184f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_489 N_A_27_47#_M1021_g N_A_1714_47#_c_1872_n 0.00935459f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_490 N_A_27_47#_c_381_n N_A_1714_47#_c_1872_n 0.00669245f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_491 N_A_27_47#_c_382_n N_A_1714_47#_c_1872_n 0.0028948f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_492 N_A_27_47#_c_361_n N_A_1714_47#_c_1875_n 0.00390894f $X=8.62 $Y=0.87
+ $X2=0 $Y2=0
cc_493 N_A_27_47#_c_362_n N_A_1714_47#_c_1875_n 0.00184507f $X=8.62 $Y=0.87
+ $X2=0 $Y2=0
cc_494 N_A_27_47#_c_363_n N_A_1714_47#_c_1875_n 0.00315233f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_495 N_A_27_47#_c_361_n N_A_1714_47#_c_1861_n 0.0117718f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_c_363_n N_A_1714_47#_c_1861_n 0.00837612f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_497 N_A_27_47#_c_371_n N_A_1714_47#_c_1861_n 6.65017e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_498 N_A_27_47#_M1021_g N_A_1714_47#_c_1867_n 0.00655877f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_499 N_A_27_47#_c_381_n N_A_1714_47#_c_1867_n 0.0359925f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_500 N_A_27_47#_c_382_n N_A_1714_47#_c_1867_n 0.00212049f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_501 N_A_27_47#_c_363_n N_A_1714_47#_c_1863_n 0.00588724f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_502 N_A_27_47#_c_381_n N_A_1714_47#_c_1863_n 0.00820578f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_503 N_A_27_47#_c_371_n N_A_1714_47#_c_1863_n 2.68785e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_504 N_A_27_47#_c_380_n N_VPWR_M1027_d 0.00165787f $X=0.605 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_505 N_A_27_47#_M1000_g N_VPWR_c_2071_n 0.00864163f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_c_380_n N_VPWR_c_2071_n 0.0171178f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_383_n N_VPWR_c_2071_n 0.0127225f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_508 N_A_27_47#_M1000_g N_VPWR_c_2072_n 0.00232641f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_c_380_n N_VPWR_c_2085_n 0.0018545f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_c_383_n N_VPWR_c_2085_n 0.0123893f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_511 N_A_27_47#_M1000_g N_VPWR_c_2086_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_512 N_A_27_47#_M1040_g N_VPWR_c_2088_n 0.00541732f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_M1021_g N_VPWR_c_2089_n 0.00367119f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_M1000_g N_VPWR_c_2070_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_515 N_A_27_47#_M1040_g N_VPWR_c_2070_n 0.00632491f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_M1021_g N_VPWR_c_2070_n 0.00567418f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_380_n N_VPWR_c_2070_n 0.00505319f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_518 N_A_27_47#_c_383_n N_VPWR_c_2070_n 0.00665993f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_519 N_A_27_47#_c_364_n N_A_453_47#_c_2297_n 0.00441112f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_520 N_A_27_47#_c_364_n N_A_453_47#_c_2298_n 0.0192062f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_c_364_n N_A_453_47#_c_2299_n 0.00519492f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_522 N_A_27_47#_c_364_n N_A_453_47#_c_2300_n 0.0879477f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_523 N_A_27_47#_c_364_n N_A_453_47#_c_2301_n 0.0279195f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_524 N_A_27_47#_c_364_n N_A_453_47#_c_2302_n 0.00691629f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_525 N_A_27_47#_c_355_n N_A_453_47#_c_2303_n 0.00125006f $X=4.665 $Y=1.32
+ $X2=0 $Y2=0
cc_526 N_A_27_47#_c_364_n N_A_453_47#_c_2303_n 0.0256464f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_527 N_A_27_47#_c_355_n N_A_453_47#_c_2304_n 0.0156881f $X=4.665 $Y=1.32 $X2=0
+ $Y2=0
cc_528 N_A_27_47#_c_364_n N_A_453_47#_c_2304_n 0.0170158f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_529 N_A_27_47#_c_374_n N_A_453_47#_c_2304_n 0.00205629f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_530 N_A_27_47#_c_359_n N_VGND_M1048_d 0.00162876f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_531 N_A_27_47#_M1028_g N_VGND_c_2475_n 0.00789067f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_532 N_A_27_47#_c_359_n N_VGND_c_2475_n 0.0154833f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_533 N_A_27_47#_c_364_n N_VGND_c_2475_n 2.30481e-19 $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_534 N_A_27_47#_c_365_n N_VGND_c_2475_n 0.00116209f $X=0.835 $Y=0.85 $X2=0
+ $Y2=0
cc_535 N_A_27_47#_c_372_n N_VGND_c_2475_n 5.88506e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_536 N_A_27_47#_M1028_g N_VGND_c_2476_n 0.00327532f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_537 N_A_27_47#_c_364_n N_VGND_c_2476_n 0.00475891f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_538 N_A_27_47#_c_364_n N_VGND_c_2477_n 0.00131319f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_539 N_A_27_47#_c_358_n N_VGND_c_2479_n 0.00174046f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_540 N_A_27_47#_M1020_g N_VGND_c_2487_n 0.00359964f $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_541 N_A_27_47#_c_358_n N_VGND_c_2491_n 0.00435972f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_542 N_A_27_47#_c_361_n N_VGND_c_2491_n 0.00288727f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_543 N_A_27_47#_c_362_n N_VGND_c_2491_n 2.15978e-19 $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_544 N_A_27_47#_c_617_p N_VGND_c_2493_n 0.00735289f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_545 N_A_27_47#_c_359_n N_VGND_c_2493_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_546 N_A_27_47#_M1028_g N_VGND_c_2494_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_547 N_A_27_47#_M1048_s N_VGND_c_2505_n 0.00358206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_548 N_A_27_47#_M1028_g N_VGND_c_2505_n 0.00581646f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_549 N_A_27_47#_M1020_g N_VGND_c_2505_n 0.00564268f $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_550 N_A_27_47#_c_358_n N_VGND_c_2505_n 0.00616197f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_551 N_A_27_47#_c_617_p N_VGND_c_2505_n 0.00626856f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_552 N_A_27_47#_c_359_n N_VGND_c_2505_n 0.00523689f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_553 N_A_27_47#_c_361_n N_VGND_c_2505_n 0.00224883f $X=8.62 $Y=0.87 $X2=0
+ $Y2=0
cc_554 N_A_27_47#_c_364_n N_VGND_c_2505_n 0.20509f $X=5.145 $Y=0.85 $X2=0 $Y2=0
cc_555 N_A_27_47#_c_365_n N_VGND_c_2505_n 0.0131302f $X=0.835 $Y=0.85 $X2=0
+ $Y2=0
cc_556 N_A_27_47#_c_370_n N_VGND_c_2505_n 0.0153531f $X=5.29 $Y=0.85 $X2=0 $Y2=0
cc_557 N_A_27_47#_c_374_n A_1041_47# 0.00109904f $X=5.19 $Y=0.93 $X2=-0.19
+ $Y2=-0.24
cc_558 N_SCD_M1034_g N_A_423_315#_c_676_n 0.0310159f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_559 N_SCD_c_636_n N_A_423_315#_c_678_n 0.0310159f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_560 N_SCD_M1006_g N_SCE_c_772_n 0.0604681f $X=1.83 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_561 N_SCD_M1006_g N_SCE_c_777_n 0.00706125f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_562 SCD N_SCE_c_777_n 0.0045361f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_563 N_SCD_M1006_g SCE 0.00375261f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_564 N_SCD_M1006_g SCE 0.0139689f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_565 SCD SCE 0.0355883f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_566 N_SCD_M1034_g N_A_193_47#_c_924_n 0.00922354f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_567 SCD N_A_193_47#_c_924_n 0.00832905f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_568 N_SCD_c_636_n N_A_193_47#_c_924_n 0.00149424f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_569 N_SCD_M1034_g N_A_193_47#_c_925_n 9.04442e-19 $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_570 N_SCD_M1006_g N_A_193_47#_c_918_n 0.00875591f $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_571 N_SCD_M1034_g N_A_193_47#_c_918_n 0.00414955f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_572 SCD N_A_193_47#_c_918_n 0.0505627f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_573 N_SCD_c_636_n N_A_193_47#_c_918_n 0.00111062f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_574 N_SCD_M1034_g N_VPWR_c_2072_n 0.0154916f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_575 SCD N_VPWR_c_2072_n 0.0161253f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_576 N_SCD_c_636_n N_VPWR_c_2072_n 0.00297773f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_577 N_SCD_M1034_g N_VPWR_c_2087_n 0.00442511f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_578 N_SCD_M1034_g N_VPWR_c_2070_n 0.00418686f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_579 N_SCD_M1006_g N_A_453_47#_c_2297_n 3.71745e-19 $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_580 N_SCD_M1034_g N_A_453_47#_c_2306_n 0.00153013f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_581 N_SCD_M1006_g N_VGND_c_2476_n 0.00528037f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_582 SCD N_VGND_c_2476_n 0.00677187f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_583 N_SCD_c_636_n N_VGND_c_2476_n 0.00111441f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_584 N_SCD_M1006_g N_VGND_c_2495_n 0.00585385f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_585 N_SCD_M1006_g N_VGND_c_2505_n 0.00755725f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_586 N_A_423_315#_c_677_n N_SCE_c_773_n 0.00548373f $X=2.695 $Y=1.65 $X2=0
+ $Y2=0
cc_587 N_A_423_315#_c_680_n N_SCE_c_773_n 4.14413e-19 $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_588 N_A_423_315#_c_669_n N_SCE_c_773_n 0.00142101f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_589 N_A_423_315#_c_670_n N_SCE_c_773_n 0.00634935f $X=3.125 $Y=0.71 $X2=0
+ $Y2=0
cc_590 N_A_423_315#_c_669_n N_SCE_c_774_n 0.00766385f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_591 N_A_423_315#_c_675_n N_SCE_c_774_n 0.0157579f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_592 N_A_423_315#_c_677_n N_SCE_c_775_n 0.0213525f $X=2.695 $Y=1.65 $X2=0
+ $Y2=0
cc_593 N_A_423_315#_c_680_n N_SCE_c_775_n 0.0110911f $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_594 N_A_423_315#_c_682_n N_SCE_c_775_n 0.0100429f $X=2.905 $Y=1.66 $X2=0
+ $Y2=0
cc_595 N_A_423_315#_c_674_n N_SCE_c_775_n 0.00669901f $X=3.622 $Y=1.095 $X2=0
+ $Y2=0
cc_596 N_A_423_315#_c_680_n N_SCE_c_783_n 0.00779447f $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_597 N_A_423_315#_c_669_n N_SCE_c_776_n 0.00574578f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_598 N_A_423_315#_c_671_n N_SCE_c_776_n 0.00669901f $X=3.685 $Y=0.93 $X2=0
+ $Y2=0
cc_599 N_A_423_315#_c_672_n N_SCE_c_776_n 0.0207451f $X=3.685 $Y=0.93 $X2=0
+ $Y2=0
cc_600 N_A_423_315#_c_675_n N_SCE_c_776_n 9.51141e-19 $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_601 N_A_423_315#_c_679_n N_SCE_c_785_n 0.0098827f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_602 N_A_423_315#_c_678_n N_SCE_c_777_n 0.0011491f $X=2.265 $Y=1.65 $X2=0
+ $Y2=0
cc_603 N_A_423_315#_c_678_n SCE 0.00459591f $X=2.265 $Y=1.65 $X2=0 $Y2=0
cc_604 N_A_423_315#_c_678_n N_SCE_c_780_n 0.00903235f $X=2.265 $Y=1.65 $X2=0
+ $Y2=0
cc_605 N_A_423_315#_c_671_n N_D_M1024_g 0.00105116f $X=3.685 $Y=0.93 $X2=0 $Y2=0
cc_606 N_A_423_315#_c_673_n N_D_M1024_g 0.00175438f $X=3.56 $Y=1.575 $X2=0 $Y2=0
cc_607 N_A_423_315#_c_675_n N_D_M1024_g 0.0616329f $X=3.685 $Y=0.765 $X2=0 $Y2=0
cc_608 N_A_423_315#_c_680_n D 0.0135689f $X=3.475 $Y=1.66 $X2=0 $Y2=0
cc_609 N_A_423_315#_c_673_n D 0.017414f $X=3.56 $Y=1.575 $X2=0 $Y2=0
cc_610 N_A_423_315#_c_680_n N_D_c_874_n 4.98039e-19 $X=3.475 $Y=1.66 $X2=0 $Y2=0
cc_611 N_A_423_315#_c_672_n N_D_c_874_n 0.00265425f $X=3.685 $Y=0.93 $X2=0 $Y2=0
cc_612 N_A_423_315#_c_673_n N_D_c_874_n 0.00200746f $X=3.56 $Y=1.575 $X2=0 $Y2=0
cc_613 N_A_423_315#_c_676_n N_A_193_47#_c_924_n 0.006798f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_614 N_A_423_315#_c_677_n N_A_193_47#_c_924_n 0.008988f $X=2.695 $Y=1.65 $X2=0
+ $Y2=0
cc_615 N_A_423_315#_c_679_n N_A_193_47#_c_924_n 0.00711261f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_616 N_A_423_315#_c_680_n N_A_193_47#_c_924_n 0.014472f $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_617 N_A_423_315#_c_682_n N_A_193_47#_c_924_n 0.0160437f $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_618 N_A_423_315#_c_676_n N_VPWR_c_2072_n 0.00275879f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_619 N_A_423_315#_c_679_n N_VPWR_c_2073_n 0.0146793f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_620 N_A_423_315#_c_680_n N_VPWR_c_2073_n 0.00517239f $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_621 N_A_423_315#_c_676_n N_VPWR_c_2087_n 0.00489197f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_622 N_A_423_315#_c_679_n N_VPWR_c_2087_n 0.0118139f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_623 N_A_423_315#_M1035_s N_VPWR_c_2070_n 0.00335142f $X=2.855 $Y=2.065 $X2=0
+ $Y2=0
cc_624 N_A_423_315#_c_676_n N_VPWR_c_2070_n 0.00669614f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_625 N_A_423_315#_c_677_n N_VPWR_c_2070_n 2.96327e-19 $X=2.695 $Y=1.65 $X2=0
+ $Y2=0
cc_626 N_A_423_315#_c_679_n N_VPWR_c_2070_n 0.00308197f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_627 N_A_423_315#_c_682_n N_VPWR_c_2070_n 0.00196684f $X=2.905 $Y=1.66 $X2=0
+ $Y2=0
cc_628 N_A_423_315#_c_677_n N_A_453_47#_c_2297_n 0.00489054f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_629 N_A_423_315#_c_732_p N_A_453_47#_c_2298_n 0.00178467f $X=3.04 $Y=0.47
+ $X2=0 $Y2=0
cc_630 N_A_423_315#_c_670_n N_A_453_47#_c_2298_n 0.0110413f $X=3.125 $Y=0.71
+ $X2=0 $Y2=0
cc_631 N_A_423_315#_c_676_n N_A_453_47#_c_2306_n 0.0101367f $X=2.19 $Y=1.725
+ $X2=0 $Y2=0
cc_632 N_A_423_315#_c_677_n N_A_453_47#_c_2306_n 0.00422041f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_633 N_A_423_315#_c_679_n N_A_453_47#_c_2306_n 0.0237696f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_634 N_A_423_315#_c_676_n N_A_453_47#_c_2307_n 0.00285053f $X=2.19 $Y=1.725
+ $X2=0 $Y2=0
cc_635 N_A_423_315#_c_677_n N_A_453_47#_c_2307_n 0.0153223f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_636 N_A_423_315#_c_682_n N_A_453_47#_c_2307_n 0.0234269f $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_637 N_A_423_315#_c_732_p N_A_453_47#_c_2299_n 0.018839f $X=3.04 $Y=0.47 $X2=0
+ $Y2=0
cc_638 N_A_423_315#_c_680_n N_A_453_47#_c_2300_n 0.00811555f $X=3.475 $Y=1.66
+ $X2=0 $Y2=0
cc_639 N_A_423_315#_c_669_n N_A_453_47#_c_2300_n 0.00315275f $X=3.475 $Y=0.71
+ $X2=0 $Y2=0
cc_640 N_A_423_315#_c_672_n N_A_453_47#_c_2300_n 3.93982e-19 $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_641 N_A_423_315#_c_673_n N_A_453_47#_c_2300_n 0.0158823f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_642 N_A_423_315#_c_674_n N_A_453_47#_c_2300_n 0.00384754f $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_643 N_A_423_315#_c_680_n N_A_453_47#_c_2301_n 0.00168869f $X=3.475 $Y=1.66
+ $X2=0 $Y2=0
cc_644 N_A_423_315#_c_670_n N_A_453_47#_c_2301_n 0.00128058f $X=3.125 $Y=0.71
+ $X2=0 $Y2=0
cc_645 N_A_423_315#_c_673_n N_A_453_47#_c_2301_n 0.0011872f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_646 N_A_423_315#_c_682_n N_A_453_47#_c_2301_n 8.39711e-19 $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_647 N_A_423_315#_c_674_n N_A_453_47#_c_2301_n 0.00120978f $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_648 N_A_423_315#_c_677_n N_A_453_47#_c_2302_n 0.0015103f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_649 N_A_423_315#_c_680_n N_A_453_47#_c_2302_n 6.94166e-19 $X=3.475 $Y=1.66
+ $X2=0 $Y2=0
cc_650 N_A_423_315#_c_670_n N_A_453_47#_c_2302_n 0.00489394f $X=3.125 $Y=0.71
+ $X2=0 $Y2=0
cc_651 N_A_423_315#_c_682_n N_A_453_47#_c_2302_n 0.0236855f $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_652 N_A_423_315#_c_674_n N_A_453_47#_c_2302_n 0.0112934f $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_653 N_A_423_315#_c_673_n N_A_453_47#_c_2303_n 0.00152543f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_654 N_A_423_315#_c_674_n N_A_453_47#_c_2303_n 4.68942e-19 $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_655 N_A_423_315#_c_669_n N_A_453_47#_c_2304_n 0.00480985f $X=3.475 $Y=0.71
+ $X2=0 $Y2=0
cc_656 N_A_423_315#_c_671_n N_A_453_47#_c_2304_n 0.00870657f $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_657 N_A_423_315#_c_673_n N_A_453_47#_c_2304_n 0.00442233f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_658 N_A_423_315#_c_669_n N_VGND_M1013_d 0.00246138f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_659 N_A_423_315#_c_669_n N_VGND_c_2477_n 0.0177928f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_660 N_A_423_315#_c_672_n N_VGND_c_2477_n 4.49423e-19 $X=3.685 $Y=0.93 $X2=0
+ $Y2=0
cc_661 N_A_423_315#_c_675_n N_VGND_c_2477_n 0.00914963f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_662 N_A_423_315#_c_675_n N_VGND_c_2487_n 0.0046653f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_663 N_A_423_315#_c_732_p N_VGND_c_2495_n 0.00857854f $X=3.04 $Y=0.47 $X2=0
+ $Y2=0
cc_664 N_A_423_315#_c_669_n N_VGND_c_2495_n 0.00345019f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_665 N_A_423_315#_M1013_s N_VGND_c_2505_n 0.00206506f $X=2.915 $Y=0.235 $X2=0
+ $Y2=0
cc_666 N_A_423_315#_c_732_p N_VGND_c_2505_n 0.00294183f $X=3.04 $Y=0.47 $X2=0
+ $Y2=0
cc_667 N_A_423_315#_c_669_n N_VGND_c_2505_n 0.00513527f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_668 N_A_423_315#_c_675_n N_VGND_c_2505_n 0.00398879f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_669 N_SCE_c_775_n N_D_M1024_g 0.00323589f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_670 N_SCE_c_775_n N_D_M1019_g 0.00214944f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_671 N_SCE_c_783_n N_D_M1019_g 0.0334116f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_672 N_SCE_c_775_n D 0.00166353f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_673 N_SCE_c_783_n D 0.0100165f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_674 N_SCE_c_775_n N_D_c_874_n 0.00552281f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_675 N_SCE_c_775_n N_A_193_47#_c_924_n 0.0020833f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_676 N_SCE_c_783_n N_A_193_47#_c_924_n 0.0106145f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_677 N_SCE_c_785_n N_A_193_47#_c_924_n 0.0038272f $X=3.265 $Y=1.91 $X2=0 $Y2=0
cc_678 SCE N_A_193_47#_c_924_n 0.0117978f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_679 N_SCE_c_782_n N_VPWR_c_2073_n 0.0105013f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_680 N_SCE_c_783_n N_VPWR_c_2073_n 0.00200314f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_681 N_SCE_c_784_n N_VPWR_c_2073_n 0.0092059f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_682 N_SCE_c_782_n N_VPWR_c_2087_n 0.00407992f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_683 N_SCE_c_784_n N_VPWR_c_2088_n 0.0046653f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_684 N_SCE_c_782_n N_VPWR_c_2070_n 0.00533244f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_685 N_SCE_c_784_n N_VPWR_c_2070_n 0.00446764f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_686 N_SCE_c_773_n N_A_453_47#_c_2297_n 5.83037e-19 $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_687 N_SCE_c_777_n N_A_453_47#_c_2297_n 0.00122047f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_688 SCE N_A_453_47#_c_2297_n 0.0175098f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_689 N_SCE_c_780_n N_A_453_47#_c_2297_n 6.70284e-19 $X=2.415 $Y=0.915 $X2=0
+ $Y2=0
cc_690 N_SCE_c_772_n N_A_453_47#_c_2298_n 0.00214969f $X=2.19 $Y=0.735 $X2=0
+ $Y2=0
cc_691 N_SCE_c_773_n N_A_453_47#_c_2298_n 0.0133696f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_692 N_SCE_c_774_n N_A_453_47#_c_2298_n 3.87637e-19 $X=3.25 $Y=0.735 $X2=0
+ $Y2=0
cc_693 N_SCE_c_775_n N_A_453_47#_c_2298_n 0.00445882f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_694 N_SCE_c_777_n N_A_453_47#_c_2298_n 0.0172138f $X=2.25 $Y=0.93 $X2=0 $Y2=0
cc_695 SCE N_A_453_47#_c_2298_n 0.00621319f $X=1.975 $Y=0.425 $X2=0 $Y2=0
cc_696 N_SCE_c_780_n N_A_453_47#_c_2298_n 0.00422791f $X=2.415 $Y=0.915 $X2=0
+ $Y2=0
cc_697 N_SCE_c_775_n N_A_453_47#_c_2307_n 0.00365885f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_698 SCE N_A_453_47#_c_2307_n 0.0160493f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_699 N_SCE_c_773_n N_A_453_47#_c_2299_n 9.34339e-19 $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_700 N_SCE_c_774_n N_A_453_47#_c_2299_n 9.21804e-19 $X=3.25 $Y=0.735 $X2=0
+ $Y2=0
cc_701 N_SCE_c_777_n N_A_453_47#_c_2299_n 0.00112761f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_702 N_SCE_c_780_n N_A_453_47#_c_2299_n 0.006857f $X=2.415 $Y=0.915 $X2=0
+ $Y2=0
cc_703 N_SCE_c_775_n N_A_453_47#_c_2300_n 0.00696234f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_704 N_SCE_c_783_n N_A_453_47#_c_2300_n 5.63442e-19 $X=3.61 $Y=1.91 $X2=0
+ $Y2=0
cc_705 N_SCE_c_773_n N_A_453_47#_c_2301_n 0.00100011f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_706 N_SCE_c_775_n N_A_453_47#_c_2301_n 0.00229563f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_707 N_SCE_c_773_n N_A_453_47#_c_2302_n 0.00673545f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_708 N_SCE_c_775_n N_A_453_47#_c_2302_n 0.00729804f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_709 N_SCE_c_774_n N_VGND_c_2477_n 0.00409489f $X=3.25 $Y=0.735 $X2=0 $Y2=0
cc_710 N_SCE_c_772_n N_VGND_c_2495_n 0.00544863f $X=2.19 $Y=0.735 $X2=0 $Y2=0
cc_711 N_SCE_c_773_n N_VGND_c_2495_n 0.00397098f $X=3.175 $Y=0.81 $X2=0 $Y2=0
cc_712 N_SCE_c_774_n N_VGND_c_2495_n 0.0042361f $X=3.25 $Y=0.735 $X2=0 $Y2=0
cc_713 SCE N_VGND_c_2495_n 0.00725411f $X=1.975 $Y=0.425 $X2=0 $Y2=0
cc_714 N_SCE_c_772_n N_VGND_c_2505_n 0.00681989f $X=2.19 $Y=0.735 $X2=0 $Y2=0
cc_715 N_SCE_c_773_n N_VGND_c_2505_n 0.00278917f $X=3.175 $Y=0.81 $X2=0 $Y2=0
cc_716 N_SCE_c_774_n N_VGND_c_2505_n 0.00704136f $X=3.25 $Y=0.735 $X2=0 $Y2=0
cc_717 N_SCE_c_777_n N_VGND_c_2505_n 0.00343181f $X=2.25 $Y=0.93 $X2=0 $Y2=0
cc_718 SCE N_VGND_c_2505_n 0.00344584f $X=1.975 $Y=0.425 $X2=0 $Y2=0
cc_719 SCE A_381_47# 0.00111272f $X=1.975 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_720 N_D_M1024_g N_A_193_47#_c_912_n 0.0212393f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_721 N_D_M1019_g N_A_193_47#_c_924_n 0.00707191f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_722 D N_A_193_47#_c_924_n 0.0200936f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_723 N_D_c_874_n N_A_193_47#_c_924_n 9.34945e-19 $X=4.105 $Y=1.49 $X2=0 $Y2=0
cc_724 N_D_M1019_g N_VPWR_c_2073_n 0.00146693f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_725 D N_VPWR_c_2073_n 0.0112394f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_726 N_D_M1019_g N_VPWR_c_2088_n 0.00585385f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_727 D N_VPWR_c_2088_n 0.00771405f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_728 N_D_M1019_g N_VPWR_c_2070_n 0.00659811f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_729 D N_VPWR_c_2070_n 0.00345538f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_730 N_D_M1024_g N_A_453_47#_c_2300_n 0.00796014f $X=4.105 $Y=0.445 $X2=0
+ $Y2=0
cc_731 D N_A_453_47#_c_2300_n 0.00855055f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_732 N_D_c_874_n N_A_453_47#_c_2300_n 5.10457e-19 $X=4.105 $Y=1.49 $X2=0 $Y2=0
cc_733 N_D_M1024_g N_A_453_47#_c_2303_n 0.00192517f $X=4.105 $Y=0.445 $X2=0
+ $Y2=0
cc_734 N_D_M1024_g N_A_453_47#_c_2304_n 0.017252f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_735 D N_A_453_47#_c_2304_n 0.0480833f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_736 D A_752_413# 0.00729005f $X=3.825 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_737 N_D_M1024_g N_VGND_c_2477_n 0.00188039f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_738 N_D_M1024_g N_VGND_c_2487_n 0.00585385f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_739 N_D_M1024_g N_VGND_c_2505_n 0.00646586f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_740 N_A_193_47#_c_916_n N_A_1107_21#_M1038_g 5.35023e-19 $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_741 N_A_193_47#_c_926_n N_A_1107_21#_M1036_g 0.00197541f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_742 N_A_193_47#_M1032_g N_A_1107_21#_M1050_g 0.0164618f $X=8.505 $Y=2.275
+ $X2=0 $Y2=0
cc_743 N_A_193_47#_c_914_n N_A_1107_21#_M1050_g 0.00557961f $X=8.58 $Y=1.32
+ $X2=0 $Y2=0
cc_744 N_A_193_47#_c_926_n N_A_1107_21#_M1050_g 0.00750594f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_745 N_A_193_47#_c_931_n N_A_1107_21#_M1050_g 0.00910409f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_746 N_A_193_47#_c_932_n N_A_1107_21#_M1050_g 0.00264318f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_747 N_A_193_47#_c_926_n N_A_1107_21#_c_1136_n 0.0240118f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_748 N_A_193_47#_c_926_n N_A_1107_21#_c_1150_n 0.0279846f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_749 N_A_193_47#_c_926_n N_A_1107_21#_c_1138_n 0.0141612f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_750 N_A_193_47#_M1010_g N_A_1107_21#_c_1139_n 0.0161827f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_751 N_A_193_47#_c_926_n N_A_1107_21#_c_1139_n 0.00193898f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_752 N_A_193_47#_c_929_n N_A_1107_21#_c_1139_n 0.00927772f $X=5.04 $Y=1.74
+ $X2=0 $Y2=0
cc_753 N_A_193_47#_c_926_n N_A_1107_21#_c_1155_n 0.00959465f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_754 N_A_193_47#_c_914_n N_A_1107_21#_c_1132_n 0.00272432f $X=8.58 $Y=1.32
+ $X2=0 $Y2=0
cc_755 N_A_193_47#_M1003_g N_SET_B_c_1278_n 0.00574501f $X=9.04 $Y=0.415 $X2=0
+ $Y2=0
cc_756 N_A_193_47#_M1010_g N_A_931_47#_c_1414_n 0.0091014f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_757 N_A_193_47#_c_924_n N_A_931_47#_c_1414_n 2.09728e-19 $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_758 N_A_193_47#_c_926_n N_A_931_47#_c_1414_n 0.00506942f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_759 N_A_193_47#_c_927_n N_A_931_47#_c_1414_n 0.00303545f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_760 N_A_193_47#_c_929_n N_A_931_47#_c_1414_n 0.00186639f $X=5.04 $Y=1.74
+ $X2=0 $Y2=0
cc_761 N_A_193_47#_c_930_n N_A_931_47#_c_1414_n 0.0152514f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_762 N_A_193_47#_c_916_n N_A_931_47#_c_1415_n 0.00676006f $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_763 N_A_193_47#_c_917_n N_A_931_47#_c_1415_n 9.25786e-19 $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_764 N_A_193_47#_M1010_g N_A_931_47#_c_1409_n 0.00650943f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_765 N_A_193_47#_c_916_n N_A_931_47#_c_1409_n 0.00666284f $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_766 N_A_193_47#_c_926_n N_A_931_47#_c_1409_n 0.013911f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_767 N_A_193_47#_c_927_n N_A_931_47#_c_1409_n 0.00149623f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_768 N_A_193_47#_c_929_n N_A_931_47#_c_1409_n 0.00203066f $X=5.04 $Y=1.74
+ $X2=0 $Y2=0
cc_769 N_A_193_47#_c_930_n N_A_931_47#_c_1409_n 0.0282877f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_770 N_A_193_47#_c_926_n N_A_931_47#_c_1405_n 0.00350894f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_771 N_A_193_47#_c_916_n N_A_931_47#_c_1406_n 0.00728915f $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_772 N_A_193_47#_c_926_n N_A_931_47#_c_1406_n 0.00456576f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_773 N_A_193_47#_c_926_n N_A_1401_21#_M1031_g 0.00576309f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_774 N_A_193_47#_c_926_n N_A_1401_21#_c_1515_n 0.00477237f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_775 N_A_193_47#_c_913_n N_A_1401_21#_c_1524_n 0.00389341f $X=8.965 $Y=1.32
+ $X2=0 $Y2=0
cc_776 N_A_193_47#_c_926_n N_A_1401_21#_c_1524_n 0.0139809f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_777 N_A_193_47#_c_928_n N_A_1401_21#_c_1524_n 0.0255925f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_778 N_A_193_47#_c_931_n N_A_1401_21#_c_1524_n 0.00176885f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_779 N_A_193_47#_c_932_n N_A_1401_21#_c_1524_n 0.00661378f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_780 N_A_193_47#_c_933_n N_A_1401_21#_c_1524_n 0.00371524f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_781 N_A_193_47#_c_926_n N_A_1401_21#_c_1525_n 0.0264578f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_782 N_A_193_47#_c_931_n N_A_1401_21#_c_1525_n 7.96394e-19 $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_783 N_A_193_47#_c_932_n N_A_1401_21#_c_1525_n 0.00130051f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_784 N_A_193_47#_c_933_n N_A_1401_21#_c_1525_n 7.27878e-19 $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_785 N_A_193_47#_c_926_n N_A_1401_21#_c_1526_n 0.020032f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_786 N_A_193_47#_c_931_n N_A_1401_21#_c_1526_n 6.45403e-19 $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_787 N_A_193_47#_c_932_n N_A_1401_21#_c_1526_n 0.00461622f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_788 N_A_193_47#_c_933_n N_A_1401_21#_c_1526_n 0.00148716f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_789 N_A_193_47#_M1003_g N_A_1888_21#_M1042_g 0.0428045f $X=9.04 $Y=0.415
+ $X2=0 $Y2=0
cc_790 N_A_193_47#_M1032_g N_A_1714_47#_c_1872_n 0.00496872f $X=8.505 $Y=2.275
+ $X2=0 $Y2=0
cc_791 N_A_193_47#_c_928_n N_A_1714_47#_c_1872_n 0.00187313f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_792 N_A_193_47#_c_932_n N_A_1714_47#_c_1872_n 0.00141396f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_793 N_A_193_47#_M1003_g N_A_1714_47#_c_1875_n 0.0096406f $X=9.04 $Y=0.415
+ $X2=0 $Y2=0
cc_794 N_A_193_47#_M1003_g N_A_1714_47#_c_1861_n 0.010696f $X=9.04 $Y=0.415
+ $X2=0 $Y2=0
cc_795 N_A_193_47#_c_928_n N_A_1714_47#_c_1867_n 0.00214622f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_796 N_A_193_47#_c_932_n N_A_1714_47#_c_1867_n 0.0013353f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_797 N_A_193_47#_M1003_g N_A_1714_47#_c_1863_n 0.00156831f $X=9.04 $Y=0.415
+ $X2=0 $Y2=0
cc_798 N_A_193_47#_c_926_n N_VPWR_M1031_d 0.00670518f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_799 N_A_193_47#_c_918_n N_VPWR_c_2071_n 0.0127345f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_800 N_A_193_47#_c_924_n N_VPWR_c_2072_n 0.0169174f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_801 N_A_193_47#_c_925_n N_VPWR_c_2072_n 0.00138261f $X=1.295 $Y=1.87 $X2=0
+ $Y2=0
cc_802 N_A_193_47#_c_918_n N_VPWR_c_2072_n 0.0415488f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_803 N_A_193_47#_c_924_n N_VPWR_c_2073_n 0.00429349f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_804 N_A_193_47#_c_926_n N_VPWR_c_2074_n 0.00160449f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_805 N_A_193_47#_c_926_n N_VPWR_c_2075_n 0.0137399f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_806 N_A_193_47#_c_918_n N_VPWR_c_2086_n 0.0156296f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_807 N_A_193_47#_M1010_g N_VPWR_c_2088_n 0.00367119f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_808 N_A_193_47#_M1032_g N_VPWR_c_2089_n 0.00424681f $X=8.505 $Y=2.275 $X2=0
+ $Y2=0
cc_809 N_A_193_47#_c_932_n N_VPWR_c_2089_n 0.00254851f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_810 N_A_193_47#_M1010_g N_VPWR_c_2070_n 0.00562272f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_811 N_A_193_47#_M1032_g N_VPWR_c_2070_n 0.0061745f $X=8.505 $Y=2.275 $X2=0
+ $Y2=0
cc_812 N_A_193_47#_c_924_n N_VPWR_c_2070_n 0.16272f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_813 N_A_193_47#_c_925_n N_VPWR_c_2070_n 0.0151864f $X=1.295 $Y=1.87 $X2=0
+ $Y2=0
cc_814 N_A_193_47#_c_926_n N_VPWR_c_2070_n 0.159156f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_815 N_A_193_47#_c_927_n N_VPWR_c_2070_n 0.0160117f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_816 N_A_193_47#_c_928_n N_VPWR_c_2070_n 0.0148451f $X=8.51 $Y=1.87 $X2=0
+ $Y2=0
cc_817 N_A_193_47#_c_930_n N_VPWR_c_2070_n 3.19863e-19 $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_818 N_A_193_47#_c_931_n N_VPWR_c_2070_n 3.05853e-19 $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_819 N_A_193_47#_c_932_n N_VPWR_c_2070_n 0.00131252f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_820 N_A_193_47#_c_918_n N_VPWR_c_2070_n 0.00381175f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_821 N_A_193_47#_c_924_n A_381_363# 0.00298073f $X=4.685 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_822 N_A_193_47#_c_924_n N_A_453_47#_c_2297_n 0.00643756f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_823 N_A_193_47#_c_924_n N_A_453_47#_c_2306_n 0.0180928f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_824 N_A_193_47#_c_924_n N_A_453_47#_c_2307_n 0.00876668f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_825 N_A_193_47#_c_924_n N_A_453_47#_c_2300_n 0.0497172f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_826 N_A_193_47#_c_924_n N_A_453_47#_c_2301_n 0.0128789f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_827 N_A_193_47#_c_924_n N_A_453_47#_c_2302_n 0.00173167f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_828 N_A_193_47#_c_916_n N_A_453_47#_c_2303_n 0.00749938f $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_829 N_A_193_47#_c_917_n N_A_453_47#_c_2303_n 2.04896e-19 $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_830 N_A_193_47#_c_924_n N_A_453_47#_c_2303_n 0.0130335f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_831 N_A_193_47#_c_912_n N_A_453_47#_c_2304_n 0.00475032f $X=4.58 $Y=0.705
+ $X2=0 $Y2=0
cc_832 N_A_193_47#_c_916_n N_A_453_47#_c_2304_n 0.0620374f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_833 N_A_193_47#_c_924_n N_A_453_47#_c_2304_n 0.0188924f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_834 N_A_193_47#_c_927_n N_A_453_47#_c_2304_n 0.00185048f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_835 N_A_193_47#_c_930_n N_A_453_47#_c_2304_n 0.0281945f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_836 N_A_193_47#_c_926_n A_1351_329# 0.00110713f $X=8.365 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_837 N_A_193_47#_c_926_n A_1572_329# 0.00532504f $X=8.365 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_838 N_A_193_47#_c_918_n N_VGND_c_2476_n 0.0209768f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_839 N_A_193_47#_M1003_g N_VGND_c_2480_n 0.00126137f $X=9.04 $Y=0.415 $X2=0
+ $Y2=0
cc_840 N_A_193_47#_c_912_n N_VGND_c_2487_n 0.00556304f $X=4.58 $Y=0.705 $X2=0
+ $Y2=0
cc_841 N_A_193_47#_c_916_n N_VGND_c_2487_n 0.00113905f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_842 N_A_193_47#_c_917_n N_VGND_c_2487_n 2.48118e-19 $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_843 N_A_193_47#_M1003_g N_VGND_c_2491_n 0.00359964f $X=9.04 $Y=0.415 $X2=0
+ $Y2=0
cc_844 N_A_193_47#_c_918_n N_VGND_c_2494_n 0.00955835f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_845 N_A_193_47#_M1028_d N_VGND_c_2505_n 0.00217251f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_846 N_A_193_47#_c_912_n N_VGND_c_2505_n 0.00678262f $X=4.58 $Y=0.705 $X2=0
+ $Y2=0
cc_847 N_A_193_47#_M1003_g N_VGND_c_2505_n 0.00564067f $X=9.04 $Y=0.415 $X2=0
+ $Y2=0
cc_848 N_A_193_47#_c_916_n N_VGND_c_2505_n 0.00122477f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_849 N_A_193_47#_c_918_n N_VGND_c_2505_n 0.0038044f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_850 N_A_1107_21#_M1038_g N_SET_B_c_1272_n 0.0189927f $X=5.61 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_851 N_A_1107_21#_M1038_g N_SET_B_M1011_g 0.0137896f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_852 N_A_1107_21#_M1036_g N_SET_B_M1011_g 0.0101628f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_853 N_A_1107_21#_c_1136_n N_SET_B_M1011_g 0.0159332f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_854 N_A_1107_21#_c_1185_p N_SET_B_M1011_g 0.00507112f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_855 N_A_1107_21#_c_1138_n N_SET_B_M1011_g 0.00473578f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_856 N_A_1107_21#_c_1139_n N_SET_B_M1011_g 0.020182f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_857 N_A_1107_21#_M1038_g N_SET_B_M1047_g 0.0145491f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_858 N_A_1107_21#_c_1128_n N_SET_B_M1047_g 6.59324e-19 $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_859 N_A_1107_21#_M1038_g SET_B 0.00110276f $X=5.61 $Y=0.445 $X2=0 $Y2=0
cc_860 N_A_1107_21#_c_1128_n SET_B 0.00825406f $X=6.9 $Y=1.065 $X2=0 $Y2=0
cc_861 N_A_1107_21#_M1016_d N_SET_B_c_1278_n 5.1491e-19 $X=6.735 $Y=0.235 $X2=0
+ $Y2=0
cc_862 N_A_1107_21#_c_1127_n N_SET_B_c_1278_n 0.00507207f $X=8.02 $Y=0.985 $X2=0
+ $Y2=0
cc_863 N_A_1107_21#_c_1128_n N_SET_B_c_1278_n 0.0208059f $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_864 N_A_1107_21#_c_1130_n N_SET_B_c_1278_n 0.0214137f $X=7.795 $Y=0.98 $X2=0
+ $Y2=0
cc_865 N_A_1107_21#_c_1131_n N_SET_B_c_1278_n 0.0108883f $X=7.96 $Y=0.98 $X2=0
+ $Y2=0
cc_866 N_A_1107_21#_c_1128_n N_SET_B_c_1279_n 0.00230334f $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_867 N_A_1107_21#_c_1128_n N_A_931_47#_M1016_g 0.00718524f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_868 N_A_1107_21#_c_1129_n N_A_931_47#_M1016_g 0.0019289f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_869 N_A_1107_21#_c_1150_n N_A_931_47#_M1037_g 0.0126303f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_870 N_A_1107_21#_M1036_g N_A_931_47#_c_1414_n 0.00191115f $X=5.61 $Y=2.275
+ $X2=0 $Y2=0
cc_871 N_A_1107_21#_M1038_g N_A_931_47#_c_1415_n 0.00854236f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_872 N_A_1107_21#_M1038_g N_A_931_47#_c_1409_n 0.0154362f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_873 N_A_1107_21#_c_1138_n N_A_931_47#_c_1409_n 0.0330453f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_874 N_A_1107_21#_M1038_g N_A_931_47#_c_1404_n 0.0188177f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_875 N_A_1107_21#_c_1136_n N_A_931_47#_c_1405_n 0.0141289f $X=6.385 $Y=1.91
+ $X2=0 $Y2=0
cc_876 N_A_1107_21#_c_1150_n N_A_931_47#_c_1405_n 0.00218253f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_877 N_A_1107_21#_c_1129_n N_A_931_47#_c_1405_n 0.0246731f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_878 N_A_1107_21#_c_1155_n N_A_931_47#_c_1405_n 0.00650509f $X=6.47 $Y=1.87
+ $X2=0 $Y2=0
cc_879 N_A_1107_21#_M1038_g N_A_931_47#_c_1406_n 0.0109165f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_880 N_A_1107_21#_c_1138_n N_A_931_47#_c_1406_n 0.0169843f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_881 N_A_1107_21#_c_1139_n N_A_931_47#_c_1406_n 0.0011995f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_882 N_A_1107_21#_c_1129_n N_A_931_47#_c_1407_n 0.00939619f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_883 N_A_1107_21#_c_1155_n N_A_931_47#_c_1407_n 9.09922e-19 $X=6.47 $Y=1.87
+ $X2=0 $Y2=0
cc_884 N_A_1107_21#_c_1128_n N_A_1401_21#_c_1509_n 0.00781955f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_885 N_A_1107_21#_c_1130_n N_A_1401_21#_c_1509_n 0.00387342f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_886 N_A_1107_21#_c_1128_n N_A_1401_21#_c_1510_n 0.001691f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_887 N_A_1107_21#_c_1129_n N_A_1401_21#_c_1510_n 0.00751117f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_888 N_A_1107_21#_c_1130_n N_A_1401_21#_c_1510_n 0.0116453f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_889 N_A_1107_21#_c_1131_n N_A_1401_21#_c_1510_n 0.00205413f $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_890 N_A_1107_21#_c_1132_n N_A_1401_21#_c_1510_n 0.0187801f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_891 N_A_1107_21#_M1050_g N_A_1401_21#_M1031_g 0.0153539f $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_892 N_A_1107_21#_c_1150_n N_A_1401_21#_M1031_g 0.00219889f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_893 N_A_1107_21#_M1050_g N_A_1401_21#_c_1515_n 2.86505e-19 $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_894 N_A_1107_21#_c_1129_n N_A_1401_21#_c_1515_n 0.0309286f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_895 N_A_1107_21#_c_1130_n N_A_1401_21#_c_1515_n 0.0205152f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_896 N_A_1107_21#_c_1132_n N_A_1401_21#_c_1515_n 0.00382982f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_897 N_A_1107_21#_c_1131_n N_A_1401_21#_c_1525_n 9.59092e-19 $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_898 N_A_1107_21#_c_1132_n N_A_1401_21#_c_1525_n 0.00358318f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_899 N_A_1107_21#_M1050_g N_A_1401_21#_c_1526_n 0.0143059f $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_900 N_A_1107_21#_c_1130_n N_A_1401_21#_c_1526_n 0.00760725f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_901 N_A_1107_21#_c_1131_n N_A_1401_21#_c_1526_n 0.0207118f $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_902 N_A_1107_21#_c_1132_n N_A_1401_21#_c_1526_n 0.00632961f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_903 N_A_1107_21#_M1050_g N_A_1714_47#_c_1872_n 7.04843e-19 $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_904 N_A_1107_21#_M1036_g N_VPWR_c_2074_n 0.00326498f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_905 N_A_1107_21#_c_1136_n N_VPWR_c_2074_n 0.0124698f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_906 N_A_1107_21#_c_1185_p N_VPWR_c_2074_n 0.00820313f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_907 N_A_1107_21#_c_1138_n N_VPWR_c_2074_n 0.0125544f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_908 N_A_1107_21#_c_1139_n N_VPWR_c_2074_n 7.62241e-19 $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_909 N_A_1107_21#_M1050_g N_VPWR_c_2075_n 0.0163458f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_910 N_A_1107_21#_c_1150_n N_VPWR_c_2075_n 0.0048929f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_911 N_A_1107_21#_c_1136_n N_VPWR_c_2081_n 0.00474052f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_912 N_A_1107_21#_c_1185_p N_VPWR_c_2081_n 0.00725778f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_913 N_A_1107_21#_c_1150_n N_VPWR_c_2081_n 0.00598455f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_914 N_A_1107_21#_M1036_g N_VPWR_c_2088_n 0.00535335f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_915 N_A_1107_21#_c_1138_n N_VPWR_c_2088_n 0.00111392f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_916 N_A_1107_21#_M1050_g N_VPWR_c_2089_n 0.00585385f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_917 N_A_1107_21#_M1011_d N_VPWR_c_2070_n 0.0031612f $X=6.215 $Y=2.065 $X2=0
+ $Y2=0
cc_918 N_A_1107_21#_M1036_g N_VPWR_c_2070_n 0.00664368f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_919 N_A_1107_21#_M1050_g N_VPWR_c_2070_n 0.00762825f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_920 N_A_1107_21#_c_1136_n N_VPWR_c_2070_n 0.00386836f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_921 N_A_1107_21#_c_1185_p N_VPWR_c_2070_n 0.0029026f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_922 N_A_1107_21#_c_1150_n N_VPWR_c_2070_n 0.00505387f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_923 N_A_1107_21#_c_1138_n N_VPWR_c_2070_n 0.00128163f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_924 N_A_1107_21#_c_1150_n A_1351_329# 0.00339576f $X=6.815 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_925 N_A_1107_21#_c_1129_n A_1351_329# 0.00178287f $X=6.9 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_926 N_A_1107_21#_M1038_g N_VGND_c_2478_n 0.00361232f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_927 N_A_1107_21#_c_1127_n N_VGND_c_2479_n 0.0111314f $X=8.02 $Y=0.985 $X2=0
+ $Y2=0
cc_928 N_A_1107_21#_c_1130_n N_VGND_c_2479_n 0.00387395f $X=7.795 $Y=0.98 $X2=0
+ $Y2=0
cc_929 N_A_1107_21#_c_1131_n N_VGND_c_2479_n 0.00379129f $X=7.96 $Y=0.98 $X2=0
+ $Y2=0
cc_930 N_A_1107_21#_c_1132_n N_VGND_c_2479_n 8.52393e-19 $X=7.96 $Y=1.15 $X2=0
+ $Y2=0
cc_931 N_A_1107_21#_M1038_g N_VGND_c_2487_n 0.0035977f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_932 N_A_1107_21#_c_1127_n N_VGND_c_2491_n 0.0046653f $X=8.02 $Y=0.985 $X2=0
+ $Y2=0
cc_933 N_A_1107_21#_M1016_d N_VGND_c_2505_n 0.00178362f $X=6.735 $Y=0.235 $X2=0
+ $Y2=0
cc_934 N_A_1107_21#_M1038_g N_VGND_c_2505_n 0.00580574f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_935 N_A_1107_21#_c_1127_n N_VGND_c_2505_n 0.00460207f $X=8.02 $Y=0.985 $X2=0
+ $Y2=0
cc_936 N_A_1107_21#_M1016_d N_A_1251_47#_c_2713_n 0.0030477f $X=6.735 $Y=0.235
+ $X2=0 $Y2=0
cc_937 N_A_1107_21#_c_1128_n N_A_1251_47#_c_2713_n 0.0147704f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_938 N_A_1107_21#_c_1130_n N_A_1251_47#_c_2713_n 0.00259503f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_939 N_A_1107_21#_c_1127_n N_A_1251_47#_c_2716_n 0.00441801f $X=8.02 $Y=0.985
+ $X2=0 $Y2=0
cc_940 N_A_1107_21#_c_1130_n N_A_1251_47#_c_2716_n 0.0106429f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_941 N_SET_B_c_1272_n N_A_931_47#_M1016_g 0.00619508f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_942 N_SET_B_M1047_g N_A_931_47#_M1016_g 0.018553f $X=6.18 $Y=0.445 $X2=0
+ $Y2=0
cc_943 SET_B N_A_931_47#_M1016_g 0.00183601f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_944 N_SET_B_c_1278_n N_A_931_47#_M1016_g 0.00491921f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_945 N_SET_B_c_1279_n N_A_931_47#_M1016_g 0.00134231f $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_946 N_SET_B_M1011_g N_A_931_47#_M1037_g 0.0228864f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_947 N_SET_B_c_1272_n N_A_931_47#_c_1404_n 0.00216489f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_948 N_SET_B_M1011_g N_A_931_47#_c_1404_n 6.04572e-19 $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_949 N_SET_B_M1047_g N_A_931_47#_c_1404_n 0.00182721f $X=6.18 $Y=0.445 $X2=0
+ $Y2=0
cc_950 SET_B N_A_931_47#_c_1404_n 0.0244028f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_951 N_SET_B_c_1279_n N_A_931_47#_c_1404_n 0.00111115f $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_952 N_SET_B_c_1272_n N_A_931_47#_c_1405_n 0.00310411f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_953 N_SET_B_M1011_g N_A_931_47#_c_1405_n 0.0131452f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_954 SET_B N_A_931_47#_c_1405_n 0.0245807f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_955 N_SET_B_c_1278_n N_A_931_47#_c_1405_n 0.00270886f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_956 N_SET_B_c_1279_n N_A_931_47#_c_1405_n 6.67689e-19 $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_957 N_SET_B_M1011_g N_A_931_47#_c_1406_n 5.20457e-19 $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_958 N_SET_B_M1011_g N_A_931_47#_c_1407_n 0.021088f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_959 N_SET_B_c_1278_n N_A_1401_21#_c_1509_n 0.00317213f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_960 N_SET_B_c_1278_n N_A_1401_21#_c_1515_n 5.29205e-19 $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_961 N_SET_B_M1007_g N_A_1401_21#_c_1524_n 0.00583258f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_962 N_SET_B_c_1278_n N_A_1401_21#_c_1524_n 0.0486538f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_963 N_SET_B_c_1280_n N_A_1401_21#_c_1524_n 0.0135087f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_964 N_SET_B_M1004_g N_A_1888_21#_M1042_g 0.0180201f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_965 N_SET_B_M1007_g N_A_1888_21#_M1042_g 0.0136409f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_966 N_SET_B_c_1278_n N_A_1888_21#_M1042_g 0.00627116f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_967 N_SET_B_c_1280_n N_A_1888_21#_M1042_g 0.00136404f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_968 N_SET_B_c_1281_n N_A_1888_21#_M1042_g 0.00227945f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_969 N_SET_B_c_1282_n N_A_1888_21#_M1042_g 0.020875f $X=9.935 $Y=0.98 $X2=0
+ $Y2=0
cc_970 N_SET_B_M1007_g N_A_1888_21#_M1043_g 0.0109753f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_971 N_SET_B_M1007_g N_A_1888_21#_c_1686_n 0.00710111f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_972 N_SET_B_M1007_g N_A_1888_21#_c_1687_n 0.019738f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_973 N_SET_B_M1007_g N_A_1888_21#_c_1688_n 0.0136222f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_974 N_SET_B_c_1281_n N_A_1888_21#_c_1676_n 0.00828511f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_975 N_SET_B_M1004_g N_A_1888_21#_c_1707_n 6.74813e-19 $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_976 N_SET_B_c_1280_n N_A_1888_21#_c_1707_n 2.37563e-19 $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_977 N_SET_B_c_1281_n N_A_1888_21#_c_1707_n 0.00144717f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_978 N_SET_B_M1004_g N_A_1714_47#_M1001_g 0.0175593f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_979 N_SET_B_c_1281_n N_A_1714_47#_M1001_g 0.00170408f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_980 N_SET_B_c_1282_n N_A_1714_47#_M1001_g 0.009306f $X=9.935 $Y=0.98 $X2=0
+ $Y2=0
cc_981 N_SET_B_M1007_g N_A_1714_47#_M1025_g 0.0325064f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_982 N_SET_B_c_1278_n N_A_1714_47#_c_1875_n 0.00883541f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_983 N_SET_B_c_1278_n N_A_1714_47#_c_1861_n 0.017797f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_984 N_SET_B_c_1280_n N_A_1714_47#_c_1861_n 0.0022902f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_985 N_SET_B_c_1281_n N_A_1714_47#_c_1861_n 0.0118231f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_986 N_SET_B_M1007_g N_A_1714_47#_c_1862_n 0.0117331f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_987 N_SET_B_c_1278_n N_A_1714_47#_c_1862_n 0.00876649f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_988 N_SET_B_c_1280_n N_A_1714_47#_c_1862_n 0.00124273f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_989 N_SET_B_c_1281_n N_A_1714_47#_c_1862_n 0.0248283f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_990 N_SET_B_c_1282_n N_A_1714_47#_c_1862_n 0.00490678f $X=9.935 $Y=0.98 $X2=0
+ $Y2=0
cc_991 N_SET_B_c_1282_n N_A_1714_47#_c_1864_n 0.00111089f $X=9.935 $Y=0.98 $X2=0
+ $Y2=0
cc_992 N_SET_B_c_1282_n N_A_1714_47#_c_1865_n 0.0212822f $X=9.935 $Y=0.98 $X2=0
+ $Y2=0
cc_993 N_SET_B_M1011_g N_VPWR_c_2074_n 0.0094739f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_994 N_SET_B_M1011_g N_VPWR_c_2081_n 0.00373914f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_995 N_SET_B_M1007_g N_VPWR_c_2084_n 0.00368415f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_996 N_SET_B_M1007_g N_VPWR_c_2097_n 0.00857728f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_997 N_SET_B_M1011_g N_VPWR_c_2070_n 0.00439789f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_998 N_SET_B_M1007_g N_VPWR_c_2070_n 0.00444663f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_999 N_SET_B_c_1278_n N_VGND_M1041_s 0.00213341f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_1000 N_SET_B_c_1272_n N_VGND_c_2478_n 8.58768e-19 $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_1001 N_SET_B_M1047_g N_VGND_c_2478_n 0.00289978f $X=6.18 $Y=0.445 $X2=0 $Y2=0
cc_1002 SET_B N_VGND_c_2478_n 0.010979f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1003 N_SET_B_c_1278_n N_VGND_c_2479_n 0.00404506f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1004 N_SET_B_M1004_g N_VGND_c_2480_n 0.00282278f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1005 N_SET_B_c_1278_n N_VGND_c_2480_n 0.00604269f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1006 N_SET_B_c_1280_n N_VGND_c_2480_n 7.41662e-19 $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1007 N_SET_B_c_1281_n N_VGND_c_2480_n 0.00350326f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1008 N_SET_B_M1047_g N_VGND_c_2489_n 0.00422832f $X=6.18 $Y=0.445 $X2=0 $Y2=0
cc_1009 SET_B N_VGND_c_2489_n 0.00221313f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1010 N_SET_B_M1004_g N_VGND_c_2496_n 0.00439071f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1011 N_SET_B_c_1281_n N_VGND_c_2496_n 0.00352663f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1012 N_SET_B_M1047_g N_VGND_c_2505_n 0.00587817f $X=6.18 $Y=0.445 $X2=0 $Y2=0
cc_1013 N_SET_B_M1004_g N_VGND_c_2505_n 0.00595177f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1014 SET_B N_VGND_c_2505_n 0.00214053f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1015 N_SET_B_c_1278_n N_VGND_c_2505_n 0.165421f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_1016 N_SET_B_c_1279_n N_VGND_c_2505_n 0.0147353f $X=6.355 $Y=0.85 $X2=0 $Y2=0
cc_1017 N_SET_B_c_1280_n N_VGND_c_2505_n 0.0141642f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1018 N_SET_B_c_1281_n N_VGND_c_2505_n 0.00284893f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1019 N_SET_B_c_1278_n N_A_1251_47#_M1047_d 0.00182666f $X=9.745 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1020 N_SET_B_c_1279_n N_A_1251_47#_M1047_d 6.40013e-19 $X=6.355 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1021 N_SET_B_c_1278_n N_A_1251_47#_M1014_d 0.00215149f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1022 N_SET_B_c_1278_n N_A_1251_47#_c_2713_n 0.00555941f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1023 N_SET_B_c_1278_n N_A_1251_47#_c_2716_n 0.00234876f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1024 N_SET_B_M1047_g N_A_1251_47#_c_2723_n 0.00335852f $X=6.18 $Y=0.445 $X2=0
+ $Y2=0
cc_1025 SET_B N_A_1251_47#_c_2723_n 0.00237046f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1026 N_SET_B_c_1278_n N_A_1251_47#_c_2723_n 0.00393563f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1027 N_SET_B_c_1279_n N_A_1251_47#_c_2723_n 0.00215379f $X=6.355 $Y=0.85
+ $X2=0 $Y2=0
cc_1028 N_SET_B_c_1278_n A_1619_47# 0.00369541f $X=9.745 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_1029 N_SET_B_M1004_g N_A_2004_47#_c_2744_n 0.00349862f $X=9.945 $Y=0.445
+ $X2=0 $Y2=0
cc_1030 N_SET_B_c_1281_n N_A_2004_47#_c_2744_n 0.00344477f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1031 N_SET_B_c_1282_n N_A_2004_47#_c_2744_n 2.8008e-19 $X=9.935 $Y=0.98 $X2=0
+ $Y2=0
cc_1032 N_A_931_47#_M1016_g N_A_1401_21#_c_1509_n 0.0281038f $X=6.66 $Y=0.555
+ $X2=0 $Y2=0
cc_1033 N_A_931_47#_M1016_g N_A_1401_21#_c_1510_n 0.00233575f $X=6.66 $Y=0.555
+ $X2=0 $Y2=0
cc_1034 N_A_931_47#_c_1407_n N_A_1401_21#_c_1510_n 0.0322452f $X=6.56 $Y=1.32
+ $X2=0 $Y2=0
cc_1035 N_A_931_47#_M1037_g N_A_1401_21#_M1031_g 0.0322452f $X=6.68 $Y=2.065
+ $X2=0 $Y2=0
cc_1036 N_A_931_47#_M1037_g N_VPWR_c_2074_n 0.00136797f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1037 N_A_931_47#_M1037_g N_VPWR_c_2081_n 0.00432313f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1038 N_A_931_47#_c_1414_n N_VPWR_c_2088_n 0.0377433f $X=5.295 $Y=2.335 $X2=0
+ $Y2=0
cc_1039 N_A_931_47#_M1040_d N_VPWR_c_2070_n 0.00173085f $X=4.665 $Y=2.065 $X2=0
+ $Y2=0
cc_1040 N_A_931_47#_M1037_g N_VPWR_c_2070_n 0.00600471f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1041 N_A_931_47#_c_1414_n N_VPWR_c_2070_n 0.0132511f $X=5.295 $Y=2.335 $X2=0
+ $Y2=0
cc_1042 N_A_931_47#_c_1414_n N_A_453_47#_c_2304_n 0.0128808f $X=5.295 $Y=2.335
+ $X2=0 $Y2=0
cc_1043 N_A_931_47#_c_1414_n A_1017_413# 0.00858887f $X=5.295 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1044 N_A_931_47#_c_1409_n A_1017_413# 0.00579571f $X=5.38 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1045 N_A_931_47#_c_1415_n N_VGND_c_2487_n 0.055608f $X=5.545 $Y=0.365 $X2=0
+ $Y2=0
cc_1046 N_A_931_47#_M1016_g N_VGND_c_2489_n 0.00357877f $X=6.66 $Y=0.555 $X2=0
+ $Y2=0
cc_1047 N_A_931_47#_M1045_d N_VGND_c_2505_n 0.00275359f $X=4.655 $Y=0.235 $X2=0
+ $Y2=0
cc_1048 N_A_931_47#_M1016_g N_VGND_c_2505_n 0.00536866f $X=6.66 $Y=0.555 $X2=0
+ $Y2=0
cc_1049 N_A_931_47#_c_1415_n N_VGND_c_2505_n 0.0218827f $X=5.545 $Y=0.365 $X2=0
+ $Y2=0
cc_1050 N_A_931_47#_c_1415_n A_1041_47# 0.00568226f $X=5.545 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1051 N_A_931_47#_M1016_g N_A_1251_47#_c_2713_n 0.00821062f $X=6.66 $Y=0.555
+ $X2=0 $Y2=0
cc_1052 N_A_931_47#_c_1405_n N_A_1251_47#_c_2723_n 0.00116076f $X=6.395 $Y=1.32
+ $X2=0 $Y2=0
cc_1053 N_A_931_47#_c_1407_n N_A_1251_47#_c_2723_n 5.81529e-19 $X=6.56 $Y=1.32
+ $X2=0 $Y2=0
cc_1054 N_A_1401_21#_c_1524_n N_A_1888_21#_M1042_g 0.00413345f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1055 N_A_1401_21#_c_1524_n N_A_1888_21#_c_1686_n 0.015309f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1056 N_A_1401_21#_c_1524_n N_A_1888_21#_c_1687_n 0.00677286f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1057 N_A_1401_21#_c_1524_n N_A_1888_21#_c_1688_n 0.010417f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1058 N_A_1401_21#_c_1524_n N_A_1888_21#_c_1714_n 0.00964432f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1059 N_A_1401_21#_M1029_g N_A_1888_21#_c_1676_n 0.0128951f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1060 N_A_1401_21#_M1017_g N_A_1888_21#_c_1676_n 0.0062981f $X=10.955 $Y=0.555
+ $X2=0 $Y2=0
cc_1061 N_A_1401_21#_c_1513_n N_A_1888_21#_c_1676_n 0.00726543f $X=11.355
+ $Y=0.84 $X2=0 $Y2=0
cc_1062 N_A_1401_21#_c_1521_n N_A_1888_21#_c_1676_n 0.0130479f $X=11.355 $Y=1.66
+ $X2=0 $Y2=0
cc_1063 N_A_1401_21#_c_1524_n N_A_1888_21#_c_1676_n 0.0270698f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1064 N_A_1401_21#_c_1527_n N_A_1888_21#_c_1676_n 5.62937e-19 $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1065 N_A_1401_21#_c_1516_n N_A_1888_21#_c_1676_n 0.00937037f $X=10.955
+ $Y=1.32 $X2=0 $Y2=0
cc_1066 N_A_1401_21#_c_1517_n N_A_1888_21#_c_1676_n 0.046128f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1067 N_A_1401_21#_M1030_s N_A_1888_21#_c_1690_n 0.00478726f $X=11.635
+ $Y=1.505 $X2=0 $Y2=0
cc_1068 N_A_1401_21#_M1029_g N_A_1888_21#_c_1690_n 0.00712539f $X=10.895
+ $Y=2.065 $X2=0 $Y2=0
cc_1069 N_A_1401_21#_c_1521_n N_A_1888_21#_c_1690_n 0.0212381f $X=11.355 $Y=1.66
+ $X2=0 $Y2=0
cc_1070 N_A_1401_21#_c_1522_n N_A_1888_21#_c_1690_n 0.0374534f $X=11.76 $Y=1.66
+ $X2=0 $Y2=0
cc_1071 N_A_1401_21#_c_1524_n N_A_1888_21#_c_1690_n 0.00648571f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1072 N_A_1401_21#_c_1527_n N_A_1888_21#_c_1690_n 0.00170504f $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1073 N_A_1401_21#_c_1516_n N_A_1888_21#_c_1690_n 0.0026574f $X=10.955 $Y=1.32
+ $X2=0 $Y2=0
cc_1074 N_A_1401_21#_c_1522_n N_A_1888_21#_c_1691_n 0.00819527f $X=11.76 $Y=1.66
+ $X2=0 $Y2=0
cc_1075 N_A_1401_21#_c_1524_n N_A_1888_21#_c_1731_n 0.00453864f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1076 N_A_1401_21#_M1017_g N_A_1888_21#_c_1707_n 0.0077182f $X=10.955 $Y=0.555
+ $X2=0 $Y2=0
cc_1077 N_A_1401_21#_M1029_g N_A_1888_21#_c_1733_n 0.00499743f $X=10.895
+ $Y=2.065 $X2=0 $Y2=0
cc_1078 N_A_1401_21#_M1017_g N_A_1714_47#_M1001_g 0.0191895f $X=10.955 $Y=0.555
+ $X2=0 $Y2=0
cc_1079 N_A_1401_21#_M1029_g N_A_1714_47#_M1025_g 0.039703f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1080 N_A_1401_21#_c_1524_n N_A_1714_47#_M1025_g 0.00713863f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1081 N_A_1401_21#_c_1524_n N_A_1714_47#_c_1867_n 0.0219541f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1082 N_A_1401_21#_c_1524_n N_A_1714_47#_c_1862_n 0.0228947f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1083 N_A_1401_21#_M1017_g N_A_1714_47#_c_1864_n 2.36981e-19 $X=10.955
+ $Y=0.555 $X2=0 $Y2=0
cc_1084 N_A_1401_21#_c_1524_n N_A_1714_47#_c_1864_n 0.00714757f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1085 N_A_1401_21#_c_1516_n N_A_1714_47#_c_1865_n 0.0588925f $X=10.955 $Y=1.32
+ $X2=0 $Y2=0
cc_1086 N_A_1401_21#_c_1512_n N_RESET_B_M1009_g 0.00684899f $X=11.62 $Y=0.84
+ $X2=0 $Y2=0
cc_1087 N_A_1401_21#_c_1514_n N_RESET_B_M1009_g 0.00289722f $X=11.76 $Y=0.43
+ $X2=0 $Y2=0
cc_1088 N_A_1401_21#_c_1517_n N_RESET_B_M1009_g 0.00219324f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1089 N_A_1401_21#_c_1522_n N_RESET_B_M1030_g 0.00322142f $X=11.76 $Y=1.66
+ $X2=0 $Y2=0
cc_1090 N_A_1401_21#_c_1527_n N_RESET_B_M1030_g 0.00254006f $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1091 N_A_1401_21#_c_1516_n N_RESET_B_M1030_g 0.00200587f $X=10.955 $Y=1.32
+ $X2=0 $Y2=0
cc_1092 N_A_1401_21#_c_1517_n N_RESET_B_M1030_g 0.00281503f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1093 N_A_1401_21#_c_1512_n RESET_B 0.0207441f $X=11.62 $Y=0.84 $X2=0 $Y2=0
cc_1094 N_A_1401_21#_c_1522_n RESET_B 0.0164254f $X=11.76 $Y=1.66 $X2=0 $Y2=0
cc_1095 N_A_1401_21#_c_1516_n RESET_B 6.20263e-19 $X=10.955 $Y=1.32 $X2=0 $Y2=0
cc_1096 N_A_1401_21#_c_1517_n RESET_B 0.0154244f $X=11.165 $Y=1.32 $X2=0 $Y2=0
cc_1097 N_A_1401_21#_M1017_g N_RESET_B_c_1961_n 0.00175075f $X=10.955 $Y=0.555
+ $X2=0 $Y2=0
cc_1098 N_A_1401_21#_c_1512_n N_RESET_B_c_1961_n 0.00576136f $X=11.62 $Y=0.84
+ $X2=0 $Y2=0
cc_1099 N_A_1401_21#_c_1522_n N_RESET_B_c_1961_n 0.00581996f $X=11.76 $Y=1.66
+ $X2=0 $Y2=0
cc_1100 N_A_1401_21#_c_1516_n N_RESET_B_c_1961_n 0.0072561f $X=10.955 $Y=1.32
+ $X2=0 $Y2=0
cc_1101 N_A_1401_21#_c_1517_n N_RESET_B_c_1961_n 0.00323603f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1102 N_A_1401_21#_c_1515_n N_VPWR_M1031_d 0.00297048f $X=7.32 $Y=1.32 $X2=0
+ $Y2=0
cc_1103 N_A_1401_21#_c_1526_n N_VPWR_M1031_d 0.00221014f $X=8.05 $Y=1.53 $X2=0
+ $Y2=0
cc_1104 N_A_1401_21#_c_1521_n N_VPWR_M1029_d 0.00311394f $X=11.355 $Y=1.66 $X2=0
+ $Y2=0
cc_1105 N_A_1401_21#_c_1510_n N_VPWR_c_2075_n 0.00111411f $X=7.1 $Y=1.485 $X2=0
+ $Y2=0
cc_1106 N_A_1401_21#_M1031_g N_VPWR_c_2075_n 0.00353361f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1107 N_A_1401_21#_c_1515_n N_VPWR_c_2075_n 0.011531f $X=7.32 $Y=1.32 $X2=0
+ $Y2=0
cc_1108 N_A_1401_21#_c_1526_n N_VPWR_c_2075_n 7.83548e-19 $X=8.05 $Y=1.53 $X2=0
+ $Y2=0
cc_1109 N_A_1401_21#_M1031_g N_VPWR_c_2081_n 0.00583607f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1110 N_A_1401_21#_M1029_g N_VPWR_c_2083_n 0.0111257f $X=10.895 $Y=2.065 $X2=0
+ $Y2=0
cc_1111 N_A_1401_21#_M1029_g N_VPWR_c_2084_n 0.00339278f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1112 N_A_1401_21#_M1031_g N_VPWR_c_2070_n 0.00670824f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1113 N_A_1401_21#_M1029_g N_VPWR_c_2070_n 0.0038354f $X=10.895 $Y=2.065 $X2=0
+ $Y2=0
cc_1114 N_A_1401_21#_c_1526_n A_1572_329# 0.00272182f $X=8.05 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_1115 N_A_1401_21#_c_1509_n N_VGND_c_2479_n 0.00318127f $X=7.08 $Y=0.95 $X2=0
+ $Y2=0
cc_1116 N_A_1401_21#_c_1512_n N_VGND_c_2481_n 0.00351875f $X=11.62 $Y=0.84 $X2=0
+ $Y2=0
cc_1117 N_A_1401_21#_c_1514_n N_VGND_c_2481_n 0.00634982f $X=11.76 $Y=0.43 $X2=0
+ $Y2=0
cc_1118 N_A_1401_21#_c_1509_n N_VGND_c_2489_n 0.00357877f $X=7.08 $Y=0.95 $X2=0
+ $Y2=0
cc_1119 N_A_1401_21#_M1017_g N_VGND_c_2496_n 0.00357877f $X=10.955 $Y=0.555
+ $X2=0 $Y2=0
cc_1120 N_A_1401_21#_c_1512_n N_VGND_c_2496_n 0.00380144f $X=11.62 $Y=0.84 $X2=0
+ $Y2=0
cc_1121 N_A_1401_21#_c_1513_n N_VGND_c_2496_n 0.00166179f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1122 N_A_1401_21#_c_1514_n N_VGND_c_2496_n 0.0145278f $X=11.76 $Y=0.43 $X2=0
+ $Y2=0
cc_1123 N_A_1401_21#_M1009_s N_VGND_c_2505_n 0.00383158f $X=11.635 $Y=0.235
+ $X2=0 $Y2=0
cc_1124 N_A_1401_21#_c_1509_n N_VGND_c_2505_n 0.00661646f $X=7.08 $Y=0.95 $X2=0
+ $Y2=0
cc_1125 N_A_1401_21#_M1017_g N_VGND_c_2505_n 0.00657041f $X=10.955 $Y=0.555
+ $X2=0 $Y2=0
cc_1126 N_A_1401_21#_c_1512_n N_VGND_c_2505_n 0.00683133f $X=11.62 $Y=0.84 $X2=0
+ $Y2=0
cc_1127 N_A_1401_21#_c_1513_n N_VGND_c_2505_n 0.00329575f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1128 N_A_1401_21#_c_1514_n N_VGND_c_2505_n 0.00854056f $X=11.76 $Y=0.43 $X2=0
+ $Y2=0
cc_1129 N_A_1401_21#_c_1509_n N_A_1251_47#_c_2713_n 0.0105472f $X=7.08 $Y=0.95
+ $X2=0 $Y2=0
cc_1130 N_A_1401_21#_c_1513_n N_A_2004_47#_M1017_d 0.0043454f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1131 N_A_1401_21#_M1017_g N_A_2004_47#_c_2748_n 0.0112006f $X=10.955 $Y=0.555
+ $X2=0 $Y2=0
cc_1132 N_A_1401_21#_c_1513_n N_A_2004_47#_c_2749_n 0.0133877f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1133 N_A_1401_21#_c_1514_n N_A_2004_47#_c_2749_n 0.0139043f $X=11.76 $Y=0.43
+ $X2=0 $Y2=0
cc_1134 N_A_1401_21#_c_1516_n N_A_2004_47#_c_2749_n 5.38954e-19 $X=10.955
+ $Y=1.32 $X2=0 $Y2=0
cc_1135 N_A_1888_21#_c_1676_n N_A_1714_47#_M1001_g 0.0153921f $X=10.82 $Y=1.915
+ $X2=0 $Y2=0
cc_1136 N_A_1888_21#_c_1707_n N_A_1714_47#_M1001_g 0.00536261f $X=10.82 $Y=0.687
+ $X2=0 $Y2=0
cc_1137 N_A_1888_21#_c_1714_n N_A_1714_47#_M1025_g 0.0118664f $X=10.73 $Y=2
+ $X2=0 $Y2=0
cc_1138 N_A_1888_21#_M1043_g N_A_1714_47#_c_1872_n 0.00204127f $X=9.515 $Y=2.275
+ $X2=0 $Y2=0
cc_1139 N_A_1888_21#_M1042_g N_A_1714_47#_c_1875_n 0.0017558f $X=9.515 $Y=0.445
+ $X2=0 $Y2=0
cc_1140 N_A_1888_21#_M1042_g N_A_1714_47#_c_1861_n 0.0128435f $X=9.515 $Y=0.445
+ $X2=0 $Y2=0
cc_1141 N_A_1888_21#_M1042_g N_A_1714_47#_c_1867_n 0.0148682f $X=9.515 $Y=0.445
+ $X2=0 $Y2=0
cc_1142 N_A_1888_21#_c_1686_n N_A_1714_47#_c_1867_n 0.0248026f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1143 N_A_1888_21#_c_1742_p N_A_1714_47#_c_1867_n 0.0135579f $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1144 N_A_1888_21#_M1042_g N_A_1714_47#_c_1862_n 0.0115171f $X=9.515 $Y=0.445
+ $X2=0 $Y2=0
cc_1145 N_A_1888_21#_c_1686_n N_A_1714_47#_c_1862_n 0.0154844f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1146 N_A_1888_21#_c_1687_n N_A_1714_47#_c_1862_n 0.00126891f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1147 N_A_1888_21#_c_1688_n N_A_1714_47#_c_1862_n 0.00635717f $X=10.24 $Y=2
+ $X2=0 $Y2=0
cc_1148 N_A_1888_21#_c_1731_n N_A_1714_47#_c_1862_n 0.00162703f $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1149 N_A_1888_21#_c_1714_n N_A_1714_47#_c_1864_n 0.00158774f $X=10.73 $Y=2
+ $X2=0 $Y2=0
cc_1150 N_A_1888_21#_c_1676_n N_A_1714_47#_c_1864_n 0.0241621f $X=10.82 $Y=1.915
+ $X2=0 $Y2=0
cc_1151 N_A_1888_21#_c_1731_n N_A_1714_47#_c_1864_n 9.97507e-19 $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1152 N_A_1888_21#_c_1731_n N_A_1714_47#_c_1865_n 4.0151e-19 $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1153 N_A_1888_21#_c_1666_n N_RESET_B_M1009_g 0.0181825f $X=12.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1154 N_A_1888_21#_c_1670_n N_RESET_B_M1009_g 0.0206659f $X=12.95 $Y=1.16
+ $X2=0 $Y2=0
cc_1155 N_A_1888_21#_c_1677_n N_RESET_B_M1009_g 0.00215032f $X=12.395 $Y=1.16
+ $X2=0 $Y2=0
cc_1156 N_A_1888_21#_c_1690_n N_RESET_B_M1030_g 0.0143706f $X=12.24 $Y=2 $X2=0
+ $Y2=0
cc_1157 N_A_1888_21#_c_1691_n N_RESET_B_M1030_g 0.00496908f $X=12.325 $Y=1.915
+ $X2=0 $Y2=0
cc_1158 N_A_1888_21#_c_1670_n RESET_B 7.65575e-19 $X=12.95 $Y=1.16 $X2=0 $Y2=0
cc_1159 N_A_1888_21#_c_1690_n RESET_B 0.00339513f $X=12.24 $Y=2 $X2=0 $Y2=0
cc_1160 N_A_1888_21#_c_1677_n RESET_B 0.0191707f $X=12.395 $Y=1.16 $X2=0 $Y2=0
cc_1161 N_A_1888_21#_M1002_g N_RESET_B_c_1961_n 0.0294515f $X=12.455 $Y=1.985
+ $X2=0 $Y2=0
cc_1162 N_A_1888_21#_c_1677_n N_RESET_B_c_1961_n 0.00563635f $X=12.395 $Y=1.16
+ $X2=0 $Y2=0
cc_1163 N_A_1888_21#_c_1671_n N_A_2696_47#_c_1995_n 0.00248624f $X=13.685
+ $Y=1.025 $X2=0 $Y2=0
cc_1164 N_A_1888_21#_c_1673_n N_A_2696_47#_c_1995_n 0.0159717f $X=13.815 $Y=0.73
+ $X2=0 $Y2=0
cc_1165 N_A_1888_21#_c_1672_n N_A_2696_47#_M1005_g 0.00455389f $X=13.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1166 N_A_1888_21#_c_1685_n N_A_2696_47#_M1005_g 0.0111821f $X=13.815 $Y=1.61
+ $X2=0 $Y2=0
cc_1167 N_A_1888_21#_M1051_g N_A_2696_47#_c_1997_n 0.00199156f $X=12.875 $Y=0.56
+ $X2=0 $Y2=0
cc_1168 N_A_1888_21#_c_1671_n N_A_2696_47#_c_1997_n 0.00383611f $X=13.685
+ $Y=1.025 $X2=0 $Y2=0
cc_1169 N_A_1888_21#_c_1673_n N_A_2696_47#_c_1997_n 0.00966775f $X=13.815
+ $Y=0.73 $X2=0 $Y2=0
cc_1170 N_A_1888_21#_c_1674_n N_A_2696_47#_c_1997_n 0.00992783f $X=13.815
+ $Y=0.805 $X2=0 $Y2=0
cc_1171 N_A_1888_21#_M1046_g N_A_2696_47#_c_2003_n 0.00294876f $X=12.875
+ $Y=1.985 $X2=0 $Y2=0
cc_1172 N_A_1888_21#_c_1672_n N_A_2696_47#_c_2003_n 0.00716207f $X=13.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1173 N_A_1888_21#_c_1684_n N_A_2696_47#_c_2003_n 0.0105544f $X=13.815
+ $Y=1.685 $X2=0 $Y2=0
cc_1174 N_A_1888_21#_c_1685_n N_A_2696_47#_c_2003_n 0.0103307f $X=13.815 $Y=1.61
+ $X2=0 $Y2=0
cc_1175 N_A_1888_21#_c_1674_n N_A_2696_47#_c_1998_n 0.00384385f $X=13.815
+ $Y=0.805 $X2=0 $Y2=0
cc_1176 N_A_1888_21#_c_1685_n N_A_2696_47#_c_1998_n 0.0033881f $X=13.815 $Y=1.61
+ $X2=0 $Y2=0
cc_1177 N_A_1888_21#_M1051_g N_A_2696_47#_c_1999_n 2.70228e-19 $X=12.875 $Y=0.56
+ $X2=0 $Y2=0
cc_1178 N_A_1888_21#_M1046_g N_A_2696_47#_c_1999_n 2.70228e-19 $X=12.875
+ $Y=1.985 $X2=0 $Y2=0
cc_1179 N_A_1888_21#_c_1669_n N_A_2696_47#_c_1999_n 0.0151191f $X=13.61 $Y=1.16
+ $X2=0 $Y2=0
cc_1180 N_A_1888_21#_c_1671_n N_A_2696_47#_c_1999_n 0.00117559f $X=13.685
+ $Y=1.025 $X2=0 $Y2=0
cc_1181 N_A_1888_21#_c_1672_n N_A_2696_47#_c_1999_n 0.00117559f $X=13.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1182 N_A_1888_21#_c_1675_n N_A_2696_47#_c_1999_n 0.00732445f $X=13.685
+ $Y=1.16 $X2=0 $Y2=0
cc_1183 N_A_1888_21#_c_1671_n N_A_2696_47#_c_2000_n 0.0132039f $X=13.685
+ $Y=1.025 $X2=0 $Y2=0
cc_1184 N_A_1888_21#_c_1688_n N_VPWR_M1043_d 0.00124767f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1185 N_A_1888_21#_c_1742_p N_VPWR_M1043_d 0.00160397f $X=9.8 $Y=2 $X2=0 $Y2=0
cc_1186 N_A_1888_21#_c_1690_n N_VPWR_M1029_d 0.0044189f $X=12.24 $Y=2 $X2=0
+ $Y2=0
cc_1187 N_A_1888_21#_c_1690_n N_VPWR_M1030_d 0.00750664f $X=12.24 $Y=2 $X2=0
+ $Y2=0
cc_1188 N_A_1888_21#_c_1691_n N_VPWR_M1030_d 0.00490342f $X=12.325 $Y=1.915
+ $X2=0 $Y2=0
cc_1189 N_A_1888_21#_M1046_g N_VPWR_c_2076_n 0.0031094f $X=12.875 $Y=1.985 $X2=0
+ $Y2=0
cc_1190 N_A_1888_21#_c_1669_n N_VPWR_c_2076_n 0.00532717f $X=13.61 $Y=1.16 $X2=0
+ $Y2=0
cc_1191 N_A_1888_21#_c_1672_n N_VPWR_c_2076_n 5.79288e-19 $X=13.685 $Y=1.535
+ $X2=0 $Y2=0
cc_1192 N_A_1888_21#_c_1684_n N_VPWR_c_2076_n 0.00385939f $X=13.815 $Y=1.685
+ $X2=0 $Y2=0
cc_1193 N_A_1888_21#_c_1684_n N_VPWR_c_2077_n 0.00471278f $X=13.815 $Y=1.685
+ $X2=0 $Y2=0
cc_1194 N_A_1888_21#_c_1684_n N_VPWR_c_2078_n 0.00513511f $X=13.815 $Y=1.685
+ $X2=0 $Y2=0
cc_1195 N_A_1888_21#_c_1690_n N_VPWR_c_2083_n 0.0907133f $X=12.24 $Y=2 $X2=0
+ $Y2=0
cc_1196 N_A_1888_21#_c_1688_n N_VPWR_c_2084_n 0.00359839f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1197 N_A_1888_21#_c_1796_p N_VPWR_c_2084_n 0.00713694f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1198 N_A_1888_21#_c_1714_n N_VPWR_c_2084_n 0.00458994f $X=10.73 $Y=2 $X2=0
+ $Y2=0
cc_1199 N_A_1888_21#_c_1690_n N_VPWR_c_2084_n 4.74543e-19 $X=12.24 $Y=2 $X2=0
+ $Y2=0
cc_1200 N_A_1888_21#_c_1733_n N_VPWR_c_2084_n 0.00279601f $X=10.82 $Y=2 $X2=0
+ $Y2=0
cc_1201 N_A_1888_21#_M1043_g N_VPWR_c_2089_n 0.00542601f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1202 N_A_1888_21#_c_1742_p N_VPWR_c_2089_n 9.91118e-19 $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1203 N_A_1888_21#_M1002_g N_VPWR_c_2091_n 0.0046653f $X=12.455 $Y=1.985 $X2=0
+ $Y2=0
cc_1204 N_A_1888_21#_M1046_g N_VPWR_c_2091_n 0.00541359f $X=12.875 $Y=1.985
+ $X2=0 $Y2=0
cc_1205 N_A_1888_21#_M1043_g N_VPWR_c_2097_n 0.00321606f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1206 N_A_1888_21#_c_1687_n N_VPWR_c_2097_n 7.01948e-19 $X=9.635 $Y=1.74 $X2=0
+ $Y2=0
cc_1207 N_A_1888_21#_c_1688_n N_VPWR_c_2097_n 0.0106677f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1208 N_A_1888_21#_c_1742_p N_VPWR_c_2097_n 0.0126362f $X=9.8 $Y=2 $X2=0 $Y2=0
cc_1209 N_A_1888_21#_c_1796_p N_VPWR_c_2097_n 0.00687131f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1210 N_A_1888_21#_M1002_g N_VPWR_c_2098_n 0.00846949f $X=12.455 $Y=1.985
+ $X2=0 $Y2=0
cc_1211 N_A_1888_21#_M1046_g N_VPWR_c_2098_n 6.53725e-19 $X=12.875 $Y=1.985
+ $X2=0 $Y2=0
cc_1212 N_A_1888_21#_c_1690_n N_VPWR_c_2098_n 0.00915613f $X=12.24 $Y=2 $X2=0
+ $Y2=0
cc_1213 N_A_1888_21#_M1007_d N_VPWR_c_2070_n 0.00327257f $X=10.13 $Y=2.065 $X2=0
+ $Y2=0
cc_1214 N_A_1888_21#_M1043_g N_VPWR_c_2070_n 0.00997697f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1215 N_A_1888_21#_M1002_g N_VPWR_c_2070_n 0.00791913f $X=12.455 $Y=1.985
+ $X2=0 $Y2=0
cc_1216 N_A_1888_21#_M1046_g N_VPWR_c_2070_n 0.0108665f $X=12.875 $Y=1.985 $X2=0
+ $Y2=0
cc_1217 N_A_1888_21#_c_1684_n N_VPWR_c_2070_n 0.00941266f $X=13.815 $Y=1.685
+ $X2=0 $Y2=0
cc_1218 N_A_1888_21#_c_1688_n N_VPWR_c_2070_n 0.00704318f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1219 N_A_1888_21#_c_1742_p N_VPWR_c_2070_n 0.00270501f $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1220 N_A_1888_21#_c_1796_p N_VPWR_c_2070_n 0.00608739f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1221 N_A_1888_21#_c_1714_n N_VPWR_c_2070_n 0.00829558f $X=10.73 $Y=2 $X2=0
+ $Y2=0
cc_1222 N_A_1888_21#_c_1690_n N_VPWR_c_2070_n 0.00725041f $X=12.24 $Y=2 $X2=0
+ $Y2=0
cc_1223 N_A_1888_21#_c_1733_n N_VPWR_c_2070_n 0.0049407f $X=10.82 $Y=2 $X2=0
+ $Y2=0
cc_1224 N_A_1888_21#_c_1714_n A_2122_329# 0.00202121f $X=10.73 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1225 N_A_1888_21#_c_1676_n A_2122_329# 0.00305059f $X=10.82 $Y=1.915
+ $X2=-0.19 $Y2=-0.24
cc_1226 N_A_1888_21#_c_1733_n A_2122_329# 5.84995e-19 $X=10.82 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1227 N_A_1888_21#_M1046_g N_Q_N_c_2432_n 0.00137437f $X=12.875 $Y=1.985 $X2=0
+ $Y2=0
cc_1228 N_A_1888_21#_c_1670_n N_Q_N_c_2432_n 0.00146072f $X=12.95 $Y=1.16 $X2=0
+ $Y2=0
cc_1229 N_A_1888_21#_c_1666_n N_Q_N_c_2430_n 0.00480728f $X=12.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1230 N_A_1888_21#_M1051_g N_Q_N_c_2430_n 0.00684428f $X=12.875 $Y=0.56 $X2=0
+ $Y2=0
cc_1231 N_A_1888_21#_M1046_g N_Q_N_c_2430_n 0.00808355f $X=12.875 $Y=1.985 $X2=0
+ $Y2=0
cc_1232 N_A_1888_21#_c_1670_n N_Q_N_c_2430_n 0.020126f $X=12.95 $Y=1.16 $X2=0
+ $Y2=0
cc_1233 N_A_1888_21#_c_1691_n N_Q_N_c_2430_n 0.0161038f $X=12.325 $Y=1.915 $X2=0
+ $Y2=0
cc_1234 N_A_1888_21#_c_1677_n N_Q_N_c_2430_n 0.0221731f $X=12.395 $Y=1.16 $X2=0
+ $Y2=0
cc_1235 N_A_1888_21#_M1051_g Q_N 0.00137437f $X=12.875 $Y=0.56 $X2=0 $Y2=0
cc_1236 N_A_1888_21#_c_1670_n Q_N 0.00141867f $X=12.95 $Y=1.16 $X2=0 $Y2=0
cc_1237 N_A_1888_21#_M1046_g Q_N 0.00905711f $X=12.875 $Y=1.985 $X2=0 $Y2=0
cc_1238 N_A_1888_21#_M1051_g N_Q_N_c_2443_n 0.00480183f $X=12.875 $Y=0.56 $X2=0
+ $Y2=0
cc_1239 N_A_1888_21#_M1042_g N_VGND_c_2480_n 0.00846638f $X=9.515 $Y=0.445 $X2=0
+ $Y2=0
cc_1240 N_A_1888_21#_c_1666_n N_VGND_c_2481_n 0.0105719f $X=12.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1241 N_A_1888_21#_M1051_g N_VGND_c_2481_n 7.66026e-19 $X=12.875 $Y=0.56 $X2=0
+ $Y2=0
cc_1242 N_A_1888_21#_c_1670_n N_VGND_c_2481_n 7.52163e-19 $X=12.95 $Y=1.16 $X2=0
+ $Y2=0
cc_1243 N_A_1888_21#_c_1677_n N_VGND_c_2481_n 0.0110684f $X=12.395 $Y=1.16 $X2=0
+ $Y2=0
cc_1244 N_A_1888_21#_M1051_g N_VGND_c_2482_n 0.00311062f $X=12.875 $Y=0.56 $X2=0
+ $Y2=0
cc_1245 N_A_1888_21#_c_1669_n N_VGND_c_2482_n 0.00576862f $X=13.61 $Y=1.16 $X2=0
+ $Y2=0
cc_1246 N_A_1888_21#_c_1673_n N_VGND_c_2482_n 0.00352378f $X=13.815 $Y=0.73
+ $X2=0 $Y2=0
cc_1247 N_A_1888_21#_c_1674_n N_VGND_c_2482_n 4.71945e-19 $X=13.815 $Y=0.805
+ $X2=0 $Y2=0
cc_1248 N_A_1888_21#_c_1673_n N_VGND_c_2483_n 0.00541359f $X=13.815 $Y=0.73
+ $X2=0 $Y2=0
cc_1249 N_A_1888_21#_c_1674_n N_VGND_c_2483_n 2.96334e-19 $X=13.815 $Y=0.805
+ $X2=0 $Y2=0
cc_1250 N_A_1888_21#_c_1673_n N_VGND_c_2484_n 0.00420958f $X=13.815 $Y=0.73
+ $X2=0 $Y2=0
cc_1251 N_A_1888_21#_M1042_g N_VGND_c_2491_n 0.0046653f $X=9.515 $Y=0.445 $X2=0
+ $Y2=0
cc_1252 N_A_1888_21#_c_1666_n N_VGND_c_2497_n 0.0046653f $X=12.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1253 N_A_1888_21#_M1051_g N_VGND_c_2497_n 0.00541359f $X=12.875 $Y=0.56 $X2=0
+ $Y2=0
cc_1254 N_A_1888_21#_M1001_d N_VGND_c_2505_n 0.00216833f $X=10.61 $Y=0.235 $X2=0
+ $Y2=0
cc_1255 N_A_1888_21#_M1042_g N_VGND_c_2505_n 0.00460207f $X=9.515 $Y=0.445 $X2=0
+ $Y2=0
cc_1256 N_A_1888_21#_c_1666_n N_VGND_c_2505_n 0.00796766f $X=12.455 $Y=0.995
+ $X2=0 $Y2=0
cc_1257 N_A_1888_21#_M1051_g N_VGND_c_2505_n 0.0108665f $X=12.875 $Y=0.56 $X2=0
+ $Y2=0
cc_1258 N_A_1888_21#_c_1673_n N_VGND_c_2505_n 0.0110992f $X=13.815 $Y=0.73 $X2=0
+ $Y2=0
cc_1259 N_A_1888_21#_M1001_d N_A_2004_47#_c_2748_n 0.00312752f $X=10.61 $Y=0.235
+ $X2=0 $Y2=0
cc_1260 N_A_1888_21#_c_1707_n N_A_2004_47#_c_2748_n 0.0145304f $X=10.82 $Y=0.687
+ $X2=0 $Y2=0
cc_1261 N_A_1714_47#_M1025_g N_VPWR_c_2083_n 0.00209073f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1262 N_A_1714_47#_M1025_g N_VPWR_c_2084_n 0.00425094f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1263 N_A_1714_47#_c_1872_n N_VPWR_c_2089_n 0.0377433f $X=9.21 $Y=2.335 $X2=0
+ $Y2=0
cc_1264 N_A_1714_47#_M1025_g N_VPWR_c_2097_n 0.00144209f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1265 N_A_1714_47#_M1032_d N_VPWR_c_2070_n 0.00205544f $X=8.58 $Y=2.065 $X2=0
+ $Y2=0
cc_1266 N_A_1714_47#_M1025_g N_VPWR_c_2070_n 0.00591666f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1267 N_A_1714_47#_c_1872_n N_VPWR_c_2070_n 0.0272797f $X=9.21 $Y=2.335 $X2=0
+ $Y2=0
cc_1268 N_A_1714_47#_c_1872_n A_1800_413# 0.0111731f $X=9.21 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1269 N_A_1714_47#_c_1867_n A_1800_413# 0.00577347f $X=9.295 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1270 N_A_1714_47#_c_1875_n N_VGND_c_2480_n 0.0155419f $X=9.21 $Y=0.365 $X2=0
+ $Y2=0
cc_1271 N_A_1714_47#_c_1861_n N_VGND_c_2480_n 0.00412668f $X=9.295 $Y=1.235
+ $X2=0 $Y2=0
cc_1272 N_A_1714_47#_c_1875_n N_VGND_c_2491_n 0.0433655f $X=9.21 $Y=0.365 $X2=0
+ $Y2=0
cc_1273 N_A_1714_47#_M1001_g N_VGND_c_2496_n 0.00357877f $X=10.535 $Y=0.555
+ $X2=0 $Y2=0
cc_1274 N_A_1714_47#_M1008_d N_VGND_c_2505_n 0.00272713f $X=8.57 $Y=0.235 $X2=0
+ $Y2=0
cc_1275 N_A_1714_47#_M1001_g N_VGND_c_2505_n 0.00569618f $X=10.535 $Y=0.555
+ $X2=0 $Y2=0
cc_1276 N_A_1714_47#_c_1875_n N_VGND_c_2505_n 0.0129183f $X=9.21 $Y=0.365 $X2=0
+ $Y2=0
cc_1277 N_A_1714_47#_c_1875_n A_1823_47# 0.0053026f $X=9.21 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1278 N_A_1714_47#_c_1861_n A_1823_47# 0.00495481f $X=9.295 $Y=1.235 $X2=-0.19
+ $Y2=-0.24
cc_1279 N_A_1714_47#_M1001_g N_A_2004_47#_c_2748_n 0.0110234f $X=10.535 $Y=0.555
+ $X2=0 $Y2=0
cc_1280 N_A_1714_47#_c_1864_n N_A_2004_47#_c_2748_n 0.00293167f $X=10.475
+ $Y=1.24 $X2=0 $Y2=0
cc_1281 N_A_1714_47#_c_1864_n N_A_2004_47#_c_2744_n 0.00206243f $X=10.475
+ $Y=1.24 $X2=0 $Y2=0
cc_1282 N_A_1714_47#_c_1865_n N_A_2004_47#_c_2744_n 3.6952e-19 $X=10.475 $Y=1.24
+ $X2=0 $Y2=0
cc_1283 N_RESET_B_M1030_g N_VPWR_c_2090_n 0.00655753f $X=11.97 $Y=1.825 $X2=0
+ $Y2=0
cc_1284 N_RESET_B_M1009_g N_VGND_c_2481_n 0.00665319f $X=11.97 $Y=0.445 $X2=0
+ $Y2=0
cc_1285 N_RESET_B_M1009_g N_VGND_c_2496_n 0.00585385f $X=11.97 $Y=0.445 $X2=0
+ $Y2=0
cc_1286 N_RESET_B_M1009_g N_VGND_c_2505_n 0.0120869f $X=11.97 $Y=0.445 $X2=0
+ $Y2=0
cc_1287 N_A_2696_47#_c_2003_n N_VPWR_c_2076_n 0.0621353f $X=13.605 $Y=1.91 $X2=0
+ $Y2=0
cc_1288 N_A_2696_47#_c_2003_n N_VPWR_c_2077_n 0.0169454f $X=13.605 $Y=1.91 $X2=0
+ $Y2=0
cc_1289 N_A_2696_47#_M1005_g N_VPWR_c_2078_n 0.0129456f $X=14.29 $Y=1.985 $X2=0
+ $Y2=0
cc_1290 N_A_2696_47#_M1018_g N_VPWR_c_2078_n 7.73813e-19 $X=14.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1291 N_A_2696_47#_c_2003_n N_VPWR_c_2078_n 0.0477132f $X=13.605 $Y=1.91 $X2=0
+ $Y2=0
cc_1292 N_A_2696_47#_c_1998_n N_VPWR_c_2078_n 0.010742f $X=14.205 $Y=1.16 $X2=0
+ $Y2=0
cc_1293 N_A_2696_47#_c_2000_n N_VPWR_c_2078_n 0.00259291f $X=14.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1294 N_A_2696_47#_M1018_g N_VPWR_c_2080_n 0.0031131f $X=14.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1295 N_A_2696_47#_M1005_g N_VPWR_c_2092_n 0.0046653f $X=14.29 $Y=1.985 $X2=0
+ $Y2=0
cc_1296 N_A_2696_47#_M1018_g N_VPWR_c_2092_n 0.00541359f $X=14.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1297 N_A_2696_47#_M1005_g N_VPWR_c_2070_n 0.00796766f $X=14.29 $Y=1.985 $X2=0
+ $Y2=0
cc_1298 N_A_2696_47#_M1018_g N_VPWR_c_2070_n 0.0104946f $X=14.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1299 N_A_2696_47#_c_2003_n N_VPWR_c_2070_n 0.0116159f $X=13.605 $Y=1.91 $X2=0
+ $Y2=0
cc_1300 N_A_2696_47#_c_1997_n N_Q_N_c_2430_n 0.00308112f $X=13.605 $Y=0.51 $X2=0
+ $Y2=0
cc_1301 N_A_2696_47#_c_2003_n N_Q_N_c_2430_n 0.00477082f $X=13.605 $Y=1.91 $X2=0
+ $Y2=0
cc_1302 N_A_2696_47#_c_1999_n N_Q_N_c_2430_n 0.0087488f $X=13.612 $Y=1.16 $X2=0
+ $Y2=0
cc_1303 N_A_2696_47#_c_1996_n N_Q_c_2457_n 0.00199113f $X=14.71 $Y=0.995 $X2=0
+ $Y2=0
cc_1304 N_A_2696_47#_M1005_g N_Q_c_2455_n 0.00156336f $X=14.29 $Y=1.985 $X2=0
+ $Y2=0
cc_1305 N_A_2696_47#_M1018_g N_Q_c_2455_n 0.00404758f $X=14.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1306 N_A_2696_47#_c_2003_n N_Q_c_2455_n 0.00487354f $X=13.605 $Y=1.91 $X2=0
+ $Y2=0
cc_1307 N_A_2696_47#_c_1995_n N_Q_c_2454_n 0.00395407f $X=14.29 $Y=0.995 $X2=0
+ $Y2=0
cc_1308 N_A_2696_47#_M1005_g N_Q_c_2454_n 0.00278423f $X=14.29 $Y=1.985 $X2=0
+ $Y2=0
cc_1309 N_A_2696_47#_c_1996_n N_Q_c_2454_n 0.00649275f $X=14.71 $Y=0.995 $X2=0
+ $Y2=0
cc_1310 N_A_2696_47#_M1018_g N_Q_c_2454_n 0.00582533f $X=14.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1311 N_A_2696_47#_c_1998_n N_Q_c_2454_n 0.0253118f $X=14.205 $Y=1.16 $X2=0
+ $Y2=0
cc_1312 N_A_2696_47#_c_2000_n N_Q_c_2454_n 0.027787f $X=14.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1313 N_A_2696_47#_c_1996_n Q 0.00609939f $X=14.71 $Y=0.995 $X2=0 $Y2=0
cc_1314 N_A_2696_47#_M1018_g Q 0.0115229f $X=14.71 $Y=1.985 $X2=0 $Y2=0
cc_1315 N_A_2696_47#_c_1997_n N_VGND_c_2482_n 0.0425491f $X=13.605 $Y=0.51 $X2=0
+ $Y2=0
cc_1316 N_A_2696_47#_c_1997_n N_VGND_c_2483_n 0.0199954f $X=13.605 $Y=0.51 $X2=0
+ $Y2=0
cc_1317 N_A_2696_47#_c_1995_n N_VGND_c_2484_n 0.00785757f $X=14.29 $Y=0.995
+ $X2=0 $Y2=0
cc_1318 N_A_2696_47#_c_1996_n N_VGND_c_2484_n 6.52632e-19 $X=14.71 $Y=0.995
+ $X2=0 $Y2=0
cc_1319 N_A_2696_47#_c_1997_n N_VGND_c_2484_n 0.0212808f $X=13.605 $Y=0.51 $X2=0
+ $Y2=0
cc_1320 N_A_2696_47#_c_1998_n N_VGND_c_2484_n 0.0104995f $X=14.205 $Y=1.16 $X2=0
+ $Y2=0
cc_1321 N_A_2696_47#_c_2000_n N_VGND_c_2484_n 0.00255976f $X=14.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1322 N_A_2696_47#_c_1996_n N_VGND_c_2486_n 0.0031131f $X=14.71 $Y=0.995 $X2=0
+ $Y2=0
cc_1323 N_A_2696_47#_c_1995_n N_VGND_c_2498_n 0.0046653f $X=14.29 $Y=0.995 $X2=0
+ $Y2=0
cc_1324 N_A_2696_47#_c_1996_n N_VGND_c_2498_n 0.00541359f $X=14.71 $Y=0.995
+ $X2=0 $Y2=0
cc_1325 N_A_2696_47#_M1044_s N_VGND_c_2505_n 0.00210122f $X=13.48 $Y=0.235 $X2=0
+ $Y2=0
cc_1326 N_A_2696_47#_c_1995_n N_VGND_c_2505_n 0.00796766f $X=14.29 $Y=0.995
+ $X2=0 $Y2=0
cc_1327 N_A_2696_47#_c_1996_n N_VGND_c_2505_n 0.0104946f $X=14.71 $Y=0.995 $X2=0
+ $Y2=0
cc_1328 N_A_2696_47#_c_1997_n N_VGND_c_2505_n 0.0119216f $X=13.605 $Y=0.51 $X2=0
+ $Y2=0
cc_1329 N_VPWR_c_2070_n N_A_453_47#_M1019_d 0.00306969f $X=14.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1330 N_VPWR_c_2072_n N_A_453_47#_c_2306_n 0.0170763f $X=1.62 $Y=1.97 $X2=0
+ $Y2=0
cc_1331 N_VPWR_c_2087_n N_A_453_47#_c_2306_n 0.0151498f $X=3.295 $Y=2.72 $X2=0
+ $Y2=0
cc_1332 N_VPWR_c_2070_n N_A_453_47#_c_2306_n 0.00610123f $X=14.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1333 N_VPWR_c_2088_n N_A_453_47#_c_2304_n 0.0154725f $X=5.705 $Y=2.72 $X2=0
+ $Y2=0
cc_1334 N_VPWR_c_2070_n N_A_453_47#_c_2304_n 0.00409094f $X=14.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1335 N_VPWR_c_2070_n A_752_413# 0.00238611f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1336 N_VPWR_c_2070_n A_1017_413# 0.00355877f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1337 N_VPWR_c_2070_n A_1351_329# 0.0026811f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1338 N_VPWR_c_2070_n A_1572_329# 0.00777501f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1339 N_VPWR_c_2070_n A_1800_413# 0.00566996f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1340 N_VPWR_c_2070_n A_2122_329# 0.00245111f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1341 N_VPWR_c_2070_n N_Q_N_M1002_d 0.00393857f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1342 N_VPWR_c_2091_n Q_N 0.0151826f $X=13 $Y=2.72 $X2=0 $Y2=0
cc_1343 N_VPWR_c_2070_n Q_N 0.00941829f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1344 N_VPWR_c_2070_n N_Q_M1005_s 0.00393857f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1345 N_VPWR_c_2092_n Q 0.0151826f $X=14.835 $Y=2.72 $X2=0 $Y2=0
cc_1346 N_VPWR_c_2070_n Q 0.00941829f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1347 N_VPWR_c_2076_n N_VGND_c_2482_n 0.00786011f $X=13.085 $Y=1.66 $X2=0
+ $Y2=0
cc_1348 N_VPWR_c_2080_n N_VGND_c_2486_n 0.00810308f $X=14.92 $Y=1.66 $X2=0 $Y2=0
cc_1349 N_A_453_47#_c_2304_n N_VGND_c_2487_n 0.0115451f $X=4.315 $Y=0.47 $X2=0
+ $Y2=0
cc_1350 N_A_453_47#_c_2299_n N_VGND_c_2495_n 0.0259189f $X=2.645 $Y=0.43 $X2=0
+ $Y2=0
cc_1351 N_A_453_47#_M1012_d N_VGND_c_2505_n 0.00187997f $X=2.265 $Y=0.235 $X2=0
+ $Y2=0
cc_1352 N_A_453_47#_M1024_d N_VGND_c_2505_n 0.00295839f $X=4.18 $Y=0.235 $X2=0
+ $Y2=0
cc_1353 N_A_453_47#_c_2299_n N_VGND_c_2505_n 0.00727734f $X=2.645 $Y=0.43 $X2=0
+ $Y2=0
cc_1354 N_A_453_47#_c_2304_n N_VGND_c_2505_n 0.00398697f $X=4.315 $Y=0.47 $X2=0
+ $Y2=0
cc_1355 N_Q_N_c_2430_n N_VGND_c_2481_n 0.00491339f $X=12.705 $Y=1.63 $X2=0 $Y2=0
cc_1356 N_Q_N_c_2443_n N_VGND_c_2497_n 0.0150393f $X=12.705 $Y=0.59 $X2=0 $Y2=0
cc_1357 N_Q_N_M1049_s N_VGND_c_2505_n 0.00393857f $X=12.53 $Y=0.235 $X2=0 $Y2=0
cc_1358 N_Q_N_c_2443_n N_VGND_c_2505_n 0.00938807f $X=12.705 $Y=0.59 $X2=0 $Y2=0
cc_1359 Q N_VGND_c_2498_n 0.0151484f $X=14.44 $Y=0.425 $X2=0 $Y2=0
cc_1360 N_Q_M1015_d N_VGND_c_2505_n 0.00393857f $X=14.365 $Y=0.235 $X2=0 $Y2=0
cc_1361 Q N_VGND_c_2505_n 0.00941054f $X=14.44 $Y=0.425 $X2=0 $Y2=0
cc_1362 N_VGND_c_2505_n A_381_47# 0.00165237f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1363 N_VGND_c_2505_n A_764_47# 0.00302076f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1364 N_VGND_c_2505_n A_1041_47# 0.0022723f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1365 N_VGND_c_2505_n N_A_1251_47#_M1047_d 0.00214379f $X=14.95 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1366 N_VGND_c_2505_n N_A_1251_47#_M1014_d 0.00204204f $X=14.95 $Y=0 $X2=0
+ $Y2=0
cc_1367 N_VGND_c_2479_n N_A_1251_47#_c_2713_n 0.010563f $X=7.81 $Y=0.38 $X2=0
+ $Y2=0
cc_1368 N_VGND_c_2489_n N_A_1251_47#_c_2713_n 0.0113927f $X=7.645 $Y=0 $X2=0
+ $Y2=0
cc_1369 N_VGND_c_2505_n N_A_1251_47#_c_2713_n 0.00305438f $X=14.95 $Y=0 $X2=0
+ $Y2=0
cc_1370 N_VGND_c_2479_n N_A_1251_47#_c_2716_n 0.0022149f $X=7.81 $Y=0.38 $X2=0
+ $Y2=0
cc_1371 N_VGND_c_2489_n N_A_1251_47#_c_2723_n 0.0540424f $X=7.645 $Y=0 $X2=0
+ $Y2=0
cc_1372 N_VGND_c_2505_n N_A_1251_47#_c_2723_n 0.0159669f $X=14.95 $Y=0 $X2=0
+ $Y2=0
cc_1373 N_VGND_c_2505_n A_1619_47# 0.00467499f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1374 N_VGND_c_2505_n A_1823_47# 0.00261578f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1375 N_VGND_c_2505_n N_A_2004_47#_M1004_d 0.00378249f $X=14.95 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1376 N_VGND_c_2505_n N_A_2004_47#_M1017_d 0.00251082f $X=14.95 $Y=0 $X2=0
+ $Y2=0
cc_1377 N_VGND_c_2496_n N_A_2004_47#_c_2748_n 0.0358653f $X=12.08 $Y=0 $X2=0
+ $Y2=0
cc_1378 N_VGND_c_2505_n N_A_2004_47#_c_2748_n 0.0235203f $X=14.95 $Y=0 $X2=0
+ $Y2=0
cc_1379 N_VGND_c_2496_n N_A_2004_47#_c_2744_n 0.0215241f $X=12.08 $Y=0 $X2=0
+ $Y2=0
cc_1380 N_VGND_c_2505_n N_A_2004_47#_c_2744_n 0.01237f $X=14.95 $Y=0 $X2=0 $Y2=0
cc_1381 N_VGND_c_2496_n N_A_2004_47#_c_2749_n 0.0110309f $X=12.08 $Y=0 $X2=0
+ $Y2=0
cc_1382 N_VGND_c_2505_n N_A_2004_47#_c_2749_n 0.0063548f $X=14.95 $Y=0 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__o2111ai_4.pxi.spice
* Created: Thu Aug 27 14:34:20 2020
* 
x_PM_SKY130_FD_SC_HD__O2111AI_4%D1 N_D1_M1016_g N_D1_c_134_n N_D1_M1003_g
+ N_D1_M1020_g N_D1_c_135_n N_D1_M1009_g N_D1_M1023_g N_D1_c_136_n N_D1_M1025_g
+ N_D1_M1039_g N_D1_c_137_n N_D1_M1036_g D1 D1 D1 N_D1_c_133_n
+ PM_SKY130_FD_SC_HD__O2111AI_4%D1
x_PM_SKY130_FD_SC_HD__O2111AI_4%C1 N_C1_M1021_g N_C1_M1001_g N_C1_M1026_g
+ N_C1_M1010_g N_C1_M1032_g N_C1_M1030_g N_C1_M1033_g N_C1_M1037_g C1 C1 C1 C1
+ N_C1_c_200_n PM_SKY130_FD_SC_HD__O2111AI_4%C1
x_PM_SKY130_FD_SC_HD__O2111AI_4%B1 N_B1_M1007_g N_B1_M1014_g N_B1_M1013_g
+ N_B1_M1017_g N_B1_M1015_g N_B1_c_270_n N_B1_M1022_g N_B1_M1038_g N_B1_c_272_n
+ N_B1_c_273_n N_B1_c_274_n N_B1_M1027_g B1 B1 B1 B1
+ PM_SKY130_FD_SC_HD__O2111AI_4%B1
x_PM_SKY130_FD_SC_HD__O2111AI_4%A2 N_A2_c_354_n N_A2_M1002_g N_A2_c_345_n
+ N_A2_c_346_n N_A2_M1024_g N_A2_c_357_n N_A2_M1008_g N_A2_M1028_g N_A2_M1011_g
+ N_A2_M1029_g N_A2_c_351_n N_A2_M1034_g N_A2_M1031_g A2 A2 A2
+ PM_SKY130_FD_SC_HD__O2111AI_4%A2
x_PM_SKY130_FD_SC_HD__O2111AI_4%A1 N_A1_M1005_g N_A1_M1000_g N_A1_M1006_g
+ N_A1_M1004_g N_A1_M1012_g N_A1_M1019_g N_A1_M1018_g N_A1_M1035_g A1 A1 A1 A1
+ N_A1_c_443_n PM_SKY130_FD_SC_HD__O2111AI_4%A1
x_PM_SKY130_FD_SC_HD__O2111AI_4%Y N_Y_M1016_s N_Y_M1023_s N_Y_M1003_s
+ N_Y_M1009_s N_Y_M1036_s N_Y_M1010_s N_Y_M1037_s N_Y_M1013_s N_Y_M1038_s
+ N_Y_M1008_d N_Y_M1034_d N_Y_c_508_n N_Y_c_514_n N_Y_c_579_p N_Y_c_518_n
+ N_Y_c_580_p N_Y_c_526_n N_Y_c_581_p N_Y_c_530_n N_Y_c_538_n N_Y_c_539_n
+ N_Y_c_583_p N_Y_c_543_n N_Y_c_552_n N_Y_c_547_n N_Y_c_608_p N_Y_c_522_n
+ N_Y_c_534_n N_Y_c_535_n N_Y_c_537_n N_Y_c_548_n N_Y_c_550_n N_Y_c_557_n
+ N_Y_c_504_n N_Y_c_561_n Y Y Y Y Y N_Y_c_502_n Y
+ PM_SKY130_FD_SC_HD__O2111AI_4%Y
x_PM_SKY130_FD_SC_HD__O2111AI_4%VPWR N_VPWR_M1003_d N_VPWR_M1025_d
+ N_VPWR_M1001_d N_VPWR_M1030_d N_VPWR_M1007_d N_VPWR_M1015_d N_VPWR_M1000_d
+ N_VPWR_M1004_d N_VPWR_M1035_d N_VPWR_c_629_n N_VPWR_c_630_n N_VPWR_c_631_n
+ N_VPWR_c_632_n N_VPWR_c_633_n N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_636_n
+ N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n N_VPWR_c_641_n
+ N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n N_VPWR_c_646_n
+ N_VPWR_c_647_n N_VPWR_c_648_n VPWR N_VPWR_c_649_n N_VPWR_c_650_n
+ N_VPWR_c_651_n N_VPWR_c_652_n N_VPWR_c_653_n N_VPWR_c_654_n N_VPWR_c_655_n
+ N_VPWR_c_628_n PM_SKY130_FD_SC_HD__O2111AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O2111AI_4%A_1163_297# N_A_1163_297#_M1002_s
+ N_A_1163_297#_M1011_s N_A_1163_297#_M1000_s N_A_1163_297#_M1019_s
+ N_A_1163_297#_c_786_n N_A_1163_297#_c_789_n N_A_1163_297#_c_792_n
+ N_A_1163_297#_c_794_n N_A_1163_297#_c_785_n N_A_1163_297#_c_797_n
+ N_A_1163_297#_c_835_n N_A_1163_297#_c_801_n N_A_1163_297#_c_805_n
+ N_A_1163_297#_c_839_n N_A_1163_297#_c_841_n
+ PM_SKY130_FD_SC_HD__O2111AI_4%A_1163_297#
x_PM_SKY130_FD_SC_HD__O2111AI_4%A_27_47# N_A_27_47#_M1016_d N_A_27_47#_M1020_d
+ N_A_27_47#_M1039_d N_A_27_47#_M1026_s N_A_27_47#_M1033_s N_A_27_47#_c_842_n
+ N_A_27_47#_c_849_n N_A_27_47#_c_843_n PM_SKY130_FD_SC_HD__O2111AI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O2111AI_4%A_445_47# N_A_445_47#_M1021_d
+ N_A_445_47#_M1032_d N_A_445_47#_M1014_d N_A_445_47#_M1022_d
+ N_A_445_47#_c_878_n PM_SKY130_FD_SC_HD__O2111AI_4%A_445_47#
x_PM_SKY130_FD_SC_HD__O2111AI_4%A_803_47# N_A_803_47#_M1014_s
+ N_A_803_47#_M1017_s N_A_803_47#_M1027_s N_A_803_47#_M1028_d
+ N_A_803_47#_M1031_d N_A_803_47#_M1006_s N_A_803_47#_M1018_s
+ N_A_803_47#_c_908_n PM_SKY130_FD_SC_HD__O2111AI_4%A_803_47#
x_PM_SKY130_FD_SC_HD__O2111AI_4%VGND N_VGND_M1024_s N_VGND_M1029_s
+ N_VGND_M1005_d N_VGND_M1012_d N_VGND_c_959_n N_VGND_c_960_n N_VGND_c_961_n
+ N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n VGND N_VGND_c_965_n
+ N_VGND_c_966_n N_VGND_c_967_n N_VGND_c_968_n N_VGND_c_969_n N_VGND_c_970_n
+ N_VGND_c_971_n N_VGND_c_972_n PM_SKY130_FD_SC_HD__O2111AI_4%VGND
cc_1 VNB N_D1_M1016_g 0.0207797f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_D1_M1020_g 0.0174986f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_D1_M1023_g 0.017506f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_4 VNB N_D1_M1039_g 0.017802f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_5 VNB N_D1_c_133_n 0.0610365f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.205
cc_6 VNB N_C1_M1021_g 0.017802f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_7 VNB N_C1_M1001_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_8 VNB N_C1_M1026_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C1_M1010_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_10 VNB N_C1_M1032_g 0.017506f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.385
cc_11 VNB N_C1_M1030_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_12 VNB N_C1_M1033_g 0.0238324f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_13 VNB N_C1_M1037_g 4.35699e-19 $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_14 VNB C1 0.0053307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_C1_c_200_n 0.0635056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_M1007_g 4.35699e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_17 VNB N_B1_M1014_g 0.0234953f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_18 VNB N_B1_M1013_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B1_M1017_g 0.017055f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_20 VNB N_B1_M1015_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.385
cc_21 VNB N_B1_c_270_n 0.0140536f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_22 VNB N_B1_M1038_g 3.36363e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.385
cc_23 VNB N_B1_c_272_n 0.0187228f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_24 VNB N_B1_c_273_n 0.0807034f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_25 VNB N_B1_c_274_n 0.0144056f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_26 VNB B1 0.00520689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A2_c_345_n 0.00530647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A2_c_346_n 0.00487696f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.385
cc_29 VNB N_A2_M1024_g 0.0176044f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_30 VNB N_A2_M1028_g 0.0173006f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_31 VNB N_A2_M1011_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.385
cc_32 VNB N_A2_M1029_g 0.0173006f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_33 VNB N_A2_c_351_n 0.0751798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A2_M1034_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_35 VNB N_A2_M1031_g 0.0176044f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_36 VNB N_A1_M1005_g 0.0176044f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_37 VNB N_A1_M1000_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_38 VNB N_A1_M1006_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A1_M1004_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_40 VNB N_A1_M1012_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.385
cc_41 VNB N_A1_M1019_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_42 VNB N_A1_M1018_g 0.0236684f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_43 VNB N_A1_M1035_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_44 VNB A1 0.0170052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A1_c_443_n 0.0832065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_502_n 0.00771117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB Y 0.0249535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_628_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_27_47#_c_842_n 0.00860317f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_50 VNB N_A_27_47#_c_843_n 0.00391512f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_51 VNB N_A_445_47#_c_878_n 0.0077648f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_52 VNB N_A_803_47#_c_908_n 0.0527475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_959_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_54 VNB N_VGND_c_960_n 3.10008e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.385
cc_55 VNB N_VGND_c_961_n 3.06325e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_56 VNB N_VGND_c_962_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_57 VNB N_VGND_c_963_n 0.011903f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_58 VNB N_VGND_c_964_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_59 VNB N_VGND_c_965_n 0.14239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_966_n 0.0124541f $X=-0.19 $Y=-0.24 $X2=1.565 $Y2=1.205
cc_61 VNB N_VGND_c_967_n 0.0125918f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.21
cc_62 VNB N_VGND_c_968_n 0.0203624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_969_n 0.455195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_970_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_971_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_972_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VPB N_D1_c_134_n 0.0184709f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.385
cc_68 VPB N_D1_c_135_n 0.0152726f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.385
cc_69 VPB N_D1_c_136_n 0.0155051f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.385
cc_70 VPB N_D1_c_137_n 0.0155605f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.385
cc_71 VPB N_D1_c_133_n 0.0219658f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.205
cc_72 VPB N_C1_M1001_g 0.0193615f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_73 VPB N_C1_M1010_g 0.0190588f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_74 VPB N_C1_M1030_g 0.0190588f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_75 VPB N_C1_M1037_g 0.0214991f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_76 VPB C1 0.00990535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_B1_M1007_g 0.0214153f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_78 VPB N_B1_M1013_g 0.0190588f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_B1_M1015_g 0.0190588f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.385
cc_80 VPB N_B1_M1038_g 0.0198354f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.385
cc_81 VPB B1 0.0103246f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A2_c_354_n 0.0146376f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.025
cc_83 VPB N_A2_c_345_n 0.00341503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A2_c_346_n 0.00478656f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.385
cc_85 VPB N_A2_c_357_n 0.0142545f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_86 VPB N_A2_M1011_g 0.0192302f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.385
cc_87 VPB N_A2_c_351_n 0.00484905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A2_M1034_g 0.0267826f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_89 VPB A2 0.00776907f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.205
cc_90 VPB N_A1_M1000_g 0.0259101f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_91 VPB N_A1_M1004_g 0.0191286f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_92 VPB N_A1_M1019_g 0.0190728f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_93 VPB N_A1_M1035_g 0.0268619f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_94 VPB A1 0.0143153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_Y_c_504_n 0.00391181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB Y 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB Y 0.0301593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB Y 0.010326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_629_n 4.01705e-19 $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_100 VPB N_VPWR_c_630_n 0.00184027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_631_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.16
cc_102 VPB N_VPWR_c_632_n 3.99007e-19 $X=-0.19 $Y=1.305 $X2=1.565 $Y2=1.205
cc_103 VPB N_VPWR_c_633_n 3.99099e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_634_n 0.0025461f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.21
cc_105 VPB N_VPWR_c_635_n 0.00635656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_636_n 3.1087e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_637_n 0.0108492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_638_n 0.0420559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_639_n 0.0145068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_640_n 0.00427244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_641_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_642_n 0.00410235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_643_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_644_n 0.00410235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_645_n 0.018986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_646_n 0.0043021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_647_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_648_n 0.00436862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_649_n 0.0153939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_650_n 0.0581754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_651_n 0.0121474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_652_n 0.0144639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_653_n 0.00416893f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_654_n 0.00507318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_655_n 0.00410235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_628_n 0.0466435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_1163_297#_c_785_n 0.0126665f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_128 N_D1_M1039_g N_C1_M1021_g 0.02306f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_129 N_D1_c_137_n N_C1_M1001_g 0.02306f $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_130 D1 C1 0.0224052f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_131 N_D1_c_133_n C1 0.00227309f $X=1.73 $Y=1.205 $X2=0 $Y2=0
cc_132 D1 N_C1_c_200_n 2.46803e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_133 N_D1_c_133_n N_C1_c_200_n 0.02306f $X=1.73 $Y=1.205 $X2=0 $Y2=0
cc_134 N_D1_M1016_g N_Y_c_508_n 0.0143719f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_135 N_D1_M1020_g N_Y_c_508_n 0.00887971f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_136 N_D1_M1023_g N_Y_c_508_n 0.00887971f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_137 N_D1_M1039_g N_Y_c_508_n 0.00264703f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_138 D1 N_Y_c_508_n 0.0498613f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_139 N_D1_c_133_n N_Y_c_508_n 0.00614247f $X=1.73 $Y=1.205 $X2=0 $Y2=0
cc_140 N_D1_c_134_n N_Y_c_514_n 0.0205647f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_141 N_D1_c_135_n N_Y_c_514_n 0.014062f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_142 D1 N_Y_c_514_n 0.0278503f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_143 N_D1_c_133_n N_Y_c_514_n 0.0021532f $X=1.73 $Y=1.205 $X2=0 $Y2=0
cc_144 N_D1_c_136_n N_Y_c_518_n 0.0149489f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_145 N_D1_c_137_n N_Y_c_518_n 0.0158507f $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_146 D1 N_Y_c_518_n 0.0345141f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_147 N_D1_c_133_n N_Y_c_518_n 0.0021532f $X=1.73 $Y=1.205 $X2=0 $Y2=0
cc_148 D1 N_Y_c_522_n 0.013582f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_149 N_D1_c_133_n N_Y_c_522_n 0.00223856f $X=1.73 $Y=1.205 $X2=0 $Y2=0
cc_150 N_D1_M1016_g Y 0.0255072f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_151 D1 Y 0.0222691f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_152 N_D1_c_134_n N_VPWR_c_629_n 0.0114522f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_153 N_D1_c_135_n N_VPWR_c_629_n 0.0109027f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_154 N_D1_c_136_n N_VPWR_c_629_n 6.40449e-19 $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_155 N_D1_c_136_n N_VPWR_c_630_n 0.00155375f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_156 N_D1_c_137_n N_VPWR_c_630_n 0.00975795f $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_157 N_D1_c_137_n N_VPWR_c_631_n 6.17924e-19 $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_158 N_D1_c_135_n N_VPWR_c_639_n 0.0046653f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_159 N_D1_c_136_n N_VPWR_c_639_n 0.00585385f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_160 N_D1_c_137_n N_VPWR_c_641_n 0.00505556f $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_161 N_D1_c_134_n N_VPWR_c_649_n 0.00525069f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_162 N_D1_c_134_n N_VPWR_c_628_n 0.00976741f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_163 N_D1_c_135_n N_VPWR_c_628_n 0.00789179f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_164 N_D1_c_136_n N_VPWR_c_628_n 0.0104242f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_165 N_D1_c_137_n N_VPWR_c_628_n 0.00853327f $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_166 N_D1_M1016_g N_A_27_47#_c_842_n 0.00834759f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_167 N_D1_M1020_g N_A_27_47#_c_842_n 0.00834759f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_168 N_D1_M1023_g N_A_27_47#_c_842_n 0.00829818f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_169 N_D1_M1039_g N_A_27_47#_c_842_n 0.0115341f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_170 D1 N_A_27_47#_c_842_n 0.00174796f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_171 N_D1_M1039_g N_A_445_47#_c_878_n 2.26e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_172 N_D1_M1016_g N_VGND_c_965_n 0.00364081f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_173 N_D1_M1020_g N_VGND_c_965_n 0.00364081f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_174 N_D1_M1023_g N_VGND_c_965_n 0.00364081f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_175 N_D1_M1039_g N_VGND_c_965_n 0.00364081f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_176 N_D1_M1016_g N_VGND_c_969_n 0.00618903f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_177 N_D1_M1020_g N_VGND_c_969_n 0.00523483f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_178 N_D1_M1023_g N_VGND_c_969_n 0.00523483f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_179 N_D1_M1039_g N_VGND_c_969_n 0.00530203f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_180 N_C1_M1037_g N_B1_M1007_g 0.0209867f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_181 N_C1_M1033_g N_B1_c_273_n 0.00887041f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_182 C1 N_B1_c_273_n 8.98283e-19 $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_183 C1 B1 0.0183754f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_184 N_C1_c_200_n B1 0.00110625f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_185 N_C1_M1001_g N_Y_c_526_n 0.0143236f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_186 N_C1_M1010_g N_Y_c_526_n 0.0143678f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_187 C1 N_Y_c_526_n 0.0408845f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_188 N_C1_c_200_n N_Y_c_526_n 5.55696e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_189 N_C1_M1030_g N_Y_c_530_n 0.0143678f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_190 N_C1_M1037_g N_Y_c_530_n 0.0152892f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_191 C1 N_Y_c_530_n 0.0408845f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_192 N_C1_c_200_n N_Y_c_530_n 5.55696e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_193 C1 N_Y_c_534_n 0.0073538f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_194 C1 N_Y_c_535_n 0.0147075f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_195 N_C1_c_200_n N_Y_c_535_n 6.26351e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_196 C1 N_Y_c_537_n 0.00137301f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_197 N_C1_M1001_g N_VPWR_c_630_n 6.16453e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_198 N_C1_M1001_g N_VPWR_c_631_n 0.0100176f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_199 N_C1_M1010_g N_VPWR_c_631_n 0.0100176f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_200 N_C1_M1030_g N_VPWR_c_631_n 6.17924e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_201 N_C1_M1010_g N_VPWR_c_632_n 6.17924e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_202 N_C1_M1030_g N_VPWR_c_632_n 0.0100176f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_203 N_C1_M1037_g N_VPWR_c_632_n 0.0113861f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_204 N_C1_M1037_g N_VPWR_c_633_n 0.00105067f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_205 N_C1_M1001_g N_VPWR_c_641_n 0.00505556f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_206 N_C1_M1010_g N_VPWR_c_643_n 0.00505556f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_207 N_C1_M1030_g N_VPWR_c_643_n 0.00505556f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_208 N_C1_M1037_g N_VPWR_c_645_n 0.00505556f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_209 N_C1_M1001_g N_VPWR_c_628_n 0.00853327f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_210 N_C1_M1010_g N_VPWR_c_628_n 0.00850607f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_211 N_C1_M1030_g N_VPWR_c_628_n 0.00850607f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_212 N_C1_M1037_g N_VPWR_c_628_n 0.00895656f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_213 C1 N_A_27_47#_c_849_n 0.00517387f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_214 N_C1_M1021_g N_A_27_47#_c_843_n 0.0115423f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_215 N_C1_M1026_g N_A_27_47#_c_843_n 0.00983161f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_216 N_C1_M1032_g N_A_27_47#_c_843_n 0.00988628f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_217 N_C1_M1033_g N_A_27_47#_c_843_n 0.00988628f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_218 C1 N_A_27_47#_c_843_n 0.0700367f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_219 N_C1_c_200_n N_A_27_47#_c_843_n 0.00588438f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_220 N_C1_M1021_g N_A_445_47#_c_878_n 0.00288225f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_221 N_C1_M1026_g N_A_445_47#_c_878_n 0.00814603f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_222 N_C1_M1032_g N_A_445_47#_c_878_n 0.00814603f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_223 N_C1_M1033_g N_A_445_47#_c_878_n 0.0104994f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_224 N_C1_M1033_g N_A_803_47#_c_908_n 0.00161288f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_225 N_C1_M1021_g N_VGND_c_965_n 0.00409265f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_226 N_C1_M1026_g N_VGND_c_965_n 0.00357877f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_227 N_C1_M1032_g N_VGND_c_965_n 0.00357877f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_228 N_C1_M1033_g N_VGND_c_965_n 0.00357877f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_229 N_C1_M1021_g N_VGND_c_969_n 0.00570536f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_230 N_C1_M1026_g N_VGND_c_969_n 0.00522516f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_231 N_C1_M1032_g N_VGND_c_969_n 0.00522516f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_232 N_C1_M1033_g N_VGND_c_969_n 0.00660224f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_233 N_B1_M1038_g N_A2_c_346_n 0.0264769f $X=5.295 $Y=1.985 $X2=0 $Y2=0
cc_234 N_B1_c_272_n N_A2_c_346_n 0.0011985f $X=5.535 $Y=1.035 $X2=0 $Y2=0
cc_235 N_B1_c_273_n N_A2_c_346_n 0.00111887f $X=5.37 $Y=1.035 $X2=0 $Y2=0
cc_236 B1 N_A2_c_346_n 0.00109941f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_237 N_B1_c_274_n N_A2_M1024_g 0.0141706f $X=5.61 $Y=0.96 $X2=0 $Y2=0
cc_238 N_B1_c_272_n N_A2_c_351_n 0.016054f $X=5.535 $Y=1.035 $X2=0 $Y2=0
cc_239 N_B1_c_273_n N_A2_c_351_n 0.00233558f $X=5.37 $Y=1.035 $X2=0 $Y2=0
cc_240 B1 N_A2_c_351_n 0.00168061f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_241 B1 A2 0.00835016f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_242 N_B1_M1007_g N_Y_c_538_n 0.00868125f $X=4.035 $Y=1.985 $X2=0 $Y2=0
cc_243 N_B1_M1007_g N_Y_c_539_n 0.0148304f $X=4.035 $Y=1.985 $X2=0 $Y2=0
cc_244 N_B1_M1013_g N_Y_c_539_n 0.0143678f $X=4.455 $Y=1.985 $X2=0 $Y2=0
cc_245 N_B1_c_273_n N_Y_c_539_n 9.34498e-19 $X=5.37 $Y=1.035 $X2=0 $Y2=0
cc_246 B1 N_Y_c_539_n 0.0483212f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_247 N_B1_M1015_g N_Y_c_543_n 0.0143678f $X=4.875 $Y=1.985 $X2=0 $Y2=0
cc_248 N_B1_M1038_g N_Y_c_543_n 0.0150519f $X=5.295 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B1_c_273_n N_Y_c_543_n 5.46557e-19 $X=5.37 $Y=1.035 $X2=0 $Y2=0
cc_250 B1 N_Y_c_543_n 0.0408845f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_251 N_B1_c_272_n N_Y_c_547_n 2.83518e-19 $X=5.535 $Y=1.035 $X2=0 $Y2=0
cc_252 N_B1_c_273_n N_Y_c_548_n 6.17186e-19 $X=5.37 $Y=1.035 $X2=0 $Y2=0
cc_253 B1 N_Y_c_548_n 0.0147075f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_254 N_B1_c_272_n N_Y_c_550_n 0.00377546f $X=5.535 $Y=1.035 $X2=0 $Y2=0
cc_255 B1 N_Y_c_550_n 0.0030818f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_256 N_B1_M1007_g N_VPWR_c_632_n 9.56803e-19 $X=4.035 $Y=1.985 $X2=0 $Y2=0
cc_257 N_B1_M1007_g N_VPWR_c_633_n 0.0154076f $X=4.035 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B1_M1013_g N_VPWR_c_633_n 0.0100176f $X=4.455 $Y=1.985 $X2=0 $Y2=0
cc_259 N_B1_M1015_g N_VPWR_c_633_n 6.1876e-19 $X=4.875 $Y=1.985 $X2=0 $Y2=0
cc_260 N_B1_M1013_g N_VPWR_c_634_n 6.16756e-19 $X=4.455 $Y=1.985 $X2=0 $Y2=0
cc_261 N_B1_M1015_g N_VPWR_c_634_n 0.00976915f $X=4.875 $Y=1.985 $X2=0 $Y2=0
cc_262 N_B1_M1038_g N_VPWR_c_634_n 0.00308779f $X=5.295 $Y=1.985 $X2=0 $Y2=0
cc_263 N_B1_M1007_g N_VPWR_c_645_n 0.00447018f $X=4.035 $Y=1.985 $X2=0 $Y2=0
cc_264 N_B1_M1013_g N_VPWR_c_647_n 0.00505556f $X=4.455 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B1_M1015_g N_VPWR_c_647_n 0.00505556f $X=4.875 $Y=1.985 $X2=0 $Y2=0
cc_266 N_B1_M1038_g N_VPWR_c_650_n 0.00583607f $X=5.295 $Y=1.985 $X2=0 $Y2=0
cc_267 N_B1_M1007_g N_VPWR_c_628_n 0.00812834f $X=4.035 $Y=1.985 $X2=0 $Y2=0
cc_268 N_B1_M1013_g N_VPWR_c_628_n 0.00850607f $X=4.455 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B1_M1015_g N_VPWR_c_628_n 0.00850607f $X=4.875 $Y=1.985 $X2=0 $Y2=0
cc_270 N_B1_M1038_g N_VPWR_c_628_n 0.0104934f $X=5.295 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B1_M1014_g N_A_445_47#_c_878_n 0.0107397f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_272 N_B1_M1017_g N_A_445_47#_c_878_n 0.00838637f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_273 N_B1_c_270_n N_A_445_47#_c_878_n 0.00838637f $X=5.19 $Y=0.96 $X2=0 $Y2=0
cc_274 N_B1_c_273_n N_A_445_47#_c_878_n 0.00190775f $X=5.37 $Y=1.035 $X2=0 $Y2=0
cc_275 N_B1_c_274_n N_A_445_47#_c_878_n 0.0040785f $X=5.61 $Y=0.96 $X2=0 $Y2=0
cc_276 B1 N_A_445_47#_c_878_n 0.00467659f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_277 N_B1_M1014_g N_A_803_47#_c_908_n 0.0110908f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_278 N_B1_M1017_g N_A_803_47#_c_908_n 0.0109368f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_279 N_B1_c_270_n N_A_803_47#_c_908_n 0.0109368f $X=5.19 $Y=0.96 $X2=0 $Y2=0
cc_280 N_B1_c_273_n N_A_803_47#_c_908_n 0.0153223f $X=5.37 $Y=1.035 $X2=0 $Y2=0
cc_281 N_B1_c_274_n N_A_803_47#_c_908_n 0.0128164f $X=5.61 $Y=0.96 $X2=0 $Y2=0
cc_282 B1 N_A_803_47#_c_908_n 0.111102f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_283 N_B1_c_274_n N_VGND_c_959_n 0.00187222f $X=5.61 $Y=0.96 $X2=0 $Y2=0
cc_284 N_B1_M1014_g N_VGND_c_965_n 0.00357877f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_285 N_B1_M1017_g N_VGND_c_965_n 0.00357877f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_286 N_B1_c_270_n N_VGND_c_965_n 0.00357877f $X=5.19 $Y=0.96 $X2=0 $Y2=0
cc_287 N_B1_c_274_n N_VGND_c_965_n 0.00413993f $X=5.61 $Y=0.96 $X2=0 $Y2=0
cc_288 N_B1_M1014_g N_VGND_c_969_n 0.00660224f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_289 N_B1_M1017_g N_VGND_c_969_n 0.00522516f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_290 N_B1_c_270_n N_VGND_c_969_n 0.00522516f $X=5.19 $Y=0.96 $X2=0 $Y2=0
cc_291 N_B1_c_274_n N_VGND_c_969_n 0.00584536f $X=5.61 $Y=0.96 $X2=0 $Y2=0
cc_292 N_A2_M1031_g N_A1_M1005_g 0.0193894f $X=7.335 $Y=0.56 $X2=0 $Y2=0
cc_293 A2 N_A1_M1000_g 4.19056e-19 $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_294 N_A2_c_351_n A1 8.61314e-19 $X=7 $Y=1.295 $X2=0 $Y2=0
cc_295 A2 A1 0.00966851f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_296 N_A2_c_351_n N_A1_c_443_n 0.0193894f $X=7 $Y=1.295 $X2=0 $Y2=0
cc_297 A2 N_A1_c_443_n 9.12663e-19 $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_298 N_A2_c_354_n N_Y_c_552_n 0.00555275f $X=5.74 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A2_c_354_n N_Y_c_547_n 0.0152484f $X=5.74 $Y=1.41 $X2=0 $Y2=0
cc_300 N_A2_c_345_n N_Y_c_547_n 0.00240394f $X=5.98 $Y=1.335 $X2=0 $Y2=0
cc_301 N_A2_c_357_n N_Y_c_547_n 0.0122883f $X=6.16 $Y=1.41 $X2=0 $Y2=0
cc_302 A2 N_Y_c_547_n 0.010804f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_303 N_A2_c_351_n N_Y_c_557_n 6.05689e-19 $X=7 $Y=1.295 $X2=0 $Y2=0
cc_304 A2 N_Y_c_557_n 0.0147558f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_305 N_A2_c_351_n N_Y_c_504_n 0.00332991f $X=7 $Y=1.295 $X2=0 $Y2=0
cc_306 N_A2_M1034_g N_Y_c_504_n 0.00188573f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A2_M1011_g N_Y_c_561_n 0.0123545f $X=6.58 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A2_c_351_n N_Y_c_561_n 5.47065e-19 $X=7 $Y=1.295 $X2=0 $Y2=0
cc_309 N_A2_M1034_g N_Y_c_561_n 0.00724892f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_310 A2 N_Y_c_561_n 0.0559298f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_311 N_A2_M1034_g N_VPWR_c_635_n 0.00644903f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A2_c_354_n N_VPWR_c_650_n 0.00539841f $X=5.74 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A2_c_357_n N_VPWR_c_650_n 0.00357835f $X=6.16 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A2_M1011_g N_VPWR_c_650_n 0.00357877f $X=6.58 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A2_M1034_g N_VPWR_c_650_n 0.00390837f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A2_c_354_n N_VPWR_c_628_n 0.00967497f $X=5.74 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A2_c_357_n N_VPWR_c_628_n 0.00522513f $X=6.16 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A2_M1011_g N_VPWR_c_628_n 0.00526405f $X=6.58 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A2_M1034_g N_VPWR_c_628_n 0.00695541f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A2_c_354_n N_A_1163_297#_c_786_n 0.0048829f $X=5.74 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A2_c_357_n N_A_1163_297#_c_786_n 0.00611592f $X=6.16 $Y=1.41 $X2=0
+ $Y2=0
cc_322 N_A2_M1011_g N_A_1163_297#_c_786_n 5.23146e-19 $X=6.58 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A2_c_357_n N_A_1163_297#_c_789_n 0.00864661f $X=6.16 $Y=1.41 $X2=0
+ $Y2=0
cc_324 N_A2_M1011_g N_A_1163_297#_c_789_n 0.0118936f $X=6.58 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A2_M1034_g N_A_1163_297#_c_789_n 0.00694404f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A2_c_354_n N_A_1163_297#_c_792_n 0.00235828f $X=5.74 $Y=1.41 $X2=0
+ $Y2=0
cc_327 N_A2_c_357_n N_A_1163_297#_c_792_n 7.72367e-19 $X=6.16 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_A2_M1034_g N_A_1163_297#_c_794_n 0.00892166f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A2_c_351_n N_A_1163_297#_c_785_n 5.99961e-19 $X=7 $Y=1.295 $X2=0 $Y2=0
cc_330 N_A2_M1034_g N_A_1163_297#_c_785_n 0.00776664f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A2_M1034_g N_A_1163_297#_c_797_n 0.00293267f $X=7 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A2_M1024_g N_A_445_47#_c_878_n 5.61217e-19 $X=6.055 $Y=0.56 $X2=0 $Y2=0
cc_333 N_A2_c_346_n N_A_803_47#_c_908_n 0.00691761f $X=5.815 $Y=1.335 $X2=0
+ $Y2=0
cc_334 N_A2_M1024_g N_A_803_47#_c_908_n 0.0136352f $X=6.055 $Y=0.56 $X2=0 $Y2=0
cc_335 N_A2_M1028_g N_A_803_47#_c_908_n 0.011851f $X=6.475 $Y=0.56 $X2=0 $Y2=0
cc_336 N_A2_M1029_g N_A_803_47#_c_908_n 0.011851f $X=6.915 $Y=0.56 $X2=0 $Y2=0
cc_337 N_A2_c_351_n N_A_803_47#_c_908_n 0.00768227f $X=7 $Y=1.295 $X2=0 $Y2=0
cc_338 N_A2_M1031_g N_A_803_47#_c_908_n 0.0130563f $X=7.335 $Y=0.56 $X2=0 $Y2=0
cc_339 A2 N_A_803_47#_c_908_n 0.0911818f $X=7.045 $Y=1.105 $X2=0 $Y2=0
cc_340 N_A2_M1024_g N_VGND_c_959_n 0.00982835f $X=6.055 $Y=0.56 $X2=0 $Y2=0
cc_341 N_A2_M1028_g N_VGND_c_959_n 0.00860636f $X=6.475 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A2_M1029_g N_VGND_c_959_n 0.00117244f $X=6.915 $Y=0.56 $X2=0 $Y2=0
cc_343 N_A2_M1028_g N_VGND_c_960_n 0.00117244f $X=6.475 $Y=0.56 $X2=0 $Y2=0
cc_344 N_A2_M1029_g N_VGND_c_960_n 0.00860636f $X=6.915 $Y=0.56 $X2=0 $Y2=0
cc_345 N_A2_M1031_g N_VGND_c_960_n 0.00864336f $X=7.335 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A2_M1031_g N_VGND_c_961_n 0.00117473f $X=7.335 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A2_M1024_g N_VGND_c_965_n 0.00341689f $X=6.055 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A2_M1028_g N_VGND_c_966_n 0.00341689f $X=6.475 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A2_M1029_g N_VGND_c_966_n 0.00341689f $X=6.915 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A2_M1031_g N_VGND_c_967_n 0.00341689f $X=7.335 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A2_M1024_g N_VGND_c_969_n 0.00411722f $X=6.055 $Y=0.56 $X2=0 $Y2=0
cc_352 N_A2_M1028_g N_VGND_c_969_n 0.00408046f $X=6.475 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A2_M1029_g N_VGND_c_969_n 0.00408046f $X=6.915 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A2_M1031_g N_VGND_c_969_n 0.00411722f $X=7.335 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A1_M1000_g N_Y_c_504_n 0.00367431f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_356 N_A1_M1000_g N_VPWR_c_635_n 0.00804316f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_357 N_A1_M1004_g N_VPWR_c_635_n 5.22478e-19 $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_358 N_A1_M1000_g N_VPWR_c_636_n 5.53443e-19 $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_359 N_A1_M1004_g N_VPWR_c_636_n 0.00962936f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A1_M1019_g N_VPWR_c_636_n 0.0104779f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A1_M1035_g N_VPWR_c_636_n 6.31999e-19 $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A1_M1035_g N_VPWR_c_638_n 0.00889532f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_363 A1 N_VPWR_c_638_n 0.0216047f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_364 N_A1_M1000_g N_VPWR_c_651_n 0.00342263f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_365 N_A1_M1004_g N_VPWR_c_651_n 0.00525069f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A1_M1019_g N_VPWR_c_652_n 0.00486043f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A1_M1035_g N_VPWR_c_652_n 0.00583607f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A1_M1000_g N_VPWR_c_628_n 0.00399267f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A1_M1004_g N_VPWR_c_628_n 0.0088132f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_370 N_A1_M1019_g N_VPWR_c_628_n 0.00819893f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_371 N_A1_M1035_g N_VPWR_c_628_n 0.0113526f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_372 N_A1_M1000_g N_A_1163_297#_c_785_n 0.0134891f $X=7.93 $Y=1.985 $X2=0
+ $Y2=0
cc_373 A1 N_A_1163_297#_c_785_n 0.0053397f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_374 N_A1_c_443_n N_A_1163_297#_c_785_n 0.00282451f $X=9.19 $Y=1.16 $X2=0
+ $Y2=0
cc_375 N_A1_M1004_g N_A_1163_297#_c_801_n 0.0140639f $X=8.35 $Y=1.985 $X2=0
+ $Y2=0
cc_376 N_A1_M1019_g N_A_1163_297#_c_801_n 0.0137743f $X=8.77 $Y=1.985 $X2=0
+ $Y2=0
cc_377 A1 N_A_1163_297#_c_801_n 0.0544992f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_378 N_A1_c_443_n N_A_1163_297#_c_801_n 0.00117541f $X=9.19 $Y=1.16 $X2=0
+ $Y2=0
cc_379 A1 N_A_1163_297#_c_805_n 0.0143788f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_380 N_A1_c_443_n N_A_1163_297#_c_805_n 6.23984e-19 $X=9.19 $Y=1.16 $X2=0
+ $Y2=0
cc_381 N_A1_M1005_g N_A_803_47#_c_908_n 0.0151591f $X=7.78 $Y=0.56 $X2=0 $Y2=0
cc_382 N_A1_M1006_g N_A_803_47#_c_908_n 0.0118378f $X=8.2 $Y=0.56 $X2=0 $Y2=0
cc_383 N_A1_M1012_g N_A_803_47#_c_908_n 0.0118378f $X=8.62 $Y=0.56 $X2=0 $Y2=0
cc_384 N_A1_M1018_g N_A_803_47#_c_908_n 0.0119986f $X=9.04 $Y=0.56 $X2=0 $Y2=0
cc_385 A1 N_A_803_47#_c_908_n 0.122197f $X=9.345 $Y=1.105 $X2=0 $Y2=0
cc_386 N_A1_c_443_n N_A_803_47#_c_908_n 0.0119451f $X=9.19 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A1_M1005_g N_VGND_c_960_n 0.00117473f $X=7.78 $Y=0.56 $X2=0 $Y2=0
cc_388 N_A1_M1005_g N_VGND_c_961_n 0.00864336f $X=7.78 $Y=0.56 $X2=0 $Y2=0
cc_389 N_A1_M1006_g N_VGND_c_961_n 0.00845732f $X=8.2 $Y=0.56 $X2=0 $Y2=0
cc_390 N_A1_M1012_g N_VGND_c_961_n 0.00116151f $X=8.62 $Y=0.56 $X2=0 $Y2=0
cc_391 N_A1_M1006_g N_VGND_c_962_n 0.00116151f $X=8.2 $Y=0.56 $X2=0 $Y2=0
cc_392 N_A1_M1012_g N_VGND_c_962_n 0.00845732f $X=8.62 $Y=0.56 $X2=0 $Y2=0
cc_393 N_A1_M1018_g N_VGND_c_962_n 0.0161007f $X=9.04 $Y=0.56 $X2=0 $Y2=0
cc_394 N_A1_M1006_g N_VGND_c_963_n 0.00341689f $X=8.2 $Y=0.56 $X2=0 $Y2=0
cc_395 N_A1_M1012_g N_VGND_c_963_n 0.00341689f $X=8.62 $Y=0.56 $X2=0 $Y2=0
cc_396 N_A1_M1005_g N_VGND_c_967_n 0.00341689f $X=7.78 $Y=0.56 $X2=0 $Y2=0
cc_397 N_A1_M1018_g N_VGND_c_968_n 0.00341689f $X=9.04 $Y=0.56 $X2=0 $Y2=0
cc_398 N_A1_M1005_g N_VGND_c_969_n 0.00411722f $X=7.78 $Y=0.56 $X2=0 $Y2=0
cc_399 N_A1_M1006_g N_VGND_c_969_n 0.0040262f $X=8.2 $Y=0.56 $X2=0 $Y2=0
cc_400 N_A1_M1012_g N_VGND_c_969_n 0.0040262f $X=8.62 $Y=0.56 $X2=0 $Y2=0
cc_401 N_A1_M1018_g N_VGND_c_969_n 0.00513758f $X=9.04 $Y=0.56 $X2=0 $Y2=0
cc_402 N_Y_c_514_n N_VPWR_M1003_d 0.00310556f $X=1.015 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_403 N_Y_c_518_n N_VPWR_M1025_d 0.00310556f $X=1.845 $Y=1.6 $X2=0 $Y2=0
cc_404 N_Y_c_526_n N_VPWR_M1001_d 0.00312854f $X=2.685 $Y=1.6 $X2=0 $Y2=0
cc_405 N_Y_c_530_n N_VPWR_M1030_d 0.00312854f $X=3.525 $Y=1.6 $X2=0 $Y2=0
cc_406 N_Y_c_539_n N_VPWR_M1007_d 0.00312854f $X=4.57 $Y=1.6 $X2=0 $Y2=0
cc_407 N_Y_c_543_n N_VPWR_M1015_d 0.00312854f $X=5.41 $Y=1.6 $X2=0 $Y2=0
cc_408 N_Y_c_514_n N_VPWR_c_629_n 0.0158832f $X=1.015 $Y=1.6 $X2=0 $Y2=0
cc_409 N_Y_c_518_n N_VPWR_c_630_n 0.0140971f $X=1.845 $Y=1.6 $X2=0 $Y2=0
cc_410 N_Y_c_526_n N_VPWR_c_631_n 0.0155023f $X=2.685 $Y=1.6 $X2=0 $Y2=0
cc_411 N_Y_c_530_n N_VPWR_c_632_n 0.0155023f $X=3.525 $Y=1.6 $X2=0 $Y2=0
cc_412 N_Y_c_538_n N_VPWR_c_633_n 0.0254721f $X=3.62 $Y=1.96 $X2=0 $Y2=0
cc_413 N_Y_c_539_n N_VPWR_c_633_n 0.016645f $X=4.57 $Y=1.6 $X2=0 $Y2=0
cc_414 N_Y_c_543_n N_VPWR_c_634_n 0.0140971f $X=5.41 $Y=1.6 $X2=0 $Y2=0
cc_415 N_Y_c_579_p N_VPWR_c_639_n 0.0117506f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_416 N_Y_c_580_p N_VPWR_c_641_n 0.0121054f $X=1.94 $Y=1.96 $X2=0 $Y2=0
cc_417 N_Y_c_581_p N_VPWR_c_643_n 0.0121054f $X=2.78 $Y=1.96 $X2=0 $Y2=0
cc_418 N_Y_c_538_n N_VPWR_c_645_n 0.0126629f $X=3.62 $Y=1.96 $X2=0 $Y2=0
cc_419 N_Y_c_583_p N_VPWR_c_647_n 0.0121054f $X=4.665 $Y=1.96 $X2=0 $Y2=0
cc_420 Y N_VPWR_c_649_n 0.0185333f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_421 N_Y_c_552_n N_VPWR_c_650_n 0.0126629f $X=5.505 $Y=1.96 $X2=0 $Y2=0
cc_422 N_Y_M1003_s N_VPWR_c_628_n 0.00330824f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_423 N_Y_M1009_s N_VPWR_c_628_n 0.00527642f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_424 N_Y_M1036_s N_VPWR_c_628_n 0.00492927f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_425 N_Y_M1010_s N_VPWR_c_628_n 0.00492927f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_426 N_Y_M1037_s N_VPWR_c_628_n 0.0137542f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_427 N_Y_M1013_s N_VPWR_c_628_n 0.00492927f $X=4.53 $Y=1.485 $X2=0 $Y2=0
cc_428 N_Y_M1038_s N_VPWR_c_628_n 0.00599791f $X=5.37 $Y=1.485 $X2=0 $Y2=0
cc_429 N_Y_M1008_d N_VPWR_c_628_n 0.00216833f $X=6.235 $Y=1.485 $X2=0 $Y2=0
cc_430 N_Y_M1034_d N_VPWR_c_628_n 0.003022f $X=7.075 $Y=1.485 $X2=0 $Y2=0
cc_431 N_Y_c_579_p N_VPWR_c_628_n 0.00685509f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_432 N_Y_c_580_p N_VPWR_c_628_n 0.00724021f $X=1.94 $Y=1.96 $X2=0 $Y2=0
cc_433 N_Y_c_581_p N_VPWR_c_628_n 0.00724021f $X=2.78 $Y=1.96 $X2=0 $Y2=0
cc_434 N_Y_c_538_n N_VPWR_c_628_n 0.00724021f $X=3.62 $Y=1.96 $X2=0 $Y2=0
cc_435 N_Y_c_583_p N_VPWR_c_628_n 0.00724021f $X=4.665 $Y=1.96 $X2=0 $Y2=0
cc_436 N_Y_c_552_n N_VPWR_c_628_n 0.00724021f $X=5.505 $Y=1.96 $X2=0 $Y2=0
cc_437 Y N_VPWR_c_628_n 0.0105137f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_438 N_Y_c_547_n N_A_1163_297#_M1002_s 0.00423749f $X=6.285 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_439 N_Y_c_561_n N_A_1163_297#_M1011_s 0.00326792f $X=7.045 $Y=1.617 $X2=0
+ $Y2=0
cc_440 N_Y_c_552_n N_A_1163_297#_c_786_n 0.0289069f $X=5.505 $Y=1.96 $X2=0 $Y2=0
cc_441 N_Y_c_547_n N_A_1163_297#_c_786_n 0.0168753f $X=6.285 $Y=1.6 $X2=0 $Y2=0
cc_442 N_Y_M1008_d N_A_1163_297#_c_789_n 0.00313673f $X=6.235 $Y=1.485 $X2=0
+ $Y2=0
cc_443 N_Y_c_547_n N_A_1163_297#_c_789_n 0.00295233f $X=6.285 $Y=1.6 $X2=0 $Y2=0
cc_444 N_Y_c_608_p N_A_1163_297#_c_789_n 0.0119291f $X=6.37 $Y=1.935 $X2=0 $Y2=0
cc_445 N_Y_c_561_n N_A_1163_297#_c_789_n 0.00369353f $X=7.045 $Y=1.617 $X2=0
+ $Y2=0
cc_446 N_Y_c_552_n N_A_1163_297#_c_792_n 0.0144619f $X=5.505 $Y=1.96 $X2=0 $Y2=0
cc_447 N_Y_M1034_d N_A_1163_297#_c_785_n 0.00599172f $X=7.075 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_Y_c_504_n N_A_1163_297#_c_785_n 0.0211973f $X=7.21 $Y=1.63 $X2=0 $Y2=0
cc_449 N_Y_c_561_n N_A_1163_297#_c_785_n 0.00227568f $X=7.045 $Y=1.617 $X2=0
+ $Y2=0
cc_450 N_Y_c_561_n N_A_1163_297#_c_797_n 0.0160594f $X=7.045 $Y=1.617 $X2=0
+ $Y2=0
cc_451 N_Y_c_502_n N_A_27_47#_M1016_d 0.00292289f $X=0.23 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_452 Y N_A_27_47#_M1016_d 3.05534e-19 $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_453 N_Y_c_508_n N_A_27_47#_M1020_d 0.00335926f $X=1.52 $Y=0.73 $X2=0 $Y2=0
cc_454 N_Y_M1016_s N_A_27_47#_c_842_n 0.00314262f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_455 N_Y_M1023_s N_A_27_47#_c_842_n 0.00314262f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_456 N_Y_c_508_n N_A_27_47#_c_842_n 0.0635866f $X=1.52 $Y=0.73 $X2=0 $Y2=0
cc_457 N_Y_c_502_n N_A_27_47#_c_842_n 0.0189726f $X=0.23 $Y=0.815 $X2=0 $Y2=0
cc_458 N_Y_c_547_n N_A_803_47#_c_908_n 0.0118232f $X=6.285 $Y=1.6 $X2=0 $Y2=0
cc_459 N_Y_c_550_n N_A_803_47#_c_908_n 0.00461686f $X=5.505 $Y=1.6 $X2=0 $Y2=0
cc_460 N_Y_c_504_n N_A_803_47#_c_908_n 0.00182057f $X=7.21 $Y=1.63 $X2=0 $Y2=0
cc_461 N_Y_M1016_s N_VGND_c_969_n 0.00218391f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_462 N_Y_M1023_s N_VGND_c_969_n 0.00218391f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_463 N_Y_c_502_n N_VGND_c_969_n 0.00100009f $X=0.23 $Y=0.815 $X2=0 $Y2=0
cc_464 N_VPWR_c_628_n N_A_1163_297#_M1002_s 0.00215201f $X=9.43 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_465 N_VPWR_c_628_n N_A_1163_297#_M1011_s 0.00216812f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_628_n N_A_1163_297#_M1000_s 0.003729f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_628_n N_A_1163_297#_M1019_s 0.00492927f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_635_n N_A_1163_297#_c_789_n 0.00671917f $X=7.72 $Y=2.34 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_650_n N_A_1163_297#_c_789_n 0.0509939f $X=7.555 $Y=2.72 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_628_n N_A_1163_297#_c_789_n 0.0319402f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_650_n N_A_1163_297#_c_792_n 0.0189234f $X=7.555 $Y=2.72 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_628_n N_A_1163_297#_c_792_n 0.0122542f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_635_n N_A_1163_297#_c_794_n 0.00128672f $X=7.72 $Y=2.34 $X2=0
+ $Y2=0
cc_474 N_VPWR_M1000_d N_A_1163_297#_c_785_n 0.00800195f $X=7.595 $Y=2.2 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_635_n N_A_1163_297#_c_785_n 0.0207773f $X=7.72 $Y=2.34 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_650_n N_A_1163_297#_c_785_n 0.00877686f $X=7.555 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_651_n N_A_1163_297#_c_785_n 0.00220527f $X=8.41 $Y=2.72 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_628_n N_A_1163_297#_c_785_n 0.0201752f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_651_n N_A_1163_297#_c_835_n 0.0117506f $X=8.41 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_628_n N_A_1163_297#_c_835_n 0.00685509f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_481 N_VPWR_M1004_d N_A_1163_297#_c_801_n 0.0031455f $X=8.425 $Y=1.485 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_636_n N_A_1163_297#_c_801_n 0.0155023f $X=8.56 $Y=2.02 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_652_n N_A_1163_297#_c_839_n 0.0121054f $X=9.265 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_628_n N_A_1163_297#_c_839_n 0.00724021f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_628_n N_A_1163_297#_c_841_n 2.92335e-19 $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_843_n N_A_445_47#_M1021_d 0.00333793f $X=3.62 $Y=0.7
+ $X2=-0.19 $Y2=-0.24
cc_487 N_A_27_47#_c_843_n N_A_445_47#_M1032_d 0.00333793f $X=3.62 $Y=0.7 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_M1026_s N_A_445_47#_c_878_n 0.00305132f $X=2.645 $Y=0.235
+ $X2=0 $Y2=0
cc_489 N_A_27_47#_M1033_s N_A_445_47#_c_878_n 0.00491625f $X=3.485 $Y=0.235
+ $X2=0 $Y2=0
cc_490 N_A_27_47#_c_843_n N_A_445_47#_c_878_n 0.0814f $X=3.62 $Y=0.7 $X2=0 $Y2=0
cc_491 N_A_27_47#_c_843_n N_A_803_47#_c_908_n 0.0145425f $X=3.62 $Y=0.7 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_842_n N_VGND_c_965_n 0.092203f $X=1.855 $Y=0.38 $X2=0 $Y2=0
cc_493 N_A_27_47#_c_843_n N_VGND_c_965_n 0.00259391f $X=3.62 $Y=0.7 $X2=0 $Y2=0
cc_494 N_A_27_47#_M1016_d N_VGND_c_969_n 0.00210839f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_M1020_d N_VGND_c_969_n 0.00216774f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_M1039_d N_VGND_c_969_n 0.00234859f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_M1026_s N_VGND_c_969_n 0.00216833f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_M1033_s N_VGND_c_969_n 0.00210147f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_842_n N_VGND_c_969_n 0.0679534f $X=1.855 $Y=0.38 $X2=0 $Y2=0
cc_500 N_A_27_47#_c_843_n N_VGND_c_969_n 0.00745687f $X=3.62 $Y=0.7 $X2=0 $Y2=0
cc_501 N_A_445_47#_c_878_n N_A_803_47#_M1014_s 0.00489431f $X=5.4 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_502 N_A_445_47#_c_878_n N_A_803_47#_M1017_s 0.003196f $X=5.4 $Y=0.36 $X2=0
+ $Y2=0
cc_503 N_A_445_47#_M1014_d N_A_803_47#_c_908_n 0.00177239f $X=4.425 $Y=0.235
+ $X2=0 $Y2=0
cc_504 N_A_445_47#_M1022_d N_A_803_47#_c_908_n 0.00177239f $X=5.265 $Y=0.235
+ $X2=0 $Y2=0
cc_505 N_A_445_47#_c_878_n N_A_803_47#_c_908_n 0.0686747f $X=5.4 $Y=0.36 $X2=0
+ $Y2=0
cc_506 N_A_445_47#_c_878_n N_VGND_c_959_n 0.00584613f $X=5.4 $Y=0.36 $X2=0 $Y2=0
cc_507 N_A_445_47#_c_878_n N_VGND_c_965_n 0.190659f $X=5.4 $Y=0.36 $X2=0 $Y2=0
cc_508 N_A_445_47#_M1021_d N_VGND_c_969_n 0.00215227f $X=2.225 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_445_47#_M1032_d N_VGND_c_969_n 0.00215227f $X=3.065 $Y=0.235 $X2=0
+ $Y2=0
cc_510 N_A_445_47#_M1014_d N_VGND_c_969_n 0.00215227f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_511 N_A_445_47#_M1022_d N_VGND_c_969_n 0.00215227f $X=5.265 $Y=0.235 $X2=0
+ $Y2=0
cc_512 N_A_445_47#_c_878_n N_VGND_c_969_n 0.120885f $X=5.4 $Y=0.36 $X2=0 $Y2=0
cc_513 N_A_803_47#_c_908_n N_VGND_M1024_s 0.00162029f $X=9.25 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_514 N_A_803_47#_c_908_n N_VGND_M1029_s 0.00162029f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_803_47#_c_908_n N_VGND_M1005_d 0.00162029f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_516 N_A_803_47#_c_908_n N_VGND_M1012_d 0.00162029f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_517 N_A_803_47#_c_908_n N_VGND_c_959_n 0.0164771f $X=9.25 $Y=0.74 $X2=0 $Y2=0
cc_518 N_A_803_47#_c_908_n N_VGND_c_960_n 0.0164771f $X=9.25 $Y=0.74 $X2=0 $Y2=0
cc_519 N_A_803_47#_c_908_n N_VGND_c_961_n 0.0164771f $X=9.25 $Y=0.74 $X2=0 $Y2=0
cc_520 N_A_803_47#_c_908_n N_VGND_c_962_n 0.0164771f $X=9.25 $Y=0.74 $X2=0 $Y2=0
cc_521 N_A_803_47#_c_908_n N_VGND_c_963_n 0.00755316f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_522 N_A_803_47#_c_908_n N_VGND_c_965_n 0.00799243f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_523 N_A_803_47#_c_908_n N_VGND_c_966_n 0.00789715f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_524 N_A_803_47#_c_908_n N_VGND_c_967_n 0.00798315f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_525 N_A_803_47#_c_908_n N_VGND_c_968_n 0.00707734f $X=9.25 $Y=0.74 $X2=0
+ $Y2=0
cc_526 N_A_803_47#_M1014_s N_VGND_c_969_n 0.00210147f $X=4.015 $Y=0.235 $X2=0
+ $Y2=0
cc_527 N_A_803_47#_M1017_s N_VGND_c_969_n 0.00216833f $X=4.845 $Y=0.235 $X2=0
+ $Y2=0
cc_528 N_A_803_47#_M1027_s N_VGND_c_969_n 0.00353055f $X=5.685 $Y=0.235 $X2=0
+ $Y2=0
cc_529 N_A_803_47#_M1028_d N_VGND_c_969_n 0.00347071f $X=6.55 $Y=0.235 $X2=0
+ $Y2=0
cc_530 N_A_803_47#_M1031_d N_VGND_c_969_n 0.00353055f $X=7.41 $Y=0.235 $X2=0
+ $Y2=0
cc_531 N_A_803_47#_M1006_s N_VGND_c_969_n 0.00323135f $X=8.275 $Y=0.235 $X2=0
+ $Y2=0
cc_532 N_A_803_47#_M1018_s N_VGND_c_969_n 0.00342852f $X=9.115 $Y=0.235 $X2=0
+ $Y2=0
cc_533 N_A_803_47#_c_908_n N_VGND_c_969_n 0.0765513f $X=9.25 $Y=0.74 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.65e+11p pd=2.73e+06u as=6.118e+11p ps=4.51e+06u
M1001 a_421_47# B a_27_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.226e+11p ps=2.74e+06u
M1002 VGND C a_421_47# VNB nshort w=420000u l=150000u
+  ad=4.082e+11p pd=3.81e+06u as=0p ps=0u
M1003 a_265_341# A VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_27_47# B a_265_341# VPB phighvt w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=0p ps=0u
M1005 VGND A a_109_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 VPWR A a_109_341# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_265_47# A VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_27_47# B a_265_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.3725e+11p pd=2.03e+06u as=0p ps=0u
M1010 a_109_341# C a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_421_341# B a_27_47# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1012 VPWR C a_421_341# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_109_47# C a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

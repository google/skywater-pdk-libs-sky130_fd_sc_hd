* File: sky130_fd_sc_hd__a41oi_4.pxi.spice
* Created: Thu Aug 27 14:06:35 2020
* 
x_PM_SKY130_FD_SC_HD__A41OI_4%B1 N_B1_c_109_n N_B1_M1021_g N_B1_M1005_g
+ N_B1_c_110_n N_B1_M1024_g N_B1_M1013_g N_B1_c_111_n N_B1_M1025_g N_B1_M1026_g
+ N_B1_c_112_n N_B1_M1036_g N_B1_M1035_g B1 B1 B1 B1 B1 B1 N_B1_c_113_n
+ N_B1_c_114_n PM_SKY130_FD_SC_HD__A41OI_4%B1
x_PM_SKY130_FD_SC_HD__A41OI_4%A1 N_A1_M1002_g N_A1_c_188_n N_A1_M1003_g
+ N_A1_c_189_n N_A1_M1004_g N_A1_M1018_g N_A1_c_190_n N_A1_M1009_g N_A1_M1022_g
+ N_A1_c_191_n N_A1_M1012_g N_A1_M1030_g A1 A1 A1 A1 N_A1_c_192_n N_A1_c_193_n
+ PM_SKY130_FD_SC_HD__A41OI_4%A1
x_PM_SKY130_FD_SC_HD__A41OI_4%A2 N_A2_c_260_n N_A2_M1006_g N_A2_M1014_g
+ N_A2_c_261_n N_A2_M1010_g N_A2_M1017_g N_A2_c_262_n N_A2_M1011_g N_A2_M1019_g
+ N_A2_c_263_n N_A2_M1039_g N_A2_M1028_g N_A2_c_264_n A2 A2 A2 A2 N_A2_c_266_n
+ PM_SKY130_FD_SC_HD__A41OI_4%A2
x_PM_SKY130_FD_SC_HD__A41OI_4%A3 N_A3_c_332_n N_A3_M1000_g N_A3_M1007_g
+ N_A3_c_333_n N_A3_M1029_g N_A3_M1027_g N_A3_c_334_n N_A3_M1033_g N_A3_M1031_g
+ N_A3_c_335_n N_A3_M1034_g N_A3_M1037_g A3 A3 A3 N_A3_c_336_n
+ PM_SKY130_FD_SC_HD__A41OI_4%A3
x_PM_SKY130_FD_SC_HD__A41OI_4%A4 N_A4_c_397_n N_A4_M1001_g N_A4_M1015_g
+ N_A4_c_398_n N_A4_M1008_g N_A4_M1020_g N_A4_c_399_n N_A4_M1016_g N_A4_M1023_g
+ N_A4_c_400_n N_A4_M1038_g N_A4_M1032_g A4 A4 A4 A4 N_A4_c_402_n
+ PM_SKY130_FD_SC_HD__A41OI_4%A4
x_PM_SKY130_FD_SC_HD__A41OI_4%A_27_297# N_A_27_297#_M1005_s N_A_27_297#_M1013_s
+ N_A_27_297#_M1035_s N_A_27_297#_M1018_d N_A_27_297#_M1030_d
+ N_A_27_297#_M1017_s N_A_27_297#_M1028_s N_A_27_297#_M1027_s
+ N_A_27_297#_M1037_s N_A_27_297#_M1020_d N_A_27_297#_M1032_d
+ N_A_27_297#_c_464_n N_A_27_297#_c_471_n N_A_27_297#_c_473_n
+ N_A_27_297#_c_472_n N_A_27_297#_c_551_p N_A_27_297#_c_477_n
+ N_A_27_297#_c_481_n N_A_27_297#_c_484_n N_A_27_297#_c_485_n
+ N_A_27_297#_c_553_p N_A_27_297#_c_489_n N_A_27_297#_c_493_n
+ N_A_27_297#_c_496_n N_A_27_297#_c_544_p N_A_27_297#_c_500_n
+ N_A_27_297#_c_554_p N_A_27_297#_c_506_n N_A_27_297#_c_555_p
+ N_A_27_297#_c_510_n N_A_27_297#_c_514_n N_A_27_297#_c_483_n
+ N_A_27_297#_c_494_n N_A_27_297#_c_504_n N_A_27_297#_c_515_n
+ PM_SKY130_FD_SC_HD__A41OI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A41OI_4%Y N_Y_M1021_s N_Y_M1025_s N_Y_M1003_d N_Y_M1009_d
+ N_Y_M1005_d N_Y_M1026_d N_Y_c_650_p N_Y_c_587_n N_Y_c_591_n N_Y_c_593_n
+ N_Y_c_653_p N_Y_c_597_n N_Y_c_599_n N_Y_c_601_n N_Y_c_607_n N_Y_c_612_n Y Y Y
+ N_Y_c_617_n Y N_Y_c_585_n PM_SKY130_FD_SC_HD__A41OI_4%Y
x_PM_SKY130_FD_SC_HD__A41OI_4%VPWR N_VPWR_M1002_s N_VPWR_M1022_s N_VPWR_M1014_d
+ N_VPWR_M1019_d N_VPWR_M1007_d N_VPWR_M1031_d N_VPWR_M1015_s N_VPWR_M1023_s
+ N_VPWR_c_674_n N_VPWR_c_675_n N_VPWR_c_676_n N_VPWR_c_677_n N_VPWR_c_678_n
+ N_VPWR_c_679_n N_VPWR_c_680_n N_VPWR_c_681_n N_VPWR_c_682_n N_VPWR_c_683_n
+ VPWR N_VPWR_c_684_n N_VPWR_c_685_n N_VPWR_c_686_n N_VPWR_c_687_n
+ N_VPWR_c_688_n N_VPWR_c_689_n N_VPWR_c_673_n N_VPWR_c_691_n N_VPWR_c_692_n
+ N_VPWR_c_693_n N_VPWR_c_694_n N_VPWR_c_695_n N_VPWR_c_696_n N_VPWR_c_697_n
+ N_VPWR_c_698_n PM_SKY130_FD_SC_HD__A41OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A41OI_4%VGND N_VGND_M1021_d N_VGND_M1024_d N_VGND_M1036_d
+ N_VGND_M1001_d N_VGND_M1016_d N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n
+ N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n VGND N_VGND_c_829_n
+ N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n
+ N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n
+ PM_SKY130_FD_SC_HD__A41OI_4%VGND
x_PM_SKY130_FD_SC_HD__A41OI_4%A_493_47# N_A_493_47#_M1003_s N_A_493_47#_M1004_s
+ N_A_493_47#_M1012_s N_A_493_47#_M1010_d N_A_493_47#_M1039_d
+ N_A_493_47#_c_959_n PM_SKY130_FD_SC_HD__A41OI_4%A_493_47#
x_PM_SKY130_FD_SC_HD__A41OI_4%A_911_47# N_A_911_47#_M1006_s N_A_911_47#_M1011_s
+ N_A_911_47#_M1000_s N_A_911_47#_M1033_s N_A_911_47#_c_989_n
+ PM_SKY130_FD_SC_HD__A41OI_4%A_911_47#
x_PM_SKY130_FD_SC_HD__A41OI_4%A_1269_47# N_A_1269_47#_M1000_d
+ N_A_1269_47#_M1029_d N_A_1269_47#_M1034_d N_A_1269_47#_M1008_s
+ N_A_1269_47#_M1038_s N_A_1269_47#_c_1020_n N_A_1269_47#_c_1043_n
+ N_A_1269_47#_c_1026_n N_A_1269_47#_c_1050_n N_A_1269_47#_c_1030_n
+ N_A_1269_47#_c_1057_n N_A_1269_47#_c_1034_n
+ PM_SKY130_FD_SC_HD__A41OI_4%A_1269_47#
cc_1 VNB N_B1_c_109_n 0.0210871f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B1_c_110_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_B1_c_111_n 0.0157754f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_B1_c_112_n 0.0183349f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_B1_c_113_n 0.0908217f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_6 VNB N_B1_c_114_n 0.00936732f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.305
cc_7 VNB N_A1_c_188_n 0.0200763f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_8 VNB N_A1_c_189_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_9 VNB N_A1_c_190_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_10 VNB N_A1_c_191_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_11 VNB N_A1_c_192_n 0.00618292f $X=-0.19 $Y=-0.24 $X2=1.29 $Y2=1.16
cc_12 VNB N_A1_c_193_n 0.0836799f $X=-0.19 $Y=-0.24 $X2=1.29 $Y2=1.16
cc_13 VNB N_A2_c_260_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_A2_c_261_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_15 VNB N_A2_c_262_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_16 VNB N_A2_c_263_n 0.0231822f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_17 VNB N_A2_c_264_n 0.0330109f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB A2 0.00294247f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_19 VNB N_A2_c_266_n 0.0577905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A3_c_332_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_21 VNB N_A3_c_333_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_22 VNB N_A3_c_334_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_23 VNB N_A3_c_335_n 0.0807748f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_24 VNB N_A3_c_336_n 0.0026648f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_25 VNB N_A4_c_397_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_26 VNB N_A4_c_398_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_27 VNB N_A4_c_399_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_28 VNB N_A4_c_400_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_29 VNB A4 0.00991795f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_30 VNB N_A4_c_402_n 0.0864272f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_31 VNB Y 0.00155789f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_32 VNB Y 0.0114849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_585_n 0.0140847f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.19
cc_34 VNB N_VPWR_c_673_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_823_n 0.0102396f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_36 VNB N_VGND_c_824_n 0.0125153f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_37 VNB N_VGND_c_825_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_38 VNB N_VGND_c_826_n 0.00595785f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_39 VNB N_VGND_c_827_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_40 VNB N_VGND_c_828_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.105
cc_41 VNB N_VGND_c_829_n 0.0117278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_830_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_43 VNB N_VGND_c_831_n 0.147433f $X=-0.19 $Y=-0.24 $X2=1.29 $Y2=1.16
cc_44 VNB N_VGND_c_832_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_833_n 0.0160953f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.19
cc_46 VNB N_VGND_c_834_n 0.474451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_835_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_836_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_837_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_838_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_493_47#_c_959_n 0.00458763f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_52 VNB N_A_911_47#_c_989_n 0.00752337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1269_47#_c_1020_n 0.00216865f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_54 VPB N_B1_M1005_g 0.0218926f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_55 VPB N_B1_M1013_g 0.0185005f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_56 VPB N_B1_M1026_g 0.0185026f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_57 VPB N_B1_M1035_g 0.0214243f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_58 VPB B1 0.0258766f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_59 VPB N_B1_c_113_n 0.0205513f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_60 VPB N_A1_M1002_g 0.0243318f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_61 VPB N_A1_M1018_g 0.0213644f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_A1_M1022_g 0.0182793f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_63 VPB N_A1_M1030_g 0.0195536f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_64 VPB N_A1_c_192_n 0.00113006f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.16
cc_65 VPB N_A1_c_193_n 0.0234857f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.16
cc_66 VPB N_A2_M1014_g 0.018515f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_A2_M1017_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_A2_M1019_g 0.0208556f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_69 VPB N_A2_M1028_g 0.0213369f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_70 VPB N_A2_c_264_n 0.00944193f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_71 VPB N_A2_c_266_n 0.0206066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A3_M1007_g 0.017785f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_73 VPB N_A3_M1027_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_74 VPB N_A3_M1031_g 0.0172788f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_75 VPB N_A3_c_335_n 0.0143946f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_76 VPB N_A3_M1037_g 0.0175748f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_77 VPB N_A4_M1015_g 0.0186099f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_78 VPB N_A4_M1020_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_79 VPB N_A4_M1023_g 0.0182793f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_80 VPB N_A4_M1032_g 0.025757f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_81 VPB N_A4_c_402_n 0.0192357f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_82 VPB N_A_27_297#_c_464_n 0.00834107f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.105
cc_83 VPB Y 0.00468314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_674_n 3.17813e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_85 VPB N_VPWR_c_675_n 3.24351e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.785
cc_86 VPB N_VPWR_c_676_n 0.00614692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_677_n 3.10683e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_678_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_89 VPB N_VPWR_c_679_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_90 VPB N_VPWR_c_680_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_91 VPB N_VPWR_c_681_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_682_n 0.0151294f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_683_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_684_n 0.0117367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_685_n 0.0156335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_686_n 0.0146009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_687_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_688_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_689_n 0.016859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_673_n 0.046594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_691_n 0.0604518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_692_n 0.0121667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_693_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_694_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_695_n 0.0128614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_696_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_697_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_698_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 N_B1_M1035_g N_A1_M1002_g 0.011481f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_110 N_B1_c_113_n N_A1_c_193_n 0.011481f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_111 B1 N_A_27_297#_M1005_s 0.0119908f $X=0.145 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_112 N_B1_M1005_g N_A_27_297#_c_464_n 0.0115553f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B1_M1013_g N_A_27_297#_c_464_n 0.00922647f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B1_M1026_g N_A_27_297#_c_464_n 0.00916955f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B1_M1035_g N_A_27_297#_c_464_n 0.0125354f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_116 B1 N_A_27_297#_c_464_n 0.0107018f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_117 N_B1_M1035_g N_A_27_297#_c_471_n 0.0039689f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_118 N_B1_M1035_g N_A_27_297#_c_472_n 0.00166962f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B1_c_110_n N_Y_c_587_n 0.0115547f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B1_c_111_n N_Y_c_587_n 0.0117424f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_121 B1 N_Y_c_587_n 0.0274913f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B1_c_113_n N_Y_c_587_n 0.00207061f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_123 B1 N_Y_c_591_n 0.0090006f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B1_c_113_n N_Y_c_591_n 0.00216182f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B1_M1013_g N_Y_c_593_n 0.00889401f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B1_M1026_g N_Y_c_593_n 0.008602f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_127 B1 N_Y_c_593_n 0.0218748f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_128 N_B1_c_113_n N_Y_c_593_n 0.00192838f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B1_c_112_n N_Y_c_597_n 0.0154902f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_130 B1 N_Y_c_597_n 0.00554203f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B1_M1035_g N_Y_c_599_n 0.0119035f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_132 B1 N_Y_c_599_n 0.00380918f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B1_M1005_g N_Y_c_601_n 0.0106465f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_134 N_B1_M1013_g N_Y_c_601_n 0.00724625f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B1_M1026_g N_Y_c_601_n 9.94965e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_136 B1 N_Y_c_601_n 0.0276407f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_137 B1 N_Y_c_601_n 0.0144995f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_138 N_B1_c_113_n N_Y_c_601_n 0.00200399f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B1_M1013_g N_Y_c_607_n 0.00140055f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B1_M1026_g N_Y_c_607_n 0.0091312f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B1_M1035_g N_Y_c_607_n 0.0131793f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_142 B1 N_Y_c_607_n 0.0196107f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_143 N_B1_c_113_n N_Y_c_607_n 0.00211284f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_144 B1 N_Y_c_612_n 0.0090006f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_145 N_B1_c_113_n N_Y_c_612_n 0.00216182f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B1_c_112_n Y 0.0170836f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_147 B1 Y 0.0170614f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_148 N_B1_M1005_g N_VPWR_c_673_n 0.00619429f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B1_M1013_g N_VPWR_c_673_n 0.00524008f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B1_M1026_g N_VPWR_c_673_n 0.00524008f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B1_M1035_g N_VPWR_c_673_n 0.00591596f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B1_M1005_g N_VPWR_c_691_n 0.00366111f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B1_M1013_g N_VPWR_c_691_n 0.00366111f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B1_M1026_g N_VPWR_c_691_n 0.00366111f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B1_M1035_g N_VPWR_c_691_n 0.00366111f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B1_M1035_g N_VPWR_c_692_n 8.92616e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_157 N_B1_c_109_n N_VGND_c_824_n 0.00816685f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B1_c_110_n N_VGND_c_824_n 5.0911e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_159 B1 N_VGND_c_824_n 0.00182093f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_160 N_B1_c_113_n N_VGND_c_824_n 0.00488836f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B1_c_114_n N_VGND_c_824_n 0.00693571f $X=0.215 $Y=1.305 $X2=0 $Y2=0
cc_162 N_B1_c_109_n N_VGND_c_825_n 5.08801e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B1_c_110_n N_VGND_c_825_n 0.00664421f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B1_c_111_n N_VGND_c_825_n 0.00664421f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_165 N_B1_c_112_n N_VGND_c_825_n 5.48314e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_166 N_B1_c_111_n N_VGND_c_826_n 5.48314e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B1_c_112_n N_VGND_c_826_n 0.00774571f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B1_c_109_n N_VGND_c_829_n 0.0046653f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B1_c_110_n N_VGND_c_829_n 0.00339367f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B1_c_111_n N_VGND_c_830_n 0.00339367f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B1_c_112_n N_VGND_c_830_n 0.00339367f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_c_109_n N_VGND_c_834_n 0.00789179f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B1_c_110_n N_VGND_c_834_n 0.00394406f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B1_c_111_n N_VGND_c_834_n 0.00398704f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B1_c_112_n N_VGND_c_834_n 0.00398704f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A1_c_191_n N_A2_c_260_n 0.0220586f $X=4.06 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_177 N_A1_M1030_g N_A2_M1014_g 0.0328195f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A1_c_192_n A2 0.0163961f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A1_c_193_n A2 2.30904e-19 $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A1_c_192_n N_A2_c_266_n 0.00419482f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A1_c_193_n N_A2_c_266_n 0.0220586f $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A1_M1002_g N_A_27_297#_c_473_n 0.0153328f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A1_M1018_g N_A_27_297#_c_473_n 0.014417f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A1_c_192_n N_A_27_297#_c_473_n 0.0239985f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A1_c_193_n N_A_27_297#_c_473_n 0.00765196f $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A1_M1022_g N_A_27_297#_c_477_n 0.014055f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A1_M1030_g N_A_27_297#_c_477_n 0.0149549f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A1_c_192_n N_A_27_297#_c_477_n 0.0304209f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A1_c_193_n N_A_27_297#_c_477_n 0.00191112f $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A1_c_192_n N_A_27_297#_c_481_n 0.00996364f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A1_c_193_n N_A_27_297#_c_481_n 0.00200701f $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A1_c_192_n N_A_27_297#_c_483_n 0.00107674f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A1_M1002_g N_Y_c_607_n 2.50203e-19 $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A1_M1002_g N_Y_c_617_n 0.00536503f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A1_c_188_n Y 0.00439884f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_192_n Y 0.021261f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A1_c_193_n Y 0.00522634f $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A1_c_188_n N_Y_c_585_n 0.010581f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_c_189_n N_Y_c_585_n 0.00847802f $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_190_n N_Y_c_585_n 0.00847802f $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_191_n N_Y_c_585_n 0.00374227f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A1_c_192_n N_Y_c_585_n 0.0959248f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A1_c_193_n N_Y_c_585_n 0.0142922f $X=4.06 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A1_M1018_g N_VPWR_c_674_n 6.83205e-19 $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A1_M1022_g N_VPWR_c_674_n 0.01018f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A1_M1030_g N_VPWR_c_674_n 0.0108578f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A1_M1030_g N_VPWR_c_675_n 7.05596e-19 $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A1_M1018_g N_VPWR_c_684_n 0.00340533f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A1_M1022_g N_VPWR_c_684_n 0.0046653f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A1_M1030_g N_VPWR_c_685_n 0.0046653f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A1_M1002_g N_VPWR_c_673_n 0.00456094f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A1_M1018_g N_VPWR_c_673_n 0.00394764f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A1_M1022_g N_VPWR_c_673_n 0.00789179f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A1_M1030_g N_VPWR_c_673_n 0.00822002f $X=4.06 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A1_M1002_g N_VPWR_c_691_n 0.00340533f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A1_M1002_g N_VPWR_c_692_n 0.00916224f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A1_M1018_g N_VPWR_c_692_n 0.00778056f $X=3.22 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A1_M1022_g N_VPWR_c_692_n 5.24369e-19 $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A1_c_188_n N_VGND_c_826_n 0.00240633f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A1_c_188_n N_VGND_c_831_n 0.00366111f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A1_c_189_n N_VGND_c_831_n 0.00366111f $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A1_c_190_n N_VGND_c_831_n 0.00366111f $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A1_c_191_n N_VGND_c_831_n 0.00366111f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A1_c_188_n N_VGND_c_834_n 0.00656615f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A1_c_189_n N_VGND_c_834_n 0.00524008f $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A1_c_190_n N_VGND_c_834_n 0.00524008f $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A1_c_191_n N_VGND_c_834_n 0.00526729f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A1_c_188_n N_A_493_47#_c_959_n 0.00789149f $X=2.8 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A1_c_189_n N_A_493_47#_c_959_n 0.00789149f $X=3.22 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A1_c_190_n N_A_493_47#_c_959_n 0.00789149f $X=3.64 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A1_c_191_n N_A_493_47#_c_959_n 0.00930387f $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A1_c_192_n N_A_493_47#_c_959_n 0.00489343f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A1_c_191_n N_A_911_47#_c_989_n 4.91085e-19 $X=4.06 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_M1028_g N_A3_M1007_g 0.0211577f $X=6.24 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A2_c_264_n N_A3_c_335_n 0.0211577f $X=6.165 $Y=1.177 $X2=0 $Y2=0
cc_236 A2 N_A3_c_335_n 2.43851e-19 $X=6.1 $Y=1.105 $X2=0 $Y2=0
cc_237 N_A2_c_264_n N_A3_c_336_n 0.00131494f $X=6.165 $Y=1.177 $X2=0 $Y2=0
cc_238 A2 N_A3_c_336_n 0.0140826f $X=6.1 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A2_M1014_g N_A_27_297#_c_484_n 0.00777966f $X=4.575 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A2_M1014_g N_A_27_297#_c_485_n 0.0152163f $X=4.575 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A2_M1017_g N_A_27_297#_c_485_n 0.0147487f $X=4.995 $Y=1.985 $X2=0 $Y2=0
cc_242 A2 N_A_27_297#_c_485_n 0.0277237f $X=6.1 $Y=1.105 $X2=0 $Y2=0
cc_243 N_A2_c_266_n N_A_27_297#_c_485_n 0.00459735f $X=5.815 $Y=1.177 $X2=0
+ $Y2=0
cc_244 N_A2_M1019_g N_A_27_297#_c_489_n 0.0171984f $X=5.415 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A2_M1028_g N_A_27_297#_c_489_n 0.0172727f $X=6.24 $Y=1.985 $X2=0 $Y2=0
cc_246 A2 N_A_27_297#_c_489_n 0.0437563f $X=6.1 $Y=1.105 $X2=0 $Y2=0
cc_247 N_A2_c_266_n N_A_27_297#_c_489_n 0.011822f $X=5.815 $Y=1.177 $X2=0 $Y2=0
cc_248 N_A2_M1028_g N_A_27_297#_c_493_n 0.00522281f $X=6.24 $Y=1.985 $X2=0 $Y2=0
cc_249 A2 N_A_27_297#_c_494_n 0.00861209f $X=6.1 $Y=1.105 $X2=0 $Y2=0
cc_250 N_A2_c_266_n N_A_27_297#_c_494_n 0.00243851f $X=5.815 $Y=1.177 $X2=0
+ $Y2=0
cc_251 N_A2_c_260_n N_Y_c_585_n 4.91085e-19 $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A2_M1014_g N_VPWR_c_674_n 7.17597e-19 $X=4.575 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A2_M1014_g N_VPWR_c_675_n 0.0119952f $X=4.575 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A2_M1017_g N_VPWR_c_675_n 0.0102769f $X=4.995 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A2_M1019_g N_VPWR_c_675_n 6.23635e-19 $X=5.415 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A2_M1019_g N_VPWR_c_676_n 0.00224235f $X=5.415 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A2_M1028_g N_VPWR_c_676_n 0.0022782f $X=6.24 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A2_M1028_g N_VPWR_c_677_n 6.10772e-19 $X=6.24 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A2_M1028_g N_VPWR_c_682_n 0.00583607f $X=6.24 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A2_M1014_g N_VPWR_c_685_n 0.0046653f $X=4.575 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A2_M1017_g N_VPWR_c_686_n 0.0046653f $X=4.995 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A2_M1019_g N_VPWR_c_686_n 0.00585385f $X=5.415 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A2_M1014_g N_VPWR_c_673_n 0.00822002f $X=4.575 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A2_M1017_g N_VPWR_c_673_n 0.00789179f $X=4.995 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A2_M1019_g N_VPWR_c_673_n 0.0111738f $X=5.415 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A2_M1028_g N_VPWR_c_673_n 0.0112254f $X=6.24 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A2_c_260_n N_VGND_c_831_n 0.00366111f $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A2_c_261_n N_VGND_c_831_n 0.00366111f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A2_c_262_n N_VGND_c_831_n 0.00366111f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A2_c_263_n N_VGND_c_831_n 0.00366111f $X=5.74 $Y=1.01 $X2=0 $Y2=0
cc_271 N_A2_c_260_n N_VGND_c_834_n 0.00526729f $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A2_c_261_n N_VGND_c_834_n 0.00524008f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A2_c_262_n N_VGND_c_834_n 0.00524008f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A2_c_263_n N_VGND_c_834_n 0.00656615f $X=5.74 $Y=1.01 $X2=0 $Y2=0
cc_275 N_A2_c_260_n N_A_493_47#_c_959_n 0.00953845f $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A2_c_261_n N_A_493_47#_c_959_n 0.00789149f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A2_c_262_n N_A_493_47#_c_959_n 0.00789149f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A2_c_263_n N_A_493_47#_c_959_n 0.00789149f $X=5.74 $Y=1.01 $X2=0 $Y2=0
cc_279 A2 N_A_493_47#_c_959_n 0.00285767f $X=6.1 $Y=1.105 $X2=0 $Y2=0
cc_280 N_A2_c_260_n N_A_911_47#_c_989_n 0.00383073f $X=4.48 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A2_c_261_n N_A_911_47#_c_989_n 0.00886233f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A2_c_262_n N_A_911_47#_c_989_n 0.00893253f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A2_c_263_n N_A_911_47#_c_989_n 0.0110355f $X=5.74 $Y=1.01 $X2=0 $Y2=0
cc_284 N_A2_c_264_n N_A_911_47#_c_989_n 0.0120065f $X=6.165 $Y=1.177 $X2=0 $Y2=0
cc_285 A2 N_A_911_47#_c_989_n 0.0782776f $X=6.1 $Y=1.105 $X2=0 $Y2=0
cc_286 N_A2_c_266_n N_A_911_47#_c_989_n 0.0072106f $X=5.815 $Y=1.177 $X2=0 $Y2=0
cc_287 N_A3_c_335_n N_A4_c_397_n 0.0238532f $X=7.94 $Y=1.01 $X2=-0.19 $Y2=-0.24
cc_288 N_A3_M1037_g N_A4_M1015_g 0.0238532f $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A3_c_335_n A4 9.3002e-19 $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_290 N_A3_c_336_n A4 0.0100551f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A3_c_335_n N_A4_c_402_n 0.0238532f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_292 N_A3_c_336_n N_A4_c_402_n 3.64284e-19 $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A3_M1007_g N_A_27_297#_c_496_n 0.0147429f $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A3_M1027_g N_A_27_297#_c_496_n 0.0146685f $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A3_c_335_n N_A_27_297#_c_496_n 0.00200188f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_296 N_A3_c_336_n N_A_27_297#_c_496_n 0.0271021f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A3_M1031_g N_A_27_297#_c_500_n 0.0146685f $X=7.52 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A3_c_335_n N_A_27_297#_c_500_n 0.00198468f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_299 N_A3_M1037_g N_A_27_297#_c_500_n 0.0162142f $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A3_c_336_n N_A_27_297#_c_500_n 0.0230062f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A3_c_335_n N_A_27_297#_c_504_n 0.00211036f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_302 N_A3_c_336_n N_A_27_297#_c_504_n 0.00901315f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A3_M1007_g N_VPWR_c_677_n 0.0103323f $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A3_M1027_g N_VPWR_c_677_n 0.0101939f $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A3_M1031_g N_VPWR_c_677_n 6.0901e-19 $X=7.52 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A3_M1027_g N_VPWR_c_678_n 0.0046653f $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A3_M1031_g N_VPWR_c_678_n 0.0046653f $X=7.52 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A3_M1027_g N_VPWR_c_679_n 6.0901e-19 $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A3_M1031_g N_VPWR_c_679_n 0.0128916f $X=7.52 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A3_M1037_g N_VPWR_c_679_n 0.0128916f $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A3_M1037_g N_VPWR_c_680_n 6.0901e-19 $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A3_M1007_g N_VPWR_c_682_n 0.0046653f $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A3_M1037_g N_VPWR_c_687_n 0.0046653f $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A3_M1007_g N_VPWR_c_673_n 0.00796757f $X=6.68 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A3_M1027_g N_VPWR_c_673_n 0.00789179f $X=7.1 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A3_M1031_g N_VPWR_c_673_n 0.00789179f $X=7.52 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A3_M1037_g N_VPWR_c_673_n 0.007919f $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A3_c_335_n N_VGND_c_827_n 0.00111179f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_319 N_A3_c_332_n N_VGND_c_831_n 0.00366111f $X=6.68 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A3_c_333_n N_VGND_c_831_n 0.00366111f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A3_c_334_n N_VGND_c_831_n 0.00366111f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A3_c_335_n N_VGND_c_831_n 0.00366111f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_323 N_A3_c_332_n N_VGND_c_834_n 0.00656615f $X=6.68 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A3_c_333_n N_VGND_c_834_n 0.00524008f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A3_c_334_n N_VGND_c_834_n 0.00524008f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A3_c_335_n N_VGND_c_834_n 0.00526729f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_327 N_A3_c_332_n N_A_911_47#_c_989_n 0.0110355f $X=6.68 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A3_c_333_n N_A_911_47#_c_989_n 0.00893253f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A3_c_334_n N_A_911_47#_c_989_n 0.00893253f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A3_c_335_n N_A_911_47#_c_989_n 0.00888656f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_331 N_A3_c_336_n N_A_911_47#_c_989_n 0.0560573f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A3_c_332_n N_A_1269_47#_c_1020_n 0.00789149f $X=6.68 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A3_c_333_n N_A_1269_47#_c_1020_n 0.00789149f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A3_c_334_n N_A_1269_47#_c_1020_n 0.00784733f $X=7.52 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A3_c_335_n N_A_1269_47#_c_1020_n 0.0105238f $X=7.94 $Y=1.01 $X2=0 $Y2=0
cc_336 N_A3_c_336_n N_A_1269_47#_c_1020_n 0.00144248f $X=7.79 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_A4_M1015_g N_A_27_297#_c_506_n 0.0147309f $X=8.36 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A4_M1020_g N_A_27_297#_c_506_n 0.0147751f $X=8.78 $Y=1.985 $X2=0 $Y2=0
cc_339 A4 N_A_27_297#_c_506_n 0.024239f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_340 N_A4_c_402_n N_A_27_297#_c_506_n 0.0019496f $X=9.62 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A4_M1023_g N_A_27_297#_c_510_n 0.0147309f $X=9.2 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A4_M1032_g N_A_27_297#_c_510_n 0.016074f $X=9.62 $Y=1.985 $X2=0 $Y2=0
cc_343 A4 N_A_27_297#_c_510_n 0.0354711f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_344 N_A4_c_402_n N_A_27_297#_c_510_n 0.00713614f $X=9.62 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A4_M1032_g N_A_27_297#_c_514_n 0.0052862f $X=9.62 $Y=1.985 $X2=0 $Y2=0
cc_346 A4 N_A_27_297#_c_515_n 0.00848579f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_347 N_A4_c_402_n N_A_27_297#_c_515_n 0.00206078f $X=9.62 $Y=1.16 $X2=0 $Y2=0
cc_348 N_A4_M1015_g N_VPWR_c_679_n 6.0901e-19 $X=8.36 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A4_M1015_g N_VPWR_c_680_n 0.0101939f $X=8.36 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A4_M1020_g N_VPWR_c_680_n 0.0101939f $X=8.78 $Y=1.985 $X2=0 $Y2=0
cc_351 N_A4_M1023_g N_VPWR_c_680_n 6.0901e-19 $X=9.2 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A4_M1020_g N_VPWR_c_681_n 6.0901e-19 $X=8.78 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A4_M1023_g N_VPWR_c_681_n 0.0101939f $X=9.2 $Y=1.985 $X2=0 $Y2=0
cc_354 N_A4_M1032_g N_VPWR_c_681_n 0.0125179f $X=9.62 $Y=1.985 $X2=0 $Y2=0
cc_355 N_A4_M1015_g N_VPWR_c_687_n 0.0046653f $X=8.36 $Y=1.985 $X2=0 $Y2=0
cc_356 N_A4_M1020_g N_VPWR_c_688_n 0.0046653f $X=8.78 $Y=1.985 $X2=0 $Y2=0
cc_357 N_A4_M1023_g N_VPWR_c_688_n 0.0046653f $X=9.2 $Y=1.985 $X2=0 $Y2=0
cc_358 N_A4_M1032_g N_VPWR_c_689_n 0.0046653f $X=9.62 $Y=1.985 $X2=0 $Y2=0
cc_359 N_A4_M1015_g N_VPWR_c_673_n 0.007919f $X=8.36 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A4_M1020_g N_VPWR_c_673_n 0.00789179f $X=8.78 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A4_M1023_g N_VPWR_c_673_n 0.00789179f $X=9.2 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A4_M1032_g N_VPWR_c_673_n 0.0088736f $X=9.62 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A4_c_397_n N_VGND_c_827_n 0.00783744f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A4_c_398_n N_VGND_c_827_n 0.00664421f $X=8.78 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A4_c_399_n N_VGND_c_827_n 5.08801e-19 $X=9.2 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A4_c_398_n N_VGND_c_828_n 5.08801e-19 $X=8.78 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A4_c_399_n N_VGND_c_828_n 0.00664421f $X=9.2 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A4_c_400_n N_VGND_c_828_n 0.00834749f $X=9.62 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A4_c_397_n N_VGND_c_831_n 0.00339367f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A4_c_398_n N_VGND_c_832_n 0.00339367f $X=8.78 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A4_c_399_n N_VGND_c_832_n 0.00339367f $X=9.2 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A4_c_400_n N_VGND_c_833_n 0.00339367f $X=9.62 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A4_c_397_n N_VGND_c_834_n 0.00397127f $X=8.36 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A4_c_398_n N_VGND_c_834_n 0.00394406f $X=8.78 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A4_c_399_n N_VGND_c_834_n 0.00394406f $X=9.2 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A4_c_400_n N_VGND_c_834_n 0.00492587f $X=9.62 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A4_c_397_n N_A_1269_47#_c_1026_n 0.0115547f $X=8.36 $Y=0.995 $X2=0
+ $Y2=0
cc_378 N_A4_c_398_n N_A_1269_47#_c_1026_n 0.0119869f $X=8.78 $Y=0.995 $X2=0
+ $Y2=0
cc_379 A4 N_A_1269_47#_c_1026_n 0.0259983f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_380 N_A4_c_402_n N_A_1269_47#_c_1026_n 0.00207061f $X=9.62 $Y=1.16 $X2=0
+ $Y2=0
cc_381 N_A4_c_399_n N_A_1269_47#_c_1030_n 0.0119869f $X=9.2 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A4_c_400_n N_A_1269_47#_c_1030_n 0.0132392f $X=9.62 $Y=0.995 $X2=0
+ $Y2=0
cc_383 A4 N_A_1269_47#_c_1030_n 0.0363475f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_384 N_A4_c_402_n N_A_1269_47#_c_1030_n 0.00593149f $X=9.62 $Y=1.16 $X2=0
+ $Y2=0
cc_385 A4 N_A_1269_47#_c_1034_n 0.00892733f $X=9.8 $Y=1.105 $X2=0 $Y2=0
cc_386 N_A4_c_402_n N_A_1269_47#_c_1034_n 0.00216182f $X=9.62 $Y=1.16 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_c_464_n N_Y_M1005_d 0.00325424f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_388 N_A_27_297#_c_464_n N_Y_M1026_d 0.00325424f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_389 N_A_27_297#_M1013_s N_Y_c_593_n 0.00465037f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_390 N_A_27_297#_c_464_n N_Y_c_593_n 0.0114593f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_391 N_A_27_297#_M1035_s N_Y_c_599_n 0.00418466f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_392 N_A_27_297#_c_464_n N_Y_c_599_n 0.00517219f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_393 N_A_27_297#_c_464_n N_Y_c_601_n 0.0157268f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_394 N_A_27_297#_c_464_n N_Y_c_607_n 0.0162597f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_395 N_A_27_297#_c_471_n N_Y_c_607_n 3.13275e-19 $X=2.25 $Y=2.255 $X2=0 $Y2=0
cc_396 N_A_27_297#_c_472_n N_Y_c_607_n 0.00628238f $X=2.335 $Y=1.99 $X2=0 $Y2=0
cc_397 N_A_27_297#_M1035_s N_Y_c_617_n 0.00893707f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_398 N_A_27_297#_c_464_n N_Y_c_617_n 0.00720722f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_399 N_A_27_297#_M1035_s Y 3.01855e-19 $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_400 N_A_27_297#_c_473_n N_VPWR_M1002_s 0.0160464f $X=3.345 $Y=1.99 $X2=-0.19
+ $Y2=1.305
cc_401 N_A_27_297#_c_477_n N_VPWR_M1022_s 0.0033993f $X=4.185 $Y=1.66 $X2=0
+ $Y2=0
cc_402 N_A_27_297#_c_485_n N_VPWR_M1014_d 0.00351323f $X=5.12 $Y=1.66 $X2=0
+ $Y2=0
cc_403 N_A_27_297#_c_489_n N_VPWR_M1019_d 0.0150542f $X=6.385 $Y=1.66 $X2=0
+ $Y2=0
cc_404 N_A_27_297#_c_496_n N_VPWR_M1007_d 0.0034684f $X=7.225 $Y=1.66 $X2=0
+ $Y2=0
cc_405 N_A_27_297#_c_500_n N_VPWR_M1031_d 0.0034684f $X=8.065 $Y=1.66 $X2=0
+ $Y2=0
cc_406 N_A_27_297#_c_506_n N_VPWR_M1015_s 0.0035361f $X=8.905 $Y=1.66 $X2=0
+ $Y2=0
cc_407 N_A_27_297#_c_510_n N_VPWR_M1023_s 0.0035361f $X=9.775 $Y=1.66 $X2=0
+ $Y2=0
cc_408 N_A_27_297#_c_477_n N_VPWR_c_674_n 0.0170259f $X=4.185 $Y=1.66 $X2=0
+ $Y2=0
cc_409 N_A_27_297#_c_484_n N_VPWR_c_675_n 0.0267757f $X=4.27 $Y=2.26 $X2=0 $Y2=0
cc_410 N_A_27_297#_c_485_n N_VPWR_c_675_n 0.0170259f $X=5.12 $Y=1.66 $X2=0 $Y2=0
cc_411 N_A_27_297#_c_489_n N_VPWR_c_676_n 0.0456421f $X=6.385 $Y=1.66 $X2=0
+ $Y2=0
cc_412 N_A_27_297#_c_493_n N_VPWR_c_676_n 0.0377548f $X=6.47 $Y=1.96 $X2=0 $Y2=0
cc_413 N_A_27_297#_c_496_n N_VPWR_c_677_n 0.0170259f $X=7.225 $Y=1.66 $X2=0
+ $Y2=0
cc_414 N_A_27_297#_c_544_p N_VPWR_c_678_n 0.0113958f $X=7.31 $Y=1.96 $X2=0 $Y2=0
cc_415 N_A_27_297#_c_500_n N_VPWR_c_679_n 0.0171101f $X=8.065 $Y=1.66 $X2=0
+ $Y2=0
cc_416 N_A_27_297#_c_506_n N_VPWR_c_680_n 0.0170259f $X=8.905 $Y=1.66 $X2=0
+ $Y2=0
cc_417 N_A_27_297#_c_510_n N_VPWR_c_681_n 0.0170259f $X=9.775 $Y=1.66 $X2=0
+ $Y2=0
cc_418 N_A_27_297#_c_514_n N_VPWR_c_681_n 0.0358254f $X=9.86 $Y=1.96 $X2=0 $Y2=0
cc_419 N_A_27_297#_c_493_n N_VPWR_c_682_n 0.0116048f $X=6.47 $Y=1.96 $X2=0 $Y2=0
cc_420 N_A_27_297#_c_473_n N_VPWR_c_684_n 0.00238578f $X=3.345 $Y=1.99 $X2=0
+ $Y2=0
cc_421 N_A_27_297#_c_551_p N_VPWR_c_684_n 0.0113958f $X=3.43 $Y=2.3 $X2=0 $Y2=0
cc_422 N_A_27_297#_c_484_n N_VPWR_c_685_n 0.00922815f $X=4.27 $Y=2.26 $X2=0
+ $Y2=0
cc_423 N_A_27_297#_c_553_p N_VPWR_c_686_n 0.0113958f $X=5.205 $Y=1.96 $X2=0
+ $Y2=0
cc_424 N_A_27_297#_c_554_p N_VPWR_c_687_n 0.0113958f $X=8.15 $Y=1.96 $X2=0 $Y2=0
cc_425 N_A_27_297#_c_555_p N_VPWR_c_688_n 0.0113958f $X=8.99 $Y=1.96 $X2=0 $Y2=0
cc_426 N_A_27_297#_c_514_n N_VPWR_c_689_n 0.0118139f $X=9.86 $Y=1.96 $X2=0 $Y2=0
cc_427 N_A_27_297#_M1005_s N_VPWR_c_673_n 0.00211652f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_428 N_A_27_297#_M1013_s N_VPWR_c_673_n 0.00217615f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_429 N_A_27_297#_M1035_s N_VPWR_c_673_n 0.00490457f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_430 N_A_27_297#_M1018_d N_VPWR_c_673_n 0.00406561f $X=3.295 $Y=1.485 $X2=0
+ $Y2=0
cc_431 N_A_27_297#_M1030_d N_VPWR_c_673_n 0.00978447f $X=4.135 $Y=1.485 $X2=0
+ $Y2=0
cc_432 N_A_27_297#_M1017_s N_VPWR_c_673_n 0.00562358f $X=5.07 $Y=1.485 $X2=0
+ $Y2=0
cc_433 N_A_27_297#_M1028_s N_VPWR_c_673_n 0.00647849f $X=6.315 $Y=1.485 $X2=0
+ $Y2=0
cc_434 N_A_27_297#_M1027_s N_VPWR_c_673_n 0.00562358f $X=7.175 $Y=1.485 $X2=0
+ $Y2=0
cc_435 N_A_27_297#_M1037_s N_VPWR_c_673_n 0.00562358f $X=8.015 $Y=1.485 $X2=0
+ $Y2=0
cc_436 N_A_27_297#_M1020_d N_VPWR_c_673_n 0.00562358f $X=8.855 $Y=1.485 $X2=0
+ $Y2=0
cc_437 N_A_27_297#_M1032_d N_VPWR_c_673_n 0.00653973f $X=9.695 $Y=1.485 $X2=0
+ $Y2=0
cc_438 N_A_27_297#_c_464_n N_VPWR_c_673_n 0.0724063f $X=2.165 $Y=2.34 $X2=0
+ $Y2=0
cc_439 N_A_27_297#_c_471_n N_VPWR_c_673_n 0.00651407f $X=2.25 $Y=2.255 $X2=0
+ $Y2=0
cc_440 N_A_27_297#_c_473_n N_VPWR_c_673_n 0.0112425f $X=3.345 $Y=1.99 $X2=0
+ $Y2=0
cc_441 N_A_27_297#_c_551_p N_VPWR_c_673_n 0.00646998f $X=3.43 $Y=2.3 $X2=0 $Y2=0
cc_442 N_A_27_297#_c_484_n N_VPWR_c_673_n 0.00634211f $X=4.27 $Y=2.26 $X2=0
+ $Y2=0
cc_443 N_A_27_297#_c_553_p N_VPWR_c_673_n 0.00646998f $X=5.205 $Y=1.96 $X2=0
+ $Y2=0
cc_444 N_A_27_297#_c_493_n N_VPWR_c_673_n 0.00646998f $X=6.47 $Y=1.96 $X2=0
+ $Y2=0
cc_445 N_A_27_297#_c_544_p N_VPWR_c_673_n 0.00646998f $X=7.31 $Y=1.96 $X2=0
+ $Y2=0
cc_446 N_A_27_297#_c_554_p N_VPWR_c_673_n 0.00646998f $X=8.15 $Y=1.96 $X2=0
+ $Y2=0
cc_447 N_A_27_297#_c_555_p N_VPWR_c_673_n 0.00646998f $X=8.99 $Y=1.96 $X2=0
+ $Y2=0
cc_448 N_A_27_297#_c_514_n N_VPWR_c_673_n 0.00646998f $X=9.86 $Y=1.96 $X2=0
+ $Y2=0
cc_449 N_A_27_297#_c_464_n N_VPWR_c_691_n 0.0938507f $X=2.165 $Y=2.34 $X2=0
+ $Y2=0
cc_450 N_A_27_297#_c_471_n N_VPWR_c_691_n 0.0115494f $X=2.25 $Y=2.255 $X2=0
+ $Y2=0
cc_451 N_A_27_297#_c_473_n N_VPWR_c_691_n 0.00238578f $X=3.345 $Y=1.99 $X2=0
+ $Y2=0
cc_452 N_A_27_297#_c_473_n N_VPWR_c_692_n 0.0398744f $X=3.345 $Y=1.99 $X2=0
+ $Y2=0
cc_453 N_Y_M1005_d N_VPWR_c_673_n 0.00219239f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_454 N_Y_M1026_d N_VPWR_c_673_n 0.00219239f $X=1.385 $Y=1.485 $X2=0 $Y2=0
cc_455 N_Y_c_587_n N_VGND_M1024_d 0.00337587f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_456 N_Y_c_597_n N_VGND_M1036_d 0.00348353f $X=1.935 $Y=0.72 $X2=0 $Y2=0
cc_457 Y N_VGND_M1036_d 0.00213667f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_458 Y N_VGND_M1036_d 0.00127255f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_459 N_Y_c_587_n N_VGND_c_825_n 0.0159625f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_460 N_Y_c_597_n N_VGND_c_826_n 0.00756697f $X=1.935 $Y=0.72 $X2=0 $Y2=0
cc_461 Y N_VGND_c_826_n 0.0143704f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_462 N_Y_c_650_p N_VGND_c_829_n 0.0112274f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_463 N_Y_c_587_n N_VGND_c_829_n 0.00244309f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_464 N_Y_c_587_n N_VGND_c_830_n 0.00243651f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_465 N_Y_c_653_p N_VGND_c_830_n 0.0112274f $X=1.52 $Y=0.46 $X2=0 $Y2=0
cc_466 N_Y_c_597_n N_VGND_c_830_n 0.00243651f $X=1.935 $Y=0.72 $X2=0 $Y2=0
cc_467 Y N_VGND_c_831_n 0.00100541f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_468 N_Y_c_585_n N_VGND_c_831_n 0.00492601f $X=3.85 $Y=0.72 $X2=0 $Y2=0
cc_469 N_Y_M1021_s N_VGND_c_834_n 0.00405853f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_470 N_Y_M1025_s N_VGND_c_834_n 0.00251683f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_471 N_Y_M1003_d N_VGND_c_834_n 0.00219239f $X=2.875 $Y=0.235 $X2=0 $Y2=0
cc_472 N_Y_M1009_d N_VGND_c_834_n 0.00219239f $X=3.715 $Y=0.235 $X2=0 $Y2=0
cc_473 N_Y_c_650_p N_VGND_c_834_n 0.00643448f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_474 N_Y_c_587_n N_VGND_c_834_n 0.00987412f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_475 N_Y_c_653_p N_VGND_c_834_n 0.00643448f $X=1.52 $Y=0.46 $X2=0 $Y2=0
cc_476 N_Y_c_597_n N_VGND_c_834_n 0.0049287f $X=1.935 $Y=0.72 $X2=0 $Y2=0
cc_477 Y N_VGND_c_834_n 0.00240358f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_478 N_Y_c_585_n N_VGND_c_834_n 0.0105479f $X=3.85 $Y=0.72 $X2=0 $Y2=0
cc_479 N_Y_c_585_n N_A_493_47#_M1003_s 0.00460975f $X=3.85 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_480 N_Y_c_585_n N_A_493_47#_M1004_s 0.00312766f $X=3.85 $Y=0.72 $X2=0 $Y2=0
cc_481 N_Y_M1003_d N_A_493_47#_c_959_n 0.00315945f $X=2.875 $Y=0.235 $X2=0 $Y2=0
cc_482 N_Y_M1009_d N_A_493_47#_c_959_n 0.00315945f $X=3.715 $Y=0.235 $X2=0 $Y2=0
cc_483 N_Y_c_585_n N_A_493_47#_c_959_n 0.0797617f $X=3.85 $Y=0.72 $X2=0 $Y2=0
cc_484 N_Y_c_585_n N_A_911_47#_c_989_n 0.00576239f $X=3.85 $Y=0.72 $X2=0 $Y2=0
cc_485 N_VGND_c_834_n N_A_493_47#_M1003_s 0.00211652f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_486 N_VGND_c_834_n N_A_493_47#_M1004_s 0.00217615f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_c_834_n N_A_493_47#_M1012_s 0.00217615f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_834_n N_A_493_47#_M1010_d 0.00217615f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_834_n N_A_493_47#_M1039_d 0.00211652f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_c_826_n N_A_493_47#_c_959_n 0.00957091f $X=1.94 $Y=0.38 $X2=0
+ $Y2=0
cc_491 N_VGND_c_831_n N_A_493_47#_c_959_n 0.164437f $X=8.405 $Y=0 $X2=0 $Y2=0
cc_492 N_VGND_c_834_n N_A_493_47#_c_959_n 0.127969f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_493 N_VGND_c_834_n N_A_911_47#_M1006_s 0.00219239f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_494 N_VGND_c_834_n N_A_911_47#_M1011_s 0.00219239f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_495 N_VGND_c_834_n N_A_911_47#_M1000_s 0.00219239f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_834_n N_A_911_47#_M1033_s 0.00219239f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_831_n N_A_911_47#_c_989_n 0.00347243f $X=8.405 $Y=0 $X2=0 $Y2=0
cc_498 N_VGND_c_834_n N_A_911_47#_c_989_n 0.0111918f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_499 N_VGND_c_834_n N_A_1269_47#_M1000_d 0.00211652f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_500 N_VGND_c_834_n N_A_1269_47#_M1029_d 0.00217615f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_501 N_VGND_c_834_n N_A_1269_47#_M1034_d 0.00233519f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_502 N_VGND_c_834_n N_A_1269_47#_M1008_s 0.00249348f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_503 N_VGND_c_834_n N_A_1269_47#_M1038_s 0.00497468f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_504 N_VGND_c_831_n N_A_1269_47#_c_1020_n 0.0780741f $X=8.405 $Y=0 $X2=0 $Y2=0
cc_505 N_VGND_c_834_n N_A_1269_47#_c_1020_n 0.0608914f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_506 N_VGND_c_831_n N_A_1269_47#_c_1043_n 0.0112984f $X=8.405 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_834_n N_A_1269_47#_c_1043_n 0.00651108f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_M1001_d N_A_1269_47#_c_1026_n 0.00337587f $X=8.435 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_VGND_c_827_n N_A_1269_47#_c_1026_n 0.0159625f $X=8.57 $Y=0.38 $X2=0
+ $Y2=0
cc_510 N_VGND_c_831_n N_A_1269_47#_c_1026_n 0.00244309f $X=8.405 $Y=0 $X2=0
+ $Y2=0
cc_511 N_VGND_c_832_n N_A_1269_47#_c_1026_n 0.00244309f $X=9.245 $Y=0 $X2=0
+ $Y2=0
cc_512 N_VGND_c_834_n N_A_1269_47#_c_1026_n 0.00984256f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_832_n N_A_1269_47#_c_1050_n 0.0112274f $X=9.245 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_834_n N_A_1269_47#_c_1050_n 0.00643448f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_M1016_d N_A_1269_47#_c_1030_n 0.00337587f $X=9.275 $Y=0.235 $X2=0
+ $Y2=0
cc_516 N_VGND_c_828_n N_A_1269_47#_c_1030_n 0.0159625f $X=9.41 $Y=0.38 $X2=0
+ $Y2=0
cc_517 N_VGND_c_832_n N_A_1269_47#_c_1030_n 0.00244309f $X=9.245 $Y=0 $X2=0
+ $Y2=0
cc_518 N_VGND_c_833_n N_A_1269_47#_c_1030_n 0.00244309f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_834_n N_A_1269_47#_c_1030_n 0.00984256f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_833_n N_A_1269_47#_c_1057_n 0.01143f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_834_n N_A_1269_47#_c_1057_n 0.00643448f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_522 N_A_493_47#_c_959_n N_A_911_47#_M1006_s 0.00315945f $X=5.95 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_523 N_A_493_47#_c_959_n N_A_911_47#_M1011_s 0.00316323f $X=5.95 $Y=0.38 $X2=0
+ $Y2=0
cc_524 N_A_493_47#_M1010_d N_A_911_47#_c_989_n 0.00337959f $X=4.975 $Y=0.235
+ $X2=0 $Y2=0
cc_525 N_A_493_47#_M1039_d N_A_911_47#_c_989_n 0.00489735f $X=5.815 $Y=0.235
+ $X2=0 $Y2=0
cc_526 N_A_493_47#_c_959_n N_A_911_47#_c_989_n 0.0797617f $X=5.95 $Y=0.38 $X2=0
+ $Y2=0
cc_527 N_A_493_47#_c_959_n N_A_1269_47#_c_1020_n 0.0145425f $X=5.95 $Y=0.38
+ $X2=0 $Y2=0
cc_528 N_A_911_47#_c_989_n N_A_1269_47#_M1000_d 0.0105704f $X=7.73 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_529 N_A_911_47#_c_989_n N_A_1269_47#_M1029_d 0.00337959f $X=7.73 $Y=0.72
+ $X2=0 $Y2=0
cc_530 N_A_911_47#_M1000_s N_A_1269_47#_c_1020_n 0.00315945f $X=6.755 $Y=0.235
+ $X2=0 $Y2=0
cc_531 N_A_911_47#_M1033_s N_A_1269_47#_c_1020_n 0.00316323f $X=7.595 $Y=0.235
+ $X2=0 $Y2=0
cc_532 N_A_911_47#_c_989_n N_A_1269_47#_c_1020_n 0.0797617f $X=7.73 $Y=0.72
+ $X2=0 $Y2=0

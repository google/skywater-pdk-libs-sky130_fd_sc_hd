* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
M1000 a_1011_297# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=1.42455e+12p ps=1.291e+07u
M1001 VPWR a_101_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.4e+11p ps=5.08e+06u
M1002 VPWR a_101_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_1011_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.6515e+11p pd=1.82e+06u as=9.453e+11p ps=9.45e+06u
M1004 VGND A a_1117_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.8275e+11p ps=3.78e+06u
M1005 X a_101_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1117_297# a_1011_297# a_631_49# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=4.5445e+11p ps=4.02e+06u
M1007 a_607_325# B a_1117_297# VNB nshort w=640000u l=150000u
+  ad=5.881e+11p pd=4.47e+06u as=0p ps=0u
M1008 a_1117_297# a_1011_297# a_607_325# VPB phighvt w=840000u l=150000u
+  ad=6.958e+11p pd=5.23e+06u as=5.646e+11p ps=4.74e+06u
M1009 a_1382_49# a_1117_297# VGND VNB nshort w=640000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=0p ps=0u
M1010 VGND a_101_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.51e+11p ps=3.68e+06u
M1011 a_101_21# C a_607_325# VPB phighvt w=840000u l=150000u
+  ad=3.059e+11p pd=2.63e+06u as=0p ps=0u
M1012 a_1382_49# a_1117_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=7.77e+11p pd=5.62e+06u as=0p ps=0u
M1013 a_607_325# B a_1382_49# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_101_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_101_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_492_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=0p ps=0u
M1017 VPWR A a_1117_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_631_49# B a_1117_297# VPB phighvt w=840000u l=150000u
+  ad=8.0855e+11p pd=5.34e+06u as=0p ps=0u
M1019 a_1382_49# a_1011_297# a_631_49# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_607_325# a_492_93# a_101_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1021 a_1382_49# a_1011_297# a_607_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_101_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_631_49# B a_1382_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_101_21# C a_631_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_492_93# C VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1026 a_631_49# a_492_93# a_101_21# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_101_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

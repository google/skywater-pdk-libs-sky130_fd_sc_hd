* File: sky130_fd_sc_hd__nand3_1.spice
* Created: Thu Aug 27 14:29:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand3_1.spice.pex"
.subckt sky130_fd_sc_hd__nand3_1  VNB VPB C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1004 A_109_47# N_C_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.1
+ A=0.0975 P=1.6 MULT=1
MM1001 A_193_47# N_B_M1001_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.08775 PD=0.98 PS=0.92 NRD=20.304 NRS=14.76 M=1 R=4.33333 SA=75000.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g A_193_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=20.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_C_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.1 A=0.15
+ P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.165 PD=2.52 PS=1.33 NRD=0 NRS=10.8153 M=1 R=6.66667 SA=75001.1 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=3.5631 P=7.65
*
.include "sky130_fd_sc_hd__nand3_1.spice.SKY130_FD_SC_HD__NAND3_1.pxi"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_hd__a21o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_386_297# VPB phighvt w=1e+06u l=150000u
+  ad=8.45e+11p pd=7.69e+06u as=5.4e+11p ps=5.08e+06u
M1001 a_80_199# B1 VGND VNB nshort w=650000u l=150000u
+  ad=3.25e+11p pd=2.3e+06u as=5.655e+11p ps=5.64e+06u
M1002 a_386_297# B1 a_80_199# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1003 X a_80_199# VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1004 X a_80_199# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1005 VGND A2 a_458_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.47e+11p ps=2.06e+06u
M1006 a_458_47# A1 a_80_199# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_80_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_386_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_80_199# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


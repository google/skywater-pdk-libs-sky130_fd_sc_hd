* File: sky130_fd_sc_hd__dfrbp_1.pex.spice
* Created: Tue Sep  1 19:02:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFRBP_1%CLK 1 2 3 5 6 8 11 13 14
c40 6 0 9.23148e-20 $X=0.47 $Y=1.74
c41 1 0 2.71124e-20 $X=0.305 $Y=1.325
r42 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=1.16
+ $X2=0.265 $Y2=1.53
r43 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r44 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r47 3 18 88.7086 $w=2.58e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r50 1 18 39.2009 $w=2.58e-07 $l=1.75656e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.327 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_27_47# 1 2 9 13 17 20 21 22 25 27 29 33 37
+ 41 42 43 46 49 50 51 52 55 61 68 71 72 77
c236 77 0 4.56546e-20 $X=6.07 $Y=1.11
c237 61 0 1.76704e-20 $X=6.11 $Y=1.19
c238 51 0 1.58851e-19 $X=5.965 $Y=1.19
c239 29 0 4.11863e-20 $X=5.845 $Y=2.275
c240 22 0 1.90473e-19 $X=2.72 $Y=1.32
r241 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=1.11 $X2=6.07 $Y2=1.11
r242 71 74 47.4498 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=1.095
r243 71 73 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=0.765
r244 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=0.93 $X2=2.585 $Y2=0.93
r245 65 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r246 61 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.19
+ $X2=6.11 $Y2=1.19
r247 59 72 8.56101 $w=3.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.56 $Y=1.19
+ $X2=2.56 $Y2=0.93
r248 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r249 55 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r250 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.19
+ $X2=0.695 $Y2=1.19
r251 52 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.19
+ $X2=2.53 $Y2=1.19
r252 51 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=6.11 $Y2=1.19
r253 51 52 4.07177 $w=1.4e-07 $l=3.29e-06 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=2.675 $Y2=1.19
r254 50 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.19
+ $X2=0.695 $Y2=1.19
r255 49 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r256 49 50 1.91213 $w=1.4e-07 $l=1.545e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.84 $Y2=1.19
r257 48 55 30.3143 $w=2.28e-07 $l=6.05e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.19
r258 47 55 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.19
r259 44 46 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r260 43 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.795
r261 43 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r262 41 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r263 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r264 35 42 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.345 $Y2=0.72
r265 35 37 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.51
r266 31 76 38.5991 $w=2.92e-07 $l=1.76125e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=5.987 $Y2=1.11
r267 31 33 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=6.01 $Y2=0.415
r268 27 76 58.4073 $w=2.92e-07 $l=3.48848e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.987 $Y2=1.11
r269 27 29 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.845 $Y2=2.275
r270 23 25 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.18 $Y=1.395
+ $X2=3.18 $Y2=2.275
r271 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=3.18 $Y2=1.395
r272 21 22 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=2.72 $Y2=1.32
r273 20 22 26.9401 $w=1.5e-07 $l=1.09243e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.72 $Y2=1.32
r274 20 74 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.642 $Y2=1.095
r275 17 73 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.64 $Y=0.415
+ $X2=2.64 $Y2=0.765
r276 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r277 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r278 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r279 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r280 2 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r281 1 37 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%D 3 7 9 10 15 19
c53 10 0 1.85993e-19 $X=2.09 $Y=1.3
c54 7 0 1.77283e-19 $X=2.225 $Y=2.275
r55 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.465 $X2=1.79 $Y2=1.465
r56 15 19 1.96287 $w=4.04e-07 $l=6.5e-08 $layer=LI1_cond $X=1.615 $Y=1.53
+ $X2=1.615 $Y2=1.465
r57 9 18 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.09 $Y=1.465 $X2=1.79
+ $Y2=1.465
r58 9 10 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.465
+ $X2=2.09 $Y2=1.3
r59 5 10 37.0704 $w=1.5e-07 $l=3.91727e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.09 $Y2=1.3
r60 5 7 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.225 $Y2=2.275
r61 1 10 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.165 $Y=1.3 $X2=2.09
+ $Y2=1.3
r62 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.165 $Y=1.3
+ $X2=2.165 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_193_47# 1 2 9 13 15 17 20 23 26 27 29 30
+ 34 35 37 38 39 40 47 49 53 65 66 70
c212 66 0 3.94709e-20 $X=6.265 $Y=1.74
c213 47 0 1.77283e-19 $X=2.99 $Y=1.87
c214 39 0 1.36782e-20 $X=5.965 $Y=1.87
c215 38 0 9.23148e-20 $X=1.245 $Y=1.87
c216 37 0 1.20979e-19 $X=2.845 $Y=1.87
c217 35 0 1.61046e-19 $X=3.095 $Y=0.9
c218 29 0 1.76704e-20 $X=5.97 $Y=1.58
c219 26 0 1.28114e-19 $X=5.59 $Y=0.87
r220 65 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.74
+ $X2=6.265 $Y2=1.905
r221 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.265
+ $Y=1.74 $X2=6.265 $Y2=1.74
r222 53 56 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.695 $Y=1.74
+ $X2=2.695 $Y2=1.875
r223 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.74 $X2=2.695 $Y2=1.74
r224 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.87
+ $X2=6.11 $Y2=1.87
r225 47 54 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=1.77
+ $X2=2.695 $Y2=1.77
r226 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.87
+ $X2=2.99 $Y2=1.87
r227 43 70 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.1 $Y=1.87
+ $X2=1.1 $Y2=0.51
r228 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=1.87 $X2=1.1
+ $Y2=1.87
r229 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.87
+ $X2=2.99 $Y2=1.87
r230 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=6.11 $Y2=1.87
r231 39 40 3.50247 $w=1.4e-07 $l=2.83e-06 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=3.135 $Y2=1.87
r232 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=1.87
+ $X2=1.1 $Y2=1.87
r233 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=2.99 $Y2=1.87
r234 37 38 1.98019 $w=1.4e-07 $l=1.6e-06 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=1.245 $Y2=1.87
r235 35 58 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.095 $Y=0.9
+ $X2=3.095 $Y2=0.765
r236 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=0.9 $X2=3.095 $Y2=0.9
r237 31 34 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.875
+ $X2=3.095 $Y2=0.875
r238 29 66 5.43733 $w=3.59e-07 $l=2.995e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=6.2 $Y2=1.74
r239 29 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=5.675 $Y2=1.58
r240 27 60 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.59 $Y=0.87
+ $X2=5.465 $Y2=0.87
r241 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=0.87 $X2=5.59 $Y2=0.87
r242 24 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.675 $Y2=1.58
r243 24 26 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.57 $Y2=0.87
r244 23 47 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.99 $Y=1.575
+ $X2=2.99 $Y2=1.77
r245 22 31 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=0.875
r246 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=1.575
r247 20 68 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.275 $Y=2.275
+ $X2=6.275 $Y2=1.905
r248 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.87
r249 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.415
r250 13 58 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.12 $Y=0.415
+ $X2=3.12 $Y2=0.765
r251 9 56 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.685 $Y=2.275
+ $X2=2.685 $Y2=1.875
r252 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r253 1 70 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_761_289# 1 2 9 13 15 18 21 23 25 26 27 30
+ 33 36 37
c109 36 0 1.00332e-19 $X=5.145 $Y=0.835
c110 23 0 4.11863e-20 $X=5.19 $Y=1.525
r111 33 35 3.58511 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.36
+ $X2=5.19 $Y2=0.445
r112 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.58 $Y=2.005
+ $X2=5.58 $Y2=2.3
r113 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.58 $Y2=2.005
r114 26 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.275 $Y2=1.92
r115 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.19 $Y=1.835
+ $X2=5.275 $Y2=1.92
r116 24 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.61
r117 24 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.835
r118 23 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=1.61
r119 23 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=0.835
r120 21 36 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.835
r121 21 35 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.445
r122 18 40 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.775
r123 18 39 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.445
r124 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.61 $X2=3.94 $Y2=1.61
r125 15 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=5.19 $Y2=1.61
r126 15 17 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=3.94 $Y2=1.61
r127 13 39 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.95 $Y=0.445
+ $X2=3.95 $Y2=1.445
r128 9 40 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.88 $Y=2.275 $X2=3.88
+ $Y2=1.775
r129 2 30 600 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.645 $X2=5.58 $Y2=2.3
r130 1 33 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.2 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%RESET_B 3 6 10 14 16 17 20 23 25 26 27 29 37
+ 39 42 57
c155 37 0 1.00332e-19 $X=4.37 $Y=0.93
c156 29 0 4.83118e-21 $X=7.19 $Y=1.165
c157 23 0 6.10372e-20 $X=4.25 $Y=0.85
c158 16 0 2.92e-20 $X=7.49 $Y=0.85
c159 14 0 1.03533e-19 $X=7.235 $Y=2.275
c160 10 0 4.70414e-20 $X=7.235 $Y=0.445
r161 49 57 3.2703 $w=2.4e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=1.035
+ $X2=7.525 $Y2=1.22
r162 42 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=1.285
r163 42 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=0.955
r164 37 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=1.095
r165 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=0.765
r166 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.27
+ $Y=1.12 $X2=7.27 $Y2=1.12
r167 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.19 $Y=1.165
+ $X2=7.19 $Y2=1.165
r168 27 34 0.181159 $w=2.07e-07 $l=3e-07 $layer=MET1_cond $X=7.19 $Y=0.85
+ $X2=7.49 $Y2=0.85
r169 27 29 0.0979621 $w=2.9e-07 $l=2e-07 $layer=MET1_cond $X=7.19 $Y=0.965
+ $X2=7.19 $Y2=1.165
r170 25 27 0.10072 $w=2.07e-07 $l=1.45e-07 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=7.19 $Y2=0.85
r171 25 26 3.2797 $w=1.4e-07 $l=2.65e-06 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=4.395 $Y2=0.85
r172 23 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=0.93 $X2=4.37 $Y2=0.93
r173 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.25 $Y=0.85
+ $X2=4.25 $Y2=0.85
r174 20 26 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.395 $Y2=0.85
r175 20 22 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.25 $Y2=0.85
r176 17 57 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.49 $Y=1.22
+ $X2=7.525 $Y2=1.22
r177 17 30 9.34413 $w=3.68e-07 $l=3e-07 $layer=LI1_cond $X=7.49 $Y=1.22 $X2=7.19
+ $Y2=1.22
r178 16 49 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=0.85
+ $X2=7.525 $Y2=1.035
r179 16 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.49 $Y=0.85
+ $X2=7.49 $Y2=0.85
r180 14 45 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=7.235 $Y=2.275
+ $X2=7.235 $Y2=1.285
r181 10 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.235 $Y=0.445
+ $X2=7.235 $Y2=0.955
r182 6 40 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=4.365 $Y=2.275
+ $X2=4.365 $Y2=1.095
r183 3 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.31 $Y=0.445
+ $X2=4.31 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_543_47# 1 2 9 11 13 15 16 20 25 27 28 29
+ 34 35
c126 35 0 6.10372e-20 $X=4.85 $Y=1.17
c127 29 0 1.61046e-19 $X=3.6 $Y=1.27
c128 11 0 1.36782e-20 $X=5.275 $Y=1.495
c129 9 0 1.28114e-19 $X=4.97 $Y=0.555
r130 34 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.85 $Y=1.17 $X2=4.85
+ $Y2=1.27
r131 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.17 $X2=4.85 $Y2=1.17
r132 30 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.33 $Y=1.27
+ $X2=3.515 $Y2=1.27
r133 29 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.27
+ $X2=3.515 $Y2=1.27
r134 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=4.85 $Y2=1.27
r135 28 29 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=3.6 $Y2=1.27
r136 27 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=1.185
+ $X2=3.515 $Y2=1.27
r137 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.515 $Y=0.475
+ $X2=3.515 $Y2=1.185
r138 24 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=1.27
r139 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=2.135
r140 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=3.515 $Y2=0.475
r141 20 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=2.91 $Y2=0.39
r142 16 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=3.33 $Y2=2.135
r143 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=2.9 $Y2=2.3
r144 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.35 $Y=1.57
+ $X2=5.35 $Y2=2.065
r145 12 35 61.4314 $w=2.55e-07 $l=3.99061e-07 $layer=POLY_cond $X=5.045 $Y=1.495
+ $X2=4.88 $Y2=1.17
r146 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.35 $Y2=1.57
r147 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.045 $Y2=1.495
r148 7 35 39.2931 $w=2.55e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.88 $Y2=1.17
r149 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.97 $Y2=0.555
r150 2 18 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.065 $X2=2.9 $Y2=2.33
r151 1 22 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.91 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_1283_21# 1 2 9 13 17 19 21 22 23 24 26 28
+ 31 33 37 38 41 45 46 47 50 52 53 54 55 57 60 65 72
c190 72 0 6.15427e-20 $X=6.695 $Y=0.98
c191 65 0 1.99375e-19 $X=8.075 $Y=1.072
c192 60 0 1.94811e-19 $X=7.15 $Y=0.78
c193 37 0 1.43777e-19 $X=9.542 $Y=1.515
c194 33 0 2.92e-20 $X=8.4 $Y=1.16
c195 13 0 2.35828e-20 $X=6.695 $Y=2.275
r196 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.27
+ $Y=1.16 $X2=8.27 $Y2=1.16
r197 65 67 5.76029 $w=4.13e-07 $l=1.95e-07 $layer=LI1_cond $X=8.075 $Y=1.072
+ $X2=8.27 $Y2=1.072
r198 64 65 2.954 $w=4.13e-07 $l=1e-07 $layer=LI1_cond $X=7.975 $Y=1.072
+ $X2=8.075 $Y2=1.072
r199 56 65 5.97325 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=8.075 $Y=1.325
+ $X2=8.075 $Y2=1.072
r200 56 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.075 $Y=1.325
+ $X2=8.075 $Y2=1.915
r201 55 64 2.23379 $w=3.2e-07 $l=2.52e-07 $layer=LI1_cond $X=7.975 $Y=0.82
+ $X2=7.975 $Y2=1.072
r202 54 63 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.975 $Y=0.465
+ $X2=7.975 $Y2=0.38
r203 54 55 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=7.975 $Y=0.465
+ $X2=7.975 $Y2=0.82
r204 52 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.99 $Y=2
+ $X2=8.075 $Y2=1.915
r205 52 53 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.99 $Y=2 $X2=7.53
+ $Y2=2
r206 48 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.53 $Y2=2
r207 48 50 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.445 $Y2=2.21
r208 46 63 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.975 $Y2=0.38
r209 46 47 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.235 $Y2=0.38
r210 45 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=0.695
+ $X2=7.15 $Y2=0.78
r211 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.235 $Y2=0.38
r212 44 45 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.15 $Y2=0.695
r213 42 72 17.8171 $w=2.57e-07 $l=9.5e-08 $layer=POLY_cond $X=6.79 $Y=0.98
+ $X2=6.695 $Y2=0.98
r214 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=0.98 $X2=6.79 $Y2=0.98
r215 39 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=0.78
+ $X2=7.15 $Y2=0.78
r216 39 41 6.02413 $w=2.18e-07 $l=1.15e-07 $layer=LI1_cond $X=6.815 $Y=0.865
+ $X2=6.815 $Y2=0.98
r217 37 38 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=9.542 $Y=1.515
+ $X2=9.542 $Y2=1.665
r218 34 35 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=8.475 $Y=1.16
+ $X2=8.63 $Y2=1.16
r219 33 68 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=8.4 $Y=1.16 $X2=8.27
+ $Y2=1.16
r220 33 34 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.4 $Y=1.16
+ $X2=8.475 $Y2=1.16
r221 31 38 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.57 $Y=2.165
+ $X2=9.57 $Y2=1.665
r222 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.57 $Y=0.73
+ $X2=9.57 $Y2=0.445
r223 24 37 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.515 $Y=1.325
+ $X2=9.515 $Y2=1.515
r224 23 35 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.705 $Y=1.16
+ $X2=8.63 $Y2=1.16
r225 22 24 49.1818 $w=1.63e-07 $l=1.77989e-07 $layer=POLY_cond $X=9.542 $Y=1.16
+ $X2=9.515 $Y2=1.325
r226 22 26 127.544 $w=1.63e-07 $l=4.43779e-07 $layer=POLY_cond $X=9.542 $Y=1.16
+ $X2=9.57 $Y2=0.73
r227 22 23 128.523 $w=3.3e-07 $l=7.35e-07 $layer=POLY_cond $X=9.44 $Y=1.16
+ $X2=8.705 $Y2=1.16
r228 19 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=0.995
+ $X2=8.63 $Y2=1.16
r229 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.63 $Y=0.995
+ $X2=8.63 $Y2=0.56
r230 15 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.475 $Y=1.325
+ $X2=8.475 $Y2=1.16
r231 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.475 $Y=1.325
+ $X2=8.475 $Y2=1.985
r232 11 72 15.359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=0.98
r233 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=2.275
r234 7 72 38.4475 $w=2.57e-07 $l=2.75409e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.695 $Y2=0.98
r235 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.49 $Y2=0.445
r236 2 50 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=2.065 $X2=7.445 $Y2=2.21
r237 1 63 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=7.765
+ $Y=0.235 $X2=7.9 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_1108_47# 1 2 9 13 15 19 24 25 26 29 30
c106 25 0 2.04429e-20 $X=6.685 $Y=1.745
c107 24 0 1.60161e-19 $X=6.45 $Y=1.315
c108 19 0 1.03533e-19 $X=6.6 $Y=2.295
c109 15 0 4.70414e-20 $X=6.365 $Y=0.395
c110 13 0 1.79199e-19 $X=7.69 $Y=0.445
r111 30 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.66
+ $X2=7.655 $Y2=1.495
r112 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.655
+ $Y=1.66 $X2=7.655 $Y2=1.66
r113 27 32 3.26844 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.77 $Y=1.66 $X2=6.6
+ $Y2=1.66
r114 27 29 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.77 $Y=1.66
+ $X2=7.655 $Y2=1.66
r115 25 32 5.45986 $w=2.62e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.6 $Y2=1.66
r116 25 26 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.685 $Y2=2.125
r117 24 32 17.5667 $w=2.62e-07 $l=4.13249e-07 $layer=LI1_cond $X=6.45 $Y=1.315
+ $X2=6.6 $Y2=1.66
r118 23 24 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.45 $Y=0.535
+ $X2=6.45 $Y2=1.315
r119 19 26 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.685 $Y2=2.125
r120 19 21 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.065 $Y2=2.295
r121 15 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=6.45 $Y2=0.535
r122 15 17 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=5.75 $Y2=0.395
r123 13 34 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=7.69 $Y=0.445
+ $X2=7.69 $Y2=1.495
r124 7 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=1.66
r125 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=2.275
r126 2 21 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=2.065 $X2=6.065 $Y2=2.335
r127 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.54
+ $Y=0.235 $X2=5.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_1847_47# 1 2 9 12 16 20 24 25 27 29
r48 25 30 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=9.982 $Y=1.16
+ $X2=9.982 $Y2=1.325
r49 25 29 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=9.982 $Y=1.16
+ $X2=9.982 $Y2=0.995
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.97
+ $Y=1.16 $X2=9.97 $Y2=1.16
r51 22 27 0.881669 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.525 $Y=1.16
+ $X2=9.36 $Y2=1.16
r52 22 24 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.525 $Y=1.16
+ $X2=9.97 $Y2=1.16
r53 18 27 5.74456 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=9.36 $Y=1.325
+ $X2=9.36 $Y2=1.16
r54 18 20 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.36 $Y=1.325
+ $X2=9.36 $Y2=2
r55 14 27 5.74456 $w=2.9e-07 $l=1.83916e-07 $layer=LI1_cond $X=9.32 $Y=0.995
+ $X2=9.36 $Y2=1.16
r56 14 16 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=9.32 $Y=0.995
+ $X2=9.32 $Y2=0.51
r57 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.055 $Y=1.985
+ $X2=10.055 $Y2=1.325
r58 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.055 $Y=0.56
+ $X2=10.055 $Y2=0.995
r59 2 20 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=9.235
+ $Y=1.845 $X2=9.36 $Y2=2
r60 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=9.235
+ $Y=0.235 $X2=9.36 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 49 50
+ 52 53 55 56 57 59 64 73 93 94 97 100 103 108 111
c156 44 0 1.43777e-19 $X=9.845 $Y=1.66
r157 110 111 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.265 $Y=2.53
+ $X2=8.43 $Y2=2.53
r158 106 110 4.67558 $w=5.48e-07 $l=2.15e-07 $layer=LI1_cond $X=8.05 $Y=2.53
+ $X2=8.265 $Y2=2.53
r159 106 108 13.6377 $w=5.48e-07 $l=3.4e-07 $layer=LI1_cond $X=8.05 $Y=2.53
+ $X2=7.71 $Y2=2.53
r160 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r161 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r162 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r163 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r164 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r165 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r166 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r167 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r168 88 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r169 87 90 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r170 87 111 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=8.51 $Y=2.72
+ $X2=8.43 $Y2=2.72
r171 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r172 84 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r173 83 108 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=7.71 $Y2=2.72
r174 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r175 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r176 80 104 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.29 $Y2=2.72
r177 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r178 77 103 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.14 $Y2=2.72
r179 77 79 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=6.67 $Y2=2.72
r180 76 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r181 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r182 73 103 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=5.14 $Y2=2.72
r183 73 75 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=4.83 $Y2=2.72
r184 72 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r185 72 101 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.07 $Y2=2.72
r186 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r187 69 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=1.975 $Y2=2.72
r188 69 71 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=3.91 $Y2=2.72
r189 68 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r190 68 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r191 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r192 65 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r193 65 67 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r194 64 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.975 $Y2=2.72
r195 64 67 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r196 59 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r197 59 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r198 57 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r199 57 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r200 55 90 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.76 $Y=2.72
+ $X2=9.43 $Y2=2.72
r201 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=2.72
+ $X2=9.845 $Y2=2.72
r202 54 93 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.93 $Y=2.72
+ $X2=10.35 $Y2=2.72
r203 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.93 $Y=2.72
+ $X2=9.845 $Y2=2.72
r204 52 79 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=6.67 $Y2=2.72
r205 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=7.065 $Y2=2.72
r206 51 83 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.19 $Y=2.72 $X2=7.59
+ $Y2=2.72
r207 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.19 $Y=2.72
+ $X2=7.065 $Y2=2.72
r208 49 71 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.99 $Y=2.72 $X2=3.91
+ $Y2=2.72
r209 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=2.72
+ $X2=4.155 $Y2=2.72
r210 48 75 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.83 $Y2=2.72
r211 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.155 $Y2=2.72
r212 44 47 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.845 $Y=1.66
+ $X2=9.845 $Y2=2.34
r213 42 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.845 $Y=2.635
+ $X2=9.845 $Y2=2.72
r214 42 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.845 $Y=2.635
+ $X2=9.845 $Y2=2.34
r215 38 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.72
r216 38 40 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.34
r217 34 103 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.72
r218 34 36 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.34
r219 30 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.72
r220 30 32 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.29
r221 26 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.72
r222 26 28 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.34
r223 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r224 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r225 7 47 400 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.845 $X2=9.845 $Y2=2.34
r226 7 44 400 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.845 $X2=9.845 $Y2=1.66
r227 6 110 300 $w=1.7e-07 $l=6.58293e-07 $layer=licon1_PDIFF $count=2 $X=7.73
+ $Y=2.065 $X2=8.265 $Y2=2.34
r228 5 40 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=2.065 $X2=7.025 $Y2=2.34
r229 4 36 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=1.645 $X2=5.14 $Y2=2.34
r230 3 32 600 $w=1.7e-07 $l=3.09233e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=2.065 $X2=4.155 $Y2=2.29
r231 2 28 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=2.065 $X2=2.015 $Y2=2.34
r232 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_448_47# 1 2 8 9 11
c34 8 0 6.94938e-20 $X=2.13 $Y=1.835
r35 9 11 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.215 $Y=0.39
+ $X2=2.375 $Y2=0.39
r36 8 14 22.5629 $w=2.72e-07 $l=5.35635e-07 $layer=LI1_cond $X=2.13 $Y=1.835
+ $X2=2.282 $Y2=2.3
r37 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.215 $Y2=0.39
r38 7 8 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.13 $Y2=1.835
r39 2 14 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.065 $X2=2.435 $Y2=2.3
r40 1 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.375 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%A_651_413# 1 2 9 11 12 15
c36 12 0 1.58851e-19 $X=3.755 $Y=1.95
r37 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.035
+ $X2=4.575 $Y2=2.21
r38 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=4.575 $Y2=2.035
r39 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=3.755 $Y2=1.95
r40 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.755 $Y2=1.95
r41 7 9 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.67 $Y2=2.21
r42 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=2.065 $X2=4.575 $Y2=2.21
r43 1 9 600 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=2.065 $X2=3.67 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%Q 1 2 9 13 15 18 22
r28 15 22 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=8.84 $Y=1.177
+ $X2=8.84 $Y2=1.18
r29 15 18 27.1348 $w=3.28e-07 $l=7.77e-07 $layer=LI1_cond $X=8.84 $Y=1.177
+ $X2=8.84 $Y2=0.4
r30 14 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.84 $Y=1.455
+ $X2=8.84 $Y2=1.18
r31 13 14 5.12431 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=8.802 $Y=1.62
+ $X2=8.802 $Y2=1.455
r32 7 13 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=8.802 $Y=1.657
+ $X2=8.802 $Y2=1.62
r33 7 9 18.2968 $w=4.03e-07 $l=6.43e-07 $layer=LI1_cond $X=8.802 $Y=1.657
+ $X2=8.802 $Y2=2.3
r34 2 13 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=8.55
+ $Y=1.485 $X2=8.685 $Y2=1.62
r35 2 9 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.55
+ $Y=1.485 $X2=8.685 $Y2=2.3
r36 1 18 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.705
+ $Y=0.235 $X2=8.84 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%Q_N 1 2 7 10 12 15 18 22
r16 18 22 0.158442 $w=2.08e-07 $l=3e-09 $layer=LI1_cond $X=10.33 $Y=1.187
+ $X2=10.33 $Y2=1.19
r17 17 22 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=10.33 $Y=1.445
+ $X2=10.33 $Y2=1.19
r18 15 18 20.703 $w=2.08e-07 $l=3.92e-07 $layer=LI1_cond $X=10.33 $Y=0.795
+ $X2=10.33 $Y2=1.187
r19 10 17 6.13261 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=10.307 $Y=1.572
+ $X2=10.307 $Y2=1.445
r20 10 12 11.2081 $w=2.53e-07 $l=2.48e-07 $layer=LI1_cond $X=10.307 $Y=1.572
+ $X2=10.307 $Y2=1.82
r21 7 15 6.13261 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=10.307 $Y=0.668
+ $X2=10.307 $Y2=0.795
r22 7 9 1.81804 $w=2.55e-07 $l=3.8e-08 $layer=LI1_cond $X=10.307 $Y=0.668
+ $X2=10.307 $Y2=0.63
r23 2 12 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=10.13
+ $Y=1.485 $X2=10.265 $Y2=1.82
r24 1 9 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=10.13
+ $Y=0.235 $X2=10.265 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_1%VGND 1 2 3 4 5 6 21 23 27 31 35 39 43 46 47
+ 49 50 52 53 55 56 57 59 90 91 94 97
c156 91 0 2.26487e-19 $X=10.35 $Y=0
r157 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r158 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r159 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r160 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r161 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r162 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r163 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r164 84 87 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r165 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r166 82 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.51
+ $Y2=0
r167 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r168 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r169 78 81 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r170 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r171 76 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r172 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r173 73 76 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.67 $Y2=0
r174 72 75 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.67
+ $Y2=0
r175 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r176 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r177 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r178 67 70 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r179 67 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r180 66 69 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r181 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r182 64 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r183 64 66 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.07 $Y2=0
r184 59 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r185 59 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r186 57 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r187 57 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r188 55 87 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.76 $Y=0 $X2=9.43
+ $Y2=0
r189 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=0 $X2=9.845
+ $Y2=0
r190 54 90 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.93 $Y=0 $X2=10.35
+ $Y2=0
r191 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.93 $Y=0 $X2=9.845
+ $Y2=0
r192 52 81 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.335 $Y=0
+ $X2=8.05 $Y2=0
r193 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=0 $X2=8.42
+ $Y2=0
r194 51 84 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=8.505 $Y=0 $X2=8.51
+ $Y2=0
r195 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.505 $Y=0 $X2=8.42
+ $Y2=0
r196 49 75 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.67
+ $Y2=0
r197 49 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.8
+ $Y2=0
r198 48 78 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.895 $Y=0
+ $X2=7.13 $Y2=0
r199 48 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.895 $Y=0 $X2=6.8
+ $Y2=0
r200 46 69 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r201 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.64
+ $Y2=0
r202 45 72 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.83
+ $Y2=0
r203 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.64
+ $Y2=0
r204 41 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.845 $Y=0.085
+ $X2=9.845 $Y2=0
r205 41 43 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.845 $Y=0.085
+ $X2=9.845 $Y2=0.48
r206 37 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0
r207 37 39 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0.575
r208 33 50 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0
r209 33 35 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0.36
r210 29 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r211 29 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.38
r212 25 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r213 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.36
r214 24 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r215 23 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r216 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=0.845
+ $Y2=0
r217 19 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r218 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r219 6 43 182 $w=1.7e-07 $l=3.30189e-07 $layer=licon1_NDIFF $count=1 $X=9.645
+ $Y=0.235 $X2=9.845 $Y2=0.48
r220 5 39 182 $w=1.7e-07 $l=3.97618e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.235 $X2=8.42 $Y2=0.575
r221 4 35 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.81 $Y2=0.36
r222 3 31 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.64 $Y2=0.38
r223 2 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.71 $Y2=0.36
r224 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


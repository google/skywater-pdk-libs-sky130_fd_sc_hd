* NGSPICE file created from sky130_fd_sc_hd__o22a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VGND A2 a_215_47# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=5.655e+11p ps=5.64e+06u
M1001 a_215_47# B2 a_78_199# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1002 a_78_199# B2 a_292_297# VPB phighvt w=1e+06u l=150000u
+  ad=4.7e+11p pd=2.94e+06u as=2.35e+11p ps=2.47e+06u
M1003 VPWR a_78_199# X VPB phighvt w=1e+06u l=150000u
+  ad=1.005e+12p pd=6.01e+06u as=2.8e+11p ps=2.56e+06u
M1004 a_78_199# B1 a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_215_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_292_297# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_493_297# A2 a_78_199# VPB phighvt w=1e+06u l=150000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1008 VGND a_78_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1009 VPWR A1 a_493_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__o311ai_1.pex.spice
* Created: Thu Aug 27 14:39:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O311AI_1%A1 1 3 6 8 9 16
r23 13 16 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.405 $Y=1.16
+ $X2=0.615 $Y2=1.16
r24 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.16 $X2=0.405 $Y2=1.16
r25 9 14 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.405 $Y2=1.16
r26 8 14 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.23 $Y=1.16
+ $X2=0.405 $Y2=1.16
r27 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=1.325
+ $X2=0.615 $Y2=1.16
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.615 $Y=1.325
+ $X2=0.615 $Y2=1.985
r29 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%A2 1 3 6 8 11
c36 6 0 1.54972e-19 $X=1.035 $Y=1.985
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r38 8 12 0.954422 $w=1.468e-06 $l=1.15e-07 $layer=LI1_cond $X=1.15 $Y=1.73
+ $X2=1.035 $Y2=1.73
r39 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.325
+ $X2=1.035 $Y2=1.16
r40 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.035 $Y=1.325
+ $X2=1.035 $Y2=1.985
r41 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=0.995
+ $X2=1.035 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.035 $Y=0.995
+ $X2=1.035 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%A3 3 6 8 11 13
r31 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.16
+ $X2=1.515 $Y2=1.325
r32 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.16
+ $X2=1.515 $Y2=0.995
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=1.16 $X2=1.515 $Y2=1.16
r34 8 12 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.61 $Y=1.16
+ $X2=1.515 $Y2=1.16
r35 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.455 $Y=1.985
+ $X2=1.455 $Y2=1.325
r36 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.455 $Y=0.56
+ $X2=1.455 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%B1 3 7 8 11 13
r35 11 14 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.16
+ $X2=2.135 $Y2=1.325
r36 11 13 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.16
+ $X2=2.135 $Y2=0.995
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=1.16 $X2=2.115 $Y2=1.16
r38 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.215 $Y=0.56
+ $X2=2.215 $Y2=0.995
r39 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.055 $Y=1.985
+ $X2=2.055 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%C1 1 3 6 8 13
r25 10 13 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.575 $Y=1.16
+ $X2=2.915 $Y2=1.16
r26 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.16 $X2=2.915 $Y2=1.16
r27 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.325
+ $X2=2.575 $Y2=1.16
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.575 $Y=1.325
+ $X2=2.575 $Y2=1.985
r29 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%VPWR 1 2 7 9 15 18 19 20 30 31
c35 9 0 2.94892e-20 $X=0.405 $Y=1.62
r36 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r37 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r38 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r39 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r40 25 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 24 27 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r44 22 34 8.12166 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=0.78 $Y=2.72 $X2=0.39
+ $Y2=2.72
r45 22 24 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.78 $Y=2.72 $X2=1.15
+ $Y2=2.72
r46 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 18 27 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.15 $Y=2.72 $X2=2.07
+ $Y2=2.72
r48 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=2.72
+ $X2=2.315 $Y2=2.72
r49 17 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.48 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=2.72
+ $X2=2.315 $Y2=2.72
r51 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=2.635
+ $X2=2.315 $Y2=2.72
r52 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.315 $Y=2.635
+ $X2=2.315 $Y2=1.96
r53 9 12 11.7026 $w=6.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.432 $Y=1.62
+ $X2=0.432 $Y2=2.3
r54 7 34 2.64475 $w=6.95e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.432 $Y=2.635
+ $X2=0.39 $Y2=2.72
r55 7 12 5.76527 $w=6.93e-07 $l=3.35e-07 $layer=LI1_cond $X=0.432 $Y=2.635
+ $X2=0.432 $Y2=2.3
r56 2 15 300 $w=1.7e-07 $l=5.59911e-07 $layer=licon1_PDIFF $count=2 $X=2.13
+ $Y=1.485 $X2=2.315 $Y2=1.96
r57 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.485 $X2=0.405 $Y2=2.3
r58 1 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.485 $X2=0.405 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%Y 1 2 3 11 14 15 16 18 19 20 21 22 45
c40 14 0 2.94892e-20 $X=1.61 $Y=1.87
c41 11 0 1.54972e-19 $X=1.705 $Y=1.665
r42 63 65 4.88923 $w=5.68e-07 $l=2.33e-07 $layer=LI1_cond $X=2.552 $Y=0.54
+ $X2=2.785 $Y2=0.54
r43 42 63 6.5206 $w=2.15e-07 $l=2.85e-07 $layer=LI1_cond $X=2.552 $Y=0.825
+ $X2=2.552 $Y2=0.54
r44 42 45 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=2.552 $Y=0.825
+ $X2=2.552 $Y2=0.85
r45 22 56 2.21953 $w=4.83e-07 $l=9e-08 $layer=LI1_cond $X=2.892 $Y=2.21
+ $X2=2.892 $Y2=2.3
r46 21 22 8.38488 $w=4.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.892 $Y=1.87
+ $X2=2.892 $Y2=2.21
r47 21 50 5.05559 $w=4.83e-07 $l=2.05e-07 $layer=LI1_cond $X=2.892 $Y=1.87
+ $X2=2.892 $Y2=1.665
r48 20 65 4.30169 $w=5.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.99 $Y=0.54
+ $X2=2.785 $Y2=0.54
r49 19 43 2.73602 $w=3.5e-07 $l=2.77262e-07 $layer=LI1_cond $X=2.79 $Y=1.58
+ $X2=2.552 $Y2=1.495
r50 19 50 2.73602 $w=3.5e-07 $l=1.38109e-07 $layer=LI1_cond $X=2.79 $Y=1.58
+ $X2=2.892 $Y2=1.665
r51 19 43 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=2.552 $Y=1.47
+ $X2=2.552 $Y2=1.495
r52 18 19 15.0086 $w=2.13e-07 $l=2.8e-07 $layer=LI1_cond $X=2.552 $Y=1.19
+ $X2=2.552 $Y2=1.47
r53 16 63 0.461644 $w=5.68e-07 $l=2.2e-08 $layer=LI1_cond $X=2.53 $Y=0.54
+ $X2=2.552 $Y2=0.54
r54 16 18 16.6166 $w=2.13e-07 $l=3.1e-07 $layer=LI1_cond $X=2.552 $Y=0.88
+ $X2=2.552 $Y2=1.19
r55 16 45 1.60806 $w=2.13e-07 $l=3e-08 $layer=LI1_cond $X=2.552 $Y=0.88
+ $X2=2.552 $Y2=0.85
r56 15 40 1.95722 $w=5.48e-07 $l=9e-08 $layer=LI1_cond $X=1.705 $Y=2.21
+ $X2=1.705 $Y2=2.3
r57 14 15 7.39394 $w=5.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.705 $Y=1.87
+ $X2=1.705 $Y2=2.21
r58 11 14 4.45811 $w=5.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=1.87
r59 11 13 2.27723 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=1.58
r60 10 19 19.7147 $w=2.88e-07 $l=4.65e-07 $layer=LI1_cond $X=1.98 $Y=1.58
+ $X2=2.445 $Y2=1.58
r61 10 13 7.3675 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=1.98 $Y=1.58
+ $X2=1.705 $Y2=1.58
r62 3 19 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.485 $X2=2.815 $Y2=1.62
r63 3 56 400 $w=1.7e-07 $l=8.937e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.485 $X2=2.815 $Y2=2.3
r64 2 40 400 $w=1.7e-07 $l=9.20652e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.485 $X2=1.755 $Y2=2.3
r65 2 13 400 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.485 $X2=1.755 $Y2=1.62
r66 1 65 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=2.65
+ $Y=0.235 $X2=2.785 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%VGND 1 2 7 9 11 15 17 24 25 31
r41 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r42 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r43 22 25 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r44 22 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r45 21 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r46 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r47 19 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.245
+ $Y2=0
r48 19 21 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.61
+ $Y2=0
r49 17 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r50 17 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r52 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.36
r53 12 28 6.29768 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.285
+ $Y2=0
r54 11 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=1.245
+ $Y2=0
r55 11 12 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.57
+ $Y2=0
r56 7 28 2.80634 $w=4.85e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.327 $Y=0.085
+ $X2=0.285 $Y2=0
r57 7 9 6.78189 $w=4.83e-07 $l=2.75e-07 $layer=LI1_cond $X=0.327 $Y=0.085
+ $X2=0.327 $Y2=0.36
r58 2 15 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.235 $X2=1.245 $Y2=0.36
r59 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.26
+ $Y=0.235 $X2=0.405 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_1%A_138_47# 1 2 7 10 11 12
r24 12 14 7.89412 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.665 $Y=0.655
+ $X2=1.665 $Y2=0.545
r25 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=0.74
+ $X2=1.665 $Y2=0.655
r26 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.58 $Y=0.74
+ $X2=0.91 $Y2=0.74
r27 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.825 $Y=0.655
+ $X2=0.91 $Y2=0.74
r28 7 9 7.89412 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.825 $Y=0.655
+ $X2=0.825 $Y2=0.545
r29 2 14 182 $w=1.7e-07 $l=3.71416e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.235 $X2=1.665 $Y2=0.545
r30 1 9 182 $w=1.7e-07 $l=3.71416e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.235 $X2=0.825 $Y2=0.545
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__lpflow_inputisolatch_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 0.765000 2.125000 1.095000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.690000 0.415000 4.975000 0.745000 ;
        RECT 4.690000 1.670000 4.975000 2.455000 ;
        RECT 4.805000 0.745000 4.975000 1.670000 ;
    END
  END Q
  PIN SLEEP_B
    ANTENNAGATEAREA  0.145500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.060000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.455000  0.085000 1.785000 0.465000 ;
        RECT 3.265000  0.085000 3.595000 0.530000 ;
        RECT 4.295000  0.085000 4.465000 0.715000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.060000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.455000 2.255000 1.850000 2.635000 ;
        RECT 3.355000 2.135000 3.525000 2.635000 ;
        RECT 4.295000 1.570000 4.465000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.780000 0.805000 ;
      RECT 0.175000 1.795000 0.780000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.610000 0.805000 0.780000 1.130000 ;
      RECT 0.610000 1.130000 0.810000 1.460000 ;
      RECT 0.610000 1.460000 0.780000 1.795000 ;
      RECT 0.980000 0.740000 1.185000 0.910000 ;
      RECT 0.980000 0.910000 1.150000 1.825000 ;
      RECT 0.980000 1.825000 1.185000 1.915000 ;
      RECT 0.980000 1.915000 2.845000 1.965000 ;
      RECT 1.015000 0.345000 1.185000 0.740000 ;
      RECT 1.015000 1.965000 2.845000 2.085000 ;
      RECT 1.015000 2.085000 1.185000 2.465000 ;
      RECT 1.320000 1.240000 1.490000 1.525000 ;
      RECT 1.320000 1.525000 2.335000 1.695000 ;
      RECT 2.050000 1.355000 2.335000 1.525000 ;
      RECT 2.295000 0.705000 2.675000 1.035000 ;
      RECT 2.310000 2.255000 3.185000 2.425000 ;
      RECT 2.380000 0.365000 3.040000 0.535000 ;
      RECT 2.505000 1.035000 2.675000 1.575000 ;
      RECT 2.505000 1.575000 2.845000 1.915000 ;
      RECT 2.870000 0.535000 3.040000 0.995000 ;
      RECT 2.870000 0.995000 3.780000 1.165000 ;
      RECT 3.015000 1.165000 3.780000 1.325000 ;
      RECT 3.015000 1.325000 3.185000 2.255000 ;
      RECT 3.420000 1.535000 4.125000 1.865000 ;
      RECT 3.835000 0.415000 4.125000 0.745000 ;
      RECT 3.835000 1.865000 4.125000 2.435000 ;
      RECT 3.950000 0.745000 4.125000 1.535000 ;
  END
END sky130_fd_sc_hd__lpflow_inputisolatch_1
END LIBRARY

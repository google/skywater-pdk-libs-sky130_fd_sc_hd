* File: sky130_fd_sc_hd__o21ba_4.pxi.spice
* Created: Tue Sep  1 19:22:02 2020
* 
x_PM_SKY130_FD_SC_HD__O21BA_4%B1_N N_B1_N_c_104_n N_B1_N_M1020_g N_B1_N_M1005_g
+ B1_N B1_N N_B1_N_c_106_n N_B1_N_c_107_n PM_SKY130_FD_SC_HD__O21BA_4%B1_N
x_PM_SKY130_FD_SC_HD__O21BA_4%A_187_21# N_A_187_21#_M1012_s N_A_187_21#_M1000_s
+ N_A_187_21#_M1001_s N_A_187_21#_c_145_n N_A_187_21#_M1003_g
+ N_A_187_21#_M1006_g N_A_187_21#_c_146_n N_A_187_21#_M1011_g
+ N_A_187_21#_M1007_g N_A_187_21#_c_147_n N_A_187_21#_M1015_g
+ N_A_187_21#_M1008_g N_A_187_21#_c_148_n N_A_187_21#_M1021_g
+ N_A_187_21#_M1018_g N_A_187_21#_c_149_n N_A_187_21#_c_150_n
+ N_A_187_21#_c_264_p N_A_187_21#_c_170_p N_A_187_21#_c_151_n
+ N_A_187_21#_c_160_n N_A_187_21#_c_279_p N_A_187_21#_c_161_n
+ N_A_187_21#_c_191_p N_A_187_21#_c_152_n N_A_187_21#_c_153_n
+ N_A_187_21#_c_162_n N_A_187_21#_c_154_n PM_SKY130_FD_SC_HD__O21BA_4%A_187_21#
x_PM_SKY130_FD_SC_HD__O21BA_4%A_27_297# N_A_27_297#_M1020_s N_A_27_297#_M1005_s
+ N_A_27_297#_M1000_g N_A_27_297#_M1002_g N_A_27_297#_c_307_n
+ N_A_27_297#_M1012_g N_A_27_297#_c_308_n N_A_27_297#_M1016_g
+ N_A_27_297#_c_314_n N_A_27_297#_c_315_n N_A_27_297#_c_322_n
+ N_A_27_297#_c_381_p N_A_27_297#_c_316_n N_A_27_297#_c_309_n
+ N_A_27_297#_c_317_n N_A_27_297#_c_310_n N_A_27_297#_c_319_n
+ N_A_27_297#_c_320_n N_A_27_297#_c_361_n N_A_27_297#_c_311_n
+ PM_SKY130_FD_SC_HD__O21BA_4%A_27_297#
x_PM_SKY130_FD_SC_HD__O21BA_4%A2 N_A2_c_417_n N_A2_M1010_g N_A2_M1001_g
+ N_A2_c_418_n N_A2_M1017_g N_A2_M1004_g A2 N_A2_c_420_n
+ PM_SKY130_FD_SC_HD__O21BA_4%A2
x_PM_SKY130_FD_SC_HD__O21BA_4%A1 N_A1_c_471_n N_A1_M1013_g N_A1_M1009_g
+ N_A1_c_472_n N_A1_M1014_g N_A1_M1019_g A1 N_A1_c_474_n
+ PM_SKY130_FD_SC_HD__O21BA_4%A1
x_PM_SKY130_FD_SC_HD__O21BA_4%VPWR N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_M1018_d
+ N_VPWR_M1002_d N_VPWR_M1009_s N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n
+ N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n
+ N_VPWR_c_518_n VPWR N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n
+ N_VPWR_c_509_n N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n
+ PM_SKY130_FD_SC_HD__O21BA_4%VPWR
x_PM_SKY130_FD_SC_HD__O21BA_4%X N_X_M1003_s N_X_M1015_s N_X_M1006_s N_X_M1008_s
+ N_X_c_621_n N_X_c_616_n N_X_c_614_n N_X_c_615_n N_X_c_644_n X N_X_c_646_n
+ PM_SKY130_FD_SC_HD__O21BA_4%X
x_PM_SKY130_FD_SC_HD__O21BA_4%A_743_297# N_A_743_297#_M1001_d
+ N_A_743_297#_M1004_d N_A_743_297#_M1019_d N_A_743_297#_c_677_n
+ N_A_743_297#_c_671_n N_A_743_297#_c_697_n N_A_743_297#_c_672_n
+ N_A_743_297#_c_673_n N_A_743_297#_c_674_n N_A_743_297#_c_675_n
+ PM_SKY130_FD_SC_HD__O21BA_4%A_743_297#
x_PM_SKY130_FD_SC_HD__O21BA_4%VGND N_VGND_M1020_d N_VGND_M1011_d N_VGND_M1021_d
+ N_VGND_M1010_d N_VGND_M1013_d N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n
+ N_VGND_c_711_n N_VGND_c_712_n N_VGND_c_713_n N_VGND_c_714_n N_VGND_c_715_n
+ N_VGND_c_716_n N_VGND_c_717_n N_VGND_c_718_n N_VGND_c_719_n VGND
+ N_VGND_c_720_n N_VGND_c_721_n N_VGND_c_722_n N_VGND_c_723_n N_VGND_c_724_n
+ PM_SKY130_FD_SC_HD__O21BA_4%VGND
x_PM_SKY130_FD_SC_HD__O21BA_4%A_575_47# N_A_575_47#_M1012_d N_A_575_47#_M1016_d
+ N_A_575_47#_M1017_s N_A_575_47#_M1014_s N_A_575_47#_c_806_n
+ N_A_575_47#_c_820_n N_A_575_47#_c_807_n N_A_575_47#_c_808_n
+ N_A_575_47#_c_828_n N_A_575_47#_c_809_n N_A_575_47#_c_810_n
+ N_A_575_47#_c_811_n PM_SKY130_FD_SC_HD__O21BA_4%A_575_47#
cc_1 VNB N_B1_N_c_104_n 0.0201252f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_2 VNB B1_N 5.70638e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_3 VNB N_B1_N_c_106_n 0.0251931f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_4 VNB N_B1_N_c_107_n 0.00578081f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.285
cc_5 VNB N_A_187_21#_c_145_n 0.0157563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_187_21#_c_146_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_187_21#_c_147_n 0.0157694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_187_21#_c_148_n 0.0190654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_187_21#_c_149_n 0.00545107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_187_21#_c_150_n 0.00384988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_187_21#_c_151_n 0.00139359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_187_21#_c_152_n 0.00944039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_187_21#_c_153_n 0.00383243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_187_21#_c_154_n 0.0630782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_297#_c_307_n 0.0198994f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.285
cc_16 VNB N_A_27_297#_c_308_n 0.0157572f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.18
cc_17 VNB N_A_27_297#_c_309_n 0.0265255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_310_n 0.021622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_311_n 0.0633313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_417_n 0.0159911f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_21 VNB N_A2_c_418_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_22 VNB A2 0.01232f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.285
cc_23 VNB N_A2_c_420_n 0.0303172f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.18
cc_24 VNB N_A1_c_471_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_25 VNB N_A1_c_472_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_26 VNB A1 0.029484f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.285
cc_27 VNB N_A1_c_474_n 0.0372858f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.18
cc_28 VNB N_VPWR_c_509_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_614_n 0.00482774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_708_n 0.00599858f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.18
cc_31 VNB N_VGND_c_709_n 0.0173082f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.18
cc_32 VNB N_VGND_c_710_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_711_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_712_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_713_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_714_n 0.0206707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_715_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_716_n 0.0380087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_717_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_718_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_719_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_720_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_721_n 0.0235448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_722_n 0.306194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_723_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_724_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_575_47#_c_806_n 0.00339908f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_48 VNB N_A_575_47#_c_807_n 0.00297087f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.18
cc_49 VNB N_A_575_47#_c_808_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_575_47#_c_809_n 0.0130752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_575_47#_c_810_n 0.0183327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_575_47#_c_811_n 0.00253348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_B1_N_M1005_g 0.0224726f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.985
cc_54 VPB B1_N 0.00104379f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_55 VPB N_B1_N_c_106_n 0.00487448f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_56 VPB N_A_187_21#_M1006_g 0.0178181f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.285
cc_57 VPB N_A_187_21#_M1007_g 0.0173952f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.18
cc_58 VPB N_A_187_21#_M1008_g 0.0178805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_187_21#_M1018_g 0.0183444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_187_21#_c_151_n 0.00753731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_187_21#_c_160_n 0.00435473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_187_21#_c_161_n 0.00282418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_187_21#_c_162_n 0.0029376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_187_21#_c_154_n 0.010536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_297#_M1000_g 0.0176165f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_66 VPB N_A_27_297#_M1002_g 0.0220732f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_67 VPB N_A_27_297#_c_314_n 0.00956215f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_297#_c_315_n 0.0168446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_297#_c_316_n 0.00143124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_297#_c_317_n 0.00982375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_297#_c_310_n 0.00715877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_297#_c_319_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_297#_c_320_n 0.00327011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_297#_c_311_n 0.0217529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A2_M1001_g 0.0226275f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.985
cc_76 VPB N_A2_M1004_g 0.0188152f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_77 VPB N_A2_c_420_n 0.00410845f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.18
cc_78 VPB N_A1_M1009_g 0.0182767f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.985
cc_79 VPB N_A1_M1019_g 0.0250431f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_80 VPB N_A1_c_474_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.18
cc_81 VPB N_VPWR_c_510_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.18
cc_82 VPB N_VPWR_c_511_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_512_n 3.09829e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_513_n 0.00751304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_514_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_515_n 0.0142092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_516_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_517_n 0.034906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_518_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_519_n 0.0119877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_520_n 0.0119877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_521_n 0.0212809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_509_n 0.0550435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_523_n 0.0215642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_524_n 0.0043639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_525_n 0.0043639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_X_c_615_n 0.0048153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_743_297#_c_671_n 0.00185659f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_99 VPB N_A_743_297#_c_672_n 0.00330301f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_100 VPB N_A_743_297#_c_673_n 0.0116465f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.53
cc_101 VPB N_A_743_297#_c_674_n 0.0307403f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.18
cc_102 VPB N_A_743_297#_c_675_n 0.00347836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 N_B1_N_c_104_n N_A_187_21#_c_145_n 0.0115065f $X=0.59 $Y=0.995 $X2=0
+ $Y2=0
cc_104 N_B1_N_M1005_g N_A_187_21#_M1006_g 0.0411668f $X=0.59 $Y=1.985 $X2=0
+ $Y2=0
cc_105 B1_N N_A_187_21#_c_154_n 0.00237504f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_106 N_B1_N_c_106_n N_A_187_21#_c_154_n 0.0219715f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B1_N_c_107_n N_A_187_21#_c_154_n 0.00171241f $X=0.745 $Y=1.285 $X2=0
+ $Y2=0
cc_108 N_B1_N_M1005_g N_A_27_297#_c_322_n 0.0107479f $X=0.59 $Y=1.985 $X2=0
+ $Y2=0
cc_109 B1_N N_A_27_297#_c_322_n 0.0165277f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_110 N_B1_N_c_106_n N_A_27_297#_c_322_n 9.55259e-19 $X=0.59 $Y=1.16 $X2=0
+ $Y2=0
cc_111 N_B1_N_c_107_n N_A_27_297#_c_322_n 0.0036428f $X=0.745 $Y=1.285 $X2=0
+ $Y2=0
cc_112 N_B1_N_c_104_n N_A_27_297#_c_309_n 0.00686851f $X=0.59 $Y=0.995 $X2=0
+ $Y2=0
cc_113 N_B1_N_c_106_n N_A_27_297#_c_309_n 0.00126681f $X=0.59 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_B1_N_c_107_n N_A_27_297#_c_309_n 0.00565721f $X=0.745 $Y=1.285 $X2=0
+ $Y2=0
cc_115 N_B1_N_M1005_g N_A_27_297#_c_317_n 0.0051502f $X=0.59 $Y=1.985 $X2=0
+ $Y2=0
cc_116 B1_N N_A_27_297#_c_317_n 0.0192667f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_117 N_B1_N_c_107_n N_A_27_297#_c_317_n 7.71248e-19 $X=0.745 $Y=1.285 $X2=0
+ $Y2=0
cc_118 N_B1_N_c_104_n N_A_27_297#_c_310_n 0.00278251f $X=0.59 $Y=0.995 $X2=0
+ $Y2=0
cc_119 N_B1_N_M1005_g N_A_27_297#_c_310_n 0.00149506f $X=0.59 $Y=1.985 $X2=0
+ $Y2=0
cc_120 B1_N N_A_27_297#_c_310_n 0.00517662f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_121 N_B1_N_c_106_n N_A_27_297#_c_310_n 0.0051685f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B1_N_c_107_n N_A_27_297#_c_310_n 0.0170112f $X=0.745 $Y=1.285 $X2=0
+ $Y2=0
cc_123 B1_N N_VPWR_M1005_d 0.00202248f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_124 N_B1_N_M1005_g N_VPWR_c_510_n 0.00894936f $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_125 N_B1_N_M1005_g N_VPWR_c_509_n 0.00507315f $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B1_N_M1005_g N_VPWR_c_523_n 0.00343969f $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B1_N_c_104_n N_X_c_616_n 4.35972e-19 $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_N_M1005_g N_X_c_616_n 2.8323e-19 $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_129 B1_N N_X_c_616_n 0.0251407f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_130 N_B1_N_c_106_n N_X_c_616_n 6.22443e-19 $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B1_N_c_107_n N_X_c_616_n 0.0172195f $X=0.745 $Y=1.285 $X2=0 $Y2=0
cc_132 N_B1_N_c_104_n N_VGND_c_708_n 0.00314514f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B1_N_c_106_n N_VGND_c_708_n 2.31083e-19 $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B1_N_c_107_n N_VGND_c_708_n 0.0143616f $X=0.745 $Y=1.285 $X2=0 $Y2=0
cc_135 N_B1_N_c_104_n N_VGND_c_714_n 0.00541763f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B1_N_c_104_n N_VGND_c_722_n 0.0105802f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_187_21#_M1018_g N_A_27_297#_M1000_g 0.0273366f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_187_21#_c_170_p N_A_27_297#_M1002_g 0.0150844f $X=3.395 $Y=1.88 $X2=0
+ $Y2=0
cc_139 N_A_187_21#_c_151_n N_A_27_297#_M1002_g 0.0121993f $X=3.49 $Y=1.795 $X2=0
+ $Y2=0
cc_140 N_A_187_21#_c_150_n N_A_27_297#_c_307_n 0.00223484f $X=2.48 $Y=1.075
+ $X2=0 $Y2=0
cc_141 N_A_187_21#_c_151_n N_A_27_297#_c_307_n 0.00225935f $X=3.49 $Y=1.795
+ $X2=0 $Y2=0
cc_142 N_A_187_21#_c_152_n N_A_27_297#_c_307_n 0.0114939f $X=3.235 $Y=0.77 $X2=0
+ $Y2=0
cc_143 N_A_187_21#_c_153_n N_A_27_297#_c_307_n 0.00731515f $X=3.49 $Y=0.77 $X2=0
+ $Y2=0
cc_144 N_A_187_21#_c_151_n N_A_27_297#_c_308_n 0.00249591f $X=3.49 $Y=1.795
+ $X2=0 $Y2=0
cc_145 N_A_187_21#_c_153_n N_A_27_297#_c_308_n 0.00317808f $X=3.49 $Y=0.77 $X2=0
+ $Y2=0
cc_146 N_A_187_21#_M1006_g N_A_27_297#_c_322_n 0.0151951f $X=1.01 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_187_21#_M1007_g N_A_27_297#_c_322_n 0.0115714f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_187_21#_M1008_g N_A_27_297#_c_322_n 0.011545f $X=1.85 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_187_21#_M1018_g N_A_27_297#_c_322_n 0.0127454f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_187_21#_c_149_n N_A_27_297#_c_322_n 0.00368939f $X=2.395 $Y=1.175
+ $X2=0 $Y2=0
cc_151 N_A_187_21#_c_154_n N_A_27_297#_c_322_n 2.8637e-19 $X=2.27 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_187_21#_c_149_n N_A_27_297#_c_316_n 0.00242013f $X=2.395 $Y=1.175
+ $X2=0 $Y2=0
cc_153 N_A_187_21#_c_151_n N_A_27_297#_c_316_n 0.00666062f $X=3.49 $Y=1.795
+ $X2=0 $Y2=0
cc_154 N_A_187_21#_c_154_n N_A_27_297#_c_316_n 9.14342e-19 $X=2.27 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_187_21#_M1000_s N_A_27_297#_c_320_n 0.00262202f $X=2.765 $Y=1.485
+ $X2=0 $Y2=0
cc_156 N_A_187_21#_M1018_g N_A_27_297#_c_320_n 8.29582e-19 $X=2.27 $Y=1.985
+ $X2=0 $Y2=0
cc_157 N_A_187_21#_c_149_n N_A_27_297#_c_320_n 0.0141093f $X=2.395 $Y=1.175
+ $X2=0 $Y2=0
cc_158 N_A_187_21#_c_151_n N_A_27_297#_c_320_n 0.0062361f $X=3.49 $Y=1.795 $X2=0
+ $Y2=0
cc_159 N_A_187_21#_c_191_p N_A_27_297#_c_320_n 0.0064623f $X=2.9 $Y=1.96 $X2=0
+ $Y2=0
cc_160 N_A_187_21#_c_152_n N_A_27_297#_c_320_n 0.00517996f $X=3.235 $Y=0.77
+ $X2=0 $Y2=0
cc_161 N_A_187_21#_c_149_n N_A_27_297#_c_361_n 0.0144242f $X=2.395 $Y=1.175
+ $X2=0 $Y2=0
cc_162 N_A_187_21#_c_170_p N_A_27_297#_c_361_n 0.00321827f $X=3.395 $Y=1.88
+ $X2=0 $Y2=0
cc_163 N_A_187_21#_c_151_n N_A_27_297#_c_361_n 0.00877872f $X=3.49 $Y=1.795
+ $X2=0 $Y2=0
cc_164 N_A_187_21#_c_191_p N_A_27_297#_c_361_n 0.00239623f $X=2.9 $Y=1.96 $X2=0
+ $Y2=0
cc_165 N_A_187_21#_c_152_n N_A_27_297#_c_361_n 0.0274042f $X=3.235 $Y=0.77 $X2=0
+ $Y2=0
cc_166 N_A_187_21#_c_149_n N_A_27_297#_c_311_n 0.00200447f $X=2.395 $Y=1.175
+ $X2=0 $Y2=0
cc_167 N_A_187_21#_c_150_n N_A_27_297#_c_311_n 0.00203264f $X=2.48 $Y=1.075
+ $X2=0 $Y2=0
cc_168 N_A_187_21#_c_170_p N_A_27_297#_c_311_n 0.00556689f $X=3.395 $Y=1.88
+ $X2=0 $Y2=0
cc_169 N_A_187_21#_c_151_n N_A_27_297#_c_311_n 0.02349f $X=3.49 $Y=1.795 $X2=0
+ $Y2=0
cc_170 N_A_187_21#_c_160_n N_A_27_297#_c_311_n 0.00362047f $X=4.135 $Y=1.88
+ $X2=0 $Y2=0
cc_171 N_A_187_21#_c_191_p N_A_27_297#_c_311_n 8.05175e-19 $X=2.9 $Y=1.96 $X2=0
+ $Y2=0
cc_172 N_A_187_21#_c_152_n N_A_27_297#_c_311_n 0.0150796f $X=3.235 $Y=0.77 $X2=0
+ $Y2=0
cc_173 N_A_187_21#_c_153_n N_A_27_297#_c_311_n 0.00133833f $X=3.49 $Y=0.77 $X2=0
+ $Y2=0
cc_174 N_A_187_21#_c_154_n N_A_27_297#_c_311_n 0.0273366f $X=2.27 $Y=1.16 $X2=0
+ $Y2=0
cc_175 N_A_187_21#_c_151_n N_A2_c_417_n 9.16473e-19 $X=3.49 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_187_21#_c_151_n N_A2_M1001_g 0.00944522f $X=3.49 $Y=1.795 $X2=0 $Y2=0
cc_177 N_A_187_21#_c_160_n N_A2_M1001_g 0.0130673f $X=4.135 $Y=1.88 $X2=0 $Y2=0
cc_178 N_A_187_21#_c_161_n N_A2_M1001_g 5.31742e-19 $X=4.26 $Y=1.62 $X2=0 $Y2=0
cc_179 N_A_187_21#_c_161_n N_A2_M1004_g 5.18373e-19 $X=4.26 $Y=1.62 $X2=0 $Y2=0
cc_180 N_A_187_21#_c_151_n A2 0.014517f $X=3.49 $Y=1.795 $X2=0 $Y2=0
cc_181 N_A_187_21#_c_160_n A2 0.00991001f $X=4.135 $Y=1.88 $X2=0 $Y2=0
cc_182 N_A_187_21#_c_161_n A2 0.0198182f $X=4.26 $Y=1.62 $X2=0 $Y2=0
cc_183 N_A_187_21#_c_151_n N_A2_c_420_n 4.47591e-19 $X=3.49 $Y=1.795 $X2=0 $Y2=0
cc_184 N_A_187_21#_c_161_n N_A2_c_420_n 0.00222344f $X=4.26 $Y=1.62 $X2=0 $Y2=0
cc_185 N_A_187_21#_c_170_p N_VPWR_M1002_d 0.00413196f $X=3.395 $Y=1.88 $X2=0
+ $Y2=0
cc_186 N_A_187_21#_c_151_n N_VPWR_M1002_d 0.00467465f $X=3.49 $Y=1.795 $X2=0
+ $Y2=0
cc_187 N_A_187_21#_c_162_n N_VPWR_M1002_d 0.00100143f $X=3.49 $Y=1.88 $X2=0
+ $Y2=0
cc_188 N_A_187_21#_M1006_g N_VPWR_c_510_n 0.00877207f $X=1.01 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_187_21#_M1007_g N_VPWR_c_510_n 0.00122022f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_187_21#_M1006_g N_VPWR_c_511_n 0.00122022f $X=1.01 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_187_21#_M1007_g N_VPWR_c_511_n 0.00880597f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_187_21#_M1008_g N_VPWR_c_511_n 0.00880597f $X=1.85 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_187_21#_M1018_g N_VPWR_c_511_n 0.00122022f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_187_21#_M1008_g N_VPWR_c_512_n 0.00122022f $X=1.85 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_187_21#_M1018_g N_VPWR_c_512_n 0.00877207f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_187_21#_c_170_p N_VPWR_c_513_n 0.0120305f $X=3.395 $Y=1.88 $X2=0
+ $Y2=0
cc_197 N_A_187_21#_c_162_n N_VPWR_c_513_n 0.00467627f $X=3.49 $Y=1.88 $X2=0
+ $Y2=0
cc_198 N_A_187_21#_c_170_p N_VPWR_c_515_n 0.00233924f $X=3.395 $Y=1.88 $X2=0
+ $Y2=0
cc_199 N_A_187_21#_c_191_p N_VPWR_c_515_n 0.0113839f $X=2.9 $Y=1.96 $X2=0 $Y2=0
cc_200 N_A_187_21#_c_160_n N_VPWR_c_517_n 0.00145432f $X=4.135 $Y=1.88 $X2=0
+ $Y2=0
cc_201 N_A_187_21#_c_162_n N_VPWR_c_517_n 0.00216841f $X=3.49 $Y=1.88 $X2=0
+ $Y2=0
cc_202 N_A_187_21#_M1006_g N_VPWR_c_519_n 0.00343969f $X=1.01 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_187_21#_M1007_g N_VPWR_c_519_n 0.00343969f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_187_21#_M1008_g N_VPWR_c_520_n 0.00343969f $X=1.85 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_187_21#_M1018_g N_VPWR_c_520_n 0.00343969f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_187_21#_M1000_s N_VPWR_c_509_n 0.00414531f $X=2.765 $Y=1.485 $X2=0
+ $Y2=0
cc_207 N_A_187_21#_M1001_s N_VPWR_c_509_n 0.00216833f $X=4.125 $Y=1.485 $X2=0
+ $Y2=0
cc_208 N_A_187_21#_M1006_g N_VPWR_c_509_n 0.00406573f $X=1.01 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_187_21#_M1007_g N_VPWR_c_509_n 0.00406573f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_187_21#_M1008_g N_VPWR_c_509_n 0.00406573f $X=1.85 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_187_21#_M1018_g N_VPWR_c_509_n 0.00406573f $X=2.27 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_187_21#_c_170_p N_VPWR_c_509_n 0.00541437f $X=3.395 $Y=1.88 $X2=0
+ $Y2=0
cc_213 N_A_187_21#_c_160_n N_VPWR_c_509_n 0.00352596f $X=4.135 $Y=1.88 $X2=0
+ $Y2=0
cc_214 N_A_187_21#_c_191_p N_VPWR_c_509_n 0.00646745f $X=2.9 $Y=1.96 $X2=0 $Y2=0
cc_215 N_A_187_21#_c_162_n N_VPWR_c_509_n 0.00397985f $X=3.49 $Y=1.88 $X2=0
+ $Y2=0
cc_216 N_A_187_21#_c_145_n N_X_c_621_n 0.00513121f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_187_21#_c_146_n N_X_c_621_n 0.00630972f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_187_21#_c_147_n N_X_c_621_n 5.22228e-19 $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_187_21#_c_145_n N_X_c_616_n 0.00268639f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_187_21#_M1006_g N_X_c_616_n 0.0061917f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_187_21#_c_146_n N_X_c_616_n 0.00314877f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_187_21#_M1007_g N_X_c_616_n 0.00852169f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_187_21#_c_147_n N_X_c_616_n 5.00581e-19 $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_187_21#_M1008_g N_X_c_616_n 6.70404e-19 $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_187_21#_c_149_n N_X_c_616_n 0.0160283f $X=2.395 $Y=1.175 $X2=0 $Y2=0
cc_226 N_A_187_21#_c_154_n N_X_c_616_n 0.0288901f $X=2.27 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_187_21#_c_146_n N_X_c_614_n 0.00535291f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_187_21#_c_147_n N_X_c_614_n 0.0098365f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_187_21#_c_148_n N_X_c_614_n 0.0026237f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_187_21#_c_149_n N_X_c_614_n 0.0456865f $X=2.395 $Y=1.175 $X2=0 $Y2=0
cc_231 N_A_187_21#_c_150_n N_X_c_614_n 7.61274e-19 $X=2.48 $Y=1.075 $X2=0 $Y2=0
cc_232 N_A_187_21#_c_264_p N_X_c_614_n 0.00761667f $X=2.565 $Y=0.81 $X2=0 $Y2=0
cc_233 N_A_187_21#_c_154_n N_X_c_614_n 0.00465913f $X=2.27 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_187_21#_M1007_g N_X_c_615_n 0.00608909f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_187_21#_M1008_g N_X_c_615_n 0.0112182f $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A_187_21#_M1018_g N_X_c_615_n 0.00395702f $X=2.27 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A_187_21#_c_149_n N_X_c_615_n 0.0442241f $X=2.395 $Y=1.175 $X2=0 $Y2=0
cc_238 N_A_187_21#_c_154_n N_X_c_615_n 0.00446399f $X=2.27 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_187_21#_c_145_n N_X_c_644_n 0.00210721f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_187_21#_c_146_n N_X_c_644_n 0.00367224f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_187_21#_c_146_n N_X_c_646_n 5.22228e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_187_21#_c_147_n N_X_c_646_n 0.00630972f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_187_21#_c_148_n N_X_c_646_n 0.0109231f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_187_21#_c_160_n N_A_743_297#_M1001_d 0.00788247f $X=4.135 $Y=1.88
+ $X2=-0.19 $Y2=-0.24
cc_245 N_A_187_21#_M1001_s N_A_743_297#_c_677_n 0.00312348f $X=4.125 $Y=1.485
+ $X2=0 $Y2=0
cc_246 N_A_187_21#_c_160_n N_A_743_297#_c_677_n 0.00520504f $X=4.135 $Y=1.88
+ $X2=0 $Y2=0
cc_247 N_A_187_21#_c_279_p N_A_743_297#_c_677_n 0.0118865f $X=4.257 $Y=1.795
+ $X2=0 $Y2=0
cc_248 N_A_187_21#_c_161_n N_A_743_297#_c_671_n 0.0021265f $X=4.26 $Y=1.62 $X2=0
+ $Y2=0
cc_249 N_A_187_21#_c_160_n N_A_743_297#_c_675_n 0.0173385f $X=4.135 $Y=1.88
+ $X2=0 $Y2=0
cc_250 N_A_187_21#_c_264_p N_VGND_M1021_d 0.00315479f $X=2.565 $Y=0.81 $X2=0
+ $Y2=0
cc_251 N_A_187_21#_c_152_n N_VGND_M1021_d 0.00109197f $X=3.235 $Y=0.77 $X2=0
+ $Y2=0
cc_252 N_A_187_21#_c_145_n N_VGND_c_708_n 0.00159991f $X=1.01 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A_187_21#_c_145_n N_VGND_c_709_n 0.00541359f $X=1.01 $Y=0.995 $X2=0
+ $Y2=0
cc_254 N_A_187_21#_c_146_n N_VGND_c_709_n 0.0042327f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_255 N_A_187_21#_c_146_n N_VGND_c_710_n 0.00146448f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_256 N_A_187_21#_c_147_n N_VGND_c_710_n 0.00146448f $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A_187_21#_c_148_n N_VGND_c_711_n 0.00316354f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A_187_21#_c_264_p N_VGND_c_711_n 0.0137999f $X=2.565 $Y=0.81 $X2=0
+ $Y2=0
cc_259 N_A_187_21#_c_152_n N_VGND_c_716_n 0.00361289f $X=3.235 $Y=0.77 $X2=0
+ $Y2=0
cc_260 N_A_187_21#_c_147_n N_VGND_c_720_n 0.00423334f $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_261 N_A_187_21#_c_148_n N_VGND_c_720_n 0.00541359f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_187_21#_M1012_s N_VGND_c_722_n 0.00216833f $X=3.285 $Y=0.235 $X2=0
+ $Y2=0
cc_263 N_A_187_21#_c_145_n N_VGND_c_722_n 0.00952874f $X=1.01 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_187_21#_c_146_n N_VGND_c_722_n 0.00571514f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_187_21#_c_147_n N_VGND_c_722_n 0.0057163f $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_266 N_A_187_21#_c_148_n N_VGND_c_722_n 0.0108276f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A_187_21#_c_264_p N_VGND_c_722_n 7.10978e-19 $X=2.565 $Y=0.81 $X2=0
+ $Y2=0
cc_268 N_A_187_21#_c_152_n N_VGND_c_722_n 0.00731837f $X=3.235 $Y=0.77 $X2=0
+ $Y2=0
cc_269 N_A_187_21#_c_152_n N_A_575_47#_M1012_d 0.00319477f $X=3.235 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_270 N_A_187_21#_M1012_s N_A_575_47#_c_806_n 0.00305026f $X=3.285 $Y=0.235
+ $X2=0 $Y2=0
cc_271 N_A_187_21#_c_152_n N_A_575_47#_c_806_n 0.0187482f $X=3.235 $Y=0.77 $X2=0
+ $Y2=0
cc_272 N_A_187_21#_c_153_n N_A_575_47#_c_806_n 0.0166477f $X=3.49 $Y=0.77 $X2=0
+ $Y2=0
cc_273 N_A_187_21#_c_151_n N_A_575_47#_c_807_n 8.1259e-19 $X=3.49 $Y=1.795 $X2=0
+ $Y2=0
cc_274 N_A_187_21#_c_153_n N_A_575_47#_c_807_n 0.00752753f $X=3.49 $Y=0.77 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_c_308_n N_A2_c_417_n 0.0145082f $X=3.63 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_276 N_A_27_297#_c_311_n A2 0.00194074f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_27_297#_c_311_n N_A2_c_420_n 0.0145082f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_278 N_A_27_297#_c_322_n N_VPWR_M1005_d 0.00323291f $X=2.395 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_279 N_A_27_297#_c_322_n N_VPWR_M1007_d 0.00317502f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_280 N_A_27_297#_c_322_n N_VPWR_M1018_d 0.00194131f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_281 N_A_27_297#_c_381_p N_VPWR_M1018_d 7.41903e-19 $X=2.48 $Y=1.875 $X2=0
+ $Y2=0
cc_282 N_A_27_297#_c_320_n N_VPWR_M1018_d 6.75483e-19 $X=2.82 $Y=1.53 $X2=0
+ $Y2=0
cc_283 N_A_27_297#_c_315_n N_VPWR_c_510_n 0.0172022f $X=0.35 $Y=2.3 $X2=0 $Y2=0
cc_284 N_A_27_297#_c_322_n N_VPWR_c_510_n 0.0161563f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_285 N_A_27_297#_c_322_n N_VPWR_c_511_n 0.0161563f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_286 N_A_27_297#_M1000_g N_VPWR_c_512_n 0.00754047f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_287 N_A_27_297#_M1002_g N_VPWR_c_512_n 5.39334e-19 $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_27_297#_c_322_n N_VPWR_c_512_n 0.0149407f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_289 N_A_27_297#_c_320_n N_VPWR_c_512_n 7.52316e-19 $X=2.82 $Y=1.53 $X2=0
+ $Y2=0
cc_290 N_A_27_297#_M1002_g N_VPWR_c_513_n 0.00329978f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_M1000_g N_VPWR_c_515_n 0.0046653f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_292 N_A_27_297#_M1002_g N_VPWR_c_515_n 0.00441875f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_293 N_A_27_297#_c_322_n N_VPWR_c_519_n 0.00707682f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_294 N_A_27_297#_c_322_n N_VPWR_c_520_n 0.00707682f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_295 N_A_27_297#_M1005_s N_VPWR_c_509_n 0.00340315f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_296 N_A_27_297#_M1000_g N_VPWR_c_509_n 0.00789179f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_A_27_297#_M1002_g N_VPWR_c_509_n 0.0071988f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_27_297#_c_315_n N_VPWR_c_509_n 0.0134021f $X=0.35 $Y=2.3 $X2=0 $Y2=0
cc_299 N_A_27_297#_c_322_n N_VPWR_c_509_n 0.0343704f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_300 N_A_27_297#_c_315_n N_VPWR_c_523_n 0.0245389f $X=0.35 $Y=2.3 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_322_n N_VPWR_c_523_n 0.00264208f $X=2.395 $Y=1.96 $X2=0
+ $Y2=0
cc_302 N_A_27_297#_c_322_n N_X_M1006_s 0.00440982f $X=2.395 $Y=1.96 $X2=0 $Y2=0
cc_303 N_A_27_297#_c_322_n N_X_M1008_s 0.00441351f $X=2.395 $Y=1.96 $X2=0 $Y2=0
cc_304 N_A_27_297#_c_322_n N_X_c_616_n 0.0224262f $X=2.395 $Y=1.96 $X2=0 $Y2=0
cc_305 N_A_27_297#_c_322_n N_X_c_615_n 0.0394127f $X=2.395 $Y=1.96 $X2=0 $Y2=0
cc_306 N_A_27_297#_c_320_n N_X_c_615_n 0.00881439f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_307 N_A_27_297#_c_307_n N_VGND_c_711_n 0.0019578f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_27_297#_c_309_n N_VGND_c_714_n 0.0283284f $X=0.38 $Y=0.39 $X2=0 $Y2=0
cc_309 N_A_27_297#_c_307_n N_VGND_c_716_n 0.00357877f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_A_27_297#_c_308_n N_VGND_c_716_n 0.00357877f $X=3.63 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_A_27_297#_M1020_s N_VGND_c_722_n 0.00246589f $X=0.21 $Y=0.235 $X2=0
+ $Y2=0
cc_312 N_A_27_297#_c_307_n N_VGND_c_722_n 0.00655123f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_A_27_297#_c_308_n N_VGND_c_722_n 0.00525237f $X=3.63 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_27_297#_c_309_n N_VGND_c_722_n 0.0173073f $X=0.38 $Y=0.39 $X2=0 $Y2=0
cc_315 N_A_27_297#_c_307_n N_A_575_47#_c_806_n 0.00924081f $X=3.21 $Y=0.995
+ $X2=0 $Y2=0
cc_316 N_A_27_297#_c_308_n N_A_575_47#_c_806_n 0.0126889f $X=3.63 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A2_c_418_n N_A1_c_471_n 0.0150516f $X=4.47 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_318 N_A2_M1004_g N_A1_M1009_g 0.0150516f $X=4.47 $Y=1.985 $X2=0 $Y2=0
cc_319 A2 A1 0.0167609f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_320 A2 N_A1_c_474_n 0.00538113f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_321 N_A2_c_420_n N_A1_c_474_n 0.0150516f $X=4.47 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A2_M1001_g N_VPWR_c_513_n 0.00216743f $X=4.05 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A2_M1004_g N_VPWR_c_514_n 0.00110007f $X=4.47 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A2_M1001_g N_VPWR_c_517_n 0.00357877f $X=4.05 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A2_M1004_g N_VPWR_c_517_n 0.00357877f $X=4.47 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A2_M1001_g N_VPWR_c_509_n 0.00655123f $X=4.05 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A2_M1004_g N_VPWR_c_509_n 0.00525237f $X=4.47 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A2_M1001_g N_A_743_297#_c_677_n 0.00846708f $X=4.05 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A2_M1004_g N_A_743_297#_c_677_n 0.0121306f $X=4.47 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A2_M1004_g N_A_743_297#_c_671_n 2.63949e-19 $X=4.47 $Y=1.985 $X2=0
+ $Y2=0
cc_331 A2 N_A_743_297#_c_671_n 0.0139423f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_332 A2 N_A_743_297#_c_672_n 0.00401644f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_333 N_A2_c_417_n N_VGND_c_712_n 0.00268723f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A2_c_418_n N_VGND_c_712_n 0.00146448f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A2_c_417_n N_VGND_c_716_n 0.00421816f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A2_c_418_n N_VGND_c_718_n 0.00423334f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A2_c_417_n N_VGND_c_722_n 0.00575258f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A2_c_418_n N_VGND_c_722_n 0.0057435f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A2_c_417_n N_A_575_47#_c_820_n 0.00255288f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A2_c_417_n N_A_575_47#_c_807_n 0.0048497f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A2_c_418_n N_A_575_47#_c_807_n 4.58193e-19 $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_342 A2 N_A_575_47#_c_807_n 0.0188951f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_343 N_A2_c_417_n N_A_575_47#_c_808_n 0.00870364f $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A2_c_418_n N_A_575_47#_c_808_n 0.00865686f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_345 A2 N_A_575_47#_c_808_n 0.036111f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_346 N_A2_c_420_n N_A_575_47#_c_808_n 0.00222133f $X=4.47 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A2_c_417_n N_A_575_47#_c_828_n 5.22228e-19 $X=4.05 $Y=0.995 $X2=0 $Y2=0
cc_348 N_A2_c_418_n N_A_575_47#_c_828_n 0.00630972f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A2_c_418_n N_A_575_47#_c_811_n 0.00112787f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_350 A2 N_A_575_47#_c_811_n 0.025661f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_351 N_A1_M1009_g N_VPWR_c_514_n 0.0122146f $X=4.89 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A1_M1019_g N_VPWR_c_514_n 0.0129691f $X=5.31 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A1_M1009_g N_VPWR_c_517_n 0.0046653f $X=4.89 $Y=1.985 $X2=0 $Y2=0
cc_354 N_A1_M1019_g N_VPWR_c_521_n 0.0046653f $X=5.31 $Y=1.985 $X2=0 $Y2=0
cc_355 N_A1_M1009_g N_VPWR_c_509_n 0.007919f $X=4.89 $Y=1.985 $X2=0 $Y2=0
cc_356 N_A1_M1019_g N_VPWR_c_509_n 0.00899032f $X=5.31 $Y=1.985 $X2=0 $Y2=0
cc_357 N_A1_M1009_g N_A_743_297#_c_672_n 0.0152988f $X=4.89 $Y=1.985 $X2=0 $Y2=0
cc_358 N_A1_M1019_g N_A_743_297#_c_672_n 0.0138201f $X=5.31 $Y=1.985 $X2=0 $Y2=0
cc_359 A1 N_A_743_297#_c_672_n 0.0309573f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_360 N_A1_c_474_n N_A_743_297#_c_672_n 0.00213789f $X=5.31 $Y=1.16 $X2=0 $Y2=0
cc_361 A1 N_A_743_297#_c_673_n 0.0225537f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_362 N_A1_c_471_n N_VGND_c_713_n 0.00146448f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_363 N_A1_c_472_n N_VGND_c_713_n 0.00268723f $X=5.31 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A1_c_471_n N_VGND_c_718_n 0.00423334f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A1_c_472_n N_VGND_c_721_n 0.00423737f $X=5.31 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A1_c_471_n N_VGND_c_722_n 0.0057435f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A1_c_472_n N_VGND_c_722_n 0.00681522f $X=5.31 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A1_c_471_n N_A_575_47#_c_828_n 0.00630972f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A1_c_472_n N_A_575_47#_c_828_n 5.22228e-19 $X=5.31 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A1_c_471_n N_A_575_47#_c_809_n 0.0101811f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A1_c_472_n N_A_575_47#_c_809_n 0.0100059f $X=5.31 $Y=0.995 $X2=0 $Y2=0
cc_372 A1 N_A_575_47#_c_809_n 0.0559741f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_373 N_A1_c_474_n N_A_575_47#_c_809_n 0.00222133f $X=5.31 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A1_c_471_n N_A_575_47#_c_810_n 5.18879e-19 $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A1_c_472_n N_A_575_47#_c_810_n 0.00621819f $X=5.31 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A1_c_471_n N_A_575_47#_c_811_n 0.00144553f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_377 N_VPWR_c_509_n N_X_M1006_s 0.00331039f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_509_n N_X_M1008_s 0.00331039f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_M1007_d N_X_c_615_n 0.00168426f $X=1.505 $Y=1.485 $X2=0 $Y2=0
cc_380 N_VPWR_c_509_n N_A_743_297#_M1001_d 0.00208521f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_381 N_VPWR_c_509_n N_A_743_297#_M1004_d 0.00385313f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_509_n N_A_743_297#_M1019_d 0.00399293f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_517_n N_A_743_297#_c_677_n 0.0358391f $X=4.935 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_509_n N_A_743_297#_c_677_n 0.0234464f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_517_n N_A_743_297#_c_697_n 0.0114668f $X=4.935 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_509_n N_A_743_297#_c_697_n 0.006547f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_M1009_s N_A_743_297#_c_672_n 0.00166915f $X=4.965 $Y=1.485 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_514_n N_A_743_297#_c_672_n 0.0172742f $X=5.1 $Y=2 $X2=0 $Y2=0
cc_389 N_VPWR_c_521_n N_A_743_297#_c_674_n 0.019049f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_509_n N_A_743_297#_c_674_n 0.0105137f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_513_n N_A_743_297#_c_675_n 0.0209524f $X=3.32 $Y=2.3 $X2=0 $Y2=0
cc_392 N_VPWR_c_517_n N_A_743_297#_c_675_n 0.0157398f $X=4.935 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_509_n N_A_743_297#_c_675_n 0.00900263f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_X_c_614_n N_VGND_M1011_d 0.00162089f $X=1.895 $Y=0.815 $X2=0 $Y2=0
cc_395 N_X_c_644_n N_VGND_c_708_n 0.00830019f $X=1.255 $Y=0.815 $X2=0 $Y2=0
cc_396 N_X_c_621_n N_VGND_c_709_n 0.0189039f $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_397 N_X_c_614_n N_VGND_c_709_n 0.00104624f $X=1.895 $Y=0.815 $X2=0 $Y2=0
cc_398 N_X_c_644_n N_VGND_c_709_n 0.00103288f $X=1.255 $Y=0.815 $X2=0 $Y2=0
cc_399 N_X_c_614_n N_VGND_c_710_n 0.0122559f $X=1.895 $Y=0.815 $X2=0 $Y2=0
cc_400 N_X_c_614_n N_VGND_c_720_n 0.00198695f $X=1.895 $Y=0.815 $X2=0 $Y2=0
cc_401 N_X_c_646_n N_VGND_c_720_n 0.0188551f $X=2.06 $Y=0.39 $X2=0 $Y2=0
cc_402 N_X_M1003_s N_VGND_c_722_n 0.00215201f $X=1.085 $Y=0.235 $X2=0 $Y2=0
cc_403 N_X_M1015_s N_VGND_c_722_n 0.00215201f $X=1.925 $Y=0.235 $X2=0 $Y2=0
cc_404 N_X_c_621_n N_VGND_c_722_n 0.0122217f $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_405 N_X_c_614_n N_VGND_c_722_n 0.00685338f $X=1.895 $Y=0.815 $X2=0 $Y2=0
cc_406 N_X_c_644_n N_VGND_c_722_n 0.00161088f $X=1.255 $Y=0.815 $X2=0 $Y2=0
cc_407 N_X_c_646_n N_VGND_c_722_n 0.0122069f $X=2.06 $Y=0.39 $X2=0 $Y2=0
cc_408 N_A_743_297#_c_672_n N_A_575_47#_c_809_n 0.00400519f $X=5.435 $Y=1.56
+ $X2=0 $Y2=0
cc_409 N_A_743_297#_c_672_n N_A_575_47#_c_811_n 7.32087e-19 $X=5.435 $Y=1.56
+ $X2=0 $Y2=0
cc_410 N_VGND_c_722_n N_A_575_47#_M1012_d 0.00209344f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_411 N_VGND_c_722_n N_A_575_47#_M1016_d 0.00215206f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_722_n N_A_575_47#_M1017_s 0.00215201f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_722_n N_A_575_47#_M1014_s 0.00226063f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_711_n N_A_575_47#_c_806_n 0.0141428f $X=2.48 $Y=0.39 $X2=0 $Y2=0
cc_415 N_VGND_c_716_n N_A_575_47#_c_806_n 0.0542601f $X=4.175 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_722_n N_A_575_47#_c_806_n 0.034069f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_716_n N_A_575_47#_c_820_n 0.0152108f $X=4.175 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_722_n N_A_575_47#_c_820_n 0.00940698f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_M1010_d N_A_575_47#_c_808_n 0.00162089f $X=4.125 $Y=0.235 $X2=0
+ $Y2=0
cc_420 N_VGND_c_712_n N_A_575_47#_c_808_n 0.0122559f $X=4.26 $Y=0.39 $X2=0 $Y2=0
cc_421 N_VGND_c_716_n N_A_575_47#_c_808_n 0.00198695f $X=4.175 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_718_n N_A_575_47#_c_808_n 0.00198695f $X=5.015 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_722_n N_A_575_47#_c_808_n 0.00835832f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_718_n N_A_575_47#_c_828_n 0.0188551f $X=5.015 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_722_n N_A_575_47#_c_828_n 0.0122069f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_M1013_d N_A_575_47#_c_809_n 0.00162089f $X=4.965 $Y=0.235 $X2=0
+ $Y2=0
cc_427 N_VGND_c_713_n N_A_575_47#_c_809_n 0.0122559f $X=5.1 $Y=0.39 $X2=0 $Y2=0
cc_428 N_VGND_c_718_n N_A_575_47#_c_809_n 0.00198695f $X=5.015 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_721_n N_A_575_47#_c_809_n 0.00198695f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_722_n N_A_575_47#_c_809_n 0.00835832f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_721_n N_A_575_47#_c_810_n 0.0213509f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_722_n N_A_575_47#_c_810_n 0.0133027f $X=5.75 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__and2b_2.spice
* Created: Tue Sep  1 18:57:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and2b_2.pex.spice"
.subckt sky130_fd_sc_hd__and2b_2  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_A_27_413#_M1008_d N_A_N_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_297_47# N_A_27_413#_M1003_g N_A_212_413#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g A_297_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0567 PD=0.777196 PS=0.69 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1002_d N_A_212_413#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.123773 AS=0.08775 PD=1.2028 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_212_413#_M1009_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.08775 PD=1.84 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_27_413#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07665 AS=0.1092 PD=0.785 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1000 N_A_212_413#_M1000_d N_A_27_413#_M1000_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0609 AS=0.07665 PD=0.71 PS=0.785 NRD=2.3443 NRS=42.1974 M=1
+ R=2.8 SA=75000.7 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_212_413#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.135435 AS=0.0609 PD=1.03225 PS=0.71 NRD=21.0987 NRS=2.3443 M=1 R=2.8
+ SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1006_d N_A_212_413#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.322465 AS=0.135 PD=2.45775 PS=1.27 NRD=15.7403 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_212_413#_M1004_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX11_noxref noxref_11 A_N A_N PROBETYPE=1
pX12_noxref noxref_12 A_N A_N PROBETYPE=1
pX13_noxref noxref_13 B B PROBETYPE=1
pX14_noxref noxref_14 X X PROBETYPE=1
pX15_noxref noxref_15 X X PROBETYPE=1
*
.include "sky130_fd_sc_hd__and2b_2.pxi.spice"
*
.ends
*
*

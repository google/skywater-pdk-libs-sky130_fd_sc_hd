* File: sky130_fd_sc_hd__ebufn_8.spice.pex
* Created: Thu Aug 27 14:19:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EBUFN_8%A 1 3 6 8 10 14 16 17
c49 14 0 3.08151e-19 $X=0.925 $Y=1.985
c50 10 0 1.1321e-20 $X=0.925 $Y=0.56
c51 8 0 1.50396e-19 $X=0.925 $Y=1.025
r52 21 23 33.74 $w=3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.295 $Y=1.16 $X2=0.505
+ $Y2=1.16
r53 16 17 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.16
+ $X2=0.257 $Y2=1.53
r54 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.295
+ $Y=1.16 $X2=0.295 $Y2=1.16
r55 8 23 67.48 $w=3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.925 $Y=1.16 $X2=0.505
+ $Y2=1.16
r56 8 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.925 $Y=1.295
+ $X2=0.925 $Y2=1.985
r57 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.925 $Y=1.025
+ $X2=0.925 $Y2=0.56
r58 4 23 18.9685 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.505 $Y2=1.16
r59 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.505 $Y2=1.985
r60 1 23 18.9685 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=0.995
+ $X2=0.505 $Y2=1.16
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.505 $Y=0.995
+ $X2=0.505 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%TE_B 1 3 6 10 12 14 15 17 19 20 22 24 25 27
+ 29 30 32 34 35 37 39 40 42 44 45 47 49 50 51 52 53 54 55 56 57 58 62 63 66 67
r172 65 67 7.05226 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=1.137 $Y=1.325
+ $X2=1.137 $Y2=1.53
r173 64 66 4.98819 $w=3.33e-07 $l=1.45e-07 $layer=LI1_cond $X=1.137 $Y=0.995
+ $X2=1.137 $Y2=0.85
r174 62 65 5.19507 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=1.16
+ $X2=1.2 $Y2=1.325
r175 62 64 5.19507 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=1.16
+ $X2=1.2 $Y2=0.995
r176 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=1.16 $X2=1.345 $Y2=1.16
r177 50 51 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.92 $Y=1.232
+ $X2=2.07 $Y2=1.232
r178 47 49 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.31 $Y=1.47
+ $X2=5.31 $Y2=2.015
r179 46 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.965 $Y=1.395
+ $X2=4.89 $Y2=1.395
r180 45 47 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.235 $Y=1.395
+ $X2=5.31 $Y2=1.47
r181 45 46 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.235 $Y=1.395
+ $X2=4.965 $Y2=1.395
r182 42 58 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.89 $Y=1.47
+ $X2=4.89 $Y2=1.395
r183 42 44 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.89 $Y=1.47
+ $X2=4.89 $Y2=2.015
r184 41 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.545 $Y=1.395
+ $X2=4.47 $Y2=1.395
r185 40 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.815 $Y=1.395
+ $X2=4.89 $Y2=1.395
r186 40 41 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.815 $Y=1.395
+ $X2=4.545 $Y2=1.395
r187 37 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.47 $Y=1.47
+ $X2=4.47 $Y2=1.395
r188 37 39 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.47 $Y=1.47
+ $X2=4.47 $Y2=2.015
r189 36 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.125 $Y=1.395
+ $X2=4.05 $Y2=1.395
r190 35 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.395 $Y=1.395
+ $X2=4.47 $Y2=1.395
r191 35 36 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.395 $Y=1.395
+ $X2=4.125 $Y2=1.395
r192 32 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.05 $Y=1.47
+ $X2=4.05 $Y2=1.395
r193 32 34 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.05 $Y=1.47
+ $X2=4.05 $Y2=2.015
r194 31 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.705 $Y=1.395
+ $X2=3.63 $Y2=1.395
r195 30 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.975 $Y=1.395
+ $X2=4.05 $Y2=1.395
r196 30 31 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.975 $Y=1.395
+ $X2=3.705 $Y2=1.395
r197 27 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.63 $Y=1.47
+ $X2=3.63 $Y2=1.395
r198 27 29 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.63 $Y=1.47
+ $X2=3.63 $Y2=2.015
r199 26 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.395
+ $X2=3.21 $Y2=1.395
r200 25 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.555 $Y=1.395
+ $X2=3.63 $Y2=1.395
r201 25 26 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.555 $Y=1.395
+ $X2=3.285 $Y2=1.395
r202 22 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.21 $Y=1.47
+ $X2=3.21 $Y2=1.395
r203 22 24 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.21 $Y=1.47
+ $X2=3.21 $Y2=2.015
r204 21 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=1.395
+ $X2=2.79 $Y2=1.395
r205 20 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.135 $Y=1.395
+ $X2=3.21 $Y2=1.395
r206 20 21 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.135 $Y=1.395
+ $X2=2.865 $Y2=1.395
r207 17 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.79 $Y=1.47
+ $X2=2.79 $Y2=1.395
r208 17 19 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.79 $Y=1.47
+ $X2=2.79 $Y2=2.015
r209 16 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.395
+ $X2=2.37 $Y2=1.395
r210 15 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.715 $Y=1.395
+ $X2=2.79 $Y2=1.395
r211 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.715 $Y=1.395
+ $X2=2.445 $Y2=1.395
r212 12 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.47
+ $X2=2.37 $Y2=1.395
r213 12 14 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.37 $Y=1.47
+ $X2=2.37 $Y2=2.015
r214 10 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.295 $Y=1.395
+ $X2=2.37 $Y2=1.395
r215 10 51 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.295 $Y=1.395
+ $X2=2.07 $Y2=1.395
r216 9 63 5.03009 $w=3.3e-07 $l=1.48e-07 $layer=POLY_cond $X=1.505 $Y=1.16
+ $X2=1.357 $Y2=1.16
r217 9 50 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=1.505 $Y=1.16
+ $X2=1.92 $Y2=1.16
r218 4 63 37.0704 $w=1.5e-07 $l=1.98167e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.357 $Y2=1.16
r219 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.43 $Y2=1.985
r220 1 63 37.0704 $w=1.5e-07 $l=1.98167e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.357 $Y2=1.16
r221 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%A_301_47# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 25 27 29 30 32 34 35 37 39 40 42 44 45 46 47 48 49 50 53 56 61 65 69 70 71
c146 71 0 1.31317e-19 $X=1.792 $Y=1.15
c147 70 0 1.90789e-20 $X=1.65 $Y=1.495
c148 69 0 1.40893e-19 $X=1.64 $Y=1.63
c149 56 0 1.1321e-20 $X=1.792 $Y=1.025
c150 42 0 7.94785e-20 $X=5.55 $Y=0.96
r151 69 70 5.91105 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.65 $Y=1.63
+ $X2=1.65 $Y2=1.495
r152 65 67 6.96131 $w=5.08e-07 $l=2.65e-07 $layer=LI1_cond $X=1.73 $Y=0.56
+ $X2=1.73 $Y2=0.825
r153 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.76
+ $Y=1.16 $X2=5.76 $Y2=1.16
r154 59 71 2.06747 $w=2.5e-07 $l=1.93e-07 $layer=LI1_cond $X=1.985 $Y=1.15
+ $X2=1.792 $Y2=1.15
r155 59 61 174.019 $w=2.48e-07 $l=3.775e-06 $layer=LI1_cond $X=1.985 $Y=1.15
+ $X2=5.76 $Y2=1.15
r156 57 71 4.36486 $w=3.05e-07 $l=1.60078e-07 $layer=LI1_cond $X=1.712 $Y=1.275
+ $X2=1.792 $Y2=1.15
r157 57 70 11.2683 $w=2.23e-07 $l=2.2e-07 $layer=LI1_cond $X=1.712 $Y=1.275
+ $X2=1.712 $Y2=1.495
r158 56 71 4.36486 $w=3.05e-07 $l=1.25e-07 $layer=LI1_cond $X=1.792 $Y=1.025
+ $X2=1.792 $Y2=1.15
r159 56 67 5.98672 $w=3.83e-07 $l=2e-07 $layer=LI1_cond $X=1.792 $Y=1.025
+ $X2=1.792 $Y2=0.825
r160 51 69 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=1.65 $Y=1.67 $X2=1.65
+ $Y2=1.63
r161 51 53 21.0732 $w=3.48e-07 $l=6.4e-07 $layer=LI1_cond $X=1.65 $Y=1.67
+ $X2=1.65 $Y2=2.31
r162 42 62 35.5158 $w=2.85e-07 $l=2.81372e-07 $layer=POLY_cond $X=5.55 $Y=0.96
+ $X2=5.76 $Y2=1.127
r163 42 44 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.55 $Y=0.96 $X2=5.55
+ $Y2=0.56
r164 41 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.205 $Y=1.035
+ $X2=5.13 $Y2=1.035
r165 40 42 23.4449 $w=2.85e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.475 $Y=1.035
+ $X2=5.55 $Y2=0.96
r166 40 41 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.475 $Y=1.035
+ $X2=5.205 $Y2=1.035
r167 37 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.13 $Y=0.96
+ $X2=5.13 $Y2=1.035
r168 37 39 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.13 $Y=0.96 $X2=5.13
+ $Y2=0.56
r169 36 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.785 $Y=1.035
+ $X2=4.71 $Y2=1.035
r170 35 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.055 $Y=1.035
+ $X2=5.13 $Y2=1.035
r171 35 36 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.055 $Y=1.035
+ $X2=4.785 $Y2=1.035
r172 32 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.71 $Y=0.96
+ $X2=4.71 $Y2=1.035
r173 32 34 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.71 $Y=0.96 $X2=4.71
+ $Y2=0.56
r174 31 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.365 $Y=1.035
+ $X2=4.29 $Y2=1.035
r175 30 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.635 $Y=1.035
+ $X2=4.71 $Y2=1.035
r176 30 31 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.635 $Y=1.035
+ $X2=4.365 $Y2=1.035
r177 27 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=0.96
+ $X2=4.29 $Y2=1.035
r178 27 29 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.29 $Y=0.96 $X2=4.29
+ $Y2=0.56
r179 26 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.945 $Y=1.035
+ $X2=3.87 $Y2=1.035
r180 25 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.215 $Y=1.035
+ $X2=4.29 $Y2=1.035
r181 25 26 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.215 $Y=1.035
+ $X2=3.945 $Y2=1.035
r182 22 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.87 $Y=0.96
+ $X2=3.87 $Y2=1.035
r183 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.87 $Y=0.96 $X2=3.87
+ $Y2=0.56
r184 21 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.525 $Y=1.035
+ $X2=3.45 $Y2=1.035
r185 20 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.795 $Y=1.035
+ $X2=3.87 $Y2=1.035
r186 20 21 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.795 $Y=1.035
+ $X2=3.525 $Y2=1.035
r187 17 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.45 $Y=0.96
+ $X2=3.45 $Y2=1.035
r188 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.45 $Y=0.96 $X2=3.45
+ $Y2=0.56
r189 16 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=1.035
+ $X2=3.03 $Y2=1.035
r190 15 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.375 $Y=1.035
+ $X2=3.45 $Y2=1.035
r191 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.375 $Y=1.035
+ $X2=3.105 $Y2=1.035
r192 12 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.03 $Y=0.96
+ $X2=3.03 $Y2=1.035
r193 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.03 $Y=0.96 $X2=3.03
+ $Y2=0.56
r194 10 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=1.035
+ $X2=3.03 $Y2=1.035
r195 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.955 $Y=1.035
+ $X2=2.685 $Y2=1.035
r196 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.61 $Y=0.96
+ $X2=2.685 $Y2=1.035
r197 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.61 $Y=0.96 $X2=2.61
+ $Y2=0.56
r198 2 69 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.485 $X2=1.64 $Y2=1.63
r199 2 53 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.485 $X2=1.64 $Y2=2.31
r200 1 65 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.64 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%A_116_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 79 83 84 87 90 105 107
c151 90 0 7.94785e-20 $X=6.665 $Y=1.19
c152 87 0 6.83439e-20 $X=0.69 $Y=1.19
c153 84 0 2.38356e-19 $X=0.835 $Y=1.19
r154 106 107 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.75 $Y=1.16
+ $X2=9.17 $Y2=1.16
r155 104 106 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=8.74 $Y=1.16
+ $X2=8.75 $Y2=1.16
r156 104 105 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=8.74
+ $Y=1.16 $X2=8.74 $Y2=1.16
r157 102 104 91.0912 $w=2.7e-07 $l=4.1e-07 $layer=POLY_cond $X=8.33 $Y=1.16
+ $X2=8.74 $Y2=1.16
r158 101 102 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.91 $Y=1.16
+ $X2=8.33 $Y2=1.16
r159 100 101 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.49 $Y=1.16
+ $X2=7.91 $Y2=1.16
r160 99 100 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.07 $Y=1.16
+ $X2=7.49 $Y2=1.16
r161 98 99 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.65 $Y=1.16
+ $X2=7.07 $Y2=1.16
r162 96 98 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=6.36 $Y=1.16
+ $X2=6.65 $Y2=1.16
r163 96 97 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=6.36
+ $Y=1.16 $X2=6.36 $Y2=1.16
r164 93 96 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=6.23 $Y=1.16
+ $X2=6.36 $Y2=1.16
r165 91 105 95.6528 $w=2.48e-07 $l=2.075e-06 $layer=LI1_cond $X=6.665 $Y=1.15
+ $X2=8.74 $Y2=1.15
r166 91 97 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=6.665 $Y=1.15
+ $X2=6.36 $Y2=1.15
r167 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.665 $Y=1.19
+ $X2=6.665 $Y2=1.19
r168 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.19
+ $X2=0.69 $Y2=1.19
r169 84 86 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.19
+ $X2=0.69 $Y2=1.19
r170 83 90 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.52 $Y=1.19
+ $X2=6.665 $Y2=1.19
r171 83 84 7.03588 $w=1.4e-07 $l=5.685e-06 $layer=MET1_cond $X=6.52 $Y=1.19
+ $X2=0.835 $Y2=1.19
r172 81 87 18.0227 $w=1.98e-07 $l=3.25e-07 $layer=LI1_cond $X=0.7 $Y=1.515
+ $X2=0.7 $Y2=1.19
r173 81 82 5.62585 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=0.7 $Y=1.515 $X2=0.7
+ $Y2=1.615
r174 79 87 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.7 $Y=1.095
+ $X2=0.7 $Y2=1.19
r175 79 80 5.62585 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=0.7 $Y=1.095 $X2=0.7
+ $Y2=0.995
r176 77 82 36.2703 $w=1.83e-07 $l=6.05e-07 $layer=LI1_cond $X=0.707 $Y=2.22
+ $X2=0.707 $Y2=1.615
r177 73 80 32.973 $w=1.83e-07 $l=5.5e-07 $layer=LI1_cond $X=0.707 $Y=0.445
+ $X2=0.707 $Y2=0.995
r178 67 107 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.17 $Y=1.295
+ $X2=9.17 $Y2=1.16
r179 67 69 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.17 $Y=1.295
+ $X2=9.17 $Y2=1.985
r180 63 107 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.17 $Y=1.025
+ $X2=9.17 $Y2=1.16
r181 63 65 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.17 $Y=1.025
+ $X2=9.17 $Y2=0.56
r182 59 106 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.75 $Y=1.295
+ $X2=8.75 $Y2=1.16
r183 59 61 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.75 $Y=1.295
+ $X2=8.75 $Y2=1.985
r184 55 106 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.75 $Y=1.025
+ $X2=8.75 $Y2=1.16
r185 55 57 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.75 $Y=1.025
+ $X2=8.75 $Y2=0.56
r186 51 102 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.33 $Y=1.295
+ $X2=8.33 $Y2=1.16
r187 51 53 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.33 $Y=1.295
+ $X2=8.33 $Y2=1.985
r188 47 102 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.33 $Y=1.025
+ $X2=8.33 $Y2=1.16
r189 47 49 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.33 $Y=1.025
+ $X2=8.33 $Y2=0.56
r190 43 101 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.91 $Y=1.295
+ $X2=7.91 $Y2=1.16
r191 43 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.91 $Y=1.295
+ $X2=7.91 $Y2=1.985
r192 39 101 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.91 $Y=1.025
+ $X2=7.91 $Y2=1.16
r193 39 41 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.91 $Y=1.025
+ $X2=7.91 $Y2=0.56
r194 35 100 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.49 $Y=1.295
+ $X2=7.49 $Y2=1.16
r195 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.49 $Y=1.295
+ $X2=7.49 $Y2=1.985
r196 31 100 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.49 $Y=1.025
+ $X2=7.49 $Y2=1.16
r197 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.49 $Y=1.025
+ $X2=7.49 $Y2=0.56
r198 27 99 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.07 $Y=1.295
+ $X2=7.07 $Y2=1.16
r199 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.07 $Y=1.295
+ $X2=7.07 $Y2=1.985
r200 23 99 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.07 $Y=1.025
+ $X2=7.07 $Y2=1.16
r201 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.07 $Y=1.025
+ $X2=7.07 $Y2=0.56
r202 19 98 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.65 $Y=1.295
+ $X2=6.65 $Y2=1.16
r203 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.65 $Y=1.295
+ $X2=6.65 $Y2=1.985
r204 15 98 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.65 $Y=1.025
+ $X2=6.65 $Y2=1.16
r205 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.65 $Y=1.025
+ $X2=6.65 $Y2=0.56
r206 11 93 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.23 $Y=1.295
+ $X2=6.23 $Y2=1.16
r207 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.23 $Y=1.295
+ $X2=6.23 $Y2=1.985
r208 7 93 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.23 $Y=1.025
+ $X2=6.23 $Y2=1.16
r209 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.23 $Y=1.025
+ $X2=6.23 $Y2=0.56
r210 2 77 600 $w=1.7e-07 $l=7.99656e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.485 $X2=0.715 $Y2=2.22
r211 1 73 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.235 $X2=0.715 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%VPWR 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 49 51 56 61 77 78 84 87 90
r137 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r138 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r139 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 77 78 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r141 75 78 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=9.43 $Y2=2.72
r142 74 77 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=9.43 $Y2=2.72
r143 74 75 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r144 72 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r145 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r146 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r147 69 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r148 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r149 66 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.42 $Y2=2.72
r150 66 68 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.91 $Y2=2.72
r151 65 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r152 65 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r153 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r154 62 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.58 $Y2=2.72
r155 62 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.99 $Y2=2.72
r156 61 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=3.42 $Y2=2.72
r157 61 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=2.72
+ $X2=2.99 $Y2=2.72
r158 60 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r159 60 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r160 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r161 57 84 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.137 $Y2=2.72
r162 57 59 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=2.07 $Y2=2.72
r163 56 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.58 $Y2=2.72
r164 56 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.07 $Y2=2.72
r165 55 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r166 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r167 52 81 5.0973 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.222 $Y2=2.72
r168 52 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.69 $Y2=2.72
r169 51 84 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.97 $Y=2.72
+ $X2=1.137 $Y2=2.72
r170 51 54 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.97 $Y=2.72
+ $X2=0.69 $Y2=2.72
r171 49 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r172 49 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r173 47 71 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=4.83 $Y2=2.72
r174 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=5.1 $Y2=2.72
r175 46 74 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.29 $Y2=2.72
r176 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.1 $Y2=2.72
r177 44 68 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=3.91 $Y2=2.72
r178 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=4.26 $Y2=2.72
r179 43 71 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.83 $Y2=2.72
r180 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.26 $Y2=2.72
r181 39 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=2.635 $X2=5.1
+ $Y2=2.72
r182 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.1 $Y=2.635
+ $X2=5.1 $Y2=2.36
r183 35 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=2.635
+ $X2=4.26 $Y2=2.72
r184 35 37 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.26 $Y=2.635
+ $X2=4.26 $Y2=2.36
r185 31 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.635
+ $X2=3.42 $Y2=2.72
r186 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.42 $Y=2.635
+ $X2=3.42 $Y2=2.36
r187 27 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.635
+ $X2=2.58 $Y2=2.72
r188 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.58 $Y=2.635
+ $X2=2.58 $Y2=2.36
r189 23 84 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.137 $Y=2.635
+ $X2=1.137 $Y2=2.72
r190 23 25 21.1568 $w=3.33e-07 $l=6.15e-07 $layer=LI1_cond $X=1.137 $Y=2.635
+ $X2=1.137 $Y2=2.02
r191 19 81 2.92581 $w=3.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.222 $Y2=2.72
r192 19 21 19.6876 $w=3.58e-07 $l=6.15e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.02
r193 6 41 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.545 $X2=5.1 $Y2=2.36
r194 5 37 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=1.545 $X2=4.26 $Y2=2.36
r195 4 33 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.545 $X2=3.42 $Y2=2.36
r196 3 29 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.545 $X2=2.58 $Y2=2.36
r197 2 25 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.485 $X2=1.135 $Y2=2.02
r198 1 21 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%A_407_309# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 52 60 62 63 64 67
r91 66 67 17.2004 $w=5.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.945 $Y=2.18
+ $X2=5.435 $Y2=2.18
r92 58 60 17.6264 $w=5.68e-07 $l=8.4e-07 $layer=LI1_cond $X=8.54 $Y=2.18
+ $X2=9.38 $Y2=2.18
r93 56 58 17.6264 $w=5.68e-07 $l=8.4e-07 $layer=LI1_cond $X=7.7 $Y=2.18 $X2=8.54
+ $Y2=2.18
r94 54 56 17.6264 $w=5.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.86 $Y=2.18 $X2=7.7
+ $Y2=2.18
r95 52 66 1.25903 $w=5.68e-07 $l=6e-08 $layer=LI1_cond $X=6.005 $Y=2.18
+ $X2=5.945 $Y2=2.18
r96 52 54 17.9412 $w=5.68e-07 $l=8.55e-07 $layer=LI1_cond $X=6.005 $Y=2.18
+ $X2=6.86 $Y2=2.18
r97 51 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=1.98
+ $X2=4.68 $Y2=1.98
r98 51 67 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.765 $Y=1.98
+ $X2=5.435 $Y2=1.98
r99 46 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.68 $Y=2.065
+ $X2=4.68 $Y2=1.98
r100 46 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.68 $Y=2.065
+ $X2=4.68 $Y2=2.3
r101 45 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=1.98
+ $X2=3.84 $Y2=1.98
r102 44 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=1.98
+ $X2=4.68 $Y2=1.98
r103 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.595 $Y=1.98
+ $X2=3.925 $Y2=1.98
r104 40 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=2.065
+ $X2=3.84 $Y2=1.98
r105 40 42 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.84 $Y=2.065
+ $X2=3.84 $Y2=2.3
r106 39 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=1.98 $X2=3
+ $Y2=1.98
r107 38 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=1.98
+ $X2=3.84 $Y2=1.98
r108 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.755 $Y=1.98
+ $X2=3.085 $Y2=1.98
r109 34 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=2.065 $X2=3
+ $Y2=1.98
r110 34 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3 $Y=2.065 $X2=3
+ $Y2=2.3
r111 32 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=1.98 $X2=3
+ $Y2=1.98
r112 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.915 $Y=1.98
+ $X2=2.245 $Y2=1.98
r113 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.12 $Y=2.065
+ $X2=2.245 $Y2=1.98
r114 28 30 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=2.12 $Y=2.065
+ $X2=2.12 $Y2=2.3
r115 9 60 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=9.245
+ $Y=1.485 $X2=9.38 $Y2=2.02
r116 8 58 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=8.405
+ $Y=1.485 $X2=8.54 $Y2=2.02
r117 7 56 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=7.565
+ $Y=1.485 $X2=7.7 $Y2=2.02
r118 6 54 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.725
+ $Y=1.485 $X2=6.86 $Y2=2.02
r119 5 66 300 $w=1.7e-07 $l=9.96406e-07 $layer=licon1_PDIFF $count=2 $X=5.385
+ $Y=1.545 $X2=5.945 $Y2=2.3
r120 4 48 600 $w=1.7e-07 $l=8.19726e-07 $layer=licon1_PDIFF $count=1 $X=4.545
+ $Y=1.545 $X2=4.68 $Y2=2.3
r121 3 42 600 $w=1.7e-07 $l=8.19726e-07 $layer=licon1_PDIFF $count=1 $X=3.705
+ $Y=1.545 $X2=3.84 $Y2=2.3
r122 2 36 600 $w=1.7e-07 $l=8.19726e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=1.545 $X2=3 $Y2=2.3
r123 1 30 600 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=1.545 $X2=2.16 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%Z 1 2 3 4 5 6 7 8 25 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 71 109
r108 51 71 3.22874 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=9.45 $Y=1.585
+ $X2=9.325 $Y2=1.585
r109 50 51 8.86994 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=9.45 $Y=1.19
+ $X2=9.45 $Y2=1.445
r110 49 109 3.3405 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=9.45 $Y=0.735
+ $X2=9.45 $Y2=0.855
r111 49 50 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.45 $Y=0.895
+ $X2=9.45 $Y2=1.19
r112 49 109 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=9.45 $Y=0.895
+ $X2=9.45 $Y2=0.855
r113 48 71 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=8.965 $Y=1.585
+ $X2=9.325 $Y2=1.585
r114 48 106 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=8.965 $Y=1.585
+ $X2=8.96 $Y2=1.585
r115 47 106 18.7272 $w=2.78e-07 $l=4.55e-07 $layer=LI1_cond $X=8.505 $Y=1.585
+ $X2=8.96 $Y2=1.585
r116 47 102 15.8461 $w=2.78e-07 $l=3.85e-07 $layer=LI1_cond $X=8.505 $Y=1.585
+ $X2=8.12 $Y2=1.585
r117 46 102 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=8.045 $Y=1.585
+ $X2=8.12 $Y2=1.585
r118 45 46 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=7.585 $Y=1.585
+ $X2=8.045 $Y2=1.585
r119 45 96 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=7.585 $Y=1.585
+ $X2=7.28 $Y2=1.585
r120 44 96 6.3796 $w=2.78e-07 $l=1.55e-07 $layer=LI1_cond $X=7.125 $Y=1.585
+ $X2=7.28 $Y2=1.585
r121 44 92 28.1937 $w=2.78e-07 $l=6.85e-07 $layer=LI1_cond $X=7.125 $Y=1.585
+ $X2=6.44 $Y2=1.585
r122 43 92 9.67229 $w=2.78e-07 $l=2.35e-07 $layer=LI1_cond $X=6.205 $Y=1.585
+ $X2=6.44 $Y2=1.585
r123 42 43 18.7272 $w=2.78e-07 $l=4.55e-07 $layer=LI1_cond $X=5.75 $Y=1.585
+ $X2=6.205 $Y2=1.585
r124 41 42 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=5.29 $Y=1.585
+ $X2=5.75 $Y2=1.585
r125 40 41 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=4.83 $Y=1.585
+ $X2=5.29 $Y2=1.585
r126 39 40 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=4.37 $Y=1.585
+ $X2=4.83 $Y2=1.585
r127 38 39 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=1.585
+ $X2=4.37 $Y2=1.585
r128 37 38 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=3.45 $Y=1.585
+ $X2=3.91 $Y2=1.585
r129 36 37 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=1.585
+ $X2=3.45 $Y2=1.585
r130 35 36 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=1.585
+ $X2=2.99 $Y2=1.585
r131 32 34 40.3355 $w=2.38e-07 $l=8.4e-07 $layer=LI1_cond $X=8.12 $Y=0.735
+ $X2=8.96 $Y2=0.735
r132 30 32 40.3355 $w=2.38e-07 $l=8.4e-07 $layer=LI1_cond $X=7.28 $Y=0.735
+ $X2=8.12 $Y2=0.735
r133 27 30 40.3355 $w=2.38e-07 $l=8.4e-07 $layer=LI1_cond $X=6.44 $Y=0.735
+ $X2=7.28 $Y2=0.735
r134 25 49 3.47969 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=9.325 $Y=0.735
+ $X2=9.45 $Y2=0.735
r135 25 34 17.5267 $w=2.38e-07 $l=3.65e-07 $layer=LI1_cond $X=9.325 $Y=0.735
+ $X2=8.96 $Y2=0.735
r136 8 106 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=8.825
+ $Y=1.485 $X2=8.96 $Y2=1.64
r137 7 102 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=7.985
+ $Y=1.485 $X2=8.12 $Y2=1.64
r138 6 96 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=7.145
+ $Y=1.485 $X2=7.28 $Y2=1.64
r139 5 92 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.485 $X2=6.44 $Y2=1.64
r140 4 34 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=8.825
+ $Y=0.235 $X2=8.96 $Y2=0.76
r141 3 32 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=7.985
+ $Y=0.235 $X2=8.12 $Y2=0.76
r142 2 30 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.235 $X2=7.28 $Y2=0.76
r143 1 27 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=6.305
+ $Y=0.235 $X2=6.44 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%VGND 1 2 3 4 5 6 19 21 25 29 33 35 39 43 46
+ 47 48 49 50 52 67 77 78 84 87 90
r134 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r135 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r136 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r137 77 78 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r138 75 78 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r139 75 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r140 74 77 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r141 74 75 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r142 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=0 $X2=5.34
+ $Y2=0
r143 72 74 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.505 $Y=0 $X2=5.75
+ $Y2=0
r144 71 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r145 71 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r146 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r147 68 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.5
+ $Y2=0
r148 68 70 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=0
+ $X2=4.83 $Y2=0
r149 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.34
+ $Y2=0
r150 67 70 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=4.83
+ $Y2=0
r151 66 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r152 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r153 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r154 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r155 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r156 60 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r157 59 62 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r158 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r159 57 84 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=1.137 $Y2=0
r160 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=1.61 $Y2=0
r161 56 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r162 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r163 53 81 5.0973 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r164 53 55 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.69
+ $Y2=0
r165 52 84 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.137
+ $Y2=0
r166 52 55 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.69
+ $Y2=0
r167 50 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r168 50 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r169 48 65 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.45
+ $Y2=0
r170 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.66
+ $Y2=0
r171 46 62 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=0
+ $X2=2.53 $Y2=0
r172 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.82
+ $Y2=0
r173 45 65 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=3.45 $Y2=0
r174 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.82
+ $Y2=0
r175 41 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0
r176 41 43 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.34 $Y=0.085
+ $X2=5.34 $Y2=0.36
r177 37 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=0.085 $X2=4.5
+ $Y2=0
r178 37 39 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.5 $Y=0.085
+ $X2=4.5 $Y2=0.36
r179 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.66
+ $Y2=0
r180 35 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.5
+ $Y2=0
r181 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=3.825 $Y2=0
r182 31 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=0.085
+ $X2=3.66 $Y2=0
r183 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.66 $Y=0.085
+ $X2=3.66 $Y2=0.36
r184 27 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0
r185 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0.36
r186 23 84 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0
r187 23 25 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0.36
r188 19 81 2.92581 $w=3.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.222 $Y2=0
r189 19 21 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.36
r190 6 43 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.205
+ $Y=0.235 $X2=5.34 $Y2=0.36
r191 5 39 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.365
+ $Y=0.235 $X2=4.5 $Y2=0.36
r192 4 33 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.525
+ $Y=0.235 $X2=3.66 $Y2=0.36
r193 3 29 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.685
+ $Y=0.235 $X2=2.82 $Y2=0.36
r194 2 25 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.135 $Y2=0.36
r195 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_8%A_455_47# 1 2 3 4 5 6 7 8 9 28 31 32 33 36
+ 38 41 43 46 56 58 59 60 61
r104 64 65 5.22619 $w=4.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.89 $Y=0.56
+ $X2=5.89 $Y2=0.755
r105 61 64 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.89 $Y=0.35
+ $X2=5.89 $Y2=0.56
r106 54 56 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=8.54 $Y=0.35
+ $X2=9.38 $Y2=0.35
r107 52 54 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=7.7 $Y=0.35
+ $X2=8.54 $Y2=0.35
r108 50 52 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=6.86 $Y=0.35
+ $X2=7.7 $Y2=0.35
r109 48 61 5.54258 $w=1.9e-07 $l=2.15e-07 $layer=LI1_cond $X=6.105 $Y=0.35
+ $X2=5.89 $Y2=0.35
r110 48 50 44.0718 $w=1.88e-07 $l=7.55e-07 $layer=LI1_cond $X=6.105 $Y=0.35
+ $X2=6.86 $Y2=0.35
r111 47 60 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=0.755
+ $X2=4.92 $Y2=0.755
r112 46 65 5.23352 $w=2e-07 $l=2.15e-07 $layer=LI1_cond $X=5.675 $Y=0.755
+ $X2=5.89 $Y2=0.755
r113 46 47 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=5.675 $Y=0.755
+ $X2=5.005 $Y2=0.755
r114 43 60 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.92 $Y=0.655 $X2=4.92
+ $Y2=0.755
r115 43 45 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.92 $Y=0.655
+ $X2=4.92 $Y2=0.56
r116 42 59 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.755
+ $X2=4.08 $Y2=0.755
r117 41 60 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=0.755
+ $X2=4.92 $Y2=0.755
r118 41 42 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=4.835 $Y=0.755
+ $X2=4.165 $Y2=0.755
r119 38 59 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.08 $Y=0.655 $X2=4.08
+ $Y2=0.755
r120 38 40 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.08 $Y=0.655
+ $X2=4.08 $Y2=0.56
r121 37 58 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=0.755
+ $X2=3.24 $Y2=0.755
r122 36 59 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0.755
+ $X2=4.08 $Y2=0.755
r123 36 37 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=3.995 $Y=0.755
+ $X2=3.325 $Y2=0.755
r124 33 58 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.24 $Y=0.655 $X2=3.24
+ $Y2=0.755
r125 33 35 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.24 $Y=0.655
+ $X2=3.24 $Y2=0.56
r126 31 58 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=0.755
+ $X2=3.24 $Y2=0.755
r127 31 32 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=3.155 $Y=0.755
+ $X2=2.485 $Y2=0.755
r128 28 32 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.32 $Y=0.655
+ $X2=2.485 $Y2=0.755
r129 28 30 3.51212 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.32 $Y=0.655
+ $X2=2.32 $Y2=0.56
r130 9 56 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=9.245
+ $Y=0.235 $X2=9.38 $Y2=0.36
r131 8 54 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=8.405
+ $Y=0.235 $X2=8.54 $Y2=0.36
r132 7 52 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.565
+ $Y=0.235 $X2=7.7 $Y2=0.36
r133 6 50 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.725
+ $Y=0.235 $X2=6.86 $Y2=0.36
r134 5 64 182 $w=1.7e-07 $l=4.39744e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.895 $Y2=0.56
r135 4 45 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.785
+ $Y=0.235 $X2=4.92 $Y2=0.56
r136 3 40 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.945
+ $Y=0.235 $X2=4.08 $Y2=0.56
r137 2 35 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.24 $Y2=0.56
r138 1 30 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.4 $Y2=0.56
.ends


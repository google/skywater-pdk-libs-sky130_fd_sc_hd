/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_TB_V
`define SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_TB_V

/**
 * lpflow_lsbuf_lh_hl_isowell_tap: Level-shift buffer, low-to-high,
 *                                 isolated well on input buffer,
 *                                 vpb/vnb taps, double-row-height
 *                                 cell.
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap.v"

module top();

    // Inputs are registered
    reg A;
    reg VPWRIN;
    reg VPWR;
    reg VGND;
    reg VPB;

    // Outputs are wires
    wire X;

    initial
    begin
        // Initial state is x for all inputs.
        A      = 1'bX;
        VGND   = 1'bX;
        VPB    = 1'bX;
        VPWR   = 1'bX;
        VPWRIN = 1'bX;

        #20   A      = 1'b0;
        #40   VGND   = 1'b0;
        #60   VPB    = 1'b0;
        #80   VPWR   = 1'b0;
        #100  VPWRIN = 1'b0;
        #120  A      = 1'b1;
        #140  VGND   = 1'b1;
        #160  VPB    = 1'b1;
        #180  VPWR   = 1'b1;
        #200  VPWRIN = 1'b1;
        #220  A      = 1'b0;
        #240  VGND   = 1'b0;
        #260  VPB    = 1'b0;
        #280  VPWR   = 1'b0;
        #300  VPWRIN = 1'b0;
        #320  VPWRIN = 1'b1;
        #340  VPWR   = 1'b1;
        #360  VPB    = 1'b1;
        #380  VGND   = 1'b1;
        #400  A      = 1'b1;
        #420  VPWRIN = 1'bx;
        #440  VPWR   = 1'bx;
        #460  VPB    = 1'bx;
        #480  VGND   = 1'bx;
        #500  A      = 1'bx;
    end

    sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap dut (.A(A), .VPWRIN(VPWRIN), .VPWR(VPWR), .VGND(VGND), .VPB(VPB), .X(X));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_TB_V

* File: sky130_fd_sc_hd__nor4_4.spice.SKY130_FD_SC_HD__NOR4_4.pxi
* Created: Thu Aug 27 14:32:55 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4_4%A N_A_c_121_n N_A_M1006_g N_A_M1003_g N_A_c_122_n
+ N_A_M1010_g N_A_M1021_g N_A_c_123_n N_A_M1018_g N_A_M1024_g N_A_c_124_n
+ N_A_M1019_g N_A_M1029_g A N_A_c_125_n N_A_c_126_n PM_SKY130_FD_SC_HD__NOR4_4%A
x_PM_SKY130_FD_SC_HD__NOR4_4%B N_B_c_195_n N_B_M1012_g N_B_M1002_g N_B_c_196_n
+ N_B_M1020_g N_B_M1014_g N_B_c_197_n N_B_M1023_g N_B_M1015_g N_B_c_198_n
+ N_B_M1027_g N_B_M1025_g B B B N_B_c_200_n PM_SKY130_FD_SC_HD__NOR4_4%B
x_PM_SKY130_FD_SC_HD__NOR4_4%C N_C_c_273_n N_C_M1004_g N_C_M1001_g N_C_c_274_n
+ N_C_M1007_g N_C_M1016_g N_C_c_275_n N_C_M1008_g N_C_M1026_g N_C_c_276_n
+ N_C_M1011_g N_C_M1030_g C N_C_c_277_n N_C_c_278_n PM_SKY130_FD_SC_HD__NOR4_4%C
x_PM_SKY130_FD_SC_HD__NOR4_4%D N_D_c_350_n N_D_M1000_g N_D_M1017_g N_D_c_351_n
+ N_D_M1005_g N_D_M1022_g N_D_c_352_n N_D_M1009_g N_D_M1028_g N_D_c_353_n
+ N_D_M1013_g N_D_M1031_g D N_D_c_354_n N_D_c_355_n PM_SKY130_FD_SC_HD__NOR4_4%D
x_PM_SKY130_FD_SC_HD__NOR4_4%A_27_297# N_A_27_297#_M1003_s N_A_27_297#_M1021_s
+ N_A_27_297#_M1029_s N_A_27_297#_M1014_d N_A_27_297#_M1025_d
+ N_A_27_297#_c_428_n N_A_27_297#_c_429_n N_A_27_297#_c_430_n
+ N_A_27_297#_c_457_p N_A_27_297#_c_431_n N_A_27_297#_c_432_n
+ N_A_27_297#_c_458_p N_A_27_297#_c_448_n N_A_27_297#_c_477_p
+ N_A_27_297#_c_433_n N_A_27_297#_c_434_n N_A_27_297#_c_435_n
+ N_A_27_297#_c_461_p PM_SKY130_FD_SC_HD__NOR4_4%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR4_4%VPWR N_VPWR_M1003_d N_VPWR_M1024_d N_VPWR_c_491_n
+ N_VPWR_c_492_n VPWR N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_490_n N_VPWR_c_497_n N_VPWR_c_498_n PM_SKY130_FD_SC_HD__NOR4_4%VPWR
x_PM_SKY130_FD_SC_HD__NOR4_4%A_449_297# N_A_449_297#_M1002_s
+ N_A_449_297#_M1015_s N_A_449_297#_M1001_d N_A_449_297#_M1026_d
+ N_A_449_297#_c_583_n N_A_449_297#_c_584_n N_A_449_297#_c_585_n
+ N_A_449_297#_c_586_n N_A_449_297#_c_587_n N_A_449_297#_c_588_n
+ N_A_449_297#_c_589_n PM_SKY130_FD_SC_HD__NOR4_4%A_449_297#
x_PM_SKY130_FD_SC_HD__NOR4_4%A_807_297# N_A_807_297#_M1001_s
+ N_A_807_297#_M1016_s N_A_807_297#_M1030_s N_A_807_297#_M1022_d
+ N_A_807_297#_M1031_d N_A_807_297#_c_641_n N_A_807_297#_c_644_n
+ N_A_807_297#_c_642_n N_A_807_297#_c_683_n N_A_807_297#_c_646_n
+ N_A_807_297#_c_648_n N_A_807_297#_c_649_n N_A_807_297#_c_691_p
+ N_A_807_297#_c_643_n N_A_807_297#_c_695_p N_A_807_297#_c_670_n
+ N_A_807_297#_c_672_n N_A_807_297#_c_674_n
+ PM_SKY130_FD_SC_HD__NOR4_4%A_807_297#
x_PM_SKY130_FD_SC_HD__NOR4_4%Y N_Y_M1006_d N_Y_M1018_d N_Y_M1012_s N_Y_M1023_s
+ N_Y_M1004_s N_Y_M1008_s N_Y_M1000_d N_Y_M1009_d N_Y_M1017_s N_Y_M1028_s
+ N_Y_c_721_n N_Y_c_698_n N_Y_c_699_n N_Y_c_732_n N_Y_c_700_n N_Y_c_737_n
+ N_Y_c_701_n N_Y_c_752_n N_Y_c_702_n N_Y_c_767_n N_Y_c_703_n N_Y_c_774_n
+ N_Y_c_704_n N_Y_c_779_n N_Y_c_716_n N_Y_c_705_n N_Y_c_802_n N_Y_c_717_n
+ N_Y_c_706_n N_Y_c_707_n N_Y_c_708_n N_Y_c_709_n N_Y_c_710_n N_Y_c_711_n
+ N_Y_c_712_n N_Y_c_718_n N_Y_c_713_n N_Y_c_719_n Y N_Y_c_715_n
+ PM_SKY130_FD_SC_HD__NOR4_4%Y
x_PM_SKY130_FD_SC_HD__NOR4_4%VGND N_VGND_M1006_s N_VGND_M1010_s N_VGND_M1019_s
+ N_VGND_M1020_d N_VGND_M1027_d N_VGND_M1007_d N_VGND_M1011_d N_VGND_M1005_s
+ N_VGND_M1013_s N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n
+ N_VGND_c_913_n N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n
+ N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_920_n N_VGND_c_921_n N_VGND_c_922_n
+ N_VGND_c_923_n N_VGND_c_924_n N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n
+ N_VGND_c_928_n N_VGND_c_929_n VGND N_VGND_c_930_n N_VGND_c_931_n
+ N_VGND_c_932_n N_VGND_c_933_n N_VGND_c_934_n PM_SKY130_FD_SC_HD__NOR4_4%VGND
cc_1 VNB N_A_c_121_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_122_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_A_c_123_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_A_c_124_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB N_A_c_125_n 0.0161158f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_6 VNB N_A_c_126_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_7 VNB N_B_c_195_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B_c_196_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_9 VNB N_B_c_197_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_10 VNB N_B_c_198_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_11 VNB B 0.0163812f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_12 VNB N_B_c_200_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.18
cc_13 VNB N_C_c_273_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_14 VNB N_C_c_274_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_15 VNB N_C_c_275_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_16 VNB N_C_c_276_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_17 VNB N_C_c_277_n 0.00349977f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_18 VNB N_C_c_278_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_19 VNB N_D_c_350_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_20 VNB N_D_c_351_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_21 VNB N_D_c_352_n 0.0157971f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_22 VNB N_D_c_353_n 0.0191578f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_23 VNB N_D_c_354_n 0.00389209f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_24 VNB N_D_c_355_n 0.0651519f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_25 VNB N_VPWR_c_490_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_698_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_27 VNB N_Y_c_699_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_28 VNB N_Y_c_700_n 0.00429924f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_29 VNB N_Y_c_701_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.18
cc_30 VNB N_Y_c_702_n 0.00892184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_703_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_704_n 0.00680092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_705_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_706_n 0.00105843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_707_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_708_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_709_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_710_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_711_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_712_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_713_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB Y 0.0207103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_715_n 0.00931661f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_909_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_910_n 0.0334957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_911_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_47 VNB N_VGND_c_912_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_48 VNB N_VGND_c_913_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_914_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_915_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_916_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_917_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_918_n 0.0118141f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_919_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_920_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_921_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_922_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_923_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_924_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_925_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_926_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_927_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_928_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_929_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_930_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_931_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_932_n 0.0197313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_933_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_934_n 0.370903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VPB N_A_M1003_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_71 VPB N_A_M1021_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_72 VPB N_A_M1024_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_73 VPB N_A_M1029_g 0.0185045f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_74 VPB N_A_c_126_n 0.0108808f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_75 VPB N_B_M1002_g 0.018818f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_76 VPB N_B_M1014_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_77 VPB N_B_M1015_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_78 VPB N_B_M1025_g 0.0252703f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_79 VPB N_B_c_200_n 0.0108798f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.18
cc_80 VPB N_C_M1001_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_81 VPB N_C_M1016_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_82 VPB N_C_M1026_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_83 VPB N_C_M1030_g 0.0188261f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_84 VPB N_C_c_278_n 0.0108798f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_85 VPB N_D_M1017_g 0.0188261f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_86 VPB N_D_M1022_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_87 VPB N_D_M1028_g 0.0182002f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_88 VPB N_D_M1031_g 0.0219116f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_89 VPB N_D_c_355_n 0.0102771f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_90 VPB N_A_27_297#_c_428_n 0.010823f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_91 VPB N_A_27_297#_c_429_n 0.0327764f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.325
cc_92 VPB N_A_27_297#_c_430_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_93 VPB N_A_27_297#_c_431_n 0.00240493f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_94 VPB N_A_27_297#_c_432_n 0.00414042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_297#_c_433_n 0.00198437f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_96 VPB N_A_27_297#_c_434_n 0.00516601f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.16
cc_97 VPB N_A_27_297#_c_435_n 0.00204609f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.18
cc_98 VPB N_VPWR_c_491_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_99 VPB N_VPWR_c_492_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_100 VPB N_VPWR_c_493_n 0.0174963f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_101 VPB N_VPWR_c_494_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.995
cc_102 VPB N_VPWR_c_495_n 0.143611f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_103 VPB N_VPWR_c_490_n 0.056284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_497_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_105 VPB N_VPWR_c_498_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_106 VPB N_A_449_297#_c_583_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.995
cc_107 VPB N_A_449_297#_c_584_n 0.0178099f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_108 VPB N_A_449_297#_c_585_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_109 VPB N_A_449_297#_c_586_n 0.00225182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_449_297#_c_587_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_449_297#_c_588_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_449_297#_c_589_n 0.00235657f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_113 VPB N_A_807_297#_c_641_n 0.00451061f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.325
cc_114 VPB N_A_807_297#_c_642_n 0.00166092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_807_297#_c_643_n 0.00692367f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.16
cc_116 VPB N_Y_c_716_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_Y_c_717_n 0.0123442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_Y_c_718_n 0.00235657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_Y_c_719_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB Y 0.00779291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 N_A_c_124_n N_B_c_195_n 0.0195974f $X=1.75 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_122 N_A_M1029_g N_B_M1002_g 0.0195974f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_c_125_n B 0.0121231f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_c_126_n B 2.62535e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_125_n N_B_c_200_n 2.62535e-19 $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_c_126_n N_B_c_200_n 0.0195974f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_c_125_n N_A_27_297#_c_428_n 0.0192812f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_M1003_g N_A_27_297#_c_430_n 0.0135215f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_M1021_g N_A_27_297#_c_430_n 0.0132714f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_c_125_n N_A_27_297#_c_430_n 0.041703f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_126_n N_A_27_297#_c_430_n 0.00211509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_M1024_g N_A_27_297#_c_431_n 0.0132273f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_M1029_g N_A_27_297#_c_431_n 0.0132131f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_c_125_n N_A_27_297#_c_431_n 0.0409754f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_126_n N_A_27_297#_c_431_n 0.00211509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_125_n N_A_27_297#_c_435_n 0.0204549f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_126_n N_A_27_297#_c_435_n 0.00220041f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_M1003_g N_VPWR_c_491_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_M1021_g N_VPWR_c_491_n 0.00157837f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1024_g N_VPWR_c_492_n 0.00157837f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1029_g N_VPWR_c_492_n 0.00302074f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1003_g N_VPWR_c_493_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1021_g N_VPWR_c_494_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1024_g N_VPWR_c_494_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1029_g N_VPWR_c_495_n 0.00585385f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1003_g N_VPWR_c_490_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1021_g N_VPWR_c_490_n 0.0104367f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1024_g N_VPWR_c_490_n 0.0104367f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1029_g N_VPWR_c_490_n 0.010464f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_c_121_n N_Y_c_721_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_122_n N_Y_c_721_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_123_n N_Y_c_721_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_122_n N_Y_c_698_n 0.00870364f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_123_n N_Y_c_698_n 0.00870364f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_125_n N_Y_c_698_n 0.0362443f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_126_n N_Y_c_698_n 0.00222133f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_c_121_n N_Y_c_699_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_122_n N_Y_c_699_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_c_125_n N_Y_c_699_n 0.0266272f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_c_126_n N_Y_c_699_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_c_122_n N_Y_c_732_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_123_n N_Y_c_732_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_124_n N_Y_c_732_n 0.00630972f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_124_n N_Y_c_700_n 0.00865686f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_125_n N_Y_c_700_n 0.00826974f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_c_124_n N_Y_c_737_n 5.22228e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_123_n N_Y_c_707_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_124_n N_Y_c_707_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_125_n N_Y_c_707_n 0.0266272f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_126_n N_Y_c_707_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_c_121_n N_VGND_c_910_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_125_n N_VGND_c_910_n 0.0157677f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_122_n N_VGND_c_911_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_c_123_n N_VGND_c_911_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_c_124_n N_VGND_c_912_n 0.00146448f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_121_n N_VGND_c_920_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_122_n N_VGND_c_920_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_123_n N_VGND_c_922_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_124_n N_VGND_c_922_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_121_n N_VGND_c_934_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_122_n N_VGND_c_934_n 0.0057163f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_c_123_n N_VGND_c_934_n 0.0057163f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_124_n N_VGND_c_934_n 0.0057435f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_184 B N_C_c_277_n 0.0150083f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_185 B N_C_c_278_n 0.00157386f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_186 N_B_M1002_g N_A_27_297#_c_432_n 2.57315e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B_M1002_g N_A_27_297#_c_448_n 0.0121747f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B_M1014_g N_A_27_297#_c_448_n 0.00984328f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B_M1015_g N_A_27_297#_c_433_n 0.00988743f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B_M1025_g N_A_27_297#_c_433_n 0.00988743f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_191 N_B_M1002_g N_VPWR_c_495_n 0.00357877f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B_M1014_g N_VPWR_c_495_n 0.00357877f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B_M1015_g N_VPWR_c_495_n 0.00357877f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B_M1025_g N_VPWR_c_495_n 0.00357877f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B_M1002_g N_VPWR_c_490_n 0.00525237f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B_M1014_g N_VPWR_c_490_n 0.00522516f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B_M1015_g N_VPWR_c_490_n 0.00522516f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B_M1025_g N_VPWR_c_490_n 0.00655123f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B_M1014_g N_A_449_297#_c_583_n 0.0109258f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B_M1015_g N_A_449_297#_c_583_n 0.01094f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_201 B N_A_449_297#_c_583_n 0.0416643f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_202 N_B_c_200_n N_A_449_297#_c_583_n 0.00211509f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B_M1025_g N_A_449_297#_c_584_n 0.0130871f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_204 B N_A_449_297#_c_584_n 0.0542632f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_205 N_B_M1002_g N_A_449_297#_c_586_n 2.57315e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_206 B N_A_449_297#_c_586_n 0.0204292f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_207 N_B_c_200_n N_A_449_297#_c_586_n 0.00219557f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_208 B N_A_449_297#_c_587_n 0.0204292f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_209 N_B_c_200_n N_A_449_297#_c_587_n 0.00219557f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B_c_195_n N_Y_c_732_n 5.22228e-19 $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B_c_195_n N_Y_c_700_n 0.00865686f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_212 B N_Y_c_700_n 0.00826974f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_213 N_B_c_195_n N_Y_c_737_n 0.00630972f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B_c_196_n N_Y_c_737_n 0.00630972f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B_c_197_n N_Y_c_737_n 5.22228e-19 $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B_c_196_n N_Y_c_701_n 0.00870364f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B_c_197_n N_Y_c_701_n 0.00870364f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_218 B N_Y_c_701_n 0.0362443f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_219 N_B_c_200_n N_Y_c_701_n 0.00222133f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B_c_196_n N_Y_c_752_n 5.22228e-19 $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B_c_197_n N_Y_c_752_n 0.00630972f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B_c_198_n N_Y_c_752_n 0.0109565f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B_c_198_n N_Y_c_702_n 0.0109318f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_224 B N_Y_c_702_n 0.0516947f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_225 N_B_c_195_n N_Y_c_708_n 0.00113286f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B_c_196_n N_Y_c_708_n 0.00113286f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_227 B N_Y_c_708_n 0.0266272f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_228 N_B_c_200_n N_Y_c_708_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_229 N_B_c_197_n N_Y_c_709_n 0.00113286f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B_c_198_n N_Y_c_709_n 0.00113286f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_231 B N_Y_c_709_n 0.0266272f $X=3.83 $Y=1.105 $X2=0 $Y2=0
cc_232 N_B_c_200_n N_Y_c_709_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_233 N_B_c_195_n N_VGND_c_912_n 0.00146448f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B_c_196_n N_VGND_c_913_n 0.00146448f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B_c_197_n N_VGND_c_913_n 0.00146339f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B_c_195_n N_VGND_c_924_n 0.00423334f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B_c_196_n N_VGND_c_924_n 0.00423334f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B_c_197_n N_VGND_c_931_n 0.00423334f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B_c_198_n N_VGND_c_931_n 0.00423334f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B_c_198_n N_VGND_c_932_n 0.00335921f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B_c_195_n N_VGND_c_934_n 0.0057435f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B_c_196_n N_VGND_c_934_n 0.0057163f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_243 N_B_c_197_n N_VGND_c_934_n 0.0057163f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_244 N_B_c_198_n N_VGND_c_934_n 0.0070399f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_245 N_C_c_276_n N_D_c_350_n 0.0236066f $X=5.63 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_246 N_C_M1030_g N_D_M1017_g 0.0236066f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_247 N_C_c_277_n N_D_c_354_n 0.0185441f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_248 N_C_c_278_n N_D_c_354_n 8.21108e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_249 N_C_c_277_n N_D_c_355_n 2.16854e-19 $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_250 N_C_c_278_n N_D_c_355_n 0.0236066f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_251 N_C_M1001_g N_VPWR_c_495_n 0.00357877f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_252 N_C_M1016_g N_VPWR_c_495_n 0.00357877f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_253 N_C_M1026_g N_VPWR_c_495_n 0.00357877f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_254 N_C_M1030_g N_VPWR_c_495_n 0.00357877f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_255 N_C_M1001_g N_VPWR_c_490_n 0.00655123f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_256 N_C_M1016_g N_VPWR_c_490_n 0.00522516f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_257 N_C_M1026_g N_VPWR_c_490_n 0.00522516f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_258 N_C_M1030_g N_VPWR_c_490_n 0.00525237f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_259 N_C_M1001_g N_A_449_297#_c_584_n 0.0130871f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_260 N_C_c_277_n N_A_449_297#_c_584_n 0.0110239f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_261 N_C_M1016_g N_A_449_297#_c_585_n 0.01094f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_262 N_C_M1026_g N_A_449_297#_c_585_n 0.0109258f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_263 N_C_c_277_n N_A_449_297#_c_585_n 0.0416643f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_264 N_C_c_278_n N_A_449_297#_c_585_n 0.00211509f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_265 N_C_c_277_n N_A_449_297#_c_588_n 0.0204292f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_266 N_C_c_278_n N_A_449_297#_c_588_n 0.00219557f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_267 N_C_M1030_g N_A_449_297#_c_589_n 4.88616e-19 $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_268 N_C_c_277_n N_A_449_297#_c_589_n 0.0204292f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_269 N_C_c_278_n N_A_449_297#_c_589_n 0.00219557f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_270 N_C_M1001_g N_A_807_297#_c_644_n 0.00988743f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_271 N_C_M1016_g N_A_807_297#_c_644_n 0.00984328f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_272 N_C_M1026_g N_A_807_297#_c_646_n 0.00988743f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_273 N_C_M1030_g N_A_807_297#_c_646_n 0.0121747f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_274 N_C_c_273_n N_Y_c_702_n 0.0109318f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_275 N_C_c_277_n N_Y_c_702_n 0.00826974f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_276 N_C_c_273_n N_Y_c_767_n 0.0109565f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_277 N_C_c_274_n N_Y_c_767_n 0.00630972f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_278 N_C_c_275_n N_Y_c_767_n 5.22228e-19 $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_279 N_C_c_274_n N_Y_c_703_n 0.00870364f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_280 N_C_c_275_n N_Y_c_703_n 0.00870364f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_281 N_C_c_277_n N_Y_c_703_n 0.0362443f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_282 N_C_c_278_n N_Y_c_703_n 0.00222133f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_283 N_C_c_274_n N_Y_c_774_n 5.22228e-19 $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_284 N_C_c_275_n N_Y_c_774_n 0.00630972f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_285 N_C_c_276_n N_Y_c_774_n 0.00630972f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_286 N_C_c_276_n N_Y_c_704_n 0.00865686f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_287 N_C_c_277_n N_Y_c_704_n 0.00826974f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_288 N_C_c_276_n N_Y_c_779_n 5.22228e-19 $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_289 N_C_c_273_n N_Y_c_710_n 0.00113286f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_290 N_C_c_274_n N_Y_c_710_n 0.00113286f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_291 N_C_c_277_n N_Y_c_710_n 0.0266272f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_292 N_C_c_278_n N_Y_c_710_n 0.00230339f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_293 N_C_c_275_n N_Y_c_711_n 0.00113286f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_294 N_C_c_276_n N_Y_c_711_n 0.00113286f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_295 N_C_c_277_n N_Y_c_711_n 0.0266272f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_296 N_C_c_278_n N_Y_c_711_n 0.00230339f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_297 N_C_c_274_n N_VGND_c_914_n 0.00146339f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_298 N_C_c_275_n N_VGND_c_914_n 0.00146448f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_299 N_C_c_276_n N_VGND_c_915_n 0.00146448f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_300 N_C_c_273_n N_VGND_c_926_n 0.00423334f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_301 N_C_c_274_n N_VGND_c_926_n 0.00423334f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_302 N_C_c_275_n N_VGND_c_928_n 0.00423334f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_303 N_C_c_276_n N_VGND_c_928_n 0.00423334f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_304 N_C_c_273_n N_VGND_c_932_n 0.00335921f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_305 N_C_c_273_n N_VGND_c_934_n 0.0070399f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_306 N_C_c_274_n N_VGND_c_934_n 0.0057163f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_307 N_C_c_275_n N_VGND_c_934_n 0.0057163f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_308 N_C_c_276_n N_VGND_c_934_n 0.0057435f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_309 N_D_M1017_g N_VPWR_c_495_n 0.00357877f $X=6.05 $Y=1.985 $X2=0 $Y2=0
cc_310 N_D_M1022_g N_VPWR_c_495_n 0.00357877f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_311 N_D_M1028_g N_VPWR_c_495_n 0.00357877f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_312 N_D_M1031_g N_VPWR_c_495_n 0.00357877f $X=7.31 $Y=1.985 $X2=0 $Y2=0
cc_313 N_D_M1017_g N_VPWR_c_490_n 0.00525237f $X=6.05 $Y=1.985 $X2=0 $Y2=0
cc_314 N_D_M1022_g N_VPWR_c_490_n 0.00522516f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_315 N_D_M1028_g N_VPWR_c_490_n 0.00522516f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_316 N_D_M1031_g N_VPWR_c_490_n 0.00621563f $X=7.31 $Y=1.985 $X2=0 $Y2=0
cc_317 N_D_c_354_n N_A_807_297#_c_648_n 0.00247046f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_318 N_D_M1017_g N_A_807_297#_c_649_n 0.0121747f $X=6.05 $Y=1.985 $X2=0 $Y2=0
cc_319 N_D_M1022_g N_A_807_297#_c_649_n 0.00988743f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_320 N_D_M1028_g N_A_807_297#_c_643_n 0.00984328f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_321 N_D_M1031_g N_A_807_297#_c_643_n 0.00988743f $X=7.31 $Y=1.985 $X2=0 $Y2=0
cc_322 N_D_c_350_n N_Y_c_774_n 5.22228e-19 $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_323 N_D_c_350_n N_Y_c_704_n 0.00865686f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_324 N_D_c_354_n N_Y_c_704_n 0.0159556f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_325 N_D_c_350_n N_Y_c_779_n 0.00630972f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_326 N_D_c_351_n N_Y_c_779_n 0.00630972f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_327 N_D_c_352_n N_Y_c_779_n 5.22228e-19 $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_328 N_D_M1022_g N_Y_c_716_n 0.0109258f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_329 N_D_M1028_g N_Y_c_716_n 0.01094f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_330 N_D_c_354_n N_Y_c_716_n 0.0416643f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_331 N_D_c_355_n N_Y_c_716_n 0.00211509f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_332 N_D_c_351_n N_Y_c_705_n 0.00870364f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_333 N_D_c_352_n N_Y_c_705_n 0.00870364f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_334 N_D_c_354_n N_Y_c_705_n 0.0362443f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_335 N_D_c_355_n N_Y_c_705_n 0.00222133f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_336 N_D_c_351_n N_Y_c_802_n 5.22228e-19 $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_337 N_D_c_352_n N_Y_c_802_n 0.00630972f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_338 N_D_c_353_n N_Y_c_802_n 0.0109314f $X=7.31 $Y=0.995 $X2=0 $Y2=0
cc_339 N_D_M1031_g N_Y_c_717_n 0.0135952f $X=7.31 $Y=1.985 $X2=0 $Y2=0
cc_340 N_D_c_354_n N_Y_c_717_n 0.00482295f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_341 N_D_c_353_n N_Y_c_706_n 0.0114045f $X=7.31 $Y=0.995 $X2=0 $Y2=0
cc_342 N_D_c_354_n N_Y_c_706_n 0.00204179f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_343 N_D_c_350_n N_Y_c_712_n 0.00113286f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_344 N_D_c_351_n N_Y_c_712_n 0.00113286f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_345 N_D_c_354_n N_Y_c_712_n 0.0266272f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_346 N_D_c_355_n N_Y_c_712_n 0.00230339f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_347 N_D_M1017_g N_Y_c_718_n 4.88616e-19 $X=6.05 $Y=1.985 $X2=0 $Y2=0
cc_348 N_D_c_354_n N_Y_c_718_n 0.0204292f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_349 N_D_c_355_n N_Y_c_718_n 0.00219557f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_350 N_D_c_352_n N_Y_c_713_n 0.00113286f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_351 N_D_c_353_n N_Y_c_713_n 0.00113286f $X=7.31 $Y=0.995 $X2=0 $Y2=0
cc_352 N_D_c_354_n N_Y_c_713_n 0.0266272f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_353 N_D_c_355_n N_Y_c_713_n 0.00230339f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_354 N_D_c_354_n N_Y_c_719_n 0.0204292f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_355 N_D_c_355_n N_Y_c_719_n 0.00219557f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_356 N_D_c_353_n Y 0.0206984f $X=7.31 $Y=0.995 $X2=0 $Y2=0
cc_357 N_D_c_354_n Y 0.0171924f $X=7.13 $Y=1.16 $X2=0 $Y2=0
cc_358 N_D_c_350_n N_VGND_c_915_n 0.00146448f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_359 N_D_c_350_n N_VGND_c_916_n 0.00423334f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_360 N_D_c_351_n N_VGND_c_916_n 0.00423334f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_361 N_D_c_351_n N_VGND_c_917_n 0.00146448f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_362 N_D_c_352_n N_VGND_c_917_n 0.00146448f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_363 N_D_c_353_n N_VGND_c_919_n 0.00316354f $X=7.31 $Y=0.995 $X2=0 $Y2=0
cc_364 N_D_c_352_n N_VGND_c_930_n 0.00423334f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_365 N_D_c_353_n N_VGND_c_930_n 0.00423334f $X=7.31 $Y=0.995 $X2=0 $Y2=0
cc_366 N_D_c_350_n N_VGND_c_934_n 0.0057435f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_367 N_D_c_351_n N_VGND_c_934_n 0.0057163f $X=6.47 $Y=0.995 $X2=0 $Y2=0
cc_368 N_D_c_352_n N_VGND_c_934_n 0.0057163f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_369 N_D_c_353_n N_VGND_c_934_n 0.00670676f $X=7.31 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A_27_297#_c_430_n N_VPWR_M1003_d 0.00165831f $X=0.995 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_371 N_A_27_297#_c_431_n N_VPWR_M1024_d 0.00165831f $X=1.835 $Y=1.54 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_430_n N_VPWR_c_491_n 0.0126919f $X=0.995 $Y=1.54 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_431_n N_VPWR_c_492_n 0.0126919f $X=1.835 $Y=1.54 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_c_429_n N_VPWR_c_493_n 0.0204682f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_375 N_A_27_297#_c_457_p N_VPWR_c_494_n 0.0142343f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_376 N_A_27_297#_c_458_p N_VPWR_c_495_n 0.0143053f $X=1.96 $Y=2.295 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_c_448_n N_VPWR_c_495_n 0.0330174f $X=2.675 $Y=2.38 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_c_433_n N_VPWR_c_495_n 0.0528834f $X=3.515 $Y=2.38 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_c_461_p N_VPWR_c_495_n 0.0142933f $X=2.8 $Y=2.38 $X2=0 $Y2=0
cc_380 N_A_27_297#_M1003_s N_VPWR_c_490_n 0.00260431f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_M1021_s N_VPWR_c_490_n 0.00284632f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_M1029_s N_VPWR_c_490_n 0.00246446f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_M1014_d N_VPWR_c_490_n 0.00215203f $X=2.665 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_M1025_d N_VPWR_c_490_n 0.0020932f $X=3.505 $Y=1.485 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_c_429_n N_VPWR_c_490_n 0.0120542f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_386 N_A_27_297#_c_457_p N_VPWR_c_490_n 0.00955092f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_387 N_A_27_297#_c_458_p N_VPWR_c_490_n 0.00962794f $X=1.96 $Y=2.295 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_c_448_n N_VPWR_c_490_n 0.0204627f $X=2.675 $Y=2.38 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_c_433_n N_VPWR_c_490_n 0.0322042f $X=3.515 $Y=2.38 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_c_461_p N_VPWR_c_490_n 0.00962421f $X=2.8 $Y=2.38 $X2=0 $Y2=0
cc_391 N_A_27_297#_c_448_n N_A_449_297#_M1002_s 0.00312348f $X=2.675 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_392 N_A_27_297#_c_433_n N_A_449_297#_M1015_s 0.00312348f $X=3.515 $Y=2.38
+ $X2=0 $Y2=0
cc_393 N_A_27_297#_M1014_d N_A_449_297#_c_583_n 0.00165831f $X=2.665 $Y=1.485
+ $X2=0 $Y2=0
cc_394 N_A_27_297#_c_448_n N_A_449_297#_c_583_n 0.00320918f $X=2.675 $Y=2.38
+ $X2=0 $Y2=0
cc_395 N_A_27_297#_c_477_p N_A_449_297#_c_583_n 0.0126766f $X=2.8 $Y=1.96 $X2=0
+ $Y2=0
cc_396 N_A_27_297#_c_433_n N_A_449_297#_c_583_n 0.00320918f $X=3.515 $Y=2.38
+ $X2=0 $Y2=0
cc_397 N_A_27_297#_M1025_d N_A_449_297#_c_584_n 0.00277342f $X=3.505 $Y=1.485
+ $X2=0 $Y2=0
cc_398 N_A_27_297#_c_433_n N_A_449_297#_c_584_n 0.00320918f $X=3.515 $Y=2.38
+ $X2=0 $Y2=0
cc_399 N_A_27_297#_c_434_n N_A_449_297#_c_584_n 0.021051f $X=3.64 $Y=1.96 $X2=0
+ $Y2=0
cc_400 N_A_27_297#_c_432_n N_A_449_297#_c_586_n 0.00271526f $X=1.96 $Y=1.625
+ $X2=0 $Y2=0
cc_401 N_A_27_297#_c_448_n N_A_449_297#_c_586_n 0.0118729f $X=2.675 $Y=2.38
+ $X2=0 $Y2=0
cc_402 N_A_27_297#_c_433_n N_A_449_297#_c_587_n 0.0118729f $X=3.515 $Y=2.38
+ $X2=0 $Y2=0
cc_403 N_A_27_297#_c_434_n N_A_807_297#_c_641_n 0.0384365f $X=3.64 $Y=1.96 $X2=0
+ $Y2=0
cc_404 N_A_27_297#_c_433_n N_A_807_297#_c_642_n 0.0149966f $X=3.515 $Y=2.38
+ $X2=0 $Y2=0
cc_405 N_A_27_297#_c_431_n N_Y_c_700_n 3.18413e-19 $X=1.835 $Y=1.54 $X2=0 $Y2=0
cc_406 N_A_27_297#_c_432_n N_Y_c_700_n 0.00936521f $X=1.96 $Y=1.625 $X2=0 $Y2=0
cc_407 N_A_27_297#_c_428_n N_VGND_c_910_n 0.00367361f $X=0.247 $Y=1.625 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_490_n N_A_449_297#_M1002_s 0.00216833f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_409 N_VPWR_c_490_n N_A_449_297#_M1015_s 0.00216833f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_490_n N_A_449_297#_M1001_d 0.00216833f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_490_n N_A_449_297#_M1026_d 0.00216833f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_490_n N_A_807_297#_M1001_s 0.0020932f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_413 N_VPWR_c_490_n N_A_807_297#_M1016_s 0.00215203f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_490_n N_A_807_297#_M1030_s 0.00215203f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_490_n N_A_807_297#_M1022_d 0.00215203f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_490_n N_A_807_297#_M1031_d 0.0020932f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_495_n N_A_807_297#_c_644_n 0.0330174f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_490_n N_A_807_297#_c_644_n 0.0204627f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_495_n N_A_807_297#_c_642_n 0.0180757f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_490_n N_A_807_297#_c_642_n 0.0107791f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_495_n N_A_807_297#_c_646_n 0.0330174f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_490_n N_A_807_297#_c_646_n 0.0204627f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_495_n N_A_807_297#_c_649_n 0.0330174f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_490_n N_A_807_297#_c_649_n 0.0204627f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_495_n N_A_807_297#_c_643_n 0.0489446f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_490_n N_A_807_297#_c_643_n 0.0300869f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_495_n N_A_807_297#_c_670_n 0.0142933f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_490_n N_A_807_297#_c_670_n 0.00962421f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_495_n N_A_807_297#_c_672_n 0.0142933f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_490_n N_A_807_297#_c_672_n 0.00962421f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_495_n N_A_807_297#_c_674_n 0.0142933f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_490_n N_A_807_297#_c_674_n 0.00962421f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_490_n N_Y_M1017_s 0.00216833f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_434 N_VPWR_c_490_n N_Y_M1028_s 0.00216833f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_435 N_A_449_297#_c_584_n N_A_807_297#_M1001_s 0.00277342f $X=4.455 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_436 N_A_449_297#_c_585_n N_A_807_297#_M1016_s 0.00165831f $X=5.295 $Y=1.54
+ $X2=0 $Y2=0
cc_437 N_A_449_297#_c_584_n N_A_807_297#_c_641_n 0.0189421f $X=4.455 $Y=1.54
+ $X2=0 $Y2=0
cc_438 N_A_449_297#_M1001_d N_A_807_297#_c_644_n 0.00312348f $X=4.445 $Y=1.485
+ $X2=0 $Y2=0
cc_439 N_A_449_297#_c_584_n N_A_807_297#_c_644_n 0.00320918f $X=4.455 $Y=1.54
+ $X2=0 $Y2=0
cc_440 N_A_449_297#_c_585_n N_A_807_297#_c_644_n 0.00320918f $X=5.295 $Y=1.54
+ $X2=0 $Y2=0
cc_441 N_A_449_297#_c_588_n N_A_807_297#_c_644_n 0.0118729f $X=4.58 $Y=1.62
+ $X2=0 $Y2=0
cc_442 N_A_449_297#_c_585_n N_A_807_297#_c_683_n 0.0126766f $X=5.295 $Y=1.54
+ $X2=0 $Y2=0
cc_443 N_A_449_297#_M1026_d N_A_807_297#_c_646_n 0.00312348f $X=5.285 $Y=1.485
+ $X2=0 $Y2=0
cc_444 N_A_449_297#_c_585_n N_A_807_297#_c_646_n 0.00320918f $X=5.295 $Y=1.54
+ $X2=0 $Y2=0
cc_445 N_A_449_297#_c_589_n N_A_807_297#_c_646_n 0.0118729f $X=5.42 $Y=1.62
+ $X2=0 $Y2=0
cc_446 N_A_449_297#_c_584_n N_Y_c_702_n 0.00753964f $X=4.455 $Y=1.54 $X2=0 $Y2=0
cc_447 N_A_449_297#_c_589_n N_Y_c_718_n 0.0011195f $X=5.42 $Y=1.62 $X2=0 $Y2=0
cc_448 N_A_807_297#_c_649_n N_Y_M1017_s 0.00312348f $X=6.555 $Y=2.38 $X2=0 $Y2=0
cc_449 N_A_807_297#_c_643_n N_Y_M1028_s 0.00312348f $X=7.395 $Y=2.38 $X2=0 $Y2=0
cc_450 N_A_807_297#_M1022_d N_Y_c_716_n 0.00165831f $X=6.545 $Y=1.485 $X2=0
+ $Y2=0
cc_451 N_A_807_297#_c_649_n N_Y_c_716_n 0.00320918f $X=6.555 $Y=2.38 $X2=0 $Y2=0
cc_452 N_A_807_297#_c_691_p N_Y_c_716_n 0.0126766f $X=6.68 $Y=1.96 $X2=0 $Y2=0
cc_453 N_A_807_297#_c_643_n N_Y_c_716_n 0.00320918f $X=7.395 $Y=2.38 $X2=0 $Y2=0
cc_454 N_A_807_297#_M1031_d N_Y_c_717_n 0.00283464f $X=7.385 $Y=1.485 $X2=0
+ $Y2=0
cc_455 N_A_807_297#_c_643_n N_Y_c_717_n 0.00320918f $X=7.395 $Y=2.38 $X2=0 $Y2=0
cc_456 N_A_807_297#_c_695_p N_Y_c_717_n 0.0179537f $X=7.52 $Y=1.96 $X2=0 $Y2=0
cc_457 N_A_807_297#_c_649_n N_Y_c_718_n 0.0118729f $X=6.555 $Y=2.38 $X2=0 $Y2=0
cc_458 N_A_807_297#_c_643_n N_Y_c_719_n 0.0118729f $X=7.395 $Y=2.38 $X2=0 $Y2=0
cc_459 N_Y_c_698_n N_VGND_M1010_s 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_460 N_Y_c_700_n N_VGND_M1019_s 0.00162089f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_461 N_Y_c_701_n N_VGND_M1020_d 0.00162089f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_462 N_Y_c_702_n N_VGND_M1027_d 0.0108248f $X=4.415 $Y=0.815 $X2=0 $Y2=0
cc_463 N_Y_c_703_n N_VGND_M1007_d 0.00162089f $X=5.255 $Y=0.815 $X2=0 $Y2=0
cc_464 N_Y_c_704_n N_VGND_M1011_d 0.00162089f $X=6.095 $Y=0.815 $X2=0 $Y2=0
cc_465 N_Y_c_705_n N_VGND_M1005_s 0.00162089f $X=6.935 $Y=0.815 $X2=0 $Y2=0
cc_466 N_Y_c_706_n N_VGND_M1013_s 2.28588e-19 $X=7.465 $Y=0.815 $X2=0 $Y2=0
cc_467 N_Y_c_715_n N_VGND_M1013_s 0.0030148f $X=7.6 $Y=0.905 $X2=0 $Y2=0
cc_468 N_Y_c_699_n N_VGND_c_910_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_469 N_Y_c_698_n N_VGND_c_911_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_470 N_Y_c_700_n N_VGND_c_912_n 0.0122559f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_471 N_Y_c_701_n N_VGND_c_913_n 0.0122559f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_472 N_Y_c_703_n N_VGND_c_914_n 0.0122559f $X=5.255 $Y=0.815 $X2=0 $Y2=0
cc_473 N_Y_c_704_n N_VGND_c_915_n 0.0122559f $X=6.095 $Y=0.815 $X2=0 $Y2=0
cc_474 N_Y_c_704_n N_VGND_c_916_n 0.00198695f $X=6.095 $Y=0.815 $X2=0 $Y2=0
cc_475 N_Y_c_779_n N_VGND_c_916_n 0.0188551f $X=6.26 $Y=0.39 $X2=0 $Y2=0
cc_476 N_Y_c_705_n N_VGND_c_916_n 0.00198695f $X=6.935 $Y=0.815 $X2=0 $Y2=0
cc_477 N_Y_c_705_n N_VGND_c_917_n 0.0122559f $X=6.935 $Y=0.815 $X2=0 $Y2=0
cc_478 N_Y_c_715_n N_VGND_c_918_n 0.00218017f $X=7.6 $Y=0.905 $X2=0 $Y2=0
cc_479 N_Y_c_706_n N_VGND_c_919_n 0.00177288f $X=7.465 $Y=0.815 $X2=0 $Y2=0
cc_480 N_Y_c_715_n N_VGND_c_919_n 0.0120207f $X=7.6 $Y=0.905 $X2=0 $Y2=0
cc_481 N_Y_c_721_n N_VGND_c_920_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_482 N_Y_c_698_n N_VGND_c_920_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_483 N_Y_c_698_n N_VGND_c_922_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_484 N_Y_c_732_n N_VGND_c_922_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_485 N_Y_c_700_n N_VGND_c_922_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_486 N_Y_c_700_n N_VGND_c_924_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_487 N_Y_c_737_n N_VGND_c_924_n 0.0188551f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_488 N_Y_c_701_n N_VGND_c_924_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_489 N_Y_c_702_n N_VGND_c_926_n 0.00198695f $X=4.415 $Y=0.815 $X2=0 $Y2=0
cc_490 N_Y_c_767_n N_VGND_c_926_n 0.0188551f $X=4.58 $Y=0.39 $X2=0 $Y2=0
cc_491 N_Y_c_703_n N_VGND_c_926_n 0.00198695f $X=5.255 $Y=0.815 $X2=0 $Y2=0
cc_492 N_Y_c_703_n N_VGND_c_928_n 0.00198695f $X=5.255 $Y=0.815 $X2=0 $Y2=0
cc_493 N_Y_c_774_n N_VGND_c_928_n 0.0188551f $X=5.42 $Y=0.39 $X2=0 $Y2=0
cc_494 N_Y_c_704_n N_VGND_c_928_n 0.00198695f $X=6.095 $Y=0.815 $X2=0 $Y2=0
cc_495 N_Y_c_705_n N_VGND_c_930_n 0.00198695f $X=6.935 $Y=0.815 $X2=0 $Y2=0
cc_496 N_Y_c_802_n N_VGND_c_930_n 0.0188551f $X=7.1 $Y=0.39 $X2=0 $Y2=0
cc_497 N_Y_c_706_n N_VGND_c_930_n 0.00198695f $X=7.465 $Y=0.815 $X2=0 $Y2=0
cc_498 N_Y_c_701_n N_VGND_c_931_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_499 N_Y_c_752_n N_VGND_c_931_n 0.0188551f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_500 N_Y_c_702_n N_VGND_c_931_n 0.00198695f $X=4.415 $Y=0.815 $X2=0 $Y2=0
cc_501 N_Y_c_702_n N_VGND_c_932_n 0.0528344f $X=4.415 $Y=0.815 $X2=0 $Y2=0
cc_502 N_Y_M1006_d N_VGND_c_934_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_503 N_Y_M1018_d N_VGND_c_934_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_504 N_Y_M1012_s N_VGND_c_934_n 0.00215201f $X=2.245 $Y=0.235 $X2=0 $Y2=0
cc_505 N_Y_M1023_s N_VGND_c_934_n 0.00215201f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_506 N_Y_M1004_s N_VGND_c_934_n 0.00215201f $X=4.445 $Y=0.235 $X2=0 $Y2=0
cc_507 N_Y_M1008_s N_VGND_c_934_n 0.00215201f $X=5.285 $Y=0.235 $X2=0 $Y2=0
cc_508 N_Y_M1000_d N_VGND_c_934_n 0.00215201f $X=6.125 $Y=0.235 $X2=0 $Y2=0
cc_509 N_Y_M1009_d N_VGND_c_934_n 0.00215201f $X=6.965 $Y=0.235 $X2=0 $Y2=0
cc_510 N_Y_c_721_n N_VGND_c_934_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_511 N_Y_c_698_n N_VGND_c_934_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_512 N_Y_c_732_n N_VGND_c_934_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_513 N_Y_c_700_n N_VGND_c_934_n 0.00835832f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_514 N_Y_c_737_n N_VGND_c_934_n 0.0122069f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_515 N_Y_c_701_n N_VGND_c_934_n 0.00835832f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_516 N_Y_c_752_n N_VGND_c_934_n 0.0122069f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_517 N_Y_c_702_n N_VGND_c_934_n 0.0103256f $X=4.415 $Y=0.815 $X2=0 $Y2=0
cc_518 N_Y_c_767_n N_VGND_c_934_n 0.0122069f $X=4.58 $Y=0.39 $X2=0 $Y2=0
cc_519 N_Y_c_703_n N_VGND_c_934_n 0.00835832f $X=5.255 $Y=0.815 $X2=0 $Y2=0
cc_520 N_Y_c_774_n N_VGND_c_934_n 0.0122069f $X=5.42 $Y=0.39 $X2=0 $Y2=0
cc_521 N_Y_c_704_n N_VGND_c_934_n 0.00835832f $X=6.095 $Y=0.815 $X2=0 $Y2=0
cc_522 N_Y_c_779_n N_VGND_c_934_n 0.0122069f $X=6.26 $Y=0.39 $X2=0 $Y2=0
cc_523 N_Y_c_705_n N_VGND_c_934_n 0.00835832f $X=6.935 $Y=0.815 $X2=0 $Y2=0
cc_524 N_Y_c_802_n N_VGND_c_934_n 0.0122069f $X=7.1 $Y=0.39 $X2=0 $Y2=0
cc_525 N_Y_c_706_n N_VGND_c_934_n 0.00396723f $X=7.465 $Y=0.815 $X2=0 $Y2=0
cc_526 N_Y_c_715_n N_VGND_c_934_n 0.00430284f $X=7.6 $Y=0.905 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o22a_2.pxi.spice
* Created: Thu Aug 27 14:37:38 2020
* 
x_PM_SKY130_FD_SC_HD__O22A_2%A_81_21# N_A_81_21#_M1004_d N_A_81_21#_M1007_d
+ N_A_81_21#_c_61_n N_A_81_21#_M1000_g N_A_81_21#_M1001_g N_A_81_21#_c_62_n
+ N_A_81_21#_M1011_g N_A_81_21#_M1010_g N_A_81_21#_c_63_n N_A_81_21#_c_64_n
+ N_A_81_21#_c_65_n N_A_81_21#_c_76_p N_A_81_21#_c_99_p N_A_81_21#_c_87_p
+ N_A_81_21#_c_77_p N_A_81_21#_c_66_n N_A_81_21#_c_67_n
+ PM_SKY130_FD_SC_HD__O22A_2%A_81_21#
x_PM_SKY130_FD_SC_HD__O22A_2%B1 N_B1_c_141_n N_B1_M1004_g N_B1_M1006_g B1
+ N_B1_c_143_n PM_SKY130_FD_SC_HD__O22A_2%B1
x_PM_SKY130_FD_SC_HD__O22A_2%B2 N_B2_M1007_g N_B2_c_173_n N_B2_M1008_g B2
+ N_B2_c_174_n N_B2_c_175_n PM_SKY130_FD_SC_HD__O22A_2%B2
x_PM_SKY130_FD_SC_HD__O22A_2%A2 N_A2_M1005_g N_A2_M1003_g N_A2_c_209_n
+ N_A2_c_210_n A2 N_A2_c_211_n PM_SKY130_FD_SC_HD__O22A_2%A2
x_PM_SKY130_FD_SC_HD__O22A_2%A1 N_A1_M1002_g N_A1_M1009_g A1 A1 N_A1_c_249_n
+ N_A1_c_250_n A1 PM_SKY130_FD_SC_HD__O22A_2%A1
x_PM_SKY130_FD_SC_HD__O22A_2%VPWR N_VPWR_M1001_s N_VPWR_M1010_s N_VPWR_M1002_d
+ N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n VPWR
+ N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_277_n VPWR
+ PM_SKY130_FD_SC_HD__O22A_2%VPWR
x_PM_SKY130_FD_SC_HD__O22A_2%X N_X_M1000_d N_X_M1001_d X N_X_c_324_n
+ PM_SKY130_FD_SC_HD__O22A_2%X
x_PM_SKY130_FD_SC_HD__O22A_2%VGND N_VGND_M1000_s N_VGND_M1011_s N_VGND_M1005_d
+ N_VGND_c_344_n N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n
+ VGND N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n
+ N_VGND_c_353_n VGND PM_SKY130_FD_SC_HD__O22A_2%VGND
x_PM_SKY130_FD_SC_HD__O22A_2%A_301_47# N_A_301_47#_M1004_s N_A_301_47#_M1008_d
+ N_A_301_47#_M1009_d N_A_301_47#_c_398_n N_A_301_47#_c_412_n
+ N_A_301_47#_c_405_n N_A_301_47#_c_399_n N_A_301_47#_c_400_n
+ PM_SKY130_FD_SC_HD__O22A_2%A_301_47#
cc_1 VNB N_A_81_21#_c_61_n 0.0219487f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_2 VNB N_A_81_21#_c_62_n 0.0191669f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_3 VNB N_A_81_21#_c_63_n 0.00193773f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.16
cc_4 VNB N_A_81_21#_c_64_n 0.0618429f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.16
cc_5 VNB N_A_81_21#_c_65_n 3.65884e-19 $X=-0.19 $Y=-0.24 $X2=1.255 $Y2=0.805
cc_6 VNB N_A_81_21#_c_66_n 0.00255278f $X=-0.19 $Y=-0.24 $X2=2.05 $Y2=0.73
cc_7 VNB N_A_81_21#_c_67_n 0.0090959f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.77
cc_8 VNB N_B1_c_141_n 0.0200556f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.235
cc_9 VNB B1 0.00192886f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_10 VNB N_B1_c_143_n 0.0293906f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_11 VNB N_B2_c_173_n 0.0173813f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B2_c_174_n 0.0195875f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_13 VNB N_B2_c_175_n 0.00461989f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_14 VNB N_A2_c_209_n 0.00324628f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_15 VNB N_A2_c_210_n 0.0202316f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_16 VNB N_A2_c_211_n 0.0174493f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.56
cc_17 VNB A1 0.00152499f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_18 VNB N_A1_c_249_n 0.0302901f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_19 VNB N_A1_c_250_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.56
cc_20 VNB A1 0.0111503f $X=-0.19 $Y=-0.24 $X2=1.255 $Y2=0.805
cc_21 VNB N_VPWR_c_277_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_324_n 0.00164538f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_23 VNB N_VGND_c_344_n 0.0113721f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_24 VNB N_VGND_c_345_n 0.00676751f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_25 VNB N_VGND_c_346_n 0.00426509f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.56
cc_26 VNB N_VGND_c_347_n 0.0416551f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_27 VNB N_VGND_c_348_n 0.0046757f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.495
cc_28 VNB N_VGND_c_349_n 0.0194554f $X=-0.19 $Y=-0.24 $X2=1.85 $Y2=0.805
cc_29 VNB N_VGND_c_350_n 0.0174149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_351_n 0.204752f $X=-0.19 $Y=-0.24 $X2=2.05 $Y2=0.77
cc_31 VNB N_VGND_c_352_n 0.00343497f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_32 VNB N_VGND_c_353_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_33 VNB N_A_301_47#_c_398_n 0.00245031f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_34 VNB N_A_301_47#_c_399_n 0.00765088f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.56
cc_35 VNB N_A_301_47#_c_400_n 0.0164654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A_81_21#_M1001_g 0.0249029f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_37 VPB N_A_81_21#_M1010_g 0.0229735f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_38 VPB N_A_81_21#_c_63_n 0.00220215f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.16
cc_39 VPB N_A_81_21#_c_64_n 0.0144495f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.16
cc_40 VPB N_B1_M1006_g 0.0217335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB B1 0.00316058f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_42 VPB N_B1_c_143_n 0.00929324f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.995
cc_43 VPB N_B2_M1007_g 0.0203739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_B2_c_174_n 0.00397859f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_45 VPB N_B2_c_175_n 0.00203056f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_46 VPB N_A2_M1003_g 0.0184111f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A2_c_209_n 0.011661f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_48 VPB N_A2_c_210_n 0.00501346f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_49 VPB N_A1_M1002_g 0.0214445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB A1 0.0133558f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_51 VPB N_A1_c_249_n 0.00746684f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.995
cc_52 VPB N_VPWR_c_278_n 0.0106521f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.325
cc_53 VPB N_VPWR_c_279_n 0.0491869f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_54 VPB N_VPWR_c_280_n 0.0112011f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.56
cc_55 VPB N_VPWR_c_281_n 0.0329646f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_56 VPB N_VPWR_c_282_n 0.0180122f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.495
cc_57 VPB N_VPWR_c_283_n 0.0404458f $X=-0.19 $Y=1.305 $X2=1.255 $Y2=0.805
cc_58 VPB N_VPWR_c_284_n 0.0189908f $X=-0.19 $Y=1.305 $X2=2.41 $Y2=1.62
cc_59 VPB N_VPWR_c_277_n 0.0438461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_X_c_324_n 0.00228298f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.325
cc_61 N_A_81_21#_c_63_n N_B1_c_141_n 0.00252022f $X=1.135 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_62 N_A_81_21#_c_66_n N_B1_c_141_n 0.0070416f $X=2.05 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_63 N_A_81_21#_c_67_n N_B1_c_141_n 0.00900801f $X=1.85 $Y=0.77 $X2=-0.19
+ $Y2=-0.24
cc_64 N_A_81_21#_c_63_n N_B1_M1006_g 0.00430219f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_81_21#_c_76_p N_B1_M1006_g 0.0193911f $X=2.19 $Y=1.6 $X2=0 $Y2=0
cc_66 N_A_81_21#_c_77_p N_B1_M1006_g 0.00272508f $X=2.41 $Y=2.3 $X2=0 $Y2=0
cc_67 N_A_81_21#_c_63_n B1 0.0188413f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_81_21#_c_64_n B1 0.00166115f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_81_21#_c_76_p B1 0.0240683f $X=2.19 $Y=1.6 $X2=0 $Y2=0
cc_70 N_A_81_21#_c_67_n B1 0.0252393f $X=1.85 $Y=0.77 $X2=0 $Y2=0
cc_71 N_A_81_21#_c_63_n N_B1_c_143_n 8.36259e-19 $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_81_21#_c_64_n N_B1_c_143_n 0.0212333f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_81_21#_c_76_p N_B1_c_143_n 0.00183798f $X=2.19 $Y=1.6 $X2=0 $Y2=0
cc_74 N_A_81_21#_c_67_n N_B1_c_143_n 0.00674077f $X=1.85 $Y=0.77 $X2=0 $Y2=0
cc_75 N_A_81_21#_c_76_p N_B2_M1007_g 0.00684637f $X=2.19 $Y=1.6 $X2=0 $Y2=0
cc_76 N_A_81_21#_c_87_p N_B2_M1007_g 0.00287872f $X=2.382 $Y=1.705 $X2=0 $Y2=0
cc_77 N_A_81_21#_c_77_p N_B2_M1007_g 0.0155164f $X=2.41 $Y=2.3 $X2=0 $Y2=0
cc_78 N_A_81_21#_c_66_n N_B2_c_173_n 0.00406178f $X=2.05 $Y=0.73 $X2=0 $Y2=0
cc_79 N_A_81_21#_c_87_p N_B2_c_174_n 0.00285844f $X=2.382 $Y=1.705 $X2=0 $Y2=0
cc_80 N_A_81_21#_c_66_n N_B2_c_174_n 0.00173935f $X=2.05 $Y=0.73 $X2=0 $Y2=0
cc_81 N_A_81_21#_c_76_p N_B2_c_175_n 0.0147636f $X=2.19 $Y=1.6 $X2=0 $Y2=0
cc_82 N_A_81_21#_c_87_p N_B2_c_175_n 0.0163217f $X=2.382 $Y=1.705 $X2=0 $Y2=0
cc_83 N_A_81_21#_c_66_n N_B2_c_175_n 0.0190747f $X=2.05 $Y=0.73 $X2=0 $Y2=0
cc_84 N_A_81_21#_c_87_p N_A2_M1003_g 0.00151222f $X=2.382 $Y=1.705 $X2=0 $Y2=0
cc_85 N_A_81_21#_c_77_p N_A2_M1003_g 0.00854089f $X=2.41 $Y=2.3 $X2=0 $Y2=0
cc_86 N_A_81_21#_c_87_p N_A2_c_209_n 0.0100102f $X=2.382 $Y=1.705 $X2=0 $Y2=0
cc_87 N_A_81_21#_c_76_p N_VPWR_M1010_s 0.0141621f $X=2.19 $Y=1.6 $X2=0 $Y2=0
cc_88 N_A_81_21#_c_99_p N_VPWR_M1010_s 0.00334235f $X=1.255 $Y=1.6 $X2=0 $Y2=0
cc_89 N_A_81_21#_M1001_g N_VPWR_c_279_n 0.00409084f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_81_21#_M1001_g N_VPWR_c_282_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_81_21#_M1010_g N_VPWR_c_282_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_81_21#_c_77_p N_VPWR_c_283_n 0.0247344f $X=2.41 $Y=2.3 $X2=0 $Y2=0
cc_93 N_A_81_21#_M1010_g N_VPWR_c_284_n 0.00359017f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_81_21#_c_64_n N_VPWR_c_284_n 8.99354e-19 $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_81_21#_c_76_p N_VPWR_c_284_n 0.0395491f $X=2.19 $Y=1.6 $X2=0 $Y2=0
cc_96 N_A_81_21#_c_99_p N_VPWR_c_284_n 0.0191594f $X=1.255 $Y=1.6 $X2=0 $Y2=0
cc_97 N_A_81_21#_c_77_p N_VPWR_c_284_n 0.0240359f $X=2.41 $Y=2.3 $X2=0 $Y2=0
cc_98 N_A_81_21#_M1007_d N_VPWR_c_277_n 0.00972089f $X=2.275 $Y=1.485 $X2=0
+ $Y2=0
cc_99 N_A_81_21#_M1001_g N_VPWR_c_277_n 0.01151f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_81_21#_M1010_g N_VPWR_c_277_n 0.0117629f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_81_21#_c_77_p N_VPWR_c_277_n 0.0142934f $X=2.41 $Y=2.3 $X2=0 $Y2=0
cc_102 N_A_81_21#_c_61_n N_X_c_324_n 0.00332776f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_81_21#_M1001_g N_X_c_324_n 0.00342089f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_81_21#_c_62_n N_X_c_324_n 0.00139262f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_81_21#_M1010_g N_X_c_324_n 0.00117471f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_81_21#_c_63_n N_X_c_324_n 0.0439327f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_81_21#_c_64_n N_X_c_324_n 0.0285698f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_81_21#_c_65_n N_X_c_324_n 0.00793472f $X=1.255 $Y=0.805 $X2=0 $Y2=0
cc_109 N_A_81_21#_c_76_p A_383_297# 0.00478751f $X=2.19 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_81_21#_c_65_n N_VGND_M1011_s 0.00357679f $X=1.255 $Y=0.805 $X2=0
+ $Y2=0
cc_111 N_A_81_21#_c_61_n N_VGND_c_345_n 0.00316354f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_81_21#_c_62_n N_VGND_c_346_n 0.00317069f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_81_21#_c_64_n N_VGND_c_346_n 7.44251e-19 $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_81_21#_c_65_n N_VGND_c_346_n 0.0148358f $X=1.255 $Y=0.805 $X2=0 $Y2=0
cc_115 N_A_81_21#_c_65_n N_VGND_c_347_n 8.30317e-19 $X=1.255 $Y=0.805 $X2=0
+ $Y2=0
cc_116 N_A_81_21#_c_67_n N_VGND_c_347_n 0.00326925f $X=1.85 $Y=0.77 $X2=0 $Y2=0
cc_117 N_A_81_21#_c_61_n N_VGND_c_349_n 0.00585385f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_81_21#_c_62_n N_VGND_c_349_n 0.00585385f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_81_21#_M1004_d N_VGND_c_351_n 0.00219239f $X=1.915 $Y=0.235 $X2=0
+ $Y2=0
cc_120 N_A_81_21#_c_61_n N_VGND_c_351_n 0.0115767f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_81_21#_c_62_n N_VGND_c_351_n 0.0119391f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_81_21#_c_65_n N_VGND_c_351_n 0.00364224f $X=1.255 $Y=0.805 $X2=0
+ $Y2=0
cc_123 N_A_81_21#_c_67_n N_VGND_c_351_n 0.00647238f $X=1.85 $Y=0.77 $X2=0 $Y2=0
cc_124 N_A_81_21#_c_67_n N_A_301_47#_M1004_s 0.0031941f $X=1.85 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_125 N_A_81_21#_M1004_d N_A_301_47#_c_398_n 0.00323205f $X=1.915 $Y=0.235
+ $X2=0 $Y2=0
cc_126 N_A_81_21#_c_66_n N_A_301_47#_c_398_n 0.0173867f $X=2.05 $Y=0.73 $X2=0
+ $Y2=0
cc_127 N_A_81_21#_c_67_n N_A_301_47#_c_398_n 0.0167975f $X=1.85 $Y=0.77 $X2=0
+ $Y2=0
cc_128 N_A_81_21#_c_87_p N_A_301_47#_c_405_n 0.00472356f $X=2.382 $Y=1.705 $X2=0
+ $Y2=0
cc_129 N_A_81_21#_c_66_n N_A_301_47#_c_405_n 0.00202176f $X=2.05 $Y=0.73 $X2=0
+ $Y2=0
cc_130 N_B1_M1006_g N_B2_M1007_g 0.0499661f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_131 N_B1_c_141_n N_B2_c_173_n 0.0270126f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_c_143_n N_B2_c_174_n 0.0499661f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_133 B1 N_B2_c_175_n 0.0203744f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B1_c_143_n N_B2_c_175_n 0.00193188f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B1_M1006_g N_VPWR_c_283_n 0.00468308f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B1_M1006_g N_VPWR_c_284_n 0.0161839f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B1_M1006_g N_VPWR_c_277_n 0.00783315f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B1_c_141_n N_VGND_c_346_n 0.0024683f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_141_n N_VGND_c_347_n 0.00366111f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_c_141_n N_VGND_c_351_n 0.0065944f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B1_c_141_n N_A_301_47#_c_398_n 0.00833791f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B2_M1007_g N_A2_M1003_g 0.0156126f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B2_M1007_g N_A2_c_209_n 8.99156e-19 $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B2_c_174_n N_A2_c_209_n 7.56644e-19 $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B2_c_175_n N_A2_c_209_n 0.021387f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B2_c_174_n N_A2_c_210_n 0.0219996f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B2_c_175_n N_A2_c_210_n 8.4425e-19 $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B2_c_173_n N_A2_c_211_n 0.0171094f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_149 N_B2_M1007_g N_VPWR_c_283_n 0.00457863f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B2_M1007_g N_VPWR_c_284_n 0.00285115f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B2_M1007_g N_VPWR_c_277_n 0.00797339f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B2_c_173_n N_VGND_c_347_n 0.00366111f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B2_c_173_n N_VGND_c_351_n 0.00559166f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B2_c_173_n N_A_301_47#_c_398_n 0.0124132f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B2_c_175_n N_A_301_47#_c_398_n 0.00366332f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B2_c_173_n N_A_301_47#_c_405_n 3.64847e-19 $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_157 N_B2_c_175_n N_A_301_47#_c_405_n 0.00212316f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A2_M1003_g N_A1_M1002_g 0.0468173f $X=2.82 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A2_c_209_n N_A1_M1002_g 7.59081e-19 $X=3 $Y=1.615 $X2=0 $Y2=0
cc_160 N_A2_c_209_n A1 0.0114464f $X=3 $Y=1.615 $X2=0 $Y2=0
cc_161 N_A2_c_209_n N_A1_c_249_n 0.00184122f $X=3 $Y=1.615 $X2=0 $Y2=0
cc_162 N_A2_c_210_n N_A1_c_249_n 0.0468173f $X=2.76 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A2_c_211_n N_A1_c_250_n 0.0275186f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_209_n A1 0.0175849f $X=3 $Y=1.615 $X2=0 $Y2=0
cc_165 N_A2_c_210_n A1 6.49721e-19 $X=2.76 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A2_M1003_g N_VPWR_c_283_n 0.00585385f $X=2.82 $Y=1.985 $X2=0 $Y2=0
cc_167 A2 N_VPWR_c_283_n 0.00754929f $X=2.9 $Y=1.785 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VPWR_c_277_n 0.011136f $X=2.82 $Y=1.985 $X2=0 $Y2=0
cc_169 A2 N_VPWR_c_277_n 0.00739369f $X=2.9 $Y=1.785 $X2=0 $Y2=0
cc_170 A2 A_579_297# 0.00430709f $X=2.9 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_171 N_A2_c_211_n N_VGND_c_347_n 0.00426936f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_211_n N_VGND_c_348_n 0.00268723f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_211_n N_VGND_c_351_n 0.00604464f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A2_c_211_n N_A_301_47#_c_412_n 0.00190722f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A2_c_209_n N_A_301_47#_c_405_n 0.00702467f $X=3 $Y=1.615 $X2=0 $Y2=0
cc_176 N_A2_c_210_n N_A_301_47#_c_405_n 0.00252674f $X=2.76 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A2_c_211_n N_A_301_47#_c_405_n 0.00373752f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A2_c_209_n N_A_301_47#_c_399_n 0.0163473f $X=3 $Y=1.615 $X2=0 $Y2=0
cc_179 N_A2_c_211_n N_A_301_47#_c_399_n 0.00935532f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_211_n N_A_301_47#_c_400_n 5.09218e-19 $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_181 A1 N_VPWR_M1002_d 0.00383293f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_182 N_A1_M1002_g N_VPWR_c_281_n 0.00485839f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_183 A1 N_VPWR_c_281_n 0.0229358f $X=3.36 $Y=1.445 $X2=0 $Y2=0
cc_184 N_A1_c_249_n N_VPWR_c_281_n 6.61872e-19 $X=3.29 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A1_M1002_g N_VPWR_c_283_n 0.00585385f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A1_M1002_g N_VPWR_c_277_n 0.0113724f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A1_c_250_n N_VGND_c_348_n 0.00268723f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_250_n N_VGND_c_350_n 0.00421028f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_250_n N_VGND_c_351_n 0.00663995f $X=3.275 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A1_c_250_n N_A_301_47#_c_405_n 4.38799e-19 $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A1_c_249_n N_A_301_47#_c_399_n 0.00377739f $X=3.29 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A1_c_250_n N_A_301_47#_c_399_n 0.00944054f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_193 A1 N_A_301_47#_c_399_n 0.0289691f $X=3.45 $Y=1.19 $X2=0 $Y2=0
cc_194 N_A1_c_250_n N_A_301_47#_c_400_n 0.00581008f $X=3.275 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_277_n N_X_M1001_d 0.00406137f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_c_279_n N_X_c_324_n 0.00252736f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_197 N_VPWR_c_282_n N_X_c_324_n 0.0129925f $X=0.995 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_277_n N_X_c_324_n 0.008203f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_277_n A_383_297# 0.00897657f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_200 N_VPWR_c_277_n A_579_297# 0.00213575f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_201 N_VPWR_c_279_n N_VGND_c_345_n 0.00641101f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_202 N_X_c_324_n N_VGND_c_349_n 0.00762694f $X=0.69 $Y=0.595 $X2=0 $Y2=0
cc_203 N_X_M1000_d N_VGND_c_351_n 0.0042453f $X=0.555 $Y=0.235 $X2=0 $Y2=0
cc_204 N_X_c_324_n N_VGND_c_351_n 0.00772384f $X=0.69 $Y=0.595 $X2=0 $Y2=0
cc_205 N_VGND_c_351_n N_A_301_47#_M1004_s 0.00211652f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_206 N_VGND_c_351_n N_A_301_47#_M1008_d 0.00307637f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_351_n N_A_301_47#_M1009_d 0.00210425f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_208 N_VGND_c_346_n N_A_301_47#_c_398_n 0.0109504f $X=1.11 $Y=0.38 $X2=0 $Y2=0
cc_209 N_VGND_c_347_n N_A_301_47#_c_398_n 0.0414486f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_351_n N_A_301_47#_c_398_n 0.0321925f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_347_n N_A_301_47#_c_412_n 0.0171071f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_351_n N_A_301_47#_c_412_n 0.0126031f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_M1005_d N_A_301_47#_c_399_n 0.0046001f $X=2.865 $Y=0.235 $X2=0
+ $Y2=0
cc_214 N_VGND_c_347_n N_A_301_47#_c_399_n 0.00233346f $X=2.915 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_348_n N_A_301_47#_c_399_n 0.012114f $X=3 $Y=0.36 $X2=0 $Y2=0
cc_216 N_VGND_c_350_n N_A_301_47#_c_399_n 0.00211912f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_351_n N_A_301_47#_c_399_n 0.00890555f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_350_n N_A_301_47#_c_400_n 0.0182739f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_351_n N_A_301_47#_c_400_n 0.0124095f $X=3.45 $Y=0 $X2=0 $Y2=0

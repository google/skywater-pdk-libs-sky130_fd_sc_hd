# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a21o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.990000 1.010000 4.515000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425000 1.010000 3.820000 1.275000 ;
        RECT 3.645000 1.275000 3.820000 1.510000 ;
        RECT 3.645000 1.510000 4.935000 1.680000 ;
        RECT 4.685000 1.055000 5.100000 1.290000 ;
        RECT 4.685000 1.290000 4.935000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 0.995000 2.705000 1.525000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 1.735000 0.785000 ;
        RECT 0.145000 0.785000 0.630000 1.585000 ;
        RECT 0.145000 1.585000 1.735000 1.755000 ;
        RECT 0.625000 1.755000 0.795000 2.185000 ;
        RECT 1.485000 1.755000 1.735000 2.185000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 0.105000  0.085000 0.445000 0.445000 ;
        RECT 0.975000  0.085000 1.305000 0.445000 ;
        RECT 1.910000  0.085000 2.685000 0.445000 ;
        RECT 3.255000  0.085000 3.585000 0.445000 ;
        RECT 4.945000  0.085000 5.225000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.115000 1.935000 0.445000 2.635000 ;
        RECT 0.975000 1.935000 1.305000 2.635000 ;
        RECT 1.915000 1.515000 2.165000 2.635000 ;
        RECT 3.635000 2.275000 3.965000 2.635000 ;
        RECT 4.475000 2.275000 4.805000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.800000 0.995000 2.205000 1.325000 ;
      RECT 2.035000 0.615000 3.045000 0.670000 ;
      RECT 2.035000 0.670000 4.365000 0.785000 ;
      RECT 2.035000 0.785000 2.205000 0.995000 ;
      RECT 2.455000 1.695000 2.625000 2.295000 ;
      RECT 2.455000 2.295000 3.465000 2.465000 ;
      RECT 2.875000 0.255000 3.045000 0.615000 ;
      RECT 2.875000 0.785000 4.365000 0.840000 ;
      RECT 2.875000 0.840000 3.045000 2.125000 ;
      RECT 3.285000 1.445000 3.465000 1.850000 ;
      RECT 3.285000 1.850000 5.360000 2.020000 ;
      RECT 3.285000 2.020000 3.465000 2.295000 ;
      RECT 4.085000 0.405000 4.365000 0.670000 ;
      RECT 4.135000 2.020000 4.305000 2.465000 ;
      RECT 5.030000 2.020000 5.360000 2.395000 ;
      RECT 5.105000 1.460000 5.360000 1.850000 ;
  END
END sky130_fd_sc_hd__a21o_4

* File: sky130_fd_sc_hd__probec_p_8.spice
* Created: Tue Sep  1 19:29:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__probec_p_8.pex.spice"
.subckt sky130_fd_sc_hd__probec_p_8  VNB VPB A VPWR VGND X
* 
* X	X
* VGND	VGND
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_A_27_47#_M1007_d N_A_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1012 N_A_27_47#_M1012_d N_A_M1012_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1021 N_A_27_47#_M1012_d N_A_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1000 N_noxref_6_M1000_d N_A_27_47#_M1000_g N_VGND_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1003 N_noxref_6_M1000_d N_A_27_47#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1009 N_noxref_6_M1009_d N_A_27_47#_M1009_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1010 N_noxref_6_M1009_d N_A_27_47#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1014 N_noxref_6_M1014_d N_A_27_47#_M1014_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1016 N_noxref_6_M1014_d N_A_27_47#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75001 A=0.0975 P=1.6 MULT=1
MM1017 N_noxref_6_M1017_d N_A_27_47#_M1017_g N_VGND_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75004 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_noxref_6_M1017_d N_A_27_47#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75004.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1002_d N_A_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1013_d N_A_27_47#_M1001_g N_noxref_6_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_27_47#_M1005_g N_noxref_6_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1005_d N_A_27_47#_M1006_g N_noxref_6_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_47#_M1008_g N_noxref_6_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1008_d N_A_27_47#_M1011_g N_noxref_6_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_27_47#_M1015_g N_noxref_6_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1015_d N_A_27_47#_M1019_g N_noxref_6_M1019_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1020_d N_A_27_47#_M1020_g N_noxref_6_M1019_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=9.4695 P=15.01
R23_noxref N_X_R23_noxref_pos N_noxref_6_R23_noxref_neg SHORT 0.01 M=1
R24_noxref noxref_9 N_VGND_R24_noxref_neg SHORT 0.01 M=1
R25_noxref noxref_10 N_VPWR_R25_noxref_neg SHORT 0.01 M=1
c_84 VNB 0 2.5355e-19 $X=0.15 $Y=-0.085
c_144 VPB 0 1.73336e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__probec_p_8.pxi.spice"
*
.ends
*
*

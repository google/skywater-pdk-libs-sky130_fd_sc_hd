* File: sky130_fd_sc_hd__o31a_4.pxi.spice
* Created: Tue Sep  1 19:25:17 2020
* 
x_PM_SKY130_FD_SC_HD__O31A_4%A_102_21# N_A_102_21#_M1016_d N_A_102_21#_M1006_s
+ N_A_102_21#_M1000_d N_A_102_21#_M1002_g N_A_102_21#_M1003_g
+ N_A_102_21#_M1007_g N_A_102_21#_M1015_g N_A_102_21#_M1008_g
+ N_A_102_21#_M1022_g N_A_102_21#_M1010_g N_A_102_21#_M1023_g
+ N_A_102_21#_c_120_n N_A_102_21#_c_121_n N_A_102_21#_c_122_n
+ N_A_102_21#_c_130_n N_A_102_21#_c_134_p N_A_102_21#_c_123_n
+ N_A_102_21#_c_138_p N_A_102_21#_c_131_n N_A_102_21#_c_139_p
+ N_A_102_21#_c_169_p N_A_102_21#_c_156_p N_A_102_21#_c_124_n
+ N_A_102_21#_c_125_n PM_SKY130_FD_SC_HD__O31A_4%A_102_21#
x_PM_SKY130_FD_SC_HD__O31A_4%B1 N_B1_M1006_g N_B1_c_237_n N_B1_c_238_n
+ N_B1_M1018_g N_B1_M1016_g N_B1_M1021_g B1 B1 B1 N_B1_c_247_n N_B1_c_243_n
+ PM_SKY130_FD_SC_HD__O31A_4%B1
x_PM_SKY130_FD_SC_HD__O31A_4%A3 N_A3_M1012_g N_A3_M1000_g N_A3_M1014_g
+ N_A3_M1020_g A3 N_A3_c_306_n PM_SKY130_FD_SC_HD__O31A_4%A3
x_PM_SKY130_FD_SC_HD__O31A_4%A2 N_A2_c_347_n N_A2_M1009_g N_A2_M1011_g
+ N_A2_M1013_g N_A2_M1017_g A2 A2 A2 A2 A2 N_A2_c_351_n N_A2_c_352_n
+ N_A2_c_353_n N_A2_c_354_n N_A2_c_372_p PM_SKY130_FD_SC_HD__O31A_4%A2
x_PM_SKY130_FD_SC_HD__O31A_4%A1 N_A1_M1004_g N_A1_M1001_g N_A1_M1005_g
+ N_A1_M1019_g A1 N_A1_c_440_n PM_SKY130_FD_SC_HD__O31A_4%A1
x_PM_SKY130_FD_SC_HD__O31A_4%VPWR N_VPWR_M1003_s N_VPWR_M1015_s N_VPWR_M1023_s
+ N_VPWR_M1018_d N_VPWR_M1001_d N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n
+ N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n VPWR N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_488_n
+ N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n VPWR
+ PM_SKY130_FD_SC_HD__O31A_4%VPWR
x_PM_SKY130_FD_SC_HD__O31A_4%X N_X_M1002_s N_X_M1008_s N_X_M1003_d N_X_M1022_d
+ N_X_c_601_n N_X_c_627_n N_X_c_611_n N_X_c_604_n N_X_c_632_n N_X_c_602_n X X X
+ N_X_c_640_p PM_SKY130_FD_SC_HD__O31A_4%X
x_PM_SKY130_FD_SC_HD__O31A_4%A_672_297# N_A_672_297#_M1000_s
+ N_A_672_297#_M1020_s N_A_672_297#_M1017_s N_A_672_297#_c_649_n
+ N_A_672_297#_c_670_n N_A_672_297#_c_656_n N_A_672_297#_c_650_n
+ N_A_672_297#_c_651_n N_A_672_297#_c_657_n
+ PM_SKY130_FD_SC_HD__O31A_4%A_672_297#
x_PM_SKY130_FD_SC_HD__O31A_4%A_926_297# N_A_926_297#_M1011_d
+ N_A_926_297#_M1019_s N_A_926_297#_c_712_n N_A_926_297#_c_714_n
+ N_A_926_297#_c_716_n PM_SKY130_FD_SC_HD__O31A_4%A_926_297#
x_PM_SKY130_FD_SC_HD__O31A_4%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_M1010_d
+ N_VGND_M1012_s N_VGND_M1009_d N_VGND_M1005_s N_VGND_c_743_n N_VGND_c_744_n
+ N_VGND_c_745_n N_VGND_c_746_n N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n
+ N_VGND_c_750_n N_VGND_c_751_n VGND N_VGND_c_752_n N_VGND_c_753_n
+ N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n
+ N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n VGND
+ PM_SKY130_FD_SC_HD__O31A_4%VGND
x_PM_SKY130_FD_SC_HD__O31A_4%A_496_47# N_A_496_47#_M1016_s N_A_496_47#_M1021_s
+ N_A_496_47#_M1014_d N_A_496_47#_M1004_d N_A_496_47#_M1013_s
+ N_A_496_47#_c_854_n N_A_496_47#_c_868_n N_A_496_47#_c_855_n
+ N_A_496_47#_c_908_n N_A_496_47#_c_875_n N_A_496_47#_c_915_n
+ N_A_496_47#_c_880_n N_A_496_47#_c_856_n N_A_496_47#_c_857_n
+ N_A_496_47#_c_858_n PM_SKY130_FD_SC_HD__O31A_4%A_496_47#
cc_1 VNB N_A_102_21#_M1002_g 0.0211452f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.56
cc_2 VNB N_A_102_21#_M1003_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.985
cc_3 VNB N_A_102_21#_M1007_g 0.0176246f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.56
cc_4 VNB N_A_102_21#_M1015_g 4.59465e-19 $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.985
cc_5 VNB N_A_102_21#_M1008_g 0.0176414f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=0.56
cc_6 VNB N_A_102_21#_M1022_g 4.61158e-19 $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.985
cc_7 VNB N_A_102_21#_M1010_g 0.0208949f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=0.56
cc_8 VNB N_A_102_21#_M1023_g 4.65423e-19 $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.985
cc_9 VNB N_A_102_21#_c_120_n 0.0282584f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.16
cc_10 VNB N_A_102_21#_c_121_n 0.00497882f $X=-0.19 $Y=-0.24 $X2=2.44 $Y2=1.172
cc_11 VNB N_A_102_21#_c_122_n 0.00308414f $X=-0.19 $Y=-0.24 $X2=2.525 $Y2=1.055
cc_12 VNB N_A_102_21#_c_123_n 0.00253506f $X=-0.19 $Y=-0.24 $X2=2.61 $Y2=0.76
cc_13 VNB N_A_102_21#_c_124_n 0.0141683f $X=-0.19 $Y=-0.24 $X2=1.38 $Y2=1.16
cc_14 VNB N_A_102_21#_c_125_n 0.0242415f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.16
cc_15 VNB N_B1_M1006_g 4.70252e-19 $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.485
cc_16 VNB N_B1_c_237_n 0.0213313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B1_c_238_n 0.0154621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B1_M1018_g 5.58873e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B1_M1016_g 0.0208485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B1_M1021_g 0.0181923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB B1 0.00471848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_B1_c_243_n 0.0428089f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.295
cc_23 VNB N_A3_M1012_g 0.0179351f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.485
cc_24 VNB N_A3_M1000_g 4.50909e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A3_M1014_g 0.017453f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.56
cc_26 VNB N_A3_M1020_g 4.04481e-19 $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.985
cc_27 VNB N_A3_c_306_n 0.0311121f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.985
cc_28 VNB N_A2_c_347_n 0.0161679f $X=-0.19 $Y=-0.24 $X2=2.91 $Y2=0.235
cc_29 VNB N_A2_M1013_g 0.0243253f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.025
cc_30 VNB N_A2_M1017_g 5.17518e-19 $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.295
cc_31 VNB A2 0.0163048f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.985
cc_32 VNB N_A2_c_351_n 0.0187919f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.025
cc_33 VNB N_A2_c_352_n 0.0308707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A2_c_353_n 0.00290978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A2_c_354_n 0.00197022f $X=-0.19 $Y=-0.24 $X2=2.44 $Y2=1.172
cc_36 VNB N_A1_M1004_g 0.0174081f $X=-0.19 $Y=-0.24 $X2=3.79 $Y2=1.485
cc_37 VNB N_A1_M1001_g 3.8603e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A1_M1005_g 0.0174782f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.56
cc_39 VNB N_A1_M1019_g 4.25865e-19 $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.985
cc_40 VNB N_A1_c_440_n 0.0291202f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.985
cc_41 VNB N_VPWR_c_488_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_X_c_601_n 0.0327538f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.985
cc_43 VNB N_X_c_602_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.295
cc_44 VNB N_VGND_c_743_n 0.0130579f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.56
cc_45 VNB N_VGND_c_744_n 0.0206934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_745_n 3.15299e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_746_n 0.0119367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_747_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_748_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_749_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_750_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_751_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.16
cc_53 VNB N_VGND_c_752_n 0.0131583f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=1.16
cc_54 VNB N_VGND_c_753_n 0.0124296f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.16
cc_55 VNB N_VGND_c_754_n 0.0352128f $X=-0.19 $Y=-0.24 $X2=2.525 $Y2=1.815
cc_56 VNB N_VGND_c_755_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_756_n 0.0177682f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=1.16
cc_58 VNB N_VGND_c_757_n 0.322593f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.16
cc_59 VNB N_VGND_c_758_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_759_n 0.00490497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_760_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_761_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_496_47#_c_854_n 0.00245154f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.985
cc_64 VNB N_A_496_47#_c_855_n 0.00171622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_496_47#_c_856_n 0.00143487f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=0.56
cc_66 VNB N_A_496_47#_c_857_n 0.00140707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_496_47#_c_858_n 0.033759f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.985
cc_68 VPB N_A_102_21#_M1003_g 0.0234995f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.985
cc_69 VPB N_A_102_21#_M1015_g 0.0195304f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.985
cc_70 VPB N_A_102_21#_M1022_g 0.0195501f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_71 VPB N_A_102_21#_M1023_g 0.0194758f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.985
cc_72 VPB N_A_102_21#_c_130_n 0.00265825f $X=-0.19 $Y=1.305 $X2=2.525 $Y2=1.815
cc_73 VPB N_A_102_21#_c_131_n 0.0081319f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.97
cc_74 VPB N_B1_M1006_g 0.019687f $X=-0.19 $Y=1.305 $X2=3.79 $Y2=1.485
cc_75 VPB N_B1_M1018_g 0.0236146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB B1 0.00543253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_B1_c_247_n 0.00483343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A3_M1000_g 0.023664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A3_M1020_g 0.0196053f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.985
cc_80 VPB A3 0.0025009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A2_M1011_g 0.0187229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A2_M1017_g 0.0236032f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.295
cc_83 VPB A2 0.00119136f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=0.56
cc_84 VPB A2 0.0216795f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.985
cc_85 VPB N_A2_c_351_n 0.0043824f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.025
cc_86 VPB N_A2_c_353_n 0.00411957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A1_M1001_g 0.0185267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A1_M1019_g 0.0194101f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.985
cc_89 VPB A1 0.00197611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_489_n 0.0130612f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.985
cc_91 VPB N_VPWR_c_490_n 0.0358276f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.025
cc_92 VPB N_VPWR_c_491_n 3.12605e-19 $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.295
cc_93 VPB N_VPWR_c_492_n 0.00284364f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.025
cc_94 VPB N_VPWR_c_493_n 0.00613061f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_95 VPB N_VPWR_c_494_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.875 $Y2=0.56
cc_96 VPB N_VPWR_c_495_n 0.0145469f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.985
cc_97 VPB N_VPWR_c_496_n 0.0128277f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.16
cc_98 VPB N_VPWR_c_497_n 0.0123863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_498_n 0.0487238f $X=-0.19 $Y=1.305 $X2=2.525 $Y2=1.055
cc_100 VPB N_VPWR_c_499_n 0.0288121f $X=-0.19 $Y=1.305 $X2=3.045 $Y2=0.76
cc_101 VPB N_VPWR_c_488_n 0.046799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_501_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.525 $Y2=1.97
cc_103 VPB N_VPWR_c_502_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.38 $Y2=1.16
cc_104 VPB N_VPWR_c_503_n 0.00507259f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.16
cc_105 VPB N_VPWR_c_504_n 0.00436244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_X_c_601_n 0.0218185f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.985
cc_107 VPB N_X_c_604_n 0.00465216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_672_297#_c_649_n 0.00216365f $X=-0.19 $Y=1.305 $X2=0.585
+ $Y2=1.025
cc_109 VPB N_A_672_297#_c_650_n 0.0091049f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.295
cc_110 VPB N_A_672_297#_c_651_n 0.024997f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.985
cc_111 N_A_102_21#_M1023_g N_B1_M1006_g 0.0143247f $X=1.875 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_102_21#_c_130_n N_B1_M1006_g 0.00577255f $X=2.525 $Y=1.815 $X2=0
+ $Y2=0
cc_113 N_A_102_21#_c_134_p N_B1_M1006_g 0.00165796f $X=2.525 $Y=2.07 $X2=0 $Y2=0
cc_114 N_A_102_21#_c_121_n N_B1_c_237_n 0.00721839f $X=2.44 $Y=1.172 $X2=0 $Y2=0
cc_115 N_A_102_21#_c_122_n N_B1_c_237_n 0.00581121f $X=2.525 $Y=1.055 $X2=0
+ $Y2=0
cc_116 N_A_102_21#_c_130_n N_B1_c_237_n 0.00275579f $X=2.525 $Y=1.815 $X2=0
+ $Y2=0
cc_117 N_A_102_21#_c_138_p N_B1_c_237_n 0.0055208f $X=3.045 $Y=0.76 $X2=0 $Y2=0
cc_118 N_A_102_21#_c_139_p N_B1_c_237_n 0.00715393f $X=2.525 $Y=1.172 $X2=0
+ $Y2=0
cc_119 N_A_102_21#_c_121_n N_B1_c_238_n 0.0167493f $X=2.44 $Y=1.172 $X2=0 $Y2=0
cc_120 N_A_102_21#_c_125_n N_B1_c_238_n 0.0143247f $X=1.875 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_102_21#_c_130_n N_B1_M1018_g 0.0019517f $X=2.525 $Y=1.815 $X2=0 $Y2=0
cc_122 N_A_102_21#_c_131_n N_B1_M1018_g 0.0165301f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_123 N_A_102_21#_c_122_n N_B1_M1016_g 0.00486303f $X=2.525 $Y=1.055 $X2=0
+ $Y2=0
cc_124 N_A_102_21#_c_138_p N_B1_M1016_g 0.0133438f $X=3.045 $Y=0.76 $X2=0 $Y2=0
cc_125 N_A_102_21#_c_138_p N_B1_M1021_g 0.00341152f $X=3.045 $Y=0.76 $X2=0 $Y2=0
cc_126 N_A_102_21#_c_138_p B1 0.00326154f $X=3.045 $Y=0.76 $X2=0 $Y2=0
cc_127 N_A_102_21#_c_131_n B1 0.00628346f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_128 N_A_102_21#_c_130_n N_B1_c_247_n 0.0226733f $X=2.525 $Y=1.815 $X2=0 $Y2=0
cc_129 N_A_102_21#_c_138_p N_B1_c_247_n 0.0260126f $X=3.045 $Y=0.76 $X2=0 $Y2=0
cc_130 N_A_102_21#_c_131_n N_B1_c_247_n 0.0249454f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_131 N_A_102_21#_c_139_p N_B1_c_247_n 0.0189153f $X=2.525 $Y=1.172 $X2=0 $Y2=0
cc_132 N_A_102_21#_c_138_p N_B1_c_243_n 0.00202434f $X=3.045 $Y=0.76 $X2=0 $Y2=0
cc_133 N_A_102_21#_c_131_n N_B1_c_243_n 0.00183926f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_134 N_A_102_21#_c_131_n N_A3_M1000_g 0.0114038f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_135 N_A_102_21#_c_156_p N_A3_M1000_g 0.0136024f $X=3.925 $Y=2.02 $X2=0 $Y2=0
cc_136 N_A_102_21#_c_156_p N_A3_M1020_g 0.00676957f $X=3.925 $Y=2.02 $X2=0 $Y2=0
cc_137 N_A_102_21#_c_131_n N_VPWR_M1018_d 0.00558372f $X=3.76 $Y=1.97 $X2=0
+ $Y2=0
cc_138 N_A_102_21#_M1003_g N_VPWR_c_490_n 0.00345571f $X=0.585 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_102_21#_M1003_g N_VPWR_c_491_n 6.6524e-19 $X=0.585 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_102_21#_M1015_g N_VPWR_c_491_n 0.00997648f $X=1.005 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_102_21#_M1022_g N_VPWR_c_491_n 0.00990792f $X=1.455 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_102_21#_M1023_g N_VPWR_c_491_n 6.53233e-19 $X=1.875 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_102_21#_M1022_g N_VPWR_c_492_n 8.61039e-19 $X=1.455 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_102_21#_M1023_g N_VPWR_c_492_n 0.0152093f $X=1.875 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_102_21#_c_121_n N_VPWR_c_492_n 0.0278378f $X=2.44 $Y=1.172 $X2=0
+ $Y2=0
cc_146 N_A_102_21#_c_130_n N_VPWR_c_492_n 0.0277815f $X=2.525 $Y=1.815 $X2=0
+ $Y2=0
cc_147 N_A_102_21#_c_134_p N_VPWR_c_492_n 0.0267314f $X=2.525 $Y=2.07 $X2=0
+ $Y2=0
cc_148 N_A_102_21#_c_169_p N_VPWR_c_492_n 0.0151539f $X=2.525 $Y=1.97 $X2=0
+ $Y2=0
cc_149 N_A_102_21#_c_131_n N_VPWR_c_493_n 0.0208649f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_150 N_A_102_21#_c_156_p N_VPWR_c_493_n 0.00642921f $X=3.925 $Y=2.02 $X2=0
+ $Y2=0
cc_151 N_A_102_21#_M1003_g N_VPWR_c_495_n 0.00583607f $X=0.585 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_102_21#_M1015_g N_VPWR_c_495_n 0.00525069f $X=1.005 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_102_21#_M1022_g N_VPWR_c_496_n 0.00525069f $X=1.455 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_102_21#_M1023_g N_VPWR_c_496_n 0.0046653f $X=1.875 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_102_21#_c_134_p N_VPWR_c_497_n 0.0116048f $X=2.525 $Y=2.07 $X2=0
+ $Y2=0
cc_156 N_A_102_21#_c_131_n N_VPWR_c_497_n 0.0023707f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_157 N_A_102_21#_c_131_n N_VPWR_c_498_n 0.0107254f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_158 N_A_102_21#_c_156_p N_VPWR_c_498_n 0.0187605f $X=3.925 $Y=2.02 $X2=0
+ $Y2=0
cc_159 N_A_102_21#_M1006_s N_VPWR_c_488_n 0.00497872f $X=2.37 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_102_21#_M1000_d N_VPWR_c_488_n 0.00215201f $X=3.79 $Y=1.485 $X2=0
+ $Y2=0
cc_161 N_A_102_21#_M1003_g N_VPWR_c_488_n 0.0115212f $X=0.585 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_102_21#_M1015_g N_VPWR_c_488_n 0.00888907f $X=1.005 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_102_21#_M1022_g N_VPWR_c_488_n 0.00888907f $X=1.455 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_102_21#_M1023_g N_VPWR_c_488_n 0.00796766f $X=1.875 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_102_21#_c_134_p N_VPWR_c_488_n 0.00646998f $X=2.525 $Y=2.07 $X2=0
+ $Y2=0
cc_166 N_A_102_21#_c_131_n N_VPWR_c_488_n 0.0233834f $X=3.76 $Y=1.97 $X2=0 $Y2=0
cc_167 N_A_102_21#_c_156_p N_VPWR_c_488_n 0.0121784f $X=3.925 $Y=2.02 $X2=0
+ $Y2=0
cc_168 N_A_102_21#_M1002_g N_X_c_601_n 0.0158361f $X=0.585 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A_102_21#_M1003_g N_X_c_601_n 0.0239943f $X=0.585 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_102_21#_M1007_g N_X_c_601_n 0.00234513f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A_102_21#_M1015_g N_X_c_601_n 0.00299741f $X=1.005 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_102_21#_c_120_n N_X_c_601_n 0.0220343f $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_102_21#_c_121_n N_X_c_601_n 0.0196562f $X=2.44 $Y=1.172 $X2=0 $Y2=0
cc_174 N_A_102_21#_M1007_g N_X_c_611_n 0.0114177f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_102_21#_M1008_g N_X_c_611_n 0.011469f $X=1.455 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_102_21#_c_121_n N_X_c_611_n 0.041085f $X=2.44 $Y=1.172 $X2=0 $Y2=0
cc_177 N_A_102_21#_c_124_n N_X_c_611_n 0.00269497f $X=1.38 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_102_21#_M1015_g N_X_c_604_n 0.0155756f $X=1.005 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_102_21#_M1022_g N_X_c_604_n 0.0151865f $X=1.455 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_102_21#_M1023_g N_X_c_604_n 7.53908e-19 $X=1.875 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_102_21#_c_121_n N_X_c_604_n 0.0630562f $X=2.44 $Y=1.172 $X2=0 $Y2=0
cc_182 N_A_102_21#_c_124_n N_X_c_604_n 0.0026088f $X=1.38 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_102_21#_c_125_n N_X_c_604_n 0.00202726f $X=1.875 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_102_21#_c_121_n N_X_c_602_n 0.0140803f $X=2.44 $Y=1.172 $X2=0 $Y2=0
cc_185 N_A_102_21#_c_125_n N_X_c_602_n 0.00208088f $X=1.875 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_102_21#_c_131_n N_A_672_297#_M1000_s 0.00746329f $X=3.76 $Y=1.97
+ $X2=-0.19 $Y2=-0.24
cc_187 N_A_102_21#_M1000_d N_A_672_297#_c_649_n 0.00312957f $X=3.79 $Y=1.485
+ $X2=0 $Y2=0
cc_188 N_A_102_21#_c_131_n N_A_672_297#_c_649_n 0.0276147f $X=3.76 $Y=1.97 $X2=0
+ $Y2=0
cc_189 N_A_102_21#_c_156_p N_A_672_297#_c_649_n 0.0169935f $X=3.925 $Y=2.02
+ $X2=0 $Y2=0
cc_190 N_A_102_21#_c_156_p N_A_672_297#_c_656_n 0.00749737f $X=3.925 $Y=2.02
+ $X2=0 $Y2=0
cc_191 N_A_102_21#_c_156_p N_A_672_297#_c_657_n 0.0171501f $X=3.925 $Y=2.02
+ $X2=0 $Y2=0
cc_192 N_A_102_21#_M1002_g N_VGND_c_744_n 0.00345571f $X=0.585 $Y=0.56 $X2=0
+ $Y2=0
cc_193 N_A_102_21#_M1002_g N_VGND_c_745_n 5.52077e-19 $X=0.585 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_A_102_21#_M1007_g N_VGND_c_745_n 0.00621536f $X=1.005 $Y=0.56 $X2=0
+ $Y2=0
cc_195 N_A_102_21#_M1008_g N_VGND_c_745_n 0.00618135f $X=1.455 $Y=0.56 $X2=0
+ $Y2=0
cc_196 N_A_102_21#_M1010_g N_VGND_c_745_n 5.46103e-19 $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_197 N_A_102_21#_M1008_g N_VGND_c_746_n 5.93577e-19 $X=1.455 $Y=0.56 $X2=0
+ $Y2=0
cc_198 N_A_102_21#_M1010_g N_VGND_c_746_n 0.0108823f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_199 N_A_102_21#_c_121_n N_VGND_c_746_n 0.023739f $X=2.44 $Y=1.172 $X2=0 $Y2=0
cc_200 N_A_102_21#_c_123_n N_VGND_c_746_n 0.0203734f $X=2.61 $Y=0.76 $X2=0 $Y2=0
cc_201 N_A_102_21#_M1002_g N_VGND_c_752_n 0.00435566f $X=0.585 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_A_102_21#_M1007_g N_VGND_c_752_n 0.00384491f $X=1.005 $Y=0.56 $X2=0
+ $Y2=0
cc_203 N_A_102_21#_M1008_g N_VGND_c_753_n 0.00384491f $X=1.455 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_102_21#_M1010_g N_VGND_c_753_n 0.00525069f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_205 N_A_102_21#_M1016_d N_VGND_c_757_n 0.00216833f $X=2.91 $Y=0.235 $X2=0
+ $Y2=0
cc_206 N_A_102_21#_M1002_g N_VGND_c_757_n 0.00681221f $X=0.585 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_102_21#_M1007_g N_VGND_c_757_n 0.004459f $X=1.005 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A_102_21#_M1008_g N_VGND_c_757_n 0.004459f $X=1.455 $Y=0.56 $X2=0 $Y2=0
cc_209 N_A_102_21#_M1010_g N_VGND_c_757_n 0.00888907f $X=1.875 $Y=0.56 $X2=0
+ $Y2=0
cc_210 N_A_102_21#_c_123_n N_A_496_47#_M1016_s 0.00254953f $X=2.61 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_211 N_A_102_21#_c_138_p N_A_496_47#_M1016_s 0.00205175f $X=3.045 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_212 N_A_102_21#_M1016_d N_A_496_47#_c_854_n 0.00305599f $X=2.91 $Y=0.235
+ $X2=0 $Y2=0
cc_213 N_A_102_21#_c_123_n N_A_496_47#_c_854_n 0.0133793f $X=2.61 $Y=0.76 $X2=0
+ $Y2=0
cc_214 N_A_102_21#_c_138_p N_A_496_47#_c_854_n 0.0299173f $X=3.045 $Y=0.76 $X2=0
+ $Y2=0
cc_215 N_B1_M1021_g N_A3_M1012_g 0.0162425f $X=3.255 $Y=0.56 $X2=0 $Y2=0
cc_216 N_B1_c_247_n N_A3_M1000_g 0.00414433f $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_217 B1 A3 0.0222004f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_218 N_B1_c_247_n A3 2.07261e-19 $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_219 B1 N_A3_c_306_n 0.00366966f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_220 N_B1_c_243_n N_A3_c_306_n 0.0162425f $X=3.255 $Y=1.16 $X2=0 $Y2=0
cc_221 N_B1_c_247_n N_VPWR_M1018_d 0.00366185f $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B1_M1006_g N_VPWR_c_492_n 0.01572f $X=2.295 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B1_M1018_g N_VPWR_c_492_n 6.08646e-19 $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_224 N_B1_M1006_g N_VPWR_c_493_n 5.48834e-19 $X=2.295 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B1_M1018_g N_VPWR_c_493_n 0.00795974f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B1_M1006_g N_VPWR_c_497_n 0.0046653f $X=2.295 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B1_M1018_g N_VPWR_c_497_n 0.00341112f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_228 N_B1_M1006_g N_VPWR_c_488_n 0.00802193f $X=2.295 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B1_M1018_g N_VPWR_c_488_n 0.00407063f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_230 N_B1_M1018_g N_A_672_297#_c_649_n 6.42245e-19 $X=2.735 $Y=1.985 $X2=0
+ $Y2=0
cc_231 B1 N_A_672_297#_c_649_n 0.0193699f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_232 N_B1_c_247_n N_A_672_297#_c_649_n 0.0146271f $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_233 N_B1_c_238_n N_VGND_c_746_n 8.18625e-19 $X=2.37 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B1_M1016_g N_VGND_c_746_n 0.00656715f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_235 N_B1_M1021_g N_VGND_c_747_n 0.00119163f $X=3.255 $Y=0.56 $X2=0 $Y2=0
cc_236 N_B1_M1016_g N_VGND_c_754_n 0.00357877f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B1_M1021_g N_VGND_c_754_n 0.00357877f $X=3.255 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B1_M1016_g N_VGND_c_757_n 0.00655123f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B1_M1021_g N_VGND_c_757_n 0.00539139f $X=3.255 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B1_c_237_n N_A_496_47#_c_854_n 6.55955e-19 $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_241 N_B1_M1016_g N_A_496_47#_c_854_n 0.00861238f $X=2.835 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B1_M1021_g N_A_496_47#_c_854_n 0.0113884f $X=3.255 $Y=0.56 $X2=0 $Y2=0
cc_243 B1 N_A_496_47#_c_854_n 0.00394331f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_244 B1 N_A_496_47#_c_868_n 3.59099e-19 $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_245 B1 N_A_496_47#_c_855_n 0.0159508f $X=3.345 $Y=1.105 $X2=0 $Y2=0
cc_246 N_A3_M1014_g N_A2_c_347_n 0.0236295f $X=4.135 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_247 N_A3_M1020_g N_A2_M1011_g 0.0265534f $X=4.135 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A3_M1014_g N_A2_c_351_n 0.0214718f $X=4.135 $Y=0.56 $X2=0 $Y2=0
cc_249 A3 N_A2_c_351_n 2.10525e-19 $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_250 A3 N_A2_c_353_n 0.0255884f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_251 N_A3_c_306_n N_A2_c_353_n 0.00245355f $X=4.135 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A3_M1000_g N_VPWR_c_493_n 0.00599992f $X=3.715 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A3_M1000_g N_VPWR_c_498_n 0.00414887f $X=3.715 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A3_M1020_g N_VPWR_c_498_n 0.00541359f $X=4.135 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A3_M1000_g N_VPWR_c_488_n 0.00711255f $X=3.715 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A3_M1020_g N_VPWR_c_488_n 0.00972842f $X=4.135 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A3_M1000_g N_A_672_297#_c_649_n 0.0102082f $X=3.715 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_A3_M1020_g N_A_672_297#_c_649_n 0.0145621f $X=4.135 $Y=1.985 $X2=0
+ $Y2=0
cc_259 A3 N_A_672_297#_c_649_n 0.0209935f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_260 N_A3_c_306_n N_A_672_297#_c_649_n 5.3419e-19 $X=4.135 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A3_M1020_g N_A_672_297#_c_657_n 7.62531e-19 $X=4.135 $Y=1.985 $X2=0
+ $Y2=0
cc_262 N_A3_M1012_g N_VGND_c_747_n 0.00776184f $X=3.715 $Y=0.56 $X2=0 $Y2=0
cc_263 N_A3_M1014_g N_VGND_c_747_n 0.00645899f $X=4.135 $Y=0.56 $X2=0 $Y2=0
cc_264 N_A3_M1014_g N_VGND_c_748_n 5.4242e-19 $X=4.135 $Y=0.56 $X2=0 $Y2=0
cc_265 N_A3_M1012_g N_VGND_c_754_n 0.00339367f $X=3.715 $Y=0.56 $X2=0 $Y2=0
cc_266 N_A3_M1014_g N_VGND_c_755_n 0.00339367f $X=4.135 $Y=0.56 $X2=0 $Y2=0
cc_267 N_A3_M1012_g N_VGND_c_757_n 0.00411438f $X=3.715 $Y=0.56 $X2=0 $Y2=0
cc_268 N_A3_M1014_g N_VGND_c_757_n 0.00401529f $X=4.135 $Y=0.56 $X2=0 $Y2=0
cc_269 N_A3_M1012_g N_A_496_47#_c_854_n 0.00181821f $X=3.715 $Y=0.56 $X2=0 $Y2=0
cc_270 N_A3_M1012_g N_A_496_47#_c_868_n 0.0148169f $X=3.715 $Y=0.56 $X2=0 $Y2=0
cc_271 N_A3_M1014_g N_A_496_47#_c_868_n 0.0147173f $X=4.135 $Y=0.56 $X2=0 $Y2=0
cc_272 A3 N_A_496_47#_c_868_n 0.0203538f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_273 N_A3_c_306_n N_A_496_47#_c_868_n 0.00202434f $X=4.135 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A2_c_347_n N_A1_M1004_g 0.027158f $X=4.555 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_c_351_n N_A1_M1004_g 0.0218346f $X=4.555 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A2_M1011_g N_A1_M1001_g 0.0397253f $X=4.555 $Y=1.985 $X2=0 $Y2=0
cc_277 A2 N_A1_M1001_g 0.00886444f $X=4.745 $Y=1.445 $X2=0 $Y2=0
cc_278 N_A2_c_354_n N_A1_M1001_g 0.00148614f $X=4.825 $Y=1.36 $X2=0 $Y2=0
cc_279 N_A2_c_372_p N_A1_M1001_g 0.00650402f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_280 N_A2_M1013_g N_A1_M1005_g 0.0281263f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A2_M1017_g N_A1_M1019_g 0.0281263f $X=5.815 $Y=1.985 $X2=0 $Y2=0
cc_282 A2 N_A1_M1019_g 5.76991e-19 $X=4.745 $Y=1.445 $X2=0 $Y2=0
cc_283 N_A2_c_372_p N_A1_M1019_g 0.0102285f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_284 A2 A1 0.025707f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_285 N_A2_c_352_n A1 3.22602e-19 $X=5.905 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A2_c_354_n A1 0.0246398f $X=4.825 $Y=1.36 $X2=0 $Y2=0
cc_287 N_A2_c_372_p A1 0.0224817f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_288 A2 N_A1_c_440_n 0.00441754f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_289 N_A2_c_352_n N_A1_c_440_n 0.0281263f $X=5.905 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A2_c_354_n N_A1_c_440_n 0.00825005f $X=4.825 $Y=1.36 $X2=0 $Y2=0
cc_291 N_A2_c_372_p N_A1_c_440_n 5.28255e-19 $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_292 N_A2_c_372_p N_VPWR_M1001_d 0.00342618f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_293 N_A2_M1011_g N_VPWR_c_494_n 0.00122089f $X=4.555 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A2_M1017_g N_VPWR_c_494_n 0.00122089f $X=5.815 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A2_M1011_g N_VPWR_c_498_n 0.00541359f $X=4.555 $Y=1.985 $X2=0 $Y2=0
cc_296 N_A2_M1017_g N_VPWR_c_499_n 0.00585385f $X=5.815 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A2_M1011_g N_VPWR_c_488_n 0.00534331f $X=4.555 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A2_M1017_g N_VPWR_c_488_n 0.00657985f $X=5.815 $Y=1.985 $X2=0 $Y2=0
cc_299 A2 N_A_672_297#_M1017_s 0.00312529f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_300 N_A2_M1011_g N_A_672_297#_c_649_n 0.00323803f $X=4.555 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A2_c_351_n N_A_672_297#_c_649_n 2.70427e-19 $X=4.555 $Y=1.16 $X2=0
+ $Y2=0
cc_302 N_A2_c_353_n N_A_672_297#_c_649_n 0.0182652f $X=4.68 $Y=1.207 $X2=0 $Y2=0
cc_303 N_A2_M1011_g N_A_672_297#_c_670_n 0.00574649f $X=4.555 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_A2_M1017_g N_A_672_297#_c_670_n 0.00318286f $X=5.815 $Y=1.985 $X2=0
+ $Y2=0
cc_305 A2 N_A_672_297#_c_670_n 8.13734e-19 $X=4.745 $Y=1.445 $X2=0 $Y2=0
cc_306 A2 N_A_672_297#_c_670_n 0.00652059f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_307 N_A2_c_372_p N_A_672_297#_c_670_n 8.94099e-19 $X=5.64 $Y=1.377 $X2=0
+ $Y2=0
cc_308 N_A2_M1011_g N_A_672_297#_c_656_n 0.00103327f $X=4.555 $Y=1.985 $X2=0
+ $Y2=0
cc_309 A2 N_A_672_297#_c_650_n 0.00149821f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_310 N_A2_M1017_g N_A_672_297#_c_651_n 0.0049333f $X=5.815 $Y=1.985 $X2=0
+ $Y2=0
cc_311 A2 N_A_672_297#_c_651_n 0.0348537f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_312 N_A2_c_352_n N_A_672_297#_c_651_n 5.35519e-19 $X=5.905 $Y=1.16 $X2=0
+ $Y2=0
cc_313 N_A2_M1011_g N_A_672_297#_c_657_n 0.00974268f $X=4.555 $Y=1.985 $X2=0
+ $Y2=0
cc_314 A2 N_A_926_297#_M1011_d 0.00193824f $X=4.745 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_315 A2 N_A_926_297#_M1019_s 0.0010921f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_316 N_A2_c_372_p N_A_926_297#_M1019_s 0.00347109f $X=5.64 $Y=1.377 $X2=0
+ $Y2=0
cc_317 A2 N_A_926_297#_c_712_n 0.00508073f $X=4.745 $Y=1.445 $X2=0 $Y2=0
cc_318 N_A2_c_372_p N_A_926_297#_c_712_n 0.0259823f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_319 N_A2_M1011_g N_A_926_297#_c_714_n 0.00110724f $X=4.555 $Y=1.985 $X2=0
+ $Y2=0
cc_320 A2 N_A_926_297#_c_714_n 0.0132767f $X=4.745 $Y=1.445 $X2=0 $Y2=0
cc_321 N_A2_M1017_g N_A_926_297#_c_716_n 0.00118947f $X=5.815 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A2_c_372_p N_A_926_297#_c_716_n 0.0123458f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_323 N_A2_c_347_n N_VGND_c_747_n 5.4242e-19 $X=4.555 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A2_c_347_n N_VGND_c_748_n 0.00642509f $X=4.555 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A2_M1013_g N_VGND_c_749_n 0.00811705f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_326 N_A2_c_347_n N_VGND_c_755_n 0.00339367f $X=4.555 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A2_M1013_g N_VGND_c_756_n 0.00339367f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_328 N_A2_c_347_n N_VGND_c_757_n 0.00401529f $X=4.555 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A2_M1013_g N_VGND_c_757_n 0.00510156f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_330 N_A2_c_347_n N_A_496_47#_c_875_n 0.0129876f $X=4.555 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A2_c_351_n N_A_496_47#_c_875_n 0.00130338f $X=4.555 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A2_c_353_n N_A_496_47#_c_875_n 0.0146249f $X=4.68 $Y=1.207 $X2=0 $Y2=0
cc_333 N_A2_c_354_n N_A_496_47#_c_875_n 0.0216203f $X=4.825 $Y=1.36 $X2=0 $Y2=0
cc_334 N_A2_c_372_p N_A_496_47#_c_875_n 0.00182971f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_335 N_A2_M1013_g N_A_496_47#_c_880_n 0.0134672f $X=5.815 $Y=0.56 $X2=0 $Y2=0
cc_336 A2 N_A_496_47#_c_880_n 0.0199693f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_337 N_A2_c_372_p N_A_496_47#_c_880_n 0.00310277f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_338 N_A2_c_351_n N_A_496_47#_c_856_n 2.26132e-19 $X=4.555 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A2_c_353_n N_A_496_47#_c_856_n 0.0136988f $X=4.68 $Y=1.207 $X2=0 $Y2=0
cc_340 N_A2_c_372_p N_A_496_47#_c_857_n 0.00100641f $X=5.64 $Y=1.377 $X2=0 $Y2=0
cc_341 A2 N_A_496_47#_c_858_n 0.0369429f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_342 N_A2_c_352_n N_A_496_47#_c_858_n 0.00296376f $X=5.905 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A1_M1001_g N_VPWR_c_494_n 0.00768198f $X=4.975 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A1_M1019_g N_VPWR_c_494_n 0.00767608f $X=5.395 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A1_M1001_g N_VPWR_c_498_n 0.00341112f $X=4.975 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A1_M1019_g N_VPWR_c_499_n 0.00341112f $X=5.395 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A1_M1001_g N_VPWR_c_488_n 0.00332143f $X=4.975 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A1_M1019_g N_VPWR_c_488_n 0.00332143f $X=5.395 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A1_M1001_g N_A_672_297#_c_670_n 0.00252193f $X=4.975 $Y=1.985 $X2=0
+ $Y2=0
cc_350 N_A1_M1019_g N_A_672_297#_c_670_n 0.00252193f $X=5.395 $Y=1.985 $X2=0
+ $Y2=0
cc_351 N_A1_M1001_g N_A_672_297#_c_657_n 7.76806e-19 $X=4.975 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A1_M1001_g N_A_926_297#_c_712_n 0.00997598f $X=4.975 $Y=1.985 $X2=0
+ $Y2=0
cc_353 N_A1_M1019_g N_A_926_297#_c_712_n 0.00997884f $X=5.395 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A1_M1001_g N_A_926_297#_c_714_n 0.00136719f $X=4.975 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A1_M1019_g N_A_926_297#_c_716_n 0.00137591f $X=5.395 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A1_M1004_g N_VGND_c_748_n 0.00642509f $X=4.975 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A1_M1005_g N_VGND_c_748_n 5.4242e-19 $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A1_M1004_g N_VGND_c_749_n 5.4242e-19 $X=4.975 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A1_M1005_g N_VGND_c_749_n 0.00642509f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A1_M1004_g N_VGND_c_750_n 0.00339367f $X=4.975 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A1_M1005_g N_VGND_c_750_n 0.00339367f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A1_M1004_g N_VGND_c_757_n 0.00398704f $X=4.975 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A1_M1005_g N_VGND_c_757_n 0.00398704f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A1_M1004_g N_A_496_47#_c_875_n 0.0142125f $X=4.975 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A1_M1005_g N_A_496_47#_c_880_n 0.0130013f $X=5.395 $Y=0.56 $X2=0 $Y2=0
cc_366 A1 N_A_496_47#_c_880_n 0.0128033f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_367 A1 N_A_496_47#_c_857_n 0.0102706f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_368 N_A1_c_440_n N_A_496_47#_c_857_n 0.00208611f $X=5.395 $Y=1.16 $X2=0 $Y2=0
cc_369 N_VPWR_c_488_n N_X_M1003_d 0.00414686f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_370 N_VPWR_c_488_n N_X_M1022_d 0.00518834f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_371 N_VPWR_M1003_s N_X_c_601_n 0.00304349f $X=0.25 $Y=1.485 $X2=0 $Y2=0
cc_372 N_VPWR_c_490_n N_X_c_601_n 0.0336692f $X=0.375 $Y=2 $X2=0 $Y2=0
cc_373 N_VPWR_c_495_n N_X_c_627_n 0.0129925f $X=1.065 $Y=2.72 $X2=0 $Y2=0
cc_374 N_VPWR_c_488_n N_X_c_627_n 0.008203f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_M1015_s N_X_c_604_n 0.00198867f $X=1.08 $Y=1.485 $X2=0 $Y2=0
cc_376 N_VPWR_c_491_n N_X_c_604_n 0.0174023f $X=1.23 $Y=2.02 $X2=0 $Y2=0
cc_377 N_VPWR_c_492_n N_X_c_604_n 0.00884749f $X=2.085 $Y=1.68 $X2=0 $Y2=0
cc_378 N_VPWR_c_496_n N_X_c_632_n 0.011928f $X=1.92 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_c_488_n N_X_c_632_n 0.00704765f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_c_488_n N_A_672_297#_M1000_s 0.00334747f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_381 N_VPWR_c_488_n N_A_672_297#_M1020_s 0.00186159f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_488_n N_A_672_297#_M1017_s 0.00116343f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_M1001_d N_A_672_297#_c_670_n 0.00196478f $X=5.05 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_494_n N_A_672_297#_c_670_n 0.00901225f $X=5.185 $Y=2.36 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_498_n N_A_672_297#_c_670_n 0.00142477f $X=5.02 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_499_n N_A_672_297#_c_670_n 0.0015755f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_488_n N_A_672_297#_c_670_n 0.131383f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_c_498_n N_A_672_297#_c_656_n 3.88714e-19 $X=5.02 $Y=2.72 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_488_n N_A_672_297#_c_656_n 0.028441f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_488_n N_A_672_297#_c_650_n 0.0284534f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_499_n N_A_672_297#_c_651_n 0.0305087f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_488_n N_A_672_297#_c_651_n 0.00464908f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_498_n N_A_672_297#_c_657_n 0.0151826f $X=5.02 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_488_n N_A_672_297#_c_657_n 0.00236942f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_488_n N_A_926_297#_M1011_d 0.00152827f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_396 N_VPWR_c_488_n N_A_926_297#_M1019_s 0.0013901f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_M1001_d N_A_926_297#_c_712_n 0.00306115f $X=5.05 $Y=1.485 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_494_n N_A_926_297#_c_712_n 0.0157356f $X=5.185 $Y=2.36 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_498_n N_A_926_297#_c_712_n 0.0021583f $X=5.02 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_499_n N_A_926_297#_c_712_n 0.0021583f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_494_n N_A_926_297#_c_714_n 0.00883474f $X=5.185 $Y=2.36 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_498_n N_A_926_297#_c_714_n 0.0112892f $X=5.02 $Y=2.72 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_488_n N_A_926_297#_c_714_n 0.00180269f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_494_n N_A_926_297#_c_716_n 0.00895573f $X=5.185 $Y=2.36 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_499_n N_A_926_297#_c_716_n 0.0123537f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_488_n N_A_926_297#_c_716_n 0.0021246f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_X_c_601_n N_VGND_M1002_d 0.00294167f $X=0.787 $Y=1.665 $X2=-0.19
+ $Y2=-0.24
cc_408 N_X_c_611_n N_VGND_M1007_d 0.00364094f $X=1.565 $Y=0.77 $X2=0 $Y2=0
cc_409 N_X_c_601_n N_VGND_c_744_n 0.0322091f $X=0.787 $Y=1.665 $X2=0 $Y2=0
cc_410 N_X_c_611_n N_VGND_c_745_n 0.0165345f $X=1.565 $Y=0.77 $X2=0 $Y2=0
cc_411 N_X_c_601_n N_VGND_c_752_n 0.00240483f $X=0.787 $Y=1.665 $X2=0 $Y2=0
cc_412 N_X_c_611_n N_VGND_c_752_n 0.0024595f $X=1.565 $Y=0.77 $X2=0 $Y2=0
cc_413 N_X_c_640_p N_VGND_c_752_n 0.0129383f $X=0.795 $Y=0.72 $X2=0 $Y2=0
cc_414 N_X_c_611_n N_VGND_c_753_n 0.0024595f $X=1.565 $Y=0.77 $X2=0 $Y2=0
cc_415 N_X_c_602_n N_VGND_c_753_n 0.012399f $X=1.665 $Y=0.72 $X2=0 $Y2=0
cc_416 N_X_M1002_s N_VGND_c_757_n 0.002386f $X=0.66 $Y=0.235 $X2=0 $Y2=0
cc_417 N_X_M1008_s N_VGND_c_757_n 0.00354764f $X=1.53 $Y=0.235 $X2=0 $Y2=0
cc_418 N_X_c_601_n N_VGND_c_757_n 0.00590041f $X=0.787 $Y=1.665 $X2=0 $Y2=0
cc_419 N_X_c_611_n N_VGND_c_757_n 0.00971057f $X=1.565 $Y=0.77 $X2=0 $Y2=0
cc_420 N_X_c_602_n N_VGND_c_757_n 0.00761007f $X=1.665 $Y=0.72 $X2=0 $Y2=0
cc_421 N_X_c_640_p N_VGND_c_757_n 0.00819075f $X=0.795 $Y=0.72 $X2=0 $Y2=0
cc_422 N_A_672_297#_c_670_n N_A_926_297#_M1011_d 0.00273286f $X=6.065 $Y=2.21
+ $X2=-0.19 $Y2=1.305
cc_423 N_A_672_297#_c_670_n N_A_926_297#_M1019_s 9.33948e-19 $X=6.065 $Y=2.21
+ $X2=0 $Y2=0
cc_424 N_A_672_297#_c_670_n N_A_926_297#_c_712_n 0.0195872f $X=6.065 $Y=2.21
+ $X2=0 $Y2=0
cc_425 N_A_672_297#_c_670_n N_A_926_297#_c_714_n 0.0116591f $X=6.065 $Y=2.21
+ $X2=0 $Y2=0
cc_426 N_A_672_297#_c_656_n N_A_926_297#_c_714_n 0.00224031f $X=4.515 $Y=2.21
+ $X2=0 $Y2=0
cc_427 N_A_672_297#_c_657_n N_A_926_297#_c_714_n 0.015889f $X=4.345 $Y=1.815
+ $X2=0 $Y2=0
cc_428 N_A_672_297#_c_670_n N_A_926_297#_c_716_n 0.01296f $X=6.065 $Y=2.21 $X2=0
+ $Y2=0
cc_429 N_A_672_297#_c_650_n N_A_926_297#_c_716_n 4.54416e-19 $X=6.21 $Y=2.21
+ $X2=0 $Y2=0
cc_430 N_A_672_297#_c_651_n N_A_926_297#_c_716_n 0.0183248f $X=6.21 $Y=2.21
+ $X2=0 $Y2=0
cc_431 N_A_672_297#_c_649_n N_A_496_47#_c_868_n 0.00577725f $X=4.26 $Y=1.615
+ $X2=0 $Y2=0
cc_432 N_VGND_c_757_n N_A_496_47#_M1016_s 0.00225742f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_433 N_VGND_c_757_n N_A_496_47#_M1021_s 0.00274469f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_757_n N_A_496_47#_M1014_d 0.00251683f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_757_n N_A_496_47#_M1004_d 0.00251683f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_757_n N_A_496_47#_M1013_s 0.0022756f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_746_n N_A_496_47#_c_854_n 0.0169507f $X=2.085 $Y=0.38 $X2=0
+ $Y2=0
cc_438 N_VGND_c_747_n N_A_496_47#_c_854_n 0.0143962f $X=3.925 $Y=0.36 $X2=0
+ $Y2=0
cc_439 N_VGND_c_754_n N_A_496_47#_c_854_n 0.0665114f $X=3.76 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_757_n N_A_496_47#_c_854_n 0.041032f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_441 N_VGND_M1012_s N_A_496_47#_c_868_n 0.0031524f $X=3.79 $Y=0.235 $X2=0
+ $Y2=0
cc_442 N_VGND_c_747_n N_A_496_47#_c_868_n 0.0147951f $X=3.925 $Y=0.36 $X2=0
+ $Y2=0
cc_443 N_VGND_c_754_n N_A_496_47#_c_868_n 0.00277814f $X=3.76 $Y=0 $X2=0 $Y2=0
cc_444 N_VGND_c_755_n N_A_496_47#_c_868_n 0.00248431f $X=4.6 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_757_n N_A_496_47#_c_868_n 0.0107423f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_755_n N_A_496_47#_c_908_n 0.0113346f $X=4.6 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_c_757_n N_A_496_47#_c_908_n 0.00645703f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_448 N_VGND_M1009_d N_A_496_47#_c_875_n 0.00333492f $X=4.63 $Y=0.235 $X2=0
+ $Y2=0
cc_449 N_VGND_c_748_n N_A_496_47#_c_875_n 0.0147951f $X=4.765 $Y=0.36 $X2=0
+ $Y2=0
cc_450 N_VGND_c_750_n N_A_496_47#_c_875_n 0.00248431f $X=5.44 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_755_n N_A_496_47#_c_875_n 0.00248431f $X=4.6 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_757_n N_A_496_47#_c_875_n 0.0101669f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_c_750_n N_A_496_47#_c_915_n 0.0113346f $X=5.44 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_757_n N_A_496_47#_c_915_n 0.00645703f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_455 N_VGND_M1005_s N_A_496_47#_c_880_n 0.00452276f $X=5.47 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_VGND_c_749_n N_A_496_47#_c_880_n 0.0147951f $X=5.605 $Y=0.36 $X2=0
+ $Y2=0
cc_457 N_VGND_c_750_n N_A_496_47#_c_880_n 0.00248431f $X=5.44 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_756_n N_A_496_47#_c_880_n 0.00248431f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_757_n N_A_496_47#_c_880_n 0.0101669f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_460 N_VGND_c_756_n N_A_496_47#_c_858_n 0.0289498f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_757_n N_A_496_47#_c_858_n 0.0158735f $X=6.21 $Y=0 $X2=0 $Y2=0

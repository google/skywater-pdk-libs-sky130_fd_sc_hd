* File: sky130_fd_sc_hd__o21ba_1.pxi.spice
* Created: Thu Aug 27 14:35:59 2020
* 
x_PM_SKY130_FD_SC_HD__O21BA_1%A_79_199# N_A_79_199#_M1009_s N_A_79_199#_M1004_d
+ N_A_79_199#_M1006_g N_A_79_199#_M1005_g N_A_79_199#_c_72_n N_A_79_199#_c_119_p
+ N_A_79_199#_c_67_n N_A_79_199#_c_68_n N_A_79_199#_c_69_n N_A_79_199#_c_76_n
+ N_A_79_199#_c_102_p N_A_79_199#_c_77_n N_A_79_199#_c_70_n
+ PM_SKY130_FD_SC_HD__O21BA_1%A_79_199#
x_PM_SKY130_FD_SC_HD__O21BA_1%B1_N N_B1_N_M1002_g N_B1_N_M1003_g B1_N
+ N_B1_N_c_148_n N_B1_N_c_149_n PM_SKY130_FD_SC_HD__O21BA_1%B1_N
x_PM_SKY130_FD_SC_HD__O21BA_1%A_222_93# N_A_222_93#_M1002_d N_A_222_93#_M1003_d
+ N_A_222_93#_c_181_n N_A_222_93#_M1009_g N_A_222_93#_M1004_g
+ N_A_222_93#_c_182_n N_A_222_93#_c_183_n N_A_222_93#_c_190_n
+ N_A_222_93#_c_184_n N_A_222_93#_c_185_n N_A_222_93#_c_186_n
+ PM_SKY130_FD_SC_HD__O21BA_1%A_222_93#
x_PM_SKY130_FD_SC_HD__O21BA_1%A2 N_A2_M1000_g N_A2_M1001_g A2 N_A2_c_236_n
+ N_A2_c_237_n PM_SKY130_FD_SC_HD__O21BA_1%A2
x_PM_SKY130_FD_SC_HD__O21BA_1%A1 N_A1_M1007_g N_A1_M1008_g A1 N_A1_c_270_n
+ N_A1_c_271_n PM_SKY130_FD_SC_HD__O21BA_1%A1
x_PM_SKY130_FD_SC_HD__O21BA_1%X N_X_M1005_s N_X_M1006_s N_X_c_295_n N_X_c_297_n
+ N_X_c_296_n X PM_SKY130_FD_SC_HD__O21BA_1%X
x_PM_SKY130_FD_SC_HD__O21BA_1%VPWR N_VPWR_M1006_d N_VPWR_M1004_s N_VPWR_M1007_d
+ N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n
+ VPWR N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_314_n
+ N_VPWR_c_324_n N_VPWR_c_325_n PM_SKY130_FD_SC_HD__O21BA_1%VPWR
x_PM_SKY130_FD_SC_HD__O21BA_1%VGND N_VGND_M1005_d N_VGND_M1000_d N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n
+ VGND N_VGND_c_372_n N_VGND_c_373_n PM_SKY130_FD_SC_HD__O21BA_1%VGND
x_PM_SKY130_FD_SC_HD__O21BA_1%A_448_47# N_A_448_47#_M1009_d N_A_448_47#_M1008_d
+ N_A_448_47#_c_416_n N_A_448_47#_c_411_n N_A_448_47#_c_412_n
+ N_A_448_47#_c_413_n PM_SKY130_FD_SC_HD__O21BA_1%A_448_47#
cc_1 VNB N_A_79_199#_c_67_n 0.00194759f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=0.57
cc_2 VNB N_A_79_199#_c_68_n 0.00672603f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_3 VNB N_A_79_199#_c_69_n 0.02763f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_4 VNB N_A_79_199#_c_70_n 0.0223891f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=0.995
cc_5 VNB B1_N 0.00557272f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_6 VNB N_B1_N_c_148_n 0.0232981f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_7 VNB N_B1_N_c_149_n 0.0215776f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_8 VNB N_A_222_93#_c_181_n 0.0199431f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_9 VNB N_A_222_93#_c_182_n 0.0474247f $X=-0.19 $Y=-0.24 $X2=0.727 $Y2=1.325
cc_10 VNB N_A_222_93#_c_183_n 0.00879111f $X=-0.19 $Y=-0.24 $X2=0.727 $Y2=1.865
cc_11 VNB N_A_222_93#_c_184_n 0.0117518f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=0.57
cc_12 VNB N_A_222_93#_c_185_n 0.00315751f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_13 VNB N_A_222_93#_c_186_n 0.0021006f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.325
cc_14 VNB A2 0.00857923f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_15 VNB N_A2_c_236_n 0.0193019f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_16 VNB N_A2_c_237_n 0.0167622f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_17 VNB A1 0.025059f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_18 VNB N_A1_c_270_n 0.0326309f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_19 VNB N_A1_c_271_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_20 VNB N_X_c_295_n 0.0172248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_296_n 0.024255f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.95
cc_22 VNB N_VPWR_c_314_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_366_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_24 VNB N_VGND_c_367_n 0.00462888f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_25 VNB N_VGND_c_368_n 0.022439f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.95
cc_26 VNB N_VGND_c_369_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.95
cc_27 VNB N_VGND_c_370_n 0.0519877f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=0.57
cc_28 VNB N_VGND_c_371_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=0.57
cc_29 VNB N_VGND_c_372_n 0.0220671f $X=-0.19 $Y=-0.24 $X2=2.435 $Y2=1.96
cc_30 VNB N_VGND_c_373_n 0.22571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_448_47#_c_411_n 0.0156132f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_32 VNB N_A_448_47#_c_412_n 0.00256586f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.56
cc_33 VNB N_A_448_47#_c_413_n 0.0181301f $X=-0.19 $Y=-0.24 $X2=0.727 $Y2=1.865
cc_34 VPB N_A_79_199#_M1006_g 0.0254413f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_35 VPB N_A_79_199#_c_72_n 0.00256842f $X=-0.19 $Y=1.305 $X2=0.727 $Y2=1.865
cc_36 VPB N_A_79_199#_c_67_n 0.00285312f $X=-0.19 $Y=1.305 $X2=1.955 $Y2=0.57
cc_37 VPB N_A_79_199#_c_68_n 0.00198329f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_38 VPB N_A_79_199#_c_69_n 0.00665208f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_39 VPB N_A_79_199#_c_76_n 0.0162918f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.745
cc_40 VPB N_A_79_199#_c_77_n 0.00384288f $X=-0.19 $Y=1.305 $X2=2.435 $Y2=1.62
cc_41 VPB N_B1_N_M1003_g 0.0233542f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB B1_N 0.00256362f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_43 VPB N_B1_N_c_148_n 0.0057822f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_44 VPB N_A_222_93#_M1004_g 0.0228293f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.56
cc_45 VPB N_A_222_93#_c_182_n 0.0190302f $X=-0.19 $Y=1.305 $X2=0.727 $Y2=1.325
cc_46 VPB N_A_222_93#_c_183_n 6.60476e-19 $X=-0.19 $Y=1.305 $X2=0.727 $Y2=1.865
cc_47 VPB N_A_222_93#_c_190_n 0.00953566f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.95
cc_48 VPB N_A_222_93#_c_185_n 0.00374886f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_49 VPB N_A2_M1001_g 0.0188916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A2_c_236_n 0.00407808f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_51 VPB N_A1_M1007_g 0.0246977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A1_c_270_n 0.00717796f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_53 VPB N_X_c_297_n 0.0075044f $X=-0.19 $Y=1.305 $X2=0.727 $Y2=1.865
cc_54 VPB N_X_c_296_n 0.00825319f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.95
cc_55 VPB X 0.0322798f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.95
cc_56 VPB N_VPWR_c_315_n 0.0187885f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.56
cc_57 VPB N_VPWR_c_316_n 0.0163315f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.95
cc_58 VPB N_VPWR_c_317_n 0.0389751f $X=-0.19 $Y=1.305 $X2=1.955 $Y2=0.57
cc_59 VPB N_VPWR_c_318_n 0.0258873f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_60 VPB N_VPWR_c_319_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_61 VPB N_VPWR_c_320_n 0.0177718f $X=-0.19 $Y=1.305 $X2=1.955 $Y2=1.745
cc_62 VPB N_VPWR_c_321_n 0.0206555f $X=-0.19 $Y=1.305 $X2=2.435 $Y2=1.96
cc_63 VPB N_VPWR_c_322_n 0.0116899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_314_n 0.0607061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_324_n 0.00785178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_325_n 0.00631679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 N_A_79_199#_M1006_g N_B1_N_M1003_g 0.0143627f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_79_199#_c_72_n N_B1_N_M1003_g 0.00552641f $X=0.727 $Y=1.865 $X2=0
+ $Y2=0
cc_69 N_A_79_199#_c_76_n N_B1_N_M1003_g 0.0153002f $X=1.87 $Y=1.745 $X2=0 $Y2=0
cc_70 N_A_79_199#_c_68_n B1_N 0.0262363f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_79_199#_c_69_n B1_N 2.92622e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_79_199#_c_76_n B1_N 0.00122077f $X=1.87 $Y=1.745 $X2=0 $Y2=0
cc_73 N_A_79_199#_c_68_n N_B1_N_c_148_n 0.00552641f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_79_199#_c_69_n N_B1_N_c_148_n 0.0181094f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_79_199#_c_70_n N_B1_N_c_149_n 0.00896998f $X=0.562 $Y=0.995 $X2=0
+ $Y2=0
cc_76 N_A_79_199#_c_76_n N_A_222_93#_M1003_d 0.00248196f $X=1.87 $Y=1.745 $X2=0
+ $Y2=0
cc_77 N_A_79_199#_c_67_n N_A_222_93#_c_181_n 0.00857073f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_78 N_A_79_199#_c_67_n N_A_222_93#_M1004_g 0.00505412f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_79 N_A_79_199#_c_77_n N_A_222_93#_M1004_g 0.0303987f $X=2.435 $Y=1.62 $X2=0
+ $Y2=0
cc_80 N_A_79_199#_c_67_n N_A_222_93#_c_182_n 0.0210961f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_81 N_A_79_199#_c_76_n N_A_222_93#_c_182_n 0.00495661f $X=1.87 $Y=1.745 $X2=0
+ $Y2=0
cc_82 N_A_79_199#_c_77_n N_A_222_93#_c_182_n 0.00323506f $X=2.435 $Y=1.62 $X2=0
+ $Y2=0
cc_83 N_A_79_199#_c_72_n N_A_222_93#_c_190_n 0.0112834f $X=0.727 $Y=1.865 $X2=0
+ $Y2=0
cc_84 N_A_79_199#_c_76_n N_A_222_93#_c_190_n 0.0433983f $X=1.87 $Y=1.745 $X2=0
+ $Y2=0
cc_85 N_A_79_199#_c_77_n N_A_222_93#_c_190_n 0.0155696f $X=2.435 $Y=1.62 $X2=0
+ $Y2=0
cc_86 N_A_79_199#_c_67_n N_A_222_93#_c_184_n 0.0134462f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_87 N_A_79_199#_c_72_n N_A_222_93#_c_185_n 0.00581423f $X=0.727 $Y=1.865 $X2=0
+ $Y2=0
cc_88 N_A_79_199#_c_67_n N_A_222_93#_c_185_n 0.0448395f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_89 N_A_79_199#_c_77_n N_A_222_93#_c_185_n 0.00573599f $X=2.435 $Y=1.62 $X2=0
+ $Y2=0
cc_90 N_A_79_199#_c_67_n N_A_222_93#_c_186_n 0.00636126f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_91 N_A_79_199#_c_102_p N_A2_M1001_g 0.00636844f $X=2.412 $Y=1.745 $X2=0 $Y2=0
cc_92 N_A_79_199#_c_77_n N_A2_M1001_g 0.00923011f $X=2.435 $Y=1.62 $X2=0 $Y2=0
cc_93 N_A_79_199#_c_67_n A2 0.0156123f $X=1.955 $Y=0.57 $X2=0 $Y2=0
cc_94 N_A_79_199#_c_77_n A2 0.029981f $X=2.435 $Y=1.62 $X2=0 $Y2=0
cc_95 N_A_79_199#_c_67_n N_A2_c_236_n 6.91749e-19 $X=1.955 $Y=0.57 $X2=0 $Y2=0
cc_96 N_A_79_199#_c_77_n N_A2_c_236_n 0.00291303f $X=2.435 $Y=1.62 $X2=0 $Y2=0
cc_97 N_A_79_199#_c_102_p N_A1_M1007_g 0.00113093f $X=2.412 $Y=1.745 $X2=0 $Y2=0
cc_98 N_A_79_199#_c_77_n N_A1_M1007_g 0.00168327f $X=2.435 $Y=1.62 $X2=0 $Y2=0
cc_99 N_A_79_199#_c_69_n N_X_c_295_n 0.00137863f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_79_199#_M1006_g N_X_c_297_n 0.00254905f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_79_199#_c_72_n N_X_c_297_n 0.0146356f $X=0.727 $Y=1.865 $X2=0 $Y2=0
cc_102 N_A_79_199#_c_72_n N_X_c_296_n 0.00930955f $X=0.727 $Y=1.865 $X2=0 $Y2=0
cc_103 N_A_79_199#_c_68_n N_X_c_296_n 0.0256987f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_79_199#_c_69_n N_X_c_296_n 0.0122262f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_79_199#_c_70_n N_X_c_296_n 0.00578113f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_79_199#_M1006_g X 0.0146289f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_79_199#_c_72_n N_VPWR_M1006_d 0.0084033f $X=0.727 $Y=1.865 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_79_199#_c_119_p N_VPWR_M1006_d 0.00441535f $X=0.86 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_79_199#_c_76_n N_VPWR_M1006_d 0.00185007f $X=1.87 $Y=1.745 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_79_199#_c_76_n N_VPWR_M1004_s 0.00282833f $X=1.87 $Y=1.745 $X2=0
+ $Y2=0
cc_111 N_A_79_199#_c_77_n N_VPWR_M1004_s 0.0129876f $X=2.435 $Y=1.62 $X2=0 $Y2=0
cc_112 N_A_79_199#_M1006_g N_VPWR_c_315_n 0.0100225f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_79_199#_c_119_p N_VPWR_c_315_n 0.0220308f $X=0.86 $Y=1.95 $X2=0 $Y2=0
cc_114 N_A_79_199#_c_76_n N_VPWR_c_315_n 0.0113161f $X=1.87 $Y=1.745 $X2=0 $Y2=0
cc_115 N_A_79_199#_c_76_n N_VPWR_c_316_n 0.0218908f $X=1.87 $Y=1.745 $X2=0 $Y2=0
cc_116 N_A_79_199#_c_102_p N_VPWR_c_317_n 0.0139781f $X=2.412 $Y=1.745 $X2=0
+ $Y2=0
cc_117 N_A_79_199#_c_77_n N_VPWR_c_317_n 0.0172574f $X=2.435 $Y=1.62 $X2=0 $Y2=0
cc_118 N_A_79_199#_c_102_p N_VPWR_c_318_n 0.0185827f $X=2.412 $Y=1.745 $X2=0
+ $Y2=0
cc_119 N_A_79_199#_c_77_n N_VPWR_c_318_n 0.00255839f $X=2.435 $Y=1.62 $X2=0
+ $Y2=0
cc_120 N_A_79_199#_M1006_g N_VPWR_c_320_n 0.00541359f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_79_199#_c_76_n N_VPWR_c_321_n 0.0120672f $X=1.87 $Y=1.745 $X2=0 $Y2=0
cc_122 N_A_79_199#_M1004_d N_VPWR_c_314_n 0.00267758f $X=2.24 $Y=1.485 $X2=0
+ $Y2=0
cc_123 N_A_79_199#_M1006_g N_VPWR_c_314_n 0.0119085f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_79_199#_c_119_p N_VPWR_c_314_n 0.00121687f $X=0.86 $Y=1.95 $X2=0
+ $Y2=0
cc_125 N_A_79_199#_c_76_n N_VPWR_c_314_n 0.0223037f $X=1.87 $Y=1.745 $X2=0 $Y2=0
cc_126 N_A_79_199#_c_102_p N_VPWR_c_314_n 0.0122055f $X=2.412 $Y=1.745 $X2=0
+ $Y2=0
cc_127 N_A_79_199#_c_77_n N_VPWR_c_314_n 0.00408517f $X=2.435 $Y=1.62 $X2=0
+ $Y2=0
cc_128 N_A_79_199#_c_68_n N_VGND_c_366_n 0.0135196f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_79_199#_c_70_n N_VGND_c_366_n 0.0120662f $X=0.562 $Y=0.995 $X2=0
+ $Y2=0
cc_130 N_A_79_199#_c_70_n N_VGND_c_368_n 0.00585385f $X=0.562 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_A_79_199#_c_67_n N_VGND_c_370_n 0.0116048f $X=1.955 $Y=0.57 $X2=0 $Y2=0
cc_132 N_A_79_199#_M1009_s N_VGND_c_373_n 0.00529506f $X=1.83 $Y=0.235 $X2=0
+ $Y2=0
cc_133 N_A_79_199#_c_67_n N_VGND_c_373_n 0.00646998f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_134 N_A_79_199#_c_70_n N_VGND_c_373_n 0.0132154f $X=0.562 $Y=0.995 $X2=0
+ $Y2=0
cc_135 N_A_79_199#_c_67_n N_A_448_47#_c_412_n 0.00129594f $X=1.955 $Y=0.57 $X2=0
+ $Y2=0
cc_136 B1_N N_A_222_93#_c_182_n 0.00227505f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_137 N_B1_N_c_148_n N_A_222_93#_c_182_n 0.0217093f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_B1_N_M1003_g N_A_222_93#_c_190_n 0.00300503f $X=1.035 $Y=1.695 $X2=0
+ $Y2=0
cc_139 B1_N N_A_222_93#_c_190_n 0.0169968f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_140 N_B1_N_c_148_n N_A_222_93#_c_190_n 9.53075e-19 $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_141 B1_N N_A_222_93#_c_184_n 0.00227139f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_142 N_B1_N_M1003_g N_A_222_93#_c_185_n 0.00297981f $X=1.035 $Y=1.695 $X2=0
+ $Y2=0
cc_143 B1_N N_A_222_93#_c_185_n 0.0249156f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_144 N_B1_N_c_148_n N_A_222_93#_c_185_n 3.20855e-19 $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_B1_N_c_149_n N_A_222_93#_c_185_n 0.00405351f $X=1.115 $Y=0.995 $X2=0
+ $Y2=0
cc_146 B1_N N_A_222_93#_c_186_n 0.0132981f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_147 N_B1_N_c_148_n N_A_222_93#_c_186_n 8.01366e-19 $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_148 N_B1_N_c_149_n N_A_222_93#_c_186_n 3.5039e-19 $X=1.115 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_B1_N_M1003_g N_VPWR_c_315_n 0.00119309f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_150 N_B1_N_M1003_g N_VPWR_c_321_n 0.00181247f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_151 N_B1_N_M1003_g N_VPWR_c_314_n 0.00295025f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_152 N_B1_N_c_149_n N_VGND_c_366_n 0.00435523f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B1_N_c_149_n N_VGND_c_370_n 0.00510437f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B1_N_c_149_n N_VGND_c_373_n 0.00512902f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_222_93#_M1004_g N_A2_M1001_g 0.0116008f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_222_93#_c_183_n A2 0.00726323f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_222_93#_c_183_n N_A2_c_236_n 0.022512f $X=2.165 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_222_93#_c_181_n N_A2_c_237_n 0.00957314f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_222_93#_M1004_g N_VPWR_c_316_n 0.00491123f $X=2.165 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_222_93#_M1004_g N_VPWR_c_318_n 0.00432313f $X=2.165 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_222_93#_M1004_g N_VPWR_c_314_n 0.00718232f $X=2.165 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_222_93#_c_186_n N_VGND_c_366_n 0.0098012f $X=1.245 $Y=0.66 $X2=0
+ $Y2=0
cc_163 N_A_222_93#_c_181_n N_VGND_c_370_n 0.00585385f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_222_93#_c_184_n N_VGND_c_370_n 0.00677941f $X=1.53 $Y=0.74 $X2=0
+ $Y2=0
cc_165 N_A_222_93#_c_186_n N_VGND_c_370_n 0.00512277f $X=1.245 $Y=0.66 $X2=0
+ $Y2=0
cc_166 N_A_222_93#_c_181_n N_VGND_c_373_n 0.0122806f $X=2.165 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_222_93#_c_184_n N_VGND_c_373_n 0.0106136f $X=1.53 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_222_93#_c_186_n N_VGND_c_373_n 0.00563626f $X=1.245 $Y=0.66 $X2=0
+ $Y2=0
cc_169 N_A_222_93#_c_181_n N_A_448_47#_c_412_n 2.04248e-19 $X=2.165 $Y=0.995
+ $X2=0 $Y2=0
cc_170 N_A2_M1001_g N_A1_M1007_g 0.0492314f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_171 A2 A1 0.0182181f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A2_c_236_n A1 2.21375e-19 $X=2.585 $Y=1.16 $X2=0 $Y2=0
cc_173 A2 N_A1_c_270_n 0.00129893f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A2_c_236_n N_A1_c_270_n 0.0492314f $X=2.585 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A2_c_237_n N_A1_c_271_n 0.0258192f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A2_M1001_g N_VPWR_c_317_n 0.00380898f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M1001_g N_VPWR_c_318_n 0.00578292f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_M1001_g N_VPWR_c_314_n 0.0105848f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_c_237_n N_VGND_c_367_n 0.00268723f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_237_n N_VGND_c_370_n 0.00424416f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A2_c_237_n N_VGND_c_373_n 0.00593107f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_c_237_n N_A_448_47#_c_416_n 0.00648375f $X=2.585 $Y=0.995 $X2=0
+ $Y2=0
cc_183 A2 N_A_448_47#_c_411_n 0.0128259f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A2_c_237_n N_A_448_47#_c_411_n 0.00845772f $X=2.585 $Y=0.995 $X2=0
+ $Y2=0
cc_185 A2 N_A_448_47#_c_412_n 0.0274572f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_186 N_A2_c_236_n N_A_448_47#_c_412_n 0.00307118f $X=2.585 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A2_c_237_n N_A_448_47#_c_412_n 0.00110465f $X=2.585 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A2_c_237_n N_A_448_47#_c_413_n 5.47159e-19 $X=2.585 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A1_M1007_g N_VPWR_c_317_n 0.022185f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_190 A1 N_VPWR_c_317_n 0.0179232f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A1_c_270_n N_VPWR_c_317_n 0.00467945f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A1_M1007_g N_VPWR_c_318_n 0.0046653f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A1_M1007_g N_VPWR_c_314_n 0.00783311f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A1_c_271_n N_VGND_c_367_n 0.00268723f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A1_c_271_n N_VGND_c_372_n 0.00425021f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_271_n N_VGND_c_373_n 0.00683108f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_271_n N_A_448_47#_c_416_n 5.5158e-19 $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_198 A1 N_A_448_47#_c_411_n 0.038466f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A1_c_270_n N_A_448_47#_c_411_n 0.00564384f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A1_c_271_n N_A_448_47#_c_411_n 0.00972538f $X=3.105 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A1_c_271_n N_A_448_47#_c_413_n 0.00634641f $X=3.105 $Y=0.995 $X2=0
+ $Y2=0
cc_202 X N_VPWR_c_320_n 0.0217551f $X=0.145 $Y=2.125 $X2=0 $Y2=0
cc_203 N_X_M1006_s N_VPWR_c_314_n 0.00209319f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_204 X N_VPWR_c_314_n 0.0128119f $X=0.145 $Y=2.125 $X2=0 $Y2=0
cc_205 N_X_c_295_n N_VGND_c_368_n 0.0106755f $X=0.34 $Y=0.66 $X2=0 $Y2=0
cc_206 N_X_M1005_s N_VGND_c_373_n 0.00346044f $X=0.215 $Y=0.235 $X2=0 $Y2=0
cc_207 N_X_c_295_n N_VGND_c_373_n 0.0122067f $X=0.34 $Y=0.66 $X2=0 $Y2=0
cc_208 N_VPWR_c_314_n A_544_297# 0.00897657f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_209 N_VGND_c_373_n N_A_448_47#_M1009_d 0.00367527f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_210 N_VGND_c_373_n N_A_448_47#_M1008_d 0.00213973f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_370_n N_A_448_47#_c_416_n 0.0200223f $X=2.77 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_373_n N_A_448_47#_c_416_n 0.0124119f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_M1000_d N_A_448_47#_c_411_n 0.00165819f $X=2.72 $Y=0.235 $X2=0
+ $Y2=0
cc_214 N_VGND_c_367_n N_A_448_47#_c_411_n 0.0116529f $X=2.855 $Y=0.39 $X2=0
+ $Y2=0
cc_215 N_VGND_c_370_n N_A_448_47#_c_411_n 0.00193763f $X=2.77 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_372_n N_A_448_47#_c_411_n 0.00193763f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_373_n N_A_448_47#_c_411_n 0.00827287f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_372_n N_A_448_47#_c_413_n 0.0191098f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_373_n N_A_448_47#_c_413_n 0.0123122f $X=3.45 $Y=0 $X2=0 $Y2=0

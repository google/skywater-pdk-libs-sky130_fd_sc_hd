* File: sky130_fd_sc_hd__o311a_4.pex.spice
* Created: Thu Aug 27 14:39:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O311A_4%A_79_21# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 41 47 49 51 52 53 54 56 60 62 66 68 70 74 75 76 77 78
c137 74 0 8.02102e-20 $X=1.78 $Y=1.16
r138 83 84 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r139 79 81 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r140 75 84 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.78 $Y=1.16 $X2=1.73
+ $Y2=1.16
r141 74 75 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=1.16 $X2=1.78 $Y2=1.16
r142 70 72 6.45882 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.92 $Y=1.725 $X2=4.92
+ $Y2=1.815
r143 69 78 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=1.605
+ $X2=3.54 $Y2=1.605
r144 68 70 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=4.835 $Y=1.605
+ $X2=4.92 $Y2=1.725
r145 68 69 58.1023 $w=2.38e-07 $l=1.21e-06 $layer=LI1_cond $X=4.835 $Y=1.605
+ $X2=3.625 $Y2=1.605
r146 64 78 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.54 $Y=1.725
+ $X2=3.54 $Y2=1.605
r147 64 66 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=1.725
+ $X2=3.54 $Y2=1.815
r148 63 77 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.605
+ $X2=2.7 $Y2=1.605
r149 62 78 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=1.605
+ $X2=3.54 $Y2=1.605
r150 62 63 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=3.455 $Y=1.605
+ $X2=2.785 $Y2=1.605
r151 58 77 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.7 $Y=1.725 $X2=2.7
+ $Y2=1.605
r152 58 60 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.7 $Y=1.725 $X2=2.7
+ $Y2=1.815
r153 54 76 5.98033 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=2.3 $Y=0.78
+ $X2=2.195 $Y2=0.78
r154 54 56 30.632 $w=2.08e-07 $l=5.8e-07 $layer=LI1_cond $X=2.3 $Y=0.78 $X2=2.88
+ $Y2=0.78
r155 52 77 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=1.605
+ $X2=2.7 $Y2=1.605
r156 52 53 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=2.615 $Y=1.605
+ $X2=1.945 $Y2=1.605
r157 51 76 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.945 $Y=0.8
+ $X2=2.195 $Y2=0.8
r158 49 53 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.86 $Y=1.485
+ $X2=1.945 $Y2=1.605
r159 48 74 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.86 $Y=1.315
+ $X2=1.86 $Y2=1.185
r160 48 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.86 $Y=1.315
+ $X2=1.86 $Y2=1.485
r161 47 74 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.86 $Y=1.055
+ $X2=1.86 $Y2=1.185
r162 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.86 $Y=0.885
+ $X2=1.945 $Y2=0.8
r163 46 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.86 $Y=0.885
+ $X2=1.86 $Y2=1.055
r164 44 83 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.1 $Y=1.16
+ $X2=1.31 $Y2=1.16
r165 44 81 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.1 $Y=1.16
+ $X2=0.89 $Y2=1.16
r166 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r167 41 74 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=1.185
+ $X2=1.86 $Y2=1.185
r168 41 43 29.9192 $w=2.58e-07 $l=6.75e-07 $layer=LI1_cond $X=1.775 $Y=1.185
+ $X2=1.1 $Y2=1.185
r169 37 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r170 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r171 34 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r172 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r173 30 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r174 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r175 27 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r176 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r177 23 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r178 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r179 20 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r180 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r181 16 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r182 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r183 13 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r184 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r185 4 72 600 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=1 $X=4.785
+ $Y=1.485 $X2=4.92 $Y2=1.815
r186 3 66 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.54 $Y2=1.815
r187 2 60 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=2.565
+ $Y=1.485 $X2=2.7 $Y2=1.815
r188 1 56 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%C1 3 5 7 10 12 14 15 16 24
c53 3 0 1.54085e-20 $X=2.49 $Y=1.985
r54 22 24 14.7051 $w=2.95e-07 $l=9e-08 $layer=POLY_cond $X=2.82 $Y=1.127
+ $X2=2.91 $Y2=1.127
r55 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.16 $X2=2.82 $Y2=1.16
r56 20 22 24.5085 $w=2.95e-07 $l=1.5e-07 $layer=POLY_cond $X=2.67 $Y=1.127
+ $X2=2.82 $Y2=1.127
r57 19 20 29.4102 $w=2.95e-07 $l=1.8e-07 $layer=POLY_cond $X=2.49 $Y=1.127
+ $X2=2.67 $Y2=1.127
r58 16 23 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=2.995 $Y=1.185
+ $X2=2.82 $Y2=1.185
r59 15 23 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.535 $Y=1.185
+ $X2=2.82 $Y2=1.185
r60 12 24 29.4102 $w=2.95e-07 $l=2.4992e-07 $layer=POLY_cond $X=3.09 $Y=0.96
+ $X2=2.91 $Y2=1.127
r61 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.09 $Y=0.96 $X2=3.09
+ $Y2=0.56
r62 8 24 18.5736 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=2.91 $Y=1.295
+ $X2=2.91 $Y2=1.127
r63 8 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.91 $Y=1.295
+ $X2=2.91 $Y2=1.985
r64 5 20 18.5736 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=2.67 $Y=0.96
+ $X2=2.67 $Y2=1.127
r65 5 7 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.67 $Y=0.96 $X2=2.67
+ $Y2=0.56
r66 1 19 18.5736 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=2.49 $Y=1.295
+ $X2=2.49 $Y2=1.127
r67 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.49 $Y=1.295 $X2=2.49
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%B1 1 3 4 6 7 9 10 12 13 14 15 24
c45 24 0 1.71287e-19 $X=3.75 $Y=1.202
r46 24 25 25.8985 $w=3.35e-07 $l=1.8e-07 $layer=POLY_cond $X=3.75 $Y=1.202
+ $X2=3.93 $Y2=1.202
r47 22 24 7.19403 $w=3.35e-07 $l=5e-08 $layer=POLY_cond $X=3.7 $Y=1.202 $X2=3.75
+ $Y2=1.202
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.7
+ $Y=1.16 $X2=3.7 $Y2=1.16
r49 20 22 27.3373 $w=3.35e-07 $l=1.9e-07 $layer=POLY_cond $X=3.51 $Y=1.202
+ $X2=3.7 $Y2=1.202
r50 14 15 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=3.915 $Y=1.185
+ $X2=4.375 $Y2=1.185
r51 14 23 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=3.915 $Y=1.185
+ $X2=3.7 $Y2=1.185
r52 13 23 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=3.455 $Y=1.185
+ $X2=3.7 $Y2=1.185
r53 10 25 21.5811 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=0.56
r55 7 24 21.5811 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.75 $Y=1.41
+ $X2=3.75 $Y2=1.202
r56 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.75 $Y=1.41 $X2=3.75
+ $Y2=1.985
r57 4 20 21.5811 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.202
r58 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995 $X2=3.51
+ $Y2=0.56
r59 1 20 25.8985 $w=3.35e-07 $l=2.84085e-07 $layer=POLY_cond $X=3.33 $Y=1.41
+ $X2=3.51 $Y2=1.202
r60 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.33 $Y=1.41 $X2=3.33
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%A3 3 7 11 15 17 18 19 20 24
c49 20 0 1.71287e-19 $X=5.755 $Y=1.19
r50 33 34 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=4.88 $Y=1.16
+ $X2=5.13 $Y2=1.16
r51 31 33 13.3304 $w=2.7e-07 $l=6e-08 $layer=POLY_cond $X=4.82 $Y=1.16 $X2=4.88
+ $Y2=1.16
r52 28 31 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=4.71 $Y=1.16
+ $X2=4.82 $Y2=1.16
r53 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.5 $Y=1.16
+ $X2=5.5 $Y2=1.16
r54 24 34 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.205 $Y=1.16
+ $X2=5.13 $Y2=1.16
r55 24 26 65.5412 $w=2.7e-07 $l=2.95e-07 $layer=POLY_cond $X=5.205 $Y=1.16
+ $X2=5.5 $Y2=1.16
r56 20 27 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=5.755 $Y=1.185
+ $X2=5.5 $Y2=1.185
r57 19 27 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=5.295 $Y=1.185
+ $X2=5.5 $Y2=1.185
r58 18 19 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=4.82 $Y=1.185
+ $X2=5.295 $Y2=1.185
r59 18 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.82
+ $Y=1.16 $X2=4.82 $Y2=1.16
r60 17 26 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.575 $Y=1.16 $X2=5.5
+ $Y2=1.16
r61 13 17 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=5.65 $Y=1.025
+ $X2=5.575 $Y2=1.16
r62 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.65 $Y=1.025
+ $X2=5.65 $Y2=0.56
r63 9 34 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.13 $Y=1.295
+ $X2=5.13 $Y2=1.16
r64 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.13 $Y=1.295
+ $X2=5.13 $Y2=1.985
r65 5 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.88 $Y=1.025
+ $X2=4.88 $Y2=1.16
r66 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.88 $Y=1.025
+ $X2=4.88 $Y2=0.56
r67 1 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.71 $Y=1.295
+ $X2=4.71 $Y2=1.16
r68 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.71 $Y=1.295 $X2=4.71
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%A2 3 7 11 15 17 18 26
c47 26 0 1.94677e-19 $X=6.49 $Y=1.16
r48 24 26 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=6.2 $Y=1.16 $X2=6.49
+ $Y2=1.16
r49 21 24 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=6.07 $Y=1.16 $X2=6.2
+ $Y2=1.16
r50 17 18 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=6.2 $Y=1.185
+ $X2=6.675 $Y2=1.185
r51 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.2
+ $Y=1.16 $X2=6.2 $Y2=1.16
r52 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.49 $Y=1.295
+ $X2=6.49 $Y2=1.16
r53 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.49 $Y=1.295
+ $X2=6.49 $Y2=1.985
r54 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.49 $Y=1.025
+ $X2=6.49 $Y2=1.16
r55 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.49 $Y=1.025
+ $X2=6.49 $Y2=0.56
r56 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.07 $Y=1.295
+ $X2=6.07 $Y2=1.16
r57 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.07 $Y=1.295 $X2=6.07
+ $Y2=1.985
r58 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.07 $Y=1.025
+ $X2=6.07 $Y2=1.16
r59 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.07 $Y=1.025
+ $X2=6.07 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%A1 3 7 11 15 17 18 25
c39 18 0 1.94677e-19 $X=7.595 $Y=1.19
r40 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.455
+ $Y=1.16 $X2=7.455 $Y2=1.16
r41 25 27 21.595 $w=2.79e-07 $l=1.25e-07 $layer=POLY_cond $X=7.33 $Y=1.16
+ $X2=7.455 $Y2=1.16
r42 23 25 37.1434 $w=2.79e-07 $l=2.15e-07 $layer=POLY_cond $X=7.115 $Y=1.16
+ $X2=7.33 $Y2=1.16
r43 18 28 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=7.595 $Y=1.185
+ $X2=7.455 $Y2=1.185
r44 17 28 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=7.115 $Y=1.185
+ $X2=7.455 $Y2=1.185
r45 17 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.115
+ $Y=1.16 $X2=7.115 $Y2=1.16
r46 13 25 17.2686 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.33 $Y=1.305
+ $X2=7.33 $Y2=1.16
r47 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.33 $Y=1.305
+ $X2=7.33 $Y2=1.985
r48 9 25 17.2686 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.33 $Y=1.015
+ $X2=7.33 $Y2=1.16
r49 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.33 $Y=1.015
+ $X2=7.33 $Y2=0.56
r50 1 23 35.4158 $w=2.79e-07 $l=2.05e-07 $layer=POLY_cond $X=6.91 $Y=1.16
+ $X2=7.115 $Y2=1.16
r51 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.91 $Y=1.295 $X2=6.91
+ $Y2=1.985
r52 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.91 $Y=1.025
+ $X2=6.91 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%VPWR 1 2 3 4 5 6 19 21 27 31 33 37 39 43 47
+ 49 51 56 61 71 72 78 81 84 87 90
r116 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r117 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r118 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r120 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r121 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r122 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r123 72 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r124 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r125 69 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=2.72
+ $X2=7.12 $Y2=2.72
r126 69 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.285 $Y=2.72
+ $X2=7.59 $Y2=2.72
r127 68 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r128 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r129 65 68 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.67 $Y2=2.72
r130 65 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r131 64 67 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.67 $Y2=2.72
r132 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 62 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.045 $Y=2.72
+ $X2=3.95 $Y2=2.72
r134 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.045 $Y=2.72
+ $X2=4.37 $Y2=2.72
r135 61 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.955 $Y=2.72
+ $X2=7.12 $Y2=2.72
r136 61 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.955 $Y=2.72
+ $X2=6.67 $Y2=2.72
r137 60 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r138 60 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.1 $Y2=2.72
r141 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.61 $Y2=2.72
r142 56 81 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=2.11 $Y2=2.72
r143 56 59 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.61 $Y2=2.72
r144 55 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r145 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 52 75 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r147 52 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.1 $Y2=2.72
r149 51 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r150 49 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 49 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r152 45 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.12 $Y=2.635
+ $X2=7.12 $Y2=2.72
r153 45 47 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=7.12 $Y=2.635
+ $X2=7.12 $Y2=2.02
r154 41 87 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=2.635
+ $X2=3.95 $Y2=2.72
r155 41 43 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=3.95 $Y=2.635
+ $X2=3.95 $Y2=2.06
r156 40 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=3.12 $Y2=2.72
r157 39 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.95 $Y2=2.72
r158 39 40 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.285 $Y2=2.72
r159 35 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.635
+ $X2=3.12 $Y2=2.72
r160 35 37 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.12 $Y=2.635
+ $X2=3.12 $Y2=2.02
r161 34 81 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.445 $Y=2.72
+ $X2=2.11 $Y2=2.72
r162 33 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=2.72
+ $X2=3.12 $Y2=2.72
r163 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.955 $Y=2.72
+ $X2=2.445 $Y2=2.72
r164 29 81 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=2.635
+ $X2=2.11 $Y2=2.72
r165 29 31 10.9789 $w=6.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.11 $Y=2.635
+ $X2=2.11 $Y2=2.02
r166 25 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r167 25 27 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2.02
r168 21 24 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=2.34
r169 19 75 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.212 $Y2=2.72
r170 19 24 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.255 $Y2=2.34
r171 6 47 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.985
+ $Y=1.485 $X2=7.12 $Y2=2.02
r172 5 43 600 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=1.485 $X2=3.96 $Y2=2.06
r173 4 37 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.485 $X2=3.12 $Y2=2.02
r174 3 31 150 $w=1.7e-07 $l=7.35085e-07 $layer=licon1_PDIFF $count=4 $X=1.805
+ $Y=1.485 $X2=2.28 $Y2=2.02
r175 2 27 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.02
r176 1 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r177 1 21 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%X 1 2 3 4 16 18 21 23 25 31 34 35 36 39 40
r46 35 40 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.595 $Y=1.185
+ $X2=0.235 $Y2=1.185
r47 35 36 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=1.185
+ $X2=0.68 $Y2=1.185
r48 29 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.52 $Y=1.725 $X2=1.52
+ $Y2=1.815
r49 26 37 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.605
+ $X2=0.68 $Y2=1.605
r50 25 29 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.435 $Y=1.605
+ $X2=1.52 $Y2=1.725
r51 25 26 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=1.605
+ $X2=0.765 $Y2=1.605
r52 24 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.8 $X2=0.68
+ $Y2=0.8
r53 23 39 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0.8 $X2=1.52
+ $Y2=0.8
r54 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=0.8
+ $X2=0.765 $Y2=0.8
r55 19 37 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.68 $Y=1.725
+ $X2=0.68 $Y2=1.605
r56 19 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.68 $Y=1.725 $X2=0.68
+ $Y2=1.815
r57 18 37 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.68 $Y=1.485
+ $X2=0.68 $Y2=1.605
r58 17 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=1.315
+ $X2=0.68 $Y2=1.185
r59 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=1.315
+ $X2=0.68 $Y2=1.485
r60 16 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=1.055
+ $X2=0.68 $Y2=1.185
r61 15 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.885
+ $X2=0.68 $Y2=0.8
r62 15 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=0.885
+ $X2=0.68 $Y2=1.055
r63 4 31 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.815
r64 3 21 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.815
r65 2 39 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.72
r66 1 34 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%A_875_297# 1 2 3 12 14 15 18 20 24 26
r46 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.28 $Y=2.295
+ $X2=6.28 $Y2=2.02
r47 21 26 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.525 $Y=2.38
+ $X2=5.39 $Y2=2.38
r48 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.115 $Y=2.38
+ $X2=6.28 $Y2=2.295
r49 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.115 $Y=2.38
+ $X2=5.525 $Y2=2.38
r50 16 26 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.39 $Y=2.295
+ $X2=5.39 $Y2=2.38
r51 16 18 20.9147 $w=2.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.39 $Y=2.295
+ $X2=5.39 $Y2=1.805
r52 14 26 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.255 $Y=2.38
+ $X2=5.39 $Y2=2.38
r53 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.255 $Y=2.38
+ $X2=4.665 $Y2=2.38
r54 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.5 $Y=2.295
+ $X2=4.665 $Y2=2.38
r55 10 12 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.5 $Y=2.295
+ $X2=4.5 $Y2=2.06
r56 3 24 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.145
+ $Y=1.485 $X2=6.28 $Y2=2.02
r57 2 18 600 $w=1.7e-07 $l=3.81576e-07 $layer=licon1_PDIFF $count=1 $X=5.205
+ $Y=1.485 $X2=5.34 $Y2=1.805
r58 1 12 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=4.375
+ $Y=1.485 $X2=4.5 $Y2=2.06
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%A_1147_297# 1 2 3 10 13 14 15 18 22 24
r36 20 22 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=7.595 $Y=1.725
+ $X2=7.595 $Y2=1.815
r37 19 24 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.785 $Y=1.605
+ $X2=6.7 $Y2=1.605
r38 18 20 6.86909 $w=2.4e-07 $l=1.90788e-07 $layer=LI1_cond $X=7.455 $Y=1.605
+ $X2=7.595 $Y2=1.725
r39 18 19 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=7.455 $Y=1.605
+ $X2=6.785 $Y2=1.605
r40 15 24 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.7 $Y=1.725 $X2=6.7
+ $Y2=1.605
r41 15 17 6.45882 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.7 $Y=1.725 $X2=6.7
+ $Y2=1.815
r42 13 24 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.615 $Y=1.605
+ $X2=6.7 $Y2=1.605
r43 13 14 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=6.615 $Y=1.605
+ $X2=5.945 $Y2=1.605
r44 10 14 6.82018 $w=2.4e-07 $l=1.75e-07 $layer=LI1_cond $X=5.82 $Y=1.725
+ $X2=5.945 $Y2=1.605
r45 10 12 4.392 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.82 $Y=1.725 $X2=5.82
+ $Y2=1.815
r46 3 22 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=7.405
+ $Y=1.485 $X2=7.54 $Y2=1.815
r47 2 17 600 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=1 $X=6.565
+ $Y=1.485 $X2=6.7 $Y2=1.815
r48 1 12 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.485 $X2=5.86 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 40 41 42
+ 44 60 65 72 73 79 84 87 89 92
r126 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r127 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r128 86 87 10.1923 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5.435 $Y=0.21
+ $X2=5.605 $Y2=0.21
r129 82 86 2.93951 $w=5.88e-07 $l=1.45e-07 $layer=LI1_cond $X=5.29 $Y=0.21
+ $X2=5.435 $Y2=0.21
r130 82 84 14.1454 $w=5.88e-07 $l=3.65e-07 $layer=LI1_cond $X=5.29 $Y=0.21
+ $X2=4.925 $Y2=0.21
r131 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r132 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r133 73 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r134 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r135 70 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=0 $X2=7.12
+ $Y2=0
r136 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.285 $Y=0
+ $X2=7.59 $Y2=0
r137 69 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r138 69 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r139 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r140 66 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.28
+ $Y2=0
r141 66 68 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=6.67 $Y2=0
r142 65 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.955 $Y=0 $X2=7.12
+ $Y2=0
r143 65 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.955 $Y=0
+ $X2=6.67 $Y2=0
r144 64 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r145 64 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r146 63 87 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=5.605 $Y2=0
r147 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r148 60 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0 $X2=6.28
+ $Y2=0
r149 60 63 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.115 $Y=0
+ $X2=5.75 $Y2=0
r150 59 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r151 58 84 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.925
+ $Y2=0
r152 58 59 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r153 56 59 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=4.83 $Y2=0
r154 55 58 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.83
+ $Y2=0
r155 55 56 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r156 52 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r157 52 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r158 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r159 49 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r160 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r161 48 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r162 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r163 45 76 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r164 45 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r165 44 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r166 44 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r167 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r168 42 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r169 40 51 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.61 $Y2=0
r170 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.9
+ $Y2=0
r171 39 55 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.07
+ $Y2=0
r172 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.9
+ $Y2=0
r173 35 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.12 $Y=0.085
+ $X2=7.12 $Y2=0
r174 35 37 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.12 $Y=0.085
+ $X2=7.12 $Y2=0.36
r175 31 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=0.085
+ $X2=6.28 $Y2=0
r176 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.28 $Y=0.085
+ $X2=6.28 $Y2=0.36
r177 27 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.9 $Y=0.085
+ $X2=1.9 $Y2=0
r178 27 29 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.9 $Y=0.085
+ $X2=1.9 $Y2=0.38
r179 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r180 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.36
r181 19 76 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.212 $Y2=0
r182 19 21 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.38
r183 6 37 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.985
+ $Y=0.235 $X2=7.12 $Y2=0.36
r184 5 33 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.145
+ $Y=0.235 $X2=6.28 $Y2=0.36
r185 4 86 91 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=2 $X=4.955
+ $Y=0.235 $X2=5.435 $Y2=0.36
r186 3 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r187 2 25 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.36
r188 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%A_467_47# 1 2 3 10 16 20 23
r28 18 23 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=0.38 $X2=3.3
+ $Y2=0.38
r29 18 20 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=3.385 $Y=0.38
+ $X2=4.14 $Y2=0.38
r30 14 23 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.3 $Y=0.505 $X2=3.3
+ $Y2=0.38
r31 14 16 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.3 $Y=0.505
+ $X2=3.3 $Y2=0.7
r32 10 23 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0.38 $X2=3.3
+ $Y2=0.38
r33 10 12 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=3.215 $Y=0.38
+ $X2=2.46 $Y2=0.38
r34 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.38
r35 2 23 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.36
r36 2 16 182 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.7
r37 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_4%A_717_47# 1 2 3 4 5 16 22 26 30 35 37 39 41
r68 31 39 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.785 $Y=0.78 $X2=6.7
+ $Y2=0.78
r69 30 41 3.99943 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=7.455 $Y=0.78
+ $X2=7.595 $Y2=0.78
r70 30 31 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=7.455 $Y=0.78
+ $X2=6.785 $Y2=0.78
r71 27 37 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.945 $Y=0.78 $X2=5.86
+ $Y2=0.78
r72 26 39 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.615 $Y=0.78 $X2=6.7
+ $Y2=0.78
r73 26 27 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=6.615 $Y=0.78
+ $X2=5.945 $Y2=0.78
r74 23 35 6.33349 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=4.755 $Y=0.78
+ $X2=4.62 $Y2=0.78
r75 22 37 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.775 $Y=0.78 $X2=5.86
+ $Y2=0.78
r76 22 23 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=5.775 $Y=0.78
+ $X2=4.755 $Y2=0.78
r77 16 35 6.33349 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=4.485 $Y=0.78
+ $X2=4.62 $Y2=0.78
r78 16 18 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=4.485 $Y=0.78
+ $X2=3.72 $Y2=0.78
r79 5 41 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=7.405
+ $Y=0.235 $X2=7.54 $Y2=0.72
r80 4 39 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.7 $Y2=0.72
r81 3 37 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.725
+ $Y=0.235 $X2=5.86 $Y2=0.72
r82 2 35 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.235 $X2=4.67 $Y2=0.72
r83 1 18 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.76
.ends


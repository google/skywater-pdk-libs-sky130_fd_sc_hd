* File: sky130_fd_sc_hd__a41oi_2.spice.SKY130_FD_SC_HD__A41OI_2.pxi
* Created: Thu Aug 27 14:06:29 2020
* 
x_PM_SKY130_FD_SC_HD__A41OI_2%B1 N_B1_c_77_n N_B1_M1000_g N_B1_c_78_n
+ N_B1_M1014_g N_B1_M1006_g N_B1_M1018_g B1 B1 N_B1_c_84_p N_B1_c_79_n
+ PM_SKY130_FD_SC_HD__A41OI_2%B1
x_PM_SKY130_FD_SC_HD__A41OI_2%A1 N_A1_c_119_n N_A1_M1008_g N_A1_M1002_g
+ N_A1_c_120_n N_A1_M1011_g N_A1_M1019_g A1 N_A1_c_121_n N_A1_c_122_n
+ PM_SKY130_FD_SC_HD__A41OI_2%A1
x_PM_SKY130_FD_SC_HD__A41OI_2%A2 N_A2_M1015_g N_A2_M1010_g N_A2_M1016_g
+ N_A2_M1017_g A2 N_A2_c_166_n N_A2_c_167_n PM_SKY130_FD_SC_HD__A41OI_2%A2
x_PM_SKY130_FD_SC_HD__A41OI_2%A3 N_A3_M1001_g N_A3_M1005_g N_A3_M1012_g
+ N_A3_M1013_g N_A3_c_209_n A3 A3 N_A3_c_211_n N_A3_c_212_n
+ PM_SKY130_FD_SC_HD__A41OI_2%A3
x_PM_SKY130_FD_SC_HD__A41OI_2%A4 N_A4_M1003_g N_A4_M1004_g N_A4_M1007_g
+ N_A4_M1009_g A4 A4 A4 N_A4_c_258_n N_A4_c_259_n PM_SKY130_FD_SC_HD__A41OI_2%A4
x_PM_SKY130_FD_SC_HD__A41OI_2%A_149_297# N_A_149_297#_M1006_d
+ N_A_149_297#_M1018_d N_A_149_297#_M1019_s N_A_149_297#_M1017_d
+ N_A_149_297#_M1013_s N_A_149_297#_M1009_d N_A_149_297#_c_321_p
+ N_A_149_297#_c_294_n N_A_149_297#_c_334_p N_A_149_297#_c_296_n
+ N_A_149_297#_c_300_n N_A_149_297#_c_335_p N_A_149_297#_c_301_n
+ N_A_149_297#_c_305_n N_A_149_297#_c_308_n N_A_149_297#_c_332_p
+ N_A_149_297#_c_293_n N_A_149_297#_c_337_p N_A_149_297#_c_306_n
+ N_A_149_297#_c_317_n PM_SKY130_FD_SC_HD__A41OI_2%A_149_297#
x_PM_SKY130_FD_SC_HD__A41OI_2%Y N_Y_M1000_d N_Y_M1008_s N_Y_M1006_s N_Y_c_392_p
+ N_Y_c_350_n N_Y_c_359_n N_Y_c_361_n N_Y_c_363_n N_Y_c_353_n Y Y Y N_Y_c_351_n
+ N_Y_c_354_n Y PM_SKY130_FD_SC_HD__A41OI_2%Y
x_PM_SKY130_FD_SC_HD__A41OI_2%VPWR N_VPWR_M1002_d N_VPWR_M1010_s N_VPWR_M1001_d
+ N_VPWR_M1004_s N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n
+ N_VPWR_c_409_n N_VPWR_c_410_n VPWR N_VPWR_c_411_n N_VPWR_c_412_n
+ N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_404_n N_VPWR_c_416_n N_VPWR_c_417_n
+ N_VPWR_c_418_n PM_SKY130_FD_SC_HD__A41OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A41OI_2%VGND N_VGND_M1000_s N_VGND_M1014_s N_VGND_M1003_s
+ N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n
+ N_VGND_c_485_n VGND N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n
+ N_VGND_c_489_n PM_SKY130_FD_SC_HD__A41OI_2%VGND
x_PM_SKY130_FD_SC_HD__A41OI_2%A_317_47# N_A_317_47#_M1008_d N_A_317_47#_M1011_d
+ N_A_317_47#_M1016_d N_A_317_47#_c_559_n N_A_317_47#_c_560_n
+ PM_SKY130_FD_SC_HD__A41OI_2%A_317_47#
x_PM_SKY130_FD_SC_HD__A41OI_2%A_567_47# N_A_567_47#_M1015_s N_A_567_47#_M1005_s
+ N_A_567_47#_c_585_n PM_SKY130_FD_SC_HD__A41OI_2%A_567_47#
x_PM_SKY130_FD_SC_HD__A41OI_2%A_757_47# N_A_757_47#_M1005_d N_A_757_47#_M1012_d
+ N_A_757_47#_M1007_d N_A_757_47#_c_604_n N_A_757_47#_c_623_n
+ PM_SKY130_FD_SC_HD__A41OI_2%A_757_47#
cc_1 VNB N_B1_c_77_n 0.0183849f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.995
cc_2 VNB N_B1_c_78_n 0.0210851f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=0.995
cc_3 VNB N_B1_c_79_n 0.0650253f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.16
cc_4 VNB N_A1_c_119_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.995
cc_5 VNB N_A1_c_120_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.985
cc_6 VNB N_A1_c_121_n 0.00307632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A1_c_122_n 0.0367159f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_8 VNB N_A2_M1015_g 0.017802f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.56
cc_9 VNB N_A2_M1010_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.325
cc_10 VNB N_A2_M1016_g 0.0243831f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.325
cc_11 VNB N_A2_M1017_g 4.72682e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_12 VNB N_A2_c_166_n 0.00193269f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_13 VNB N_A2_c_167_n 0.0362021f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.16
cc_14 VNB N_A3_M1001_g 7.42991e-19 $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.56
cc_15 VNB N_A3_M1005_g 0.0243831f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.325
cc_16 VNB N_A3_M1012_g 0.017802f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.325
cc_17 VNB N_A3_M1013_g 7.36106e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_18 VNB N_A3_c_209_n 0.0124857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB A3 0.00143625f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_20 VNB N_A3_c_211_n 0.0254321f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_21 VNB N_A3_c_212_n 0.0318748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A4_M1003_g 0.0175748f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.56
cc_23 VNB N_A4_M1004_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.325
cc_24 VNB N_A4_M1007_g 0.0233553f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.325
cc_25 VNB A4 0.0131271f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_26 VNB N_A4_c_258_n 0.0291497f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_27 VNB N_A4_c_259_n 0.0384045f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.16
cc_28 VNB N_Y_c_350_n 0.0069295f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_29 VNB N_Y_c_351_n 0.00829952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB Y 0.022997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_404_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_480_n 0.0129989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_481_n 0.0118776f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.985
cc_34 VNB N_VGND_c_482_n 0.00580922f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_35 VNB N_VGND_c_483_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_484_n 0.0865679f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_37 VNB N_VGND_c_485_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.16
cc_38 VNB N_VGND_c_486_n 0.0109937f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.16
cc_39 VNB N_VGND_c_487_n 0.0192923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_488_n 0.308768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_489_n 0.00545594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_317_47#_c_559_n 0.00209378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_317_47#_c_560_n 0.00295274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_567_47#_c_585_n 0.00667811f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.325
cc_45 VNB N_A_757_47#_c_604_n 0.00213317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_B1_M1006_g 0.0232539f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.985
cc_47 VPB N_B1_M1018_g 0.0186953f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.985
cc_48 VPB N_B1_c_79_n 0.0185114f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.16
cc_49 VPB N_A1_M1002_g 0.0186075f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=0.56
cc_50 VPB N_A1_M1019_g 0.0186099f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.985
cc_51 VPB N_A1_c_122_n 0.00421932f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.16
cc_52 VPB N_A2_M1010_g 0.0196968f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.325
cc_53 VPB N_A2_M1017_g 0.0199383f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_54 VPB N_A3_M1001_g 0.028274f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.56
cc_55 VPB N_A3_M1013_g 0.0280325f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_56 VPB N_A4_M1004_g 0.0196968f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.325
cc_57 VPB N_A4_M1009_g 0.0273582f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_58 VPB N_A4_c_259_n 0.013317f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.16
cc_59 VPB N_A_149_297#_c_293_n 0.00906529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_Y_c_353_n 0.0254464f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.16
cc_61 VPB N_Y_c_354_n 0.0148348f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.177
cc_62 VPB Y 0.00817771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_405_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_64 VPB N_VPWR_c_406_n 3.20298e-19 $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_65 VPB N_VPWR_c_407_n 0.00628023f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.16
cc_66 VPB N_VPWR_c_408_n 4.07719e-19 $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.16
cc_67 VPB N_VPWR_c_409_n 0.0157658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_410_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.177
cc_69 VPB N_VPWR_c_411_n 0.0538627f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.177
cc_70 VPB N_VPWR_c_412_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_413_n 0.0170387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_414_n 0.0200412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_404_n 0.0777827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_416_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_417_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_418_n 0.0128614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 N_B1_M1018_g N_A1_M1002_g 0.0143305f $X=1.5 $Y=1.985 $X2=0 $Y2=0
cc_78 N_B1_c_84_p N_A1_c_121_n 0.0134465f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B1_c_79_n N_A1_c_121_n 9.43542e-19 $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B1_c_84_p N_A1_c_122_n 2.44182e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B1_c_79_n N_A1_c_122_n 0.0352126f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B1_M1006_g N_A_149_297#_c_294_n 0.00937268f $X=1.08 $Y=1.985 $X2=0 $Y2=0
cc_83 N_B1_M1018_g N_A_149_297#_c_294_n 0.0112437f $X=1.5 $Y=1.985 $X2=0 $Y2=0
cc_84 N_B1_c_78_n N_Y_c_350_n 0.0141261f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B1_c_84_p N_Y_c_350_n 0.0331142f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B1_c_79_n N_Y_c_350_n 0.0138267f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B1_M1006_g N_Y_c_359_n 0.011421f $X=1.08 $Y=1.985 $X2=0 $Y2=0
cc_88 N_B1_M1018_g N_Y_c_359_n 0.00559427f $X=1.5 $Y=1.985 $X2=0 $Y2=0
cc_89 N_B1_c_77_n N_Y_c_361_n 0.0140556f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B1_c_84_p N_Y_c_361_n 0.00564987f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B1_c_84_p N_Y_c_363_n 0.00920238f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_92 N_B1_c_79_n N_Y_c_363_n 0.00217728f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B1_M1006_g N_Y_c_353_n 0.0124935f $X=1.08 $Y=1.985 $X2=0 $Y2=0
cc_94 N_B1_M1018_g N_Y_c_353_n 0.00354125f $X=1.5 $Y=1.985 $X2=0 $Y2=0
cc_95 N_B1_c_84_p N_Y_c_353_n 0.0667357f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B1_c_79_n N_Y_c_353_n 0.0165242f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B1_c_77_n Y 0.0168902f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B1_M1006_g Y 0.00258743f $X=1.08 $Y=1.985 $X2=0 $Y2=0
cc_99 N_B1_c_84_p Y 0.0129089f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B1_M1018_g N_VPWR_c_405_n 0.00110007f $X=1.5 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B1_M1006_g N_VPWR_c_411_n 0.00357877f $X=1.08 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B1_M1018_g N_VPWR_c_411_n 0.00357877f $X=1.5 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_M1006_g N_VPWR_c_404_n 0.00655123f $X=1.08 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B1_M1018_g N_VPWR_c_404_n 0.00525237f $X=1.5 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B1_c_77_n N_VGND_c_481_n 0.00775781f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B1_c_78_n N_VGND_c_481_n 5.08801e-19 $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_c_77_n N_VGND_c_482_n 5.10011e-19 $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B1_c_78_n N_VGND_c_482_n 0.00779688f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B1_c_77_n N_VGND_c_486_n 0.00340533f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B1_c_78_n N_VGND_c_486_n 0.00340533f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B1_c_77_n N_VGND_c_488_n 0.00396343f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B1_c_78_n N_VGND_c_488_n 0.00396343f $X=0.98 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A1_c_120_n N_A2_M1015_g 0.0262473f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A1_c_122_n N_A2_M1010_g 0.0297623f $X=2.34 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A1_c_121_n N_A2_c_166_n 0.0148685f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_c_122_n N_A2_c_166_n 2.59194e-19 $X=2.34 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A1_c_121_n N_A2_c_167_n 8.99392e-19 $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A1_c_122_n N_A2_c_167_n 0.0188157f $X=2.34 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A1_M1002_g N_A_149_297#_c_296_n 0.0140455f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A1_M1019_g N_A_149_297#_c_296_n 0.0144336f $X=2.34 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A1_c_121_n N_A_149_297#_c_296_n 0.0297787f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A1_c_122_n N_A_149_297#_c_296_n 0.00199384f $X=2.34 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A1_c_121_n N_A_149_297#_c_300_n 3.72838e-19 $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A1_c_119_n N_Y_c_350_n 0.0110418f $X=1.92 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A1_c_120_n N_Y_c_350_n 0.00265854f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A1_c_121_n N_Y_c_350_n 0.0213252f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A1_c_122_n N_Y_c_350_n 0.00320521f $X=2.34 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A1_M1002_g N_Y_c_353_n 4.60615e-19 $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A1_M1002_g N_VPWR_c_405_n 0.0114282f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A1_M1019_g N_VPWR_c_405_n 0.0102418f $X=2.34 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A1_M1019_g N_VPWR_c_406_n 6.0901e-19 $X=2.34 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A1_M1002_g N_VPWR_c_411_n 0.0046653f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A1_M1019_g N_VPWR_c_412_n 0.0046653f $X=2.34 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A1_M1002_g N_VPWR_c_404_n 0.007919f $X=1.92 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A1_M1019_g N_VPWR_c_404_n 0.007919f $X=2.34 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A1_c_119_n N_VGND_c_482_n 0.0030548f $X=1.92 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A1_c_119_n N_VGND_c_484_n 0.00366111f $X=1.92 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A1_c_120_n N_VGND_c_484_n 0.00366111f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_c_119_n N_VGND_c_488_n 0.00656615f $X=1.92 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_c_120_n N_VGND_c_488_n 0.00530732f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A1_c_119_n N_A_317_47#_c_559_n 0.00790826f $X=1.92 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_120_n N_A_317_47#_c_559_n 0.0109652f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_c_121_n N_A_317_47#_c_559_n 0.00335763f $X=2.29 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A2_M1017_g N_A3_M1001_g 0.0273833f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A2_c_166_n N_A3_c_209_n 7.97919e-19 $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A2_c_167_n N_A3_c_209_n 0.0185804f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A2_c_166_n A3 0.0178028f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_167_n A3 3.10946e-19 $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A2_M1010_g N_A_149_297#_c_301_n 0.0145283f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A2_M1017_g N_A_149_297#_c_301_n 0.0146468f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A2_c_166_n N_A_149_297#_c_301_n 0.0291326f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A2_c_167_n N_A_149_297#_c_301_n 0.00314431f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A2_M1017_g N_A_149_297#_c_305_n 0.00593237f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A2_c_166_n N_A_149_297#_c_306_n 0.00244642f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A2_c_167_n N_A_149_297#_c_306_n 2.17164e-19 $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A2_M1010_g N_VPWR_c_405_n 6.0901e-19 $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A2_M1010_g N_VPWR_c_406_n 0.0102418f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A2_M1017_g N_VPWR_c_406_n 0.0107671f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A2_M1010_g N_VPWR_c_412_n 0.0046653f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A2_M1017_g N_VPWR_c_413_n 0.0046653f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A2_M1010_g N_VPWR_c_404_n 0.007919f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A2_M1017_g N_VPWR_c_404_n 0.00796757f $X=3.18 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_M1015_g N_VGND_c_484_n 0.00414474f $X=2.76 $Y=0.56 $X2=0 $Y2=0
cc_164 N_A2_M1016_g N_VGND_c_484_n 0.00366111f $X=3.18 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A2_M1015_g N_VGND_c_488_n 0.00576602f $X=2.76 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A2_M1016_g N_VGND_c_488_n 0.00661716f $X=3.18 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A2_M1015_g N_A_317_47#_c_560_n 0.0100324f $X=2.76 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A2_M1016_g N_A_317_47#_c_560_n 0.00888921f $X=3.18 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A2_c_166_n N_A_317_47#_c_560_n 0.030352f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A2_c_167_n N_A_317_47#_c_560_n 0.00348263f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A2_M1015_g N_A_567_47#_c_585_n 0.00246655f $X=2.76 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A2_M1016_g N_A_567_47#_c_585_n 0.0100554f $X=3.18 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A3_M1012_g N_A4_M1003_g 0.0278108f $X=4.54 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A3_M1013_g N_A4_M1004_g 0.0295861f $X=4.54 $Y=1.985 $X2=0 $Y2=0
cc_175 A3 A4 0.0186079f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A3_c_212_n A4 0.00159327f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_177 A3 N_A4_c_258_n 2.18232e-19 $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A3_c_212_n N_A4_c_258_n 0.0187866f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A3_M1001_g N_A_149_297#_c_308_n 0.0175396f $X=3.62 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A3_M1013_g N_A_149_297#_c_308_n 0.0185325f $X=4.54 $Y=1.985 $X2=0 $Y2=0
cc_181 A3 N_A_149_297#_c_308_n 0.0526793f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A3_c_211_n N_A_149_297#_c_308_n 0.0131832f $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A3_M1001_g N_VPWR_c_406_n 6.50547e-19 $X=3.62 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A3_M1001_g N_VPWR_c_407_n 0.0172927f $X=3.62 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A3_M1013_g N_VPWR_c_407_n 0.0143821f $X=4.54 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A3_M1013_g N_VPWR_c_408_n 6.37932e-19 $X=4.54 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A3_M1013_g N_VPWR_c_409_n 0.00585385f $X=4.54 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A3_M1001_g N_VPWR_c_413_n 0.00585385f $X=3.62 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A3_M1001_g N_VPWR_c_404_n 0.0120907f $X=3.62 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A3_M1013_g N_VPWR_c_404_n 0.0119919f $X=4.54 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A3_M1012_g N_VGND_c_483_n 0.0018398f $X=4.54 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A3_M1005_g N_VGND_c_484_n 0.00366111f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A3_M1012_g N_VGND_c_484_n 0.00414474f $X=4.54 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A3_M1005_g N_VGND_c_488_n 0.00661716f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A3_M1012_g N_VGND_c_488_n 0.00576602f $X=4.54 $Y=0.56 $X2=0 $Y2=0
cc_196 N_A3_c_209_n N_A_317_47#_c_560_n 2.61353e-19 $X=3.695 $Y=1.16 $X2=0 $Y2=0
cc_197 A3 N_A_317_47#_c_560_n 5.30975e-19 $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_198 N_A3_M1005_g N_A_567_47#_c_585_n 0.0100554f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A3_M1012_g N_A_567_47#_c_585_n 0.0036428f $X=4.54 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A3_c_209_n N_A_567_47#_c_585_n 0.00397513f $X=3.695 $Y=1.16 $X2=0 $Y2=0
cc_201 A3 N_A_567_47#_c_585_n 0.00525016f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A3_M1005_g N_A_757_47#_c_604_n 0.00893883f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A3_M1012_g N_A_757_47#_c_604_n 0.0110926f $X=4.54 $Y=0.56 $X2=0 $Y2=0
cc_204 A3 N_A_757_47#_c_604_n 0.0377211f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_205 N_A3_c_211_n N_A_757_47#_c_604_n 0.00644521f $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A3_c_212_n N_A_757_47#_c_604_n 0.00193451f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A4_M1004_g N_A_149_297#_c_293_n 0.0144777f $X=4.96 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A4_M1009_g N_A_149_297#_c_293_n 0.0159719f $X=5.38 $Y=1.985 $X2=0 $Y2=0
cc_209 A4 N_A_149_297#_c_293_n 0.0450021f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_210 N_A4_c_258_n N_A_149_297#_c_293_n 0.0018492f $X=5.455 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A4_c_259_n N_A_149_297#_c_293_n 0.00553433f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_212 A4 N_A_149_297#_c_317_n 0.00496679f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_213 N_A4_M1004_g N_VPWR_c_408_n 0.0104049f $X=4.96 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A4_M1009_g N_VPWR_c_408_n 0.0121374f $X=5.38 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A4_M1004_g N_VPWR_c_409_n 0.0046653f $X=4.96 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A4_M1009_g N_VPWR_c_414_n 0.0046653f $X=5.38 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A4_M1004_g N_VPWR_c_404_n 0.007919f $X=4.96 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A4_M1009_g N_VPWR_c_404_n 0.00894942f $X=5.38 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A4_M1003_g N_VGND_c_483_n 0.0093539f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A4_M1007_g N_VGND_c_483_n 0.00835959f $X=5.38 $Y=0.56 $X2=0 $Y2=0
cc_221 N_A4_M1003_g N_VGND_c_484_n 0.00340533f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A4_M1007_g N_VGND_c_487_n 0.00340533f $X=5.38 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A4_M1003_g N_VGND_c_488_n 0.00403482f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A4_M1007_g N_VGND_c_488_n 0.00502106f $X=5.38 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A4_M1003_g N_A_567_47#_c_585_n 4.913e-19 $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A4_M1003_g N_A_757_47#_c_604_n 0.00997866f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A4_M1007_g N_A_757_47#_c_604_n 0.0132313f $X=5.38 $Y=0.56 $X2=0 $Y2=0
cc_228 A4 N_A_757_47#_c_604_n 0.04186f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_229 N_A4_c_258_n N_A_757_47#_c_604_n 0.0030539f $X=5.455 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A4_c_259_n N_A_757_47#_c_604_n 0.00388852f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_149_297#_c_294_n N_Y_M1006_s 0.00312348f $X=1.625 $Y=2.38 $X2=0 $Y2=0
cc_232 N_A_149_297#_c_294_n N_Y_c_359_n 0.0159307f $X=1.625 $Y=2.38 $X2=0 $Y2=0
cc_233 N_A_149_297#_M1006_d N_Y_c_353_n 0.00390196f $X=0.745 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_A_149_297#_c_321_p N_Y_c_353_n 0.0131641f $X=0.87 $Y=1.96 $X2=0 $Y2=0
cc_235 N_A_149_297#_c_294_n N_Y_c_353_n 0.00256303f $X=1.625 $Y=2.38 $X2=0 $Y2=0
cc_236 N_A_149_297#_c_296_n N_VPWR_M1002_d 0.00351266f $X=2.465 $Y=1.62
+ $X2=-0.19 $Y2=1.305
cc_237 N_A_149_297#_c_301_n N_VPWR_M1010_s 0.0035514f $X=3.325 $Y=1.62 $X2=0
+ $Y2=0
cc_238 N_A_149_297#_c_308_n N_VPWR_M1001_d 0.0180393f $X=4.665 $Y=1.62 $X2=0
+ $Y2=0
cc_239 N_A_149_297#_c_293_n N_VPWR_M1004_s 0.0035232f $X=5.505 $Y=1.62 $X2=0
+ $Y2=0
cc_240 N_A_149_297#_c_296_n N_VPWR_c_405_n 0.0145016f $X=2.465 $Y=1.62 $X2=0
+ $Y2=0
cc_241 N_A_149_297#_c_301_n N_VPWR_c_406_n 0.0145016f $X=3.325 $Y=1.62 $X2=0
+ $Y2=0
cc_242 N_A_149_297#_c_305_n N_VPWR_c_406_n 0.0372674f $X=3.41 $Y=1.96 $X2=0
+ $Y2=0
cc_243 N_A_149_297#_c_308_n N_VPWR_c_407_n 0.045327f $X=4.665 $Y=1.62 $X2=0
+ $Y2=0
cc_244 N_A_149_297#_c_293_n N_VPWR_c_408_n 0.0145016f $X=5.505 $Y=1.62 $X2=0
+ $Y2=0
cc_245 N_A_149_297#_c_332_p N_VPWR_c_409_n 0.0113958f $X=4.75 $Y=1.96 $X2=0
+ $Y2=0
cc_246 N_A_149_297#_c_294_n N_VPWR_c_411_n 0.0473059f $X=1.625 $Y=2.38 $X2=0
+ $Y2=0
cc_247 N_A_149_297#_c_334_p N_VPWR_c_411_n 0.0116982f $X=0.955 $Y=2.38 $X2=0
+ $Y2=0
cc_248 N_A_149_297#_c_335_p N_VPWR_c_412_n 0.0113958f $X=2.55 $Y=1.96 $X2=0
+ $Y2=0
cc_249 N_A_149_297#_c_305_n N_VPWR_c_413_n 0.0116048f $X=3.41 $Y=1.96 $X2=0
+ $Y2=0
cc_250 N_A_149_297#_c_337_p N_VPWR_c_414_n 0.0116048f $X=5.59 $Y=1.96 $X2=0
+ $Y2=0
cc_251 N_A_149_297#_M1006_d N_VPWR_c_404_n 0.00348186f $X=0.745 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_149_297#_M1018_d N_VPWR_c_404_n 0.00385313f $X=1.575 $Y=1.485 $X2=0
+ $Y2=0
cc_253 N_A_149_297#_M1019_s N_VPWR_c_404_n 0.00562358f $X=2.415 $Y=1.485 $X2=0
+ $Y2=0
cc_254 N_A_149_297#_M1017_d N_VPWR_c_404_n 0.00647849f $X=3.255 $Y=1.485 $X2=0
+ $Y2=0
cc_255 N_A_149_297#_M1013_s N_VPWR_c_404_n 0.00562358f $X=4.615 $Y=1.485 $X2=0
+ $Y2=0
cc_256 N_A_149_297#_M1009_d N_VPWR_c_404_n 0.00525232f $X=5.455 $Y=1.485 $X2=0
+ $Y2=0
cc_257 N_A_149_297#_c_294_n N_VPWR_c_404_n 0.0299894f $X=1.625 $Y=2.38 $X2=0
+ $Y2=0
cc_258 N_A_149_297#_c_334_p N_VPWR_c_404_n 0.00654447f $X=0.955 $Y=2.38 $X2=0
+ $Y2=0
cc_259 N_A_149_297#_c_335_p N_VPWR_c_404_n 0.00646998f $X=2.55 $Y=1.96 $X2=0
+ $Y2=0
cc_260 N_A_149_297#_c_305_n N_VPWR_c_404_n 0.00646998f $X=3.41 $Y=1.96 $X2=0
+ $Y2=0
cc_261 N_A_149_297#_c_332_p N_VPWR_c_404_n 0.00646998f $X=4.75 $Y=1.96 $X2=0
+ $Y2=0
cc_262 N_A_149_297#_c_337_p N_VPWR_c_404_n 0.00646998f $X=5.59 $Y=1.96 $X2=0
+ $Y2=0
cc_263 N_Y_M1006_s N_VPWR_c_404_n 0.00216833f $X=1.155 $Y=1.485 $X2=0 $Y2=0
cc_264 N_Y_c_361_n N_VGND_M1000_s 0.00335579f $X=0.685 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_265 N_Y_c_351_n N_VGND_M1000_s 0.00173515f $X=0.23 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_266 Y N_VGND_M1000_s 0.00110582f $X=0.23 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_267 N_Y_c_350_n N_VGND_M1014_s 0.00489262f $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_268 N_Y_c_351_n N_VGND_c_480_n 7.9782e-19 $X=0.23 $Y=0.815 $X2=0 $Y2=0
cc_269 N_Y_c_361_n N_VGND_c_481_n 0.0101191f $X=0.685 $Y=0.73 $X2=0 $Y2=0
cc_270 N_Y_c_351_n N_VGND_c_481_n 0.0104868f $X=0.23 $Y=0.815 $X2=0 $Y2=0
cc_271 N_Y_c_350_n N_VGND_c_482_n 0.021163f $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_272 N_Y_c_350_n N_VGND_c_484_n 0.00303246f $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_273 N_Y_c_392_p N_VGND_c_486_n 0.0112415f $X=0.77 $Y=0.42 $X2=0 $Y2=0
cc_274 N_Y_c_350_n N_VGND_c_486_n 0.00238578f $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_275 N_Y_c_361_n N_VGND_c_486_n 0.00238578f $X=0.685 $Y=0.73 $X2=0 $Y2=0
cc_276 N_Y_M1000_d N_VGND_c_488_n 0.00250764f $X=0.635 $Y=0.235 $X2=0 $Y2=0
cc_277 N_Y_M1008_s N_VGND_c_488_n 0.00219239f $X=1.995 $Y=0.235 $X2=0 $Y2=0
cc_278 N_Y_c_392_p N_VGND_c_488_n 0.00643744f $X=0.77 $Y=0.42 $X2=0 $Y2=0
cc_279 N_Y_c_350_n N_VGND_c_488_n 0.0119676f $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_280 N_Y_c_361_n N_VGND_c_488_n 0.00504221f $X=0.685 $Y=0.73 $X2=0 $Y2=0
cc_281 N_Y_c_351_n N_VGND_c_488_n 0.00189762f $X=0.23 $Y=0.815 $X2=0 $Y2=0
cc_282 N_Y_c_350_n N_A_317_47#_M1008_d 0.010508f $X=2.13 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_283 N_Y_M1008_s N_A_317_47#_c_559_n 0.003196f $X=1.995 $Y=0.235 $X2=0 $Y2=0
cc_284 N_Y_c_350_n N_A_317_47#_c_559_n 0.0372327f $X=2.13 $Y=0.73 $X2=0 $Y2=0
cc_285 N_VGND_c_488_n N_A_317_47#_M1008_d 0.00211652f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_286 N_VGND_c_488_n N_A_317_47#_M1011_d 0.00237695f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_488_n N_A_317_47#_M1016_d 0.00212464f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_288 N_VGND_c_482_n N_A_317_47#_c_559_n 0.014924f $X=1.19 $Y=0.38 $X2=0 $Y2=0
cc_289 N_VGND_c_484_n N_A_317_47#_c_559_n 0.0501343f $X=5.005 $Y=0 $X2=0 $Y2=0
cc_290 N_VGND_c_488_n N_A_317_47#_c_559_n 0.0383323f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_291 N_VGND_c_484_n N_A_317_47#_c_560_n 0.00238885f $X=5.005 $Y=0 $X2=0 $Y2=0
cc_292 N_VGND_c_488_n N_A_317_47#_c_560_n 0.00560614f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_293 N_VGND_c_488_n N_A_567_47#_M1015_s 0.00217615f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_294 N_VGND_c_488_n N_A_567_47#_M1005_s 0.00217615f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_295 N_VGND_c_483_n N_A_567_47#_c_585_n 0.00545039f $X=5.17 $Y=0.38 $X2=0
+ $Y2=0
cc_296 N_VGND_c_484_n N_A_567_47#_c_585_n 0.0775216f $X=5.005 $Y=0 $X2=0 $Y2=0
cc_297 N_VGND_c_488_n N_A_567_47#_c_585_n 0.0594678f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_298 N_VGND_c_488_n N_A_757_47#_M1005_d 0.00212464f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_299 N_VGND_c_488_n N_A_757_47#_M1012_d 0.00319211f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_300 N_VGND_c_488_n N_A_757_47#_M1007_d 0.00369435f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_M1003_s N_A_757_47#_c_604_n 0.00339267f $X=5.035 $Y=0.235 $X2=0
+ $Y2=0
cc_302 N_VGND_c_483_n N_A_757_47#_c_604_n 0.0152077f $X=5.17 $Y=0.38 $X2=0 $Y2=0
cc_303 N_VGND_c_484_n N_A_757_47#_c_604_n 0.00757283f $X=5.005 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_487_n N_A_757_47#_c_604_n 0.00238578f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_488_n N_A_757_47#_c_604_n 0.020203f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_487_n N_A_757_47#_c_623_n 0.0114446f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_488_n N_A_757_47#_c_623_n 0.00643744f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_308 N_A_317_47#_c_560_n N_A_567_47#_M1015_s 0.0033933f $X=3.39 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_309 N_A_317_47#_M1016_d N_A_567_47#_c_585_n 0.00501197f $X=3.255 $Y=0.235
+ $X2=0 $Y2=0
cc_310 N_A_317_47#_c_560_n N_A_567_47#_c_585_n 0.0372291f $X=3.39 $Y=0.73 $X2=0
+ $Y2=0
cc_311 N_A_317_47#_c_560_n N_A_757_47#_c_604_n 0.0145425f $X=3.39 $Y=0.73 $X2=0
+ $Y2=0
cc_312 N_A_567_47#_c_585_n N_A_757_47#_M1005_d 0.00482233f $X=4.33 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_313 N_A_567_47#_M1005_s N_A_757_47#_c_604_n 0.00339635f $X=4.195 $Y=0.235
+ $X2=0 $Y2=0
cc_314 N_A_567_47#_c_585_n N_A_757_47#_c_604_n 0.0372291f $X=4.33 $Y=0.38 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__o31a_4.spice
* Created: Tue Sep  1 19:25:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o31a_4.pex.spice"
.subckt sky130_fd_sc_hd__o31a_4  VNB VPB B1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_102_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_102_21#_M1007_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.0975 AS=0.08775 PD=0.95 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1007_d N_A_102_21#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.0975 AS=0.08775 PD=0.95 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_102_21#_M1010_g N_X_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1016 N_A_102_21#_M1016_d N_B1_M1016_g N_A_496_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1021 N_A_102_21#_M1016_d N_B1_M1021_g N_A_496_47#_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.10075 PD=0.92 PS=0.96 NRD=0 NRS=0.912 M=1 R=4.33333
+ SA=75000.6 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1012 N_A_496_47#_M1021_s N_A3_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.08775 PD=0.96 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1014 N_A_496_47#_M1014_d N_A3_M1014_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_496_47#_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_A_496_47#_M1004_d N_A1_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_A_496_47#_M1004_d N_A1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1005_s N_A2_M1013_g N_A_496_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_102_21#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1015 N_X_M1003_d N_A_102_21#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.15 PD=1.27 PS=1.3 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1022 N_X_M1022_d N_A_102_21#_M1022_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.15 PD=1.27 PS=1.3 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1023 N_X_M1022_d N_A_102_21#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1023_s N_B1_M1006_g N_A_102_21#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1018_d N_B1_M1018_g N_A_102_21#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.145 PD=2.56 PS=1.29 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_102_21#_M1000_d N_A3_M1000_g N_A_672_297#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1020 N_A_102_21#_M1000_d N_A3_M1020_g N_A_672_297#_M1020_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1011 N_A_926_297#_M1011_d N_A2_M1011_g N_A_672_297#_M1020_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_926_297#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1001_d N_A1_M1019_g N_A_926_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_A_926_297#_M1019_s N_A2_M1017_g N_A_672_297#_M1017_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.9461 P=16.85
c_68 VNB 0 2.30751e-19 $X=0.125 $Y=-0.085
*
.include "sky130_fd_sc_hd__o31a_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a22o_4.spice.pex
* Created: Thu Aug 27 14:02:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A22O_4%A_96_21# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 41 50 52 54 55 56 57 59 60 65 66 71 72 73 79 80 88
c166 79 0 1.20852e-19 $X=5.145 $Y=0.73
c167 73 0 1.24618e-19 $X=3.805 $Y=1.87
c168 66 0 1.24618e-19 $X=2.965 $Y=1.87
c169 55 0 1.50675e-19 $X=2.84 $Y=1.87
r170 85 86 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.975 $Y=1.16
+ $X2=1.395 $Y2=1.16
r171 79 80 10.6882 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=5.145 $Y=0.775
+ $X2=4.935 $Y2=0.775
r172 73 76 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.805 $Y=1.87
+ $X2=3.805 $Y2=1.96
r173 72 80 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.605 $Y=0.82
+ $X2=4.935 $Y2=0.82
r174 66 69 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.965 $Y=1.87
+ $X2=2.965 $Y2=1.96
r175 60 71 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.3 $Y=0.775
+ $X2=3.17 $Y2=0.775
r176 60 62 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.775
+ $X2=3.385 $Y2=0.775
r177 59 72 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.475 $Y=0.775
+ $X2=3.605 $Y2=0.775
r178 59 62 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=3.475 $Y=0.775
+ $X2=3.385 $Y2=0.775
r179 58 66 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=1.87
+ $X2=2.965 $Y2=1.87
r180 57 73 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.68 $Y=1.87
+ $X2=3.805 $Y2=1.87
r181 57 58 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.68 $Y=1.87
+ $X2=3.09 $Y2=1.87
r182 55 66 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.84 $Y=1.87
+ $X2=2.965 $Y2=1.87
r183 55 56 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.84 $Y=1.87
+ $X2=2.23 $Y2=1.87
r184 54 71 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.23 $Y=0.82
+ $X2=3.17 $Y2=0.82
r185 52 65 3.53812 $w=3.1e-07 $l=1.09545e-07 $layer=LI1_cond $X=2.085 $Y=1.075
+ $X2=2.065 $Y2=1.175
r186 51 54 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.085 $Y=0.905
+ $X2=2.23 $Y2=0.82
r187 51 52 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.085 $Y=0.905
+ $X2=2.085 $Y2=1.075
r188 50 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.065 $Y=1.785
+ $X2=2.23 $Y2=1.87
r189 49 65 3.53812 $w=3.1e-07 $l=1e-07 $layer=LI1_cond $X=2.065 $Y=1.275
+ $X2=2.065 $Y2=1.175
r190 49 50 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.065 $Y=1.275
+ $X2=2.065 $Y2=1.785
r191 48 88 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.725 $Y=1.16
+ $X2=1.815 $Y2=1.16
r192 48 86 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.725 $Y=1.16
+ $X2=1.395 $Y2=1.16
r193 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.725
+ $Y=1.16 $X2=1.725 $Y2=1.16
r194 44 85 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.705 $Y=1.16
+ $X2=0.975 $Y2=1.16
r195 44 82 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.705 $Y=1.16
+ $X2=0.555 $Y2=1.16
r196 43 47 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=1.725 $Y2=1.175
r197 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=1.16 $X2=0.705 $Y2=1.16
r198 41 65 2.95888 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=1.175
+ $X2=2.065 $Y2=1.175
r199 41 47 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=1.9 $Y=1.175
+ $X2=1.725 $Y2=1.175
r200 37 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.16
r201 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.985
r202 34 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=1.16
r203 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=0.56
r204 30 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.16
r205 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.395 $Y=1.325
+ $X2=1.395 $Y2=1.985
r206 27 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=1.16
r207 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=0.56
r208 23 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.16
r209 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.985
r210 20 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=1.16
r211 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=0.56
r212 16 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.325
+ $X2=0.555 $Y2=1.16
r213 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.555 $Y=1.325
+ $X2=0.555 $Y2=1.985
r214 13 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=1.16
r215 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=0.56
r216 4 76 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=1.485 $X2=3.805 $Y2=1.96
r217 3 69 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.485 $X2=2.965 $Y2=1.96
r218 2 79 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.235 $X2=5.145 $Y2=0.73
r219 1 62 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.235 $X2=3.385 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%B2 1 3 6 8 10 13 15 19 20 22 25 26
c85 26 0 1.81811e-19 $X=2.755 $Y=1.16
c86 25 0 2.75292e-19 $X=2.755 $Y=1.16
c87 20 0 2.52452e-19 $X=4.015 $Y=1.16
r88 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.16 $X2=2.755 $Y2=1.16
r89 22 32 7.60125 $w=5.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.687 $Y=1.19
+ $X2=2.687 $Y2=1.53
r90 22 26 0.670698 $w=5.33e-07 $l=3e-08 $layer=LI1_cond $X=2.687 $Y=1.19
+ $X2=2.687 $Y2=1.16
r91 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.015
+ $Y=1.16 $X2=4.015 $Y2=1.16
r92 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.015 $Y=1.445
+ $X2=4.015 $Y2=1.16
r93 16 32 7.58357 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=2.955 $Y=1.53
+ $X2=2.687 $Y2=1.53
r94 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.85 $Y=1.53
+ $X2=4.015 $Y2=1.445
r95 15 16 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.85 $Y=1.53
+ $X2=2.955 $Y2=1.53
r96 11 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=1.16
r97 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=1.985
r98 8 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=1.16
r99 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=0.56
r100 4 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.325
+ $X2=2.755 $Y2=1.16
r101 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.755 $Y=1.325
+ $X2=2.755 $Y2=1.985
r102 1 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=0.995
+ $X2=2.755 $Y2=1.16
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.755 $Y=0.995
+ $X2=2.755 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%B1 1 3 6 8 10 13 15 22
c43 6 0 1.81811e-19 $X=3.175 $Y=1.985
r44 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.385 $Y=1.16
+ $X2=3.595 $Y2=1.16
r45 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.175 $Y=1.16
+ $X2=3.385 $Y2=1.16
r46 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.16 $X2=3.385 $Y2=1.16
r47 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.325
+ $X2=3.595 $Y2=1.16
r48 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.595 $Y=1.325
+ $X2=3.595 $Y2=1.985
r49 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=0.995
+ $X2=3.595 $Y2=1.16
r50 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.595 $Y=0.995
+ $X2=3.595 $Y2=0.56
r51 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=1.325
+ $X2=3.175 $Y2=1.16
r52 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.175 $Y=1.325
+ $X2=3.175 $Y2=1.985
r53 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=0.995
+ $X2=3.175 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.175 $Y=0.995
+ $X2=3.175 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%A2 1 3 6 8 10 13 17 18 20 21 23 24 25 29 34
c85 29 0 1.50675e-19 $X=5.775 $Y=1.16
c86 18 0 2.78509e-19 $X=4.515 $Y=1.16
c87 8 0 1.20852e-19 $X=5.775 $Y=0.995
r88 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.775
+ $Y=1.16 $X2=5.775 $Y2=1.16
r89 25 34 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=6.21 $Y=1.175 $X2=6.23
+ $Y2=1.175
r90 25 30 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=6.21 $Y=1.175
+ $X2=5.775 $Y2=1.175
r91 24 30 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=5.735 $Y=1.175
+ $X2=5.775 $Y2=1.175
r92 22 24 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.65 $Y=1.275
+ $X2=5.735 $Y2=1.175
r93 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.65 $Y=1.275
+ $X2=5.65 $Y2=1.445
r94 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.565 $Y=1.53
+ $X2=5.65 $Y2=1.445
r95 20 21 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=5.565 $Y=1.53
+ $X2=4.68 $Y2=1.53
r96 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.515
+ $Y=1.16 $X2=4.515 $Y2=1.16
r97 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.515 $Y=1.445
+ $X2=4.68 $Y2=1.53
r98 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.515 $Y=1.445
+ $X2=4.515 $Y2=1.16
r99 11 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.775 $Y=1.325
+ $X2=5.775 $Y2=1.16
r100 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.775 $Y=1.325
+ $X2=5.775 $Y2=1.985
r101 8 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.775 $Y=0.995
+ $X2=5.775 $Y2=1.16
r102 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.775 $Y=0.995
+ $X2=5.775 $Y2=0.56
r103 4 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.515 $Y=1.325
+ $X2=4.515 $Y2=1.16
r104 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.515 $Y=1.325
+ $X2=4.515 $Y2=1.985
r105 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.515 $Y=0.995
+ $X2=4.515 $Y2=1.16
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.515 $Y=0.995
+ $X2=4.515 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%A1 1 3 6 8 10 13 15 22
c43 8 0 6.86556e-20 $X=5.355 $Y=0.995
r44 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.145 $Y=1.16
+ $X2=5.355 $Y2=1.16
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.145
+ $Y=1.16 $X2=5.145 $Y2=1.16
r46 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.935 $Y=1.16
+ $X2=5.145 $Y2=1.16
r47 15 21 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.31 $Y=1.175
+ $X2=5.145 $Y2=1.175
r48 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.355 $Y=1.325
+ $X2=5.355 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.355 $Y=1.325
+ $X2=5.355 $Y2=1.985
r50 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.355 $Y=0.995
+ $X2=5.355 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.355 $Y=0.995
+ $X2=5.355 $Y2=0.56
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.325
+ $X2=4.935 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.935 $Y=1.325
+ $X2=4.935 $Y2=1.985
r54 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=0.995
+ $X2=4.935 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.935 $Y=0.995
+ $X2=4.935 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 42 44 49 62 63 69 72
r97 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r98 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r99 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r100 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r101 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r102 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r103 57 73 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=2.07 $Y2=2.72
r104 56 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r105 54 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.15 $Y=2.72
+ $X2=2.025 $Y2=2.72
r106 54 56 144.834 $w=1.68e-07 $l=2.22e-06 $layer=LI1_cond $X=2.15 $Y=2.72
+ $X2=4.37 $Y2=2.72
r107 53 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r108 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r109 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r110 50 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.31 $Y=2.72
+ $X2=1.185 $Y2=2.72
r111 50 52 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.31 $Y=2.72 $X2=1.61
+ $Y2=2.72
r112 49 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.9 $Y=2.72
+ $X2=2.025 $Y2=2.72
r113 49 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.9 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 48 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r115 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r116 45 66 3.90382 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=0.235 $Y2=2.72
r117 45 47 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 44 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.06 $Y=2.72
+ $X2=1.185 $Y2=2.72
r119 44 47 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 42 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r122 40 59 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.44 $Y=2.72
+ $X2=5.29 $Y2=2.72
r123 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.44 $Y=2.72
+ $X2=5.565 $Y2=2.72
r124 39 62 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.69 $Y=2.72
+ $X2=6.21 $Y2=2.72
r125 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.69 $Y=2.72
+ $X2=5.565 $Y2=2.72
r126 37 56 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.6 $Y=2.72
+ $X2=4.37 $Y2=2.72
r127 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.6 $Y=2.72
+ $X2=4.725 $Y2=2.72
r128 36 59 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.85 $Y=2.72
+ $X2=5.29 $Y2=2.72
r129 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.85 $Y=2.72
+ $X2=4.725 $Y2=2.72
r130 32 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.635
+ $X2=5.565 $Y2=2.72
r131 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.565 $Y=2.635
+ $X2=5.565 $Y2=2.3
r132 28 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.725 $Y=2.635
+ $X2=4.725 $Y2=2.72
r133 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.725 $Y=2.635
+ $X2=4.725 $Y2=2.3
r134 24 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.635
+ $X2=2.025 $Y2=2.72
r135 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.025 $Y=2.635
+ $X2=2.025 $Y2=2.3
r136 20 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=2.72
r137 20 22 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.185 $Y=2.635
+ $X2=1.185 $Y2=1.99
r138 16 66 3.23934 $w=2.5e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.235 $Y2=2.72
r139 16 18 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.345 $Y2=1.99
r140 5 34 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.485 $X2=5.565 $Y2=2.3
r141 4 30 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=1.485 $X2=4.725 $Y2=2.3
r142 3 26 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.485 $X2=2.025 $Y2=2.3
r143 2 22 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=1.05
+ $Y=1.485 $X2=1.185 $Y2=1.99
r144 1 18 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=1.485 $X2=0.345 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43 44
+ 45
r71 42 45 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.227 $Y=1.445
+ $X2=0.227 $Y2=1.19
r72 41 45 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=0.227 $Y=0.905
+ $X2=0.227 $Y2=1.19
r73 37 39 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=1.62
+ $X2=1.605 $Y2=2.3
r74 35 37 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=1.615
+ $X2=1.605 $Y2=1.62
r75 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.605 $Y=0.725
+ $X2=1.605 $Y2=0.39
r76 30 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=0.815
+ $X2=0.765 $Y2=0.815
r77 29 31 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.44 $Y=0.815
+ $X2=1.605 $Y2=0.725
r78 29 30 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.44 $Y=0.815
+ $X2=0.93 $Y2=0.815
r79 28 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.89 $Y=1.53
+ $X2=0.765 $Y2=1.53
r80 27 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.48 $Y=1.53
+ $X2=1.605 $Y2=1.615
r81 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.48 $Y=1.53 $X2=0.89
+ $Y2=1.53
r82 23 25 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.765 $Y=1.62
+ $X2=0.765 $Y2=2.3
r83 21 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.615
+ $X2=0.765 $Y2=1.53
r84 21 23 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.765 $Y=1.615
+ $X2=0.765 $Y2=1.62
r85 17 43 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.765 $Y=0.725
+ $X2=0.765 $Y2=0.815
r86 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.765 $Y=0.725
+ $X2=0.765 $Y2=0.39
r87 16 42 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.37 $Y=1.53
+ $X2=0.227 $Y2=1.445
r88 15 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.64 $Y=1.53
+ $X2=0.765 $Y2=1.53
r89 15 16 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.64 $Y=1.53 $X2=0.37
+ $Y2=1.53
r90 14 41 7.27854 $w=1.8e-07 $l=1.82535e-07 $layer=LI1_cond $X=0.37 $Y=0.815
+ $X2=0.227 $Y2=0.905
r91 13 43 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=0.815
+ $X2=0.765 $Y2=0.815
r92 13 14 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.6 $Y=0.815
+ $X2=0.37 $Y2=0.815
r93 4 39 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.485 $X2=1.605 $Y2=2.3
r94 4 37 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.485 $X2=1.605 $Y2=1.62
r95 3 25 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.485 $X2=0.765 $Y2=2.3
r96 3 23 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.485 $X2=0.765 $Y2=1.62
r97 2 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.47
+ $Y=0.235 $X2=1.605 $Y2=0.39
r98 1 19 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.235 $X2=0.765 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%A_484_297# 1 2 3 4 5 16 18 24 25 28 30 34 38
+ 41 46 50
c59 30 0 1.50675e-19 $X=5.905 $Y=1.87
c60 25 0 2.55669e-19 $X=4.43 $Y=1.87
c61 24 0 1.50675e-19 $X=5.02 $Y=1.87
r62 46 48 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.385 $Y=2.3 $X2=3.385
+ $Y2=2.38
r63 41 43 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.545 $Y=2.3 $X2=2.545
+ $Y2=2.38
r64 36 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.007 $Y=1.955
+ $X2=6.007 $Y2=1.87
r65 36 38 0.27051 $w=2.03e-07 $l=5e-09 $layer=LI1_cond $X=6.007 $Y=1.955
+ $X2=6.007 $Y2=1.96
r66 32 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.007 $Y=1.785
+ $X2=6.007 $Y2=1.87
r67 32 34 8.92683 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=6.007 $Y=1.785
+ $X2=6.007 $Y2=1.62
r68 31 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.27 $Y=1.87
+ $X2=5.145 $Y2=1.87
r69 30 51 2.0246 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.905 $Y=1.87
+ $X2=6.007 $Y2=1.87
r70 30 31 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.905 $Y=1.87
+ $X2=5.27 $Y2=1.87
r71 26 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=1.955
+ $X2=5.145 $Y2=1.87
r72 26 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.145 $Y=1.955
+ $X2=5.145 $Y2=1.96
r73 24 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.02 $Y=1.87
+ $X2=5.145 $Y2=1.87
r74 24 25 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.02 $Y=1.87 $X2=4.43
+ $Y2=1.87
r75 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.265 $Y=2.295
+ $X2=4.265 $Y2=1.96
r76 20 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.265 $Y=1.955
+ $X2=4.43 $Y2=1.87
r77 20 23 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=4.265 $Y=1.955
+ $X2=4.265 $Y2=1.96
r78 19 48 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.51 $Y=2.38
+ $X2=3.385 $Y2=2.38
r79 18 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.1 $Y=2.38
+ $X2=4.265 $Y2=2.295
r80 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.1 $Y=2.38 $X2=3.51
+ $Y2=2.38
r81 17 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.67 $Y=2.38
+ $X2=2.545 $Y2=2.38
r82 16 48 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.26 $Y=2.38
+ $X2=3.385 $Y2=2.38
r83 16 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.26 $Y=2.38 $X2=2.67
+ $Y2=2.38
r84 5 38 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=5.85
+ $Y=1.485 $X2=5.99 $Y2=1.96
r85 5 34 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=5.85
+ $Y=1.485 $X2=5.99 $Y2=1.62
r86 4 28 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.01
+ $Y=1.485 $X2=5.145 $Y2=1.96
r87 3 23 300 $w=1.7e-07 $l=5.53512e-07 $layer=licon1_PDIFF $count=2 $X=4.09
+ $Y=1.485 $X2=4.26 $Y2=1.96
r88 2 46 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.25
+ $Y=1.485 $X2=3.385 $Y2=2.3
r89 1 41 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.485 $X2=2.545 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%VGND 1 2 3 4 5 18 20 21 24 28 32 35 36 38 39
+ 40 61 62 70 75 81
r95 80 81 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0.235
+ $X2=2.63 $Y2=0.235
r96 77 80 0.280331 $w=6.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.545 $Y2=0.235
r97 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r98 74 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r99 73 77 8.59681 $w=6.38e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.53 $Y2=0.235
r100 73 75 9.76276 $w=6.38e-07 $l=1.3e-07 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=1.94 $Y2=0.235
r101 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r102 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r103 65 68 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.345 $Y2=0
r104 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r105 59 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r106 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r107 56 59 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.75 $Y2=0
r108 55 58 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.75
+ $Y2=0
r109 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r110 53 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r111 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r112 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r113 50 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r114 49 52 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r115 49 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.63
+ $Y2=0
r116 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r117 46 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r118 46 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r119 45 75 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.94
+ $Y2=0
r120 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r121 43 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.185
+ $Y2=0
r122 43 45 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.61
+ $Y2=0
r123 40 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r124 40 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r125 38 58 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.9 $Y=0 $X2=5.75
+ $Y2=0
r126 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0 $X2=5.985
+ $Y2=0
r127 37 61 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.07 $Y=0 $X2=6.21
+ $Y2=0
r128 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=0 $X2=5.985
+ $Y2=0
r129 35 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=3.91 $Y2=0
r130 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.27
+ $Y2=0
r131 34 55 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.37
+ $Y2=0
r132 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.27
+ $Y2=0
r133 30 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=0.085
+ $X2=5.985 $Y2=0
r134 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.985 $Y=0.085
+ $X2=5.985 $Y2=0.39
r135 26 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r136 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.39
r137 22 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r138 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.39
r139 21 68 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.345
+ $Y2=0
r140 20 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0 $X2=1.185
+ $Y2=0
r141 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=0.43
+ $Y2=0
r142 16 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0
r143 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.39
r144 5 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.85
+ $Y=0.235 $X2=5.985 $Y2=0.39
r145 4 28 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.235 $X2=4.27 $Y2=0.39
r146 3 80 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=1.89
+ $Y=0.235 $X2=2.545 $Y2=0.39
r147 2 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.235 $X2=1.185 $Y2=0.39
r148 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.235 $X2=0.345 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%A_566_47# 1 2 11
r15 8 11 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=2.965 $Y=0.365
+ $X2=3.805 $Y2=0.365
r16 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.235 $X2=3.805 $Y2=0.39
r17 1 8 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.235 $X2=2.965 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_4%A_918_47# 1 2 7 11 13
c23 13 0 6.86556e-20 $X=5.565 $Y=0.73
r24 11 16 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=5.605 $Y=0.475
+ $X2=5.605 $Y2=0.365
r25 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.605 $Y=0.475
+ $X2=5.605 $Y2=0.73
r26 7 16 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.48 $Y=0.365
+ $X2=5.605 $Y2=0.365
r27 7 9 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=5.48 $Y=0.365
+ $X2=4.725 $Y2=0.365
r28 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.43
+ $Y=0.235 $X2=5.565 $Y2=0.39
r29 2 13 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.43
+ $Y=0.235 $X2=5.565 $Y2=0.73
r30 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.59
+ $Y=0.235 $X2=4.725 $Y2=0.39
.ends


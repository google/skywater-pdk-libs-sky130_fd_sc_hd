* File: sky130_fd_sc_hd__a2111oi_2.pxi.spice
* Created: Thu Aug 27 13:59:04 2020
* 
x_PM_SKY130_FD_SC_HD__A2111OI_2%C1 N_C1_c_85_n N_C1_M1014_g N_C1_M1001_g
+ N_C1_M1013_g N_C1_M1018_g N_C1_c_93_n N_C1_c_94_n N_C1_c_86_n N_C1_c_87_n C1
+ N_C1_c_89_n N_C1_c_90_n N_C1_c_98_n C1 PM_SKY130_FD_SC_HD__A2111OI_2%C1
x_PM_SKY130_FD_SC_HD__A2111OI_2%D1 N_D1_c_169_n N_D1_M1009_g N_D1_M1007_g
+ N_D1_c_170_n N_D1_M1017_g N_D1_M1002_g D1 N_D1_c_171_n N_D1_c_172_n
+ PM_SKY130_FD_SC_HD__A2111OI_2%D1
x_PM_SKY130_FD_SC_HD__A2111OI_2%B1 N_B1_M1005_g N_B1_c_220_n N_B1_M1003_g
+ N_B1_M1010_g N_B1_c_221_n N_B1_M1012_g B1 N_B1_c_228_n N_B1_c_222_n
+ PM_SKY130_FD_SC_HD__A2111OI_2%B1
x_PM_SKY130_FD_SC_HD__A2111OI_2%A1 N_A1_c_269_n N_A1_M1000_g N_A1_M1006_g
+ N_A1_M1015_g N_A1_M1011_g N_A1_c_270_n N_A1_c_271_n N_A1_c_272_n N_A1_c_280_n
+ N_A1_c_281_n A1 N_A1_c_273_n N_A1_c_274_n PM_SKY130_FD_SC_HD__A2111OI_2%A1
x_PM_SKY130_FD_SC_HD__A2111OI_2%A2 N_A2_c_344_n N_A2_M1019_g N_A2_M1008_g
+ N_A2_M1016_g N_A2_c_345_n N_A2_M1004_g A2 N_A2_c_346_n
+ PM_SKY130_FD_SC_HD__A2111OI_2%A2
x_PM_SKY130_FD_SC_HD__A2111OI_2%A_28_297# N_A_28_297#_M1001_d
+ N_A_28_297#_M1013_d N_A_28_297#_M1010_d N_A_28_297#_c_389_n
+ N_A_28_297#_c_395_n N_A_28_297#_c_390_n N_A_28_297#_c_402_n
+ N_A_28_297#_c_417_p PM_SKY130_FD_SC_HD__A2111OI_2%A_28_297#
x_PM_SKY130_FD_SC_HD__A2111OI_2%Y N_Y_M1014_d N_Y_M1009_s N_Y_M1018_d
+ N_Y_M1012_s N_Y_M1015_d N_Y_M1007_s N_Y_c_432_n N_Y_c_433_n N_Y_c_442_n
+ N_Y_c_445_n N_Y_c_451_n N_Y_c_452_n N_Y_c_456_n N_Y_c_457_n N_Y_c_475_n
+ N_Y_c_479_n N_Y_c_492_n N_Y_c_472_n N_Y_c_459_n N_Y_c_436_n N_Y_c_483_n
+ N_Y_c_434_n Y N_Y_c_438_n Y PM_SKY130_FD_SC_HD__A2111OI_2%Y
x_PM_SKY130_FD_SC_HD__A2111OI_2%A_467_297# N_A_467_297#_M1005_s
+ N_A_467_297#_M1006_d N_A_467_297#_M1008_s N_A_467_297#_M1011_d
+ N_A_467_297#_c_568_n N_A_467_297#_c_569_n N_A_467_297#_c_581_n
+ N_A_467_297#_c_609_p N_A_467_297#_c_584_n N_A_467_297#_c_570_n
+ N_A_467_297#_c_571_n N_A_467_297#_c_575_n N_A_467_297#_c_572_n
+ N_A_467_297#_c_590_n PM_SKY130_FD_SC_HD__A2111OI_2%A_467_297#
x_PM_SKY130_FD_SC_HD__A2111OI_2%VPWR N_VPWR_M1006_s N_VPWR_M1016_d
+ N_VPWR_c_627_n N_VPWR_c_628_n N_VPWR_c_629_n N_VPWR_c_630_n VPWR
+ N_VPWR_c_631_n N_VPWR_c_632_n N_VPWR_c_626_n N_VPWR_c_634_n
+ PM_SKY130_FD_SC_HD__A2111OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A2111OI_2%VGND N_VGND_M1014_s N_VGND_M1017_d
+ N_VGND_M1003_d N_VGND_M1019_s N_VGND_c_697_n N_VGND_c_698_n N_VGND_c_699_n
+ N_VGND_c_700_n N_VGND_c_701_n VGND N_VGND_c_702_n N_VGND_c_703_n
+ N_VGND_c_704_n N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n N_VGND_c_708_n
+ N_VGND_c_709_n N_VGND_c_710_n PM_SKY130_FD_SC_HD__A2111OI_2%VGND
cc_1 VNB N_C1_c_85_n 0.022077f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_2 VNB N_C1_c_86_n 0.0037005f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_3 VNB N_C1_c_87_n 0.0223517f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_4 VNB C1 3.75757e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.445
cc_5 VNB N_C1_c_89_n 0.0435065f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_6 VNB N_C1_c_90_n 0.0180289f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=0.995
cc_7 VNB N_D1_c_169_n 0.016201f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_8 VNB N_D1_c_170_n 0.0173848f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=1.325
cc_9 VNB N_D1_c_171_n 0.00206513f $X=-0.19 $Y=-0.24 $X2=1.707 $Y2=1.152
cc_10 VNB N_D1_c_172_n 0.034592f $X=-0.19 $Y=-0.24 $X2=1.707 $Y2=1.275
cc_11 VNB N_B1_c_220_n 0.017838f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.985
cc_12 VNB N_B1_c_221_n 0.0174003f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_13 VNB N_B1_c_222_n 0.0462487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_269_n 0.0186686f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_15 VNB N_A1_c_270_n 0.00254493f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.16
cc_16 VNB N_A1_c_271_n 0.0141872f $X=-0.19 $Y=-0.24 $X2=1.707 $Y2=1.275
cc_17 VNB N_A1_c_272_n 0.0300122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_c_273_n 0.0346418f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.16
cc_19 VNB N_A1_c_274_n 0.0222431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_344_n 0.0186611f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_21 VNB N_A2_c_345_n 0.0561117f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.995
cc_22 VNB N_A2_c_346_n 0.00234832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_432_n 0.00962673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_433_n 0.0133844f $X=-0.19 $Y=-0.24 $X2=1.707 $Y2=1.152
cc_25 VNB N_Y_c_434_n 0.0219444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB Y 0.00836469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_626_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_28 VNB N_VGND_c_697_n 4.08532e-19 $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.445
cc_29 VNB N_VGND_c_698_n 0.00437091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_699_n 0.016464f $X=-0.19 $Y=-0.24 $X2=1.707 $Y2=1.152
cc_31 VNB N_VGND_c_700_n 0.00504533f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_32 VNB N_VGND_c_701_n 0.00561423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_702_n 0.0153773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_703_n 0.013512f $X=-0.19 $Y=-0.24 $X2=1.81 $Y2=1.325
cc_35 VNB N_VGND_c_704_n 0.03462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_705_n 0.0305163f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_706_n 0.280387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_707_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_708_n 0.00630653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_709_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_710_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_C1_M1001_g 0.0231823f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_43 VPB N_C1_M1013_g 0.0188557f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.985
cc_44 VPB N_C1_c_93_n 0.00443496f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_45 VPB N_C1_c_94_n 0.00980426f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.562
cc_46 VPB N_C1_c_87_n 0.00690834f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_47 VPB C1 0.00135737f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.445
cc_48 VPB N_C1_c_89_n 0.0108944f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.16
cc_49 VPB N_C1_c_98_n 0.00869034f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.562
cc_50 VPB N_D1_M1007_g 0.0185909f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_51 VPB N_D1_M1002_g 0.0185899f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_52 VPB N_D1_c_172_n 0.00606292f $X=-0.19 $Y=1.305 $X2=1.707 $Y2=1.275
cc_53 VPB N_B1_M1005_g 0.0190232f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=0.56
cc_54 VPB N_B1_M1010_g 0.0223279f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.985
cc_55 VPB N_B1_c_222_n 0.0107364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A1_M1006_g 0.0229337f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_57 VPB N_A1_M1011_g 0.023371f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_58 VPB N_A1_c_270_n 0.0011856f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_59 VPB N_A1_c_271_n 0.00529561f $X=-0.19 $Y=1.305 $X2=1.707 $Y2=1.275
cc_60 VPB N_A1_c_272_n 0.00675287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A1_c_280_n 3.32596e-19 $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_62 VPB N_A1_c_281_n 0.0120374f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_63 VPB N_A1_c_273_n 0.0109269f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_64 VPB N_A2_M1008_g 0.0183579f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_65 VPB N_A2_M1016_g 0.0187917f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.985
cc_66 VPB N_A2_c_345_n 0.00790452f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.995
cc_67 VPB N_A_28_297#_c_389_n 0.0168703f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.995
cc_68 VPB N_A_28_297#_c_390_n 0.00830264f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.445
cc_69 VPB N_Y_c_436_n 0.00262475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB Y 0.00847791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_Y_c_438_n 0.00508259f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_467_297#_c_568_n 0.0038642f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_73 VPB N_A_467_297#_c_569_n 0.0058696f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_74 VPB N_A_467_297#_c_570_n 0.0115466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_467_297#_c_571_n 0.0137698f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_467_297#_c_572_n 0.00503203f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=0.995
cc_77 VPB N_VPWR_c_627_n 4.02668e-19 $X=-0.19 $Y=1.305 $X2=1.79 $Y2=1.985
cc_78 VPB N_VPWR_c_628_n 4.02668e-19 $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_79 VPB N_VPWR_c_629_n 0.0118152f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_80 VPB N_VPWR_c_630_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_81 VPB N_VPWR_c_631_n 0.0858071f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.562
cc_82 VPB N_VPWR_c_632_n 0.0169463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_626_n 0.0488908f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.16
cc_84 VPB N_VPWR_c_634_n 0.00436029f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=0.995
cc_85 N_C1_c_85_n N_D1_c_169_n 0.0262916f $X=0.5 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_86 N_C1_M1001_g N_D1_M1007_g 0.058711f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_87 N_C1_c_93_n N_D1_M1007_g 5.82991e-19 $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_88 N_C1_c_98_n N_D1_M1007_g 0.0135738f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_89 N_C1_c_90_n N_D1_c_170_n 0.0183741f $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C1_M1013_g N_D1_M1002_g 0.0596244f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_91 N_C1_c_98_n N_D1_M1002_g 0.0130954f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_92 N_C1_c_93_n N_D1_c_171_n 0.0109239f $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_93 N_C1_c_86_n N_D1_c_171_n 0.0154251f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_94 N_C1_c_87_n N_D1_c_171_n 2.28589e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_95 N_C1_c_89_n N_D1_c_171_n 0.00161792f $X=0.5 $Y=1.16 $X2=0 $Y2=0
cc_96 N_C1_c_98_n N_D1_c_171_n 0.0487509f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_97 N_C1_c_93_n N_D1_c_172_n 6.75681e-19 $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_98 N_C1_c_86_n N_D1_c_172_n 0.00233451f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_99 N_C1_c_87_n N_D1_c_172_n 0.0221936f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_100 C1 N_D1_c_172_n 0.003522f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_101 N_C1_c_89_n N_D1_c_172_n 0.0228162f $X=0.5 $Y=1.16 $X2=0 $Y2=0
cc_102 N_C1_c_98_n N_D1_c_172_n 0.00407476f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_103 N_C1_M1013_g N_B1_M1005_g 0.0340456f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_104 N_C1_c_90_n N_B1_c_220_n 0.0103831f $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C1_c_86_n N_B1_c_228_n 0.0164523f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_106 N_C1_c_87_n N_B1_c_228_n 3.04216e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_107 N_C1_c_86_n N_B1_c_222_n 9.82276e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_108 N_C1_c_87_n N_B1_c_222_n 0.0228177f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_109 C1 N_B1_c_222_n 9.05002e-19 $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_110 N_C1_c_94_n N_A_28_297#_M1001_d 0.00365777f $X=0.455 $Y=1.562 $X2=-0.19
+ $Y2=-0.24
cc_111 N_C1_M1001_g N_A_28_297#_c_389_n 0.00755431f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_112 N_C1_c_94_n N_A_28_297#_c_389_n 0.0221169f $X=0.455 $Y=1.562 $X2=0 $Y2=0
cc_113 N_C1_c_89_n N_A_28_297#_c_389_n 0.00102472f $X=0.5 $Y=1.16 $X2=0 $Y2=0
cc_114 N_C1_M1001_g N_A_28_297#_c_395_n 0.0083072f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_115 N_C1_M1013_g N_A_28_297#_c_395_n 0.00815006f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_116 N_C1_c_98_n N_A_28_297#_c_395_n 0.00885661f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_117 N_C1_M1001_g N_A_28_297#_c_390_n 8.91003e-19 $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_118 N_C1_c_98_n A_115_297# 0.00332787f $X=1.615 $Y=1.562 $X2=-0.19 $Y2=-0.24
cc_119 N_C1_c_98_n N_Y_M1007_s 0.00178666f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_120 N_C1_c_93_n N_Y_c_432_n 0.0188083f $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C1_c_89_n N_Y_c_432_n 0.0061482f $X=0.5 $Y=1.16 $X2=0 $Y2=0
cc_122 N_C1_c_85_n N_Y_c_442_n 0.0126933f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_123 N_C1_c_93_n N_Y_c_442_n 0.0035829f $X=0.29 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C1_c_98_n N_Y_c_442_n 0.00777808f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_125 N_C1_M1001_g N_Y_c_445_n 8.83703e-19 $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C1_M1013_g N_Y_c_445_n 0.0142794f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_127 N_C1_c_86_n N_Y_c_445_n 0.00385267f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_128 N_C1_c_87_n N_Y_c_445_n 0.00209598f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_129 C1 N_Y_c_445_n 0.00980769f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_130 N_C1_c_98_n N_Y_c_445_n 0.0403401f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_131 N_C1_c_90_n N_Y_c_451_n 2.99967e-19 $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_132 N_C1_c_86_n N_Y_c_452_n 0.0219158f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_133 N_C1_c_87_n N_Y_c_452_n 0.00448883f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_134 N_C1_c_90_n N_Y_c_452_n 0.0115254f $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_135 N_C1_c_98_n N_Y_c_452_n 0.00501729f $X=1.615 $Y=1.562 $X2=0 $Y2=0
cc_136 N_C1_c_90_n N_Y_c_456_n 0.0050662f $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_137 N_C1_M1013_g N_Y_c_457_n 0.0042407f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_138 C1 N_Y_c_457_n 0.00428644f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_139 N_C1_c_86_n N_Y_c_459_n 6.83854e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_140 N_C1_M1013_g N_Y_c_436_n 0.00139311f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_141 N_C1_c_86_n N_Y_c_436_n 4.12181e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_142 C1 N_Y_c_436_n 0.0158024f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_143 C1 A_287_297# 4.58617e-19 $X=1.525 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_144 N_C1_c_98_n A_287_297# 0.00131309f $X=1.615 $Y=1.562 $X2=-0.19 $Y2=-0.24
cc_145 N_C1_M1001_g N_VPWR_c_631_n 0.00357828f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_146 N_C1_M1013_g N_VPWR_c_631_n 0.00357877f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_147 N_C1_M1001_g N_VPWR_c_626_n 0.00626064f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_148 N_C1_M1013_g N_VPWR_c_626_n 0.00542429f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_149 N_C1_c_85_n N_VGND_c_697_n 0.00785369f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_150 N_C1_c_90_n N_VGND_c_698_n 0.00181538f $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C1_c_90_n N_VGND_c_699_n 0.00419334f $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_152 N_C1_c_85_n N_VGND_c_702_n 0.00351072f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_153 N_C1_c_85_n N_VGND_c_706_n 0.00502853f $X=0.5 $Y=0.995 $X2=0 $Y2=0
cc_154 N_C1_c_90_n N_VGND_c_706_n 0.00597828f $X=1.81 $Y=0.995 $X2=0 $Y2=0
cc_155 N_D1_M1007_g N_A_28_297#_c_389_n 0.00152045f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_156 N_D1_M1007_g N_A_28_297#_c_395_n 0.0110596f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_157 N_D1_M1002_g N_A_28_297#_c_395_n 0.0104494f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_158 N_D1_c_169_n N_Y_c_442_n 0.011376f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_159 N_D1_c_171_n N_Y_c_442_n 0.013631f $X=1.26 $Y=1.16 $X2=0 $Y2=0
cc_160 N_D1_c_172_n N_Y_c_442_n 0.00148879f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_161 N_D1_M1007_g N_Y_c_445_n 0.00832762f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_162 N_D1_M1002_g N_Y_c_445_n 0.0106262f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_163 N_D1_c_170_n N_Y_c_451_n 0.0050662f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_164 N_D1_c_170_n N_Y_c_452_n 0.0118882f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_165 N_D1_c_171_n N_Y_c_452_n 0.00714467f $X=1.26 $Y=1.16 $X2=0 $Y2=0
cc_166 N_D1_c_170_n N_Y_c_456_n 2.9878e-19 $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_167 N_D1_c_170_n N_Y_c_472_n 3.30347e-19 $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_168 N_D1_c_171_n N_Y_c_472_n 0.0128296f $X=1.26 $Y=1.16 $X2=0 $Y2=0
cc_169 N_D1_c_172_n N_Y_c_472_n 0.00246912f $X=1.36 $Y=1.16 $X2=0 $Y2=0
cc_170 N_D1_M1007_g N_VPWR_c_631_n 0.00357877f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_171 N_D1_M1002_g N_VPWR_c_631_n 0.00357877f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_172 N_D1_M1007_g N_VPWR_c_626_n 0.00534514f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_173 N_D1_M1002_g N_VPWR_c_626_n 0.00534514f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_174 N_D1_c_169_n N_VGND_c_697_n 0.00634459f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_175 N_D1_c_170_n N_VGND_c_697_n 4.66587e-19 $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_176 N_D1_c_170_n N_VGND_c_698_n 0.00170614f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_177 N_D1_c_169_n N_VGND_c_703_n 0.00351072f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_178 N_D1_c_170_n N_VGND_c_703_n 0.00419334f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_179 N_D1_c_169_n N_VGND_c_706_n 0.0040731f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_180 N_D1_c_170_n N_VGND_c_706_n 0.005848f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B1_c_221_n N_A1_c_269_n 0.0122004f $X=2.915 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_182 N_B1_M1010_g N_A1_c_280_n 0.00176157f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_c_222_n N_A1_c_273_n 0.0122004f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_184 N_B1_M1005_g N_A_28_297#_c_402_n 0.00959945f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_M1010_g N_A_28_297#_c_402_n 0.00847184f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_c_220_n N_Y_c_475_n 0.0121925f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_c_221_n N_Y_c_475_n 0.0118361f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_228_n N_Y_c_475_n 0.0341506f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B1_c_222_n N_Y_c_475_n 0.00573899f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B1_c_220_n N_Y_c_479_n 3.03663e-19 $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B1_c_221_n N_Y_c_479_n 0.00537883f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B1_c_228_n N_Y_c_459_n 0.00604885f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B1_c_222_n N_Y_c_459_n 0.00291437f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B1_c_221_n N_Y_c_483_n 0.0010812f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B1_M1010_g Y 0.00383456f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B1_c_221_n Y 0.00749037f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B1_c_228_n Y 0.0198946f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B1_M1005_g N_Y_c_438_n 0.0123956f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B1_M1010_g N_Y_c_438_n 0.0126795f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B1_c_228_n N_Y_c_438_n 0.0484304f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B1_c_222_n N_Y_c_438_n 0.00974323f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_M1010_g N_A_467_297#_c_568_n 0.0110892f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B1_M1010_g N_A_467_297#_c_569_n 0.00105011f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_B1_M1005_g N_A_467_297#_c_575_n 0.00337819f $X=2.26 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_B1_M1010_g N_A_467_297#_c_575_n 0.00341091f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_B1_M1010_g N_A_467_297#_c_572_n 0.00292952f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_B1_M1005_g N_VPWR_c_631_n 0.00357877f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_M1010_g N_VPWR_c_631_n 0.00357877f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1005_g N_VPWR_c_626_n 0.00539798f $X=2.26 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_M1010_g N_VPWR_c_626_n 0.00656955f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_c_220_n N_VGND_c_699_n 0.00422112f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_c_220_n N_VGND_c_700_n 0.00188851f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_c_221_n N_VGND_c_700_n 0.00427574f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B1_c_221_n N_VGND_c_704_n 0.00413555f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B1_c_220_n N_VGND_c_706_n 0.00597519f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_221_n N_VGND_c_706_n 0.00590023f $X=2.915 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A1_c_269_n N_A2_c_344_n 0.0198188f $X=3.345 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A1_c_270_n N_A2_c_344_n 2.29569e-19 $X=3.55 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_219 N_A1_M1006_g N_A2_M1008_g 0.0441679f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A1_c_270_n N_A2_M1008_g 7.4519e-19 $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A1_c_281_n N_A2_M1008_g 0.0127584f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_222 N_A1_M1011_g N_A2_M1016_g 0.0378814f $X=4.97 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A1_c_271_n N_A2_M1016_g 7.18528e-19 $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A1_c_281_n N_A2_M1016_g 0.0130084f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_225 N_A1_c_270_n N_A2_c_345_n 0.00166459f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A1_c_271_n N_A2_c_345_n 8.32748e-19 $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A1_c_281_n N_A2_c_345_n 0.00591476f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_228 N_A1_c_273_n N_A2_c_345_n 0.0177289f $X=3.64 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A1_c_274_n N_A2_c_345_n 0.0627816f $X=5.06 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A1_c_270_n N_A2_c_346_n 0.0146466f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A1_c_271_n N_A2_c_346_n 0.022102f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A1_c_272_n N_A2_c_346_n 0.00159562f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A1_c_281_n N_A2_c_346_n 0.0561855f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_234 N_A1_c_273_n N_A2_c_346_n 0.0010332f $X=3.64 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A1_c_269_n N_Y_c_479_n 0.00778295f $X=3.345 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A1_c_269_n N_Y_c_492_n 0.0136994f $X=3.345 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A1_c_270_n N_Y_c_492_n 0.0195568f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A1_c_271_n N_Y_c_492_n 0.00870266f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A1_c_281_n N_Y_c_492_n 0.0109197f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_240 N_A1_c_273_n N_Y_c_492_n 0.00165483f $X=3.64 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A1_c_274_n N_Y_c_492_n 0.00958675f $X=5.06 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A1_c_269_n N_Y_c_483_n 0.00152448f $X=3.345 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A1_c_271_n N_Y_c_434_n 0.018942f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A1_c_272_n N_Y_c_434_n 0.00119026f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A1_c_274_n N_Y_c_434_n 0.00739389f $X=5.06 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A1_c_269_n Y 0.0059507f $X=3.345 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A1_M1006_g Y 0.00179111f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A1_c_270_n Y 0.0300505f $X=3.55 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A1_c_280_n Y 0.0142595f $X=3.715 $Y=1.56 $X2=0 $Y2=0
cc_250 N_A1_c_280_n N_A_467_297#_M1006_d 0.00310617f $X=3.715 $Y=1.56 $X2=0
+ $Y2=0
cc_251 N_A1_c_281_n N_A_467_297#_M1008_s 0.00178113f $X=4.895 $Y=1.56 $X2=0
+ $Y2=0
cc_252 N_A1_c_281_n N_A_467_297#_M1011_d 0.011252f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_253 N_A1_M1006_g N_A_467_297#_c_581_n 0.0115524f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A1_c_280_n N_A_467_297#_c_581_n 0.0116377f $X=3.715 $Y=1.56 $X2=0 $Y2=0
cc_255 N_A1_c_281_n N_A_467_297#_c_581_n 0.0233782f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_256 N_A1_M1011_g N_A_467_297#_c_584_n 0.0122425f $X=4.97 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A1_c_281_n N_A_467_297#_c_584_n 0.0381722f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_258 N_A1_c_272_n N_A_467_297#_c_570_n 5.30976e-19 $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A1_c_281_n N_A_467_297#_c_570_n 0.0168351f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_260 N_A1_c_280_n N_A_467_297#_c_572_n 0.00385468f $X=3.715 $Y=1.56 $X2=0
+ $Y2=0
cc_261 N_A1_c_273_n N_A_467_297#_c_572_n 0.00663912f $X=3.64 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A1_c_281_n N_A_467_297#_c_590_n 0.0136847f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_263 N_A1_c_281_n N_VPWR_M1006_s 0.00178548f $X=4.895 $Y=1.56 $X2=-0.19
+ $Y2=-0.24
cc_264 N_A1_c_281_n N_VPWR_M1016_d 0.00221571f $X=4.895 $Y=1.56 $X2=0 $Y2=0
cc_265 N_A1_M1006_g N_VPWR_c_627_n 0.00786361f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A1_M1011_g N_VPWR_c_628_n 0.00676393f $X=4.97 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A1_M1006_g N_VPWR_c_631_n 0.0035231f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A1_M1011_g N_VPWR_c_632_n 0.00407353f $X=4.97 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A1_M1006_g N_VPWR_c_626_n 0.00539272f $X=3.64 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A1_M1011_g N_VPWR_c_626_n 0.00563351f $X=4.97 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A1_c_269_n N_VGND_c_704_n 0.00413555f $X=3.345 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A1_c_274_n N_VGND_c_705_n 0.00414208f $X=5.06 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A1_c_269_n N_VGND_c_706_n 0.00633119f $X=3.345 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A1_c_274_n N_VGND_c_706_n 0.00676537f $X=5.06 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_c_344_n N_Y_c_479_n 0.00144014f $X=4.045 $Y=0.99 $X2=0 $Y2=0
cc_276 N_A2_c_344_n N_Y_c_492_n 0.0144173f $X=4.045 $Y=0.99 $X2=0 $Y2=0
cc_277 N_A2_c_345_n N_Y_c_492_n 0.0185587f $X=4.54 $Y=0.99 $X2=0 $Y2=0
cc_278 N_A2_c_346_n N_Y_c_492_n 0.0409856f $X=4.52 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A2_c_345_n N_Y_c_434_n 0.0013673f $X=4.54 $Y=0.99 $X2=0 $Y2=0
cc_280 N_A2_M1008_g N_A_467_297#_c_581_n 0.0115866f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A2_M1016_g N_A_467_297#_c_584_n 0.0122627f $X=4.5 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A2_M1008_g N_VPWR_c_627_n 0.00627551f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A2_M1016_g N_VPWR_c_627_n 5.06577e-19 $X=4.5 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A2_M1008_g N_VPWR_c_628_n 4.81945e-19 $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A2_M1016_g N_VPWR_c_628_n 0.00519775f $X=4.5 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A2_M1008_g N_VPWR_c_629_n 0.0035231f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A2_M1016_g N_VPWR_c_629_n 0.00407353f $X=4.5 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A2_M1008_g N_VPWR_c_626_n 0.00409303f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A2_M1016_g N_VPWR_c_626_n 0.0046373f $X=4.5 $Y=1.985 $X2=0 $Y2=0
cc_290 N_A2_c_344_n N_VGND_c_701_n 0.00326182f $X=4.045 $Y=0.99 $X2=0 $Y2=0
cc_291 N_A2_c_345_n N_VGND_c_701_n 0.00323006f $X=4.54 $Y=0.99 $X2=0 $Y2=0
cc_292 N_A2_c_344_n N_VGND_c_704_n 0.00422112f $X=4.045 $Y=0.99 $X2=0 $Y2=0
cc_293 N_A2_c_345_n N_VGND_c_705_n 0.00422112f $X=4.54 $Y=0.99 $X2=0 $Y2=0
cc_294 N_A2_c_344_n N_VGND_c_706_n 0.00632851f $X=4.045 $Y=0.99 $X2=0 $Y2=0
cc_295 N_A2_c_345_n N_VGND_c_706_n 0.00580292f $X=4.54 $Y=0.99 $X2=0 $Y2=0
cc_296 N_A_28_297#_c_395_n A_115_297# 0.00486744f $X=2.09 $Y=2.37 $X2=-0.19
+ $Y2=1.305
cc_297 N_A_28_297#_c_395_n N_Y_M1007_s 0.00333945f $X=2.09 $Y=2.37 $X2=0 $Y2=0
cc_298 N_A_28_297#_M1013_d N_Y_c_445_n 0.00411626f $X=1.865 $Y=1.485 $X2=0 $Y2=0
cc_299 N_A_28_297#_c_389_n N_Y_c_445_n 0.00868085f $X=0.285 $Y=2.02 $X2=0 $Y2=0
cc_300 N_A_28_297#_c_395_n N_Y_c_445_n 0.0660674f $X=2.09 $Y=2.37 $X2=0 $Y2=0
cc_301 N_A_28_297#_M1013_d N_Y_c_457_n 0.002593f $X=1.865 $Y=1.485 $X2=0 $Y2=0
cc_302 N_A_28_297#_M1013_d N_Y_c_436_n 0.00138807f $X=1.865 $Y=1.485 $X2=0 $Y2=0
cc_303 N_A_28_297#_M1010_d N_Y_c_438_n 0.00276414f $X=2.765 $Y=1.485 $X2=0 $Y2=0
cc_304 N_A_28_297#_c_402_n N_Y_c_438_n 0.00273666f $X=2.815 $Y=2.38 $X2=0 $Y2=0
cc_305 N_A_28_297#_c_395_n A_287_297# 0.00333945f $X=2.09 $Y=2.37 $X2=-0.19
+ $Y2=1.305
cc_306 N_A_28_297#_c_402_n N_A_467_297#_M1005_s 0.00359552f $X=2.815 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_307 N_A_28_297#_M1010_d N_A_467_297#_c_568_n 0.00518878f $X=2.765 $Y=1.485
+ $X2=0 $Y2=0
cc_308 N_A_28_297#_c_402_n N_A_467_297#_c_568_n 0.00434673f $X=2.815 $Y=2.38
+ $X2=0 $Y2=0
cc_309 N_A_28_297#_c_417_p N_A_467_297#_c_568_n 0.0120509f $X=2.9 $Y=2.3 $X2=0
+ $Y2=0
cc_310 N_A_28_297#_c_417_p N_A_467_297#_c_569_n 0.0259343f $X=2.9 $Y=2.3 $X2=0
+ $Y2=0
cc_311 N_A_28_297#_c_402_n N_A_467_297#_c_575_n 0.0112705f $X=2.815 $Y=2.38
+ $X2=0 $Y2=0
cc_312 N_A_28_297#_c_395_n N_VPWR_c_631_n 0.130684f $X=2.09 $Y=2.37 $X2=0 $Y2=0
cc_313 N_A_28_297#_c_390_n N_VPWR_c_631_n 0.0230714f $X=0.46 $Y=2.37 $X2=0 $Y2=0
cc_314 N_A_28_297#_c_417_p N_VPWR_c_631_n 0.0110309f $X=2.9 $Y=2.3 $X2=0 $Y2=0
cc_315 N_A_28_297#_M1001_d N_VPWR_c_626_n 0.00229814f $X=0.14 $Y=1.485 $X2=0
+ $Y2=0
cc_316 N_A_28_297#_M1013_d N_VPWR_c_626_n 0.00255381f $X=1.865 $Y=1.485 $X2=0
+ $Y2=0
cc_317 N_A_28_297#_M1010_d N_VPWR_c_626_n 0.0023074f $X=2.765 $Y=1.485 $X2=0
+ $Y2=0
cc_318 N_A_28_297#_c_395_n N_VPWR_c_626_n 0.0837084f $X=2.09 $Y=2.37 $X2=0 $Y2=0
cc_319 N_A_28_297#_c_390_n N_VPWR_c_626_n 0.0135841f $X=0.46 $Y=2.37 $X2=0 $Y2=0
cc_320 N_A_28_297#_c_417_p N_VPWR_c_626_n 0.0063548f $X=2.9 $Y=2.3 $X2=0 $Y2=0
cc_321 A_115_297# N_VPWR_c_626_n 0.00224864f $X=0.575 $Y=1.485 $X2=0.5 $Y2=1.16
cc_322 N_Y_c_445_n A_287_297# 0.00349173f $X=1.97 $Y=1.977 $X2=-0.19 $Y2=-0.24
cc_323 N_Y_c_438_n N_A_467_297#_M1005_s 0.00176773f $X=3.025 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_324 Y N_A_467_297#_c_568_n 0.0108576f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_325 N_Y_c_438_n N_A_467_297#_c_568_n 0.0232814f $X=3.025 $Y=1.535 $X2=0 $Y2=0
cc_326 N_Y_c_438_n N_A_467_297#_c_575_n 0.0159136f $X=3.025 $Y=1.535 $X2=0 $Y2=0
cc_327 Y N_A_467_297#_c_572_n 0.00931259f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_328 N_Y_M1007_s N_VPWR_c_626_n 0.00224864f $X=1.005 $Y=1.485 $X2=0 $Y2=0
cc_329 N_Y_c_442_n N_VGND_M1014_s 0.00467331f $X=1.05 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_330 N_Y_c_452_n N_VGND_M1017_d 0.00708074f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_331 N_Y_c_475_n N_VGND_M1003_d 0.00576665f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_332 N_Y_c_492_n N_VGND_M1019_s 0.00464181f $X=5.02 $Y=0.71 $X2=0 $Y2=0
cc_333 N_Y_c_442_n N_VGND_c_697_n 0.0162283f $X=1.05 $Y=0.73 $X2=0 $Y2=0
cc_334 N_Y_c_452_n N_VGND_c_698_n 0.0213394f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_335 N_Y_c_452_n N_VGND_c_699_n 0.00273863f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_336 N_Y_c_456_n N_VGND_c_699_n 0.0190918f $X=2.13 $Y=0.4 $X2=0 $Y2=0
cc_337 N_Y_c_475_n N_VGND_c_699_n 0.00281024f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_338 N_Y_c_475_n N_VGND_c_700_n 0.0213394f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_339 N_Y_c_492_n N_VGND_c_701_n 0.0176382f $X=5.02 $Y=0.71 $X2=0 $Y2=0
cc_340 N_Y_c_433_n N_VGND_c_702_n 0.0176056f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_341 N_Y_c_442_n N_VGND_c_702_n 0.00263122f $X=1.05 $Y=0.73 $X2=0 $Y2=0
cc_342 N_Y_c_442_n N_VGND_c_703_n 0.00263122f $X=1.05 $Y=0.73 $X2=0 $Y2=0
cc_343 N_Y_c_451_n N_VGND_c_703_n 0.0145408f $X=1.145 $Y=0.42 $X2=0 $Y2=0
cc_344 N_Y_c_452_n N_VGND_c_703_n 0.00273863f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_345 N_Y_c_475_n N_VGND_c_704_n 0.00263122f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_346 N_Y_c_479_n N_VGND_c_704_n 0.0167556f $X=3.13 $Y=0.375 $X2=0 $Y2=0
cc_347 N_Y_c_492_n N_VGND_c_704_n 0.0139982f $X=5.02 $Y=0.71 $X2=0 $Y2=0
cc_348 N_Y_c_492_n N_VGND_c_705_n 0.00907844f $X=5.02 $Y=0.71 $X2=0 $Y2=0
cc_349 N_Y_c_434_n N_VGND_c_705_n 0.0167396f $X=5.185 $Y=0.38 $X2=0 $Y2=0
cc_350 N_Y_M1014_d N_VGND_c_706_n 0.00243803f $X=0.14 $Y=0.235 $X2=0 $Y2=0
cc_351 N_Y_M1009_s N_VGND_c_706_n 0.0023722f $X=1.005 $Y=0.235 $X2=0 $Y2=0
cc_352 N_Y_M1018_d N_VGND_c_706_n 0.0025535f $X=1.975 $Y=0.235 $X2=0 $Y2=0
cc_353 N_Y_M1012_s N_VGND_c_706_n 0.00224096f $X=2.99 $Y=0.235 $X2=0 $Y2=0
cc_354 N_Y_M1015_d N_VGND_c_706_n 0.00215706f $X=5.045 $Y=0.235 $X2=0 $Y2=0
cc_355 N_Y_c_433_n N_VGND_c_706_n 0.00989931f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_356 N_Y_c_442_n N_VGND_c_706_n 0.0101289f $X=1.05 $Y=0.73 $X2=0 $Y2=0
cc_357 N_Y_c_451_n N_VGND_c_706_n 0.00921046f $X=1.145 $Y=0.42 $X2=0 $Y2=0
cc_358 N_Y_c_452_n N_VGND_c_706_n 0.00994312f $X=1.965 $Y=0.73 $X2=0 $Y2=0
cc_359 N_Y_c_456_n N_VGND_c_706_n 0.0124719f $X=2.13 $Y=0.4 $X2=0 $Y2=0
cc_360 N_Y_c_475_n N_VGND_c_706_n 0.00995639f $X=2.965 $Y=0.73 $X2=0 $Y2=0
cc_361 N_Y_c_479_n N_VGND_c_706_n 0.0121246f $X=3.13 $Y=0.375 $X2=0 $Y2=0
cc_362 N_Y_c_492_n N_VGND_c_706_n 0.038985f $X=5.02 $Y=0.71 $X2=0 $Y2=0
cc_363 N_Y_c_434_n N_VGND_c_706_n 0.0122828f $X=5.185 $Y=0.38 $X2=0 $Y2=0
cc_364 N_Y_c_492_n A_684_47# 0.0155718f $X=5.02 $Y=0.71 $X2=-0.19 $Y2=-0.24
cc_365 N_Y_c_492_n A_923_47# 0.00577135f $X=5.02 $Y=0.71 $X2=-0.19 $Y2=-0.24
cc_366 A_287_297# N_VPWR_c_626_n 0.00224864f $X=1.435 $Y=1.485 $X2=0.5 $Y2=1.16
cc_367 N_A_467_297#_c_581_n N_VPWR_M1006_s 0.00354452f $X=4.19 $Y=1.97 $X2=-0.19
+ $Y2=1.305
cc_368 N_A_467_297#_c_584_n N_VPWR_M1016_d 0.00428976f $X=5.07 $Y=1.975 $X2=0
+ $Y2=0
cc_369 N_A_467_297#_c_581_n N_VPWR_c_627_n 0.0155135f $X=4.19 $Y=1.97 $X2=0
+ $Y2=0
cc_370 N_A_467_297#_c_584_n N_VPWR_c_628_n 0.0165275f $X=5.07 $Y=1.975 $X2=0
+ $Y2=0
cc_371 N_A_467_297#_c_581_n N_VPWR_c_629_n 0.00257989f $X=4.19 $Y=1.97 $X2=0
+ $Y2=0
cc_372 N_A_467_297#_c_609_p N_VPWR_c_629_n 0.0130847f $X=4.285 $Y=2.3 $X2=0
+ $Y2=0
cc_373 N_A_467_297#_c_584_n N_VPWR_c_629_n 0.00279402f $X=5.07 $Y=1.975 $X2=0
+ $Y2=0
cc_374 N_A_467_297#_c_568_n N_VPWR_c_631_n 0.00242398f $X=3.155 $Y=1.88 $X2=0
+ $Y2=0
cc_375 N_A_467_297#_c_569_n N_VPWR_c_631_n 0.0252517f $X=3.43 $Y=2.3 $X2=0 $Y2=0
cc_376 N_A_467_297#_c_581_n N_VPWR_c_631_n 0.00257989f $X=4.19 $Y=1.97 $X2=0
+ $Y2=0
cc_377 N_A_467_297#_c_584_n N_VPWR_c_632_n 0.00279402f $X=5.07 $Y=1.975 $X2=0
+ $Y2=0
cc_378 N_A_467_297#_c_571_n N_VPWR_c_632_n 0.02187f $X=5.235 $Y=2.36 $X2=0 $Y2=0
cc_379 N_A_467_297#_M1005_s N_VPWR_c_626_n 0.00224864f $X=2.335 $Y=1.485 $X2=0
+ $Y2=0
cc_380 N_A_467_297#_M1006_d N_VPWR_c_626_n 0.00223936f $X=3.305 $Y=1.485 $X2=0
+ $Y2=0
cc_381 N_A_467_297#_M1008_s N_VPWR_c_626_n 0.00245113f $X=4.145 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_A_467_297#_M1011_d N_VPWR_c_626_n 0.00278069f $X=5.045 $Y=1.485 $X2=0
+ $Y2=0
cc_383 N_A_467_297#_c_568_n N_VPWR_c_626_n 0.00513688f $X=3.155 $Y=1.88 $X2=0
+ $Y2=0
cc_384 N_A_467_297#_c_569_n N_VPWR_c_626_n 0.01396f $X=3.43 $Y=2.3 $X2=0 $Y2=0
cc_385 N_A_467_297#_c_581_n N_VPWR_c_626_n 0.0101026f $X=4.19 $Y=1.97 $X2=0
+ $Y2=0
cc_386 N_A_467_297#_c_609_p N_VPWR_c_626_n 0.00799109f $X=4.285 $Y=2.3 $X2=0
+ $Y2=0
cc_387 N_A_467_297#_c_584_n N_VPWR_c_626_n 0.0100043f $X=5.07 $Y=1.975 $X2=0
+ $Y2=0
cc_388 N_A_467_297#_c_571_n N_VPWR_c_626_n 0.0126013f $X=5.235 $Y=2.36 $X2=0
+ $Y2=0
cc_389 N_VGND_c_706_n A_684_47# 0.0062974f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24
cc_390 N_VGND_c_706_n A_923_47# 0.00318969f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_2.pxi.spice
* Created: Tue Sep  1 19:11:14 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%A N_A_M1000_g N_A_M1001_g N_A_M1002_g
+ N_A_c_37_n N_A_M1003_g N_A_M1004_g A A A
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%Y N_Y_M1002_d N_Y_M1000_s N_Y_M1001_s
+ N_Y_c_102_n N_Y_c_96_n N_Y_c_97_n N_Y_c_91_n N_Y_c_111_n N_Y_c_98_n N_Y_c_92_n
+ N_Y_c_93_n N_Y_c_99_n Y Y Y N_Y_c_95_n N_Y_c_101_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%Y
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%KAPWR N_KAPWR_M1000_d N_KAPWR_M1003_d
+ N_KAPWR_c_159_n N_KAPWR_c_160_n N_KAPWR_c_165_n KAPWR N_KAPWR_c_166_n
+ N_KAPWR_c_161_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%VGND N_VGND_M1002_s N_VGND_M1004_s
+ N_VGND_c_198_n N_VGND_c_199_n N_VGND_c_200_n VGND N_VGND_c_201_n
+ N_VGND_c_202_n N_VGND_c_203_n N_VGND_c_204_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%VPWR VPWR N_VPWR_c_223_n
+ N_VPWR_c_222_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_2%VPWR
cc_1 VNB N_A_M1001_g 4.57292e-19 $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_2 VNB N_A_M1002_g 0.0421156f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.445
cc_3 VNB N_A_c_37_n 0.0934495f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.295
cc_4 VNB N_A_M1003_g 4.91581e-19 $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.985
cc_5 VNB N_A_M1004_g 0.0349086f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=0.445
cc_6 VNB A 0.0140604f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_7 VNB N_Y_c_91_n 0.00149799f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=0.445
cc_8 VNB N_Y_c_92_n 0.00167495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_Y_c_93_n 0.00410962f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_10 VNB Y 0.0210583f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_11 VNB N_Y_c_95_n 0.0101921f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.16
cc_12 VNB N_VGND_c_198_n 0.0193788f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.015
cc_13 VNB N_VGND_c_199_n 0.0101596f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.445
cc_14 VNB N_VGND_c_200_n 0.0154987f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.295
cc_15 VNB N_VGND_c_201_n 0.0199636f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.025
cc_16 VNB N_VGND_c_202_n 0.0142308f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_17 VNB N_VGND_c_203_n 0.00564902f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_18 VNB N_VGND_c_204_n 0.141662f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_19 VNB N_VPWR_c_222_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.015
cc_20 VPB N_A_M1000_g 0.0271137f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_21 VPB N_A_M1001_g 0.0195484f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_22 VPB N_A_c_37_n 0.00626529f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.295
cc_23 VPB N_A_M1003_g 0.0231397f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.985
cc_24 VPB N_Y_c_96_n 0.00291986f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.985
cc_25 VPB N_Y_c_97_n 0.00831597f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.985
cc_26 VPB N_Y_c_98_n 9.22346e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_Y_c_99_n 0.00145777f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_28 VPB Y 0.00792875f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_29 VPB N_Y_c_101_n 0.00805732f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.177
cc_30 VPB N_KAPWR_c_159_n 0.00903021f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_31 VPB N_KAPWR_c_160_n 0.011566f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.295
cc_32 VPB N_KAPWR_c_161_n 0.0215128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_223_n 0.0527727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_222_n 0.0424642f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.015
cc_35 N_A_M1000_g N_Y_c_102_n 0.00131597f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_36 N_A_M1000_g N_Y_c_96_n 0.0128484f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_37 N_A_M1001_g N_Y_c_96_n 0.0115307f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_38 N_A_c_37_n N_Y_c_96_n 0.0031781f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_39 A N_Y_c_96_n 0.0477264f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_40 N_A_c_37_n N_Y_c_97_n 0.00508687f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_41 A N_Y_c_97_n 0.0180799f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_42 N_A_M1002_g N_Y_c_91_n 0.00189162f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_43 N_A_M1004_g N_Y_c_91_n 0.00180689f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_44 N_A_M1001_g N_Y_c_111_n 4.82584e-19 $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_45 N_A_M1003_g N_Y_c_111_n 4.82584e-19 $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_46 N_A_c_37_n N_Y_c_98_n 4.58912e-19 $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_47 N_A_M1003_g N_Y_c_98_n 0.0145268f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_48 A N_Y_c_98_n 0.00498066f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_49 N_A_M1004_g N_Y_c_92_n 0.0146405f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_50 A N_Y_c_92_n 0.00394157f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_51 N_A_M1002_g N_Y_c_93_n 0.00568793f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_52 N_A_c_37_n N_Y_c_93_n 0.00241459f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_53 A N_Y_c_93_n 0.0183373f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A_c_37_n N_Y_c_99_n 0.00232565f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_55 A N_Y_c_99_n 0.0156166f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_M1003_g Y 0.00683246f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A_M1004_g Y 0.0148622f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_58 A Y 0.0184815f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_KAPWR_c_159_n 0.00247485f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_60 N_A_M1003_g N_KAPWR_c_159_n 0.00247485f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_M1000_g N_KAPWR_c_160_n 0.00233626f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_KAPWR_c_165_n 6.07575e-19 $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_M1000_g N_KAPWR_c_166_n 0.00761429f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_64 N_A_M1001_g N_KAPWR_c_166_n 0.00682379f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_KAPWR_c_161_n 0.00682391f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1002_g N_VGND_c_198_n 0.00365907f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_67 N_A_c_37_n N_VGND_c_198_n 0.00633207f $X=1.355 $Y=1.295 $X2=0 $Y2=0
cc_68 A N_VGND_c_198_n 0.0101104f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A_M1002_g N_VGND_c_200_n 5.86108e-19 $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_M1004_g N_VGND_c_200_n 0.00871096f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1002_g N_VGND_c_202_n 0.00585385f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_M1004_g N_VGND_c_202_n 0.00364083f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_73 N_A_M1002_g N_VGND_c_204_n 0.0119927f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_M1004_g N_VGND_c_204_n 0.00434306f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_VPWR_c_223_n 0.0054895f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_VPWR_c_223_n 0.0054895f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_VPWR_c_223_n 0.0054895f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1000_g N_VPWR_c_222_n 0.00615194f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_VPWR_c_222_n 0.00516436f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_M1003_g N_VPWR_c_222_n 0.0061063f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_81 N_Y_c_96_n N_KAPWR_M1000_d 0.00171343f $X=1.045 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_82 N_Y_c_101_n N_KAPWR_M1003_d 0.00291707f $X=1.615 $Y=1.46 $X2=0 $Y2=0
cc_83 N_Y_M1001_s N_KAPWR_c_159_n 0.00147741f $X=1 $Y=1.485 $X2=0 $Y2=0
cc_84 N_Y_c_96_n N_KAPWR_c_159_n 0.00502158f $X=1.045 $Y=1.545 $X2=0 $Y2=0
cc_85 N_Y_c_111_n N_KAPWR_c_159_n 0.0203024f $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_86 N_Y_c_98_n N_KAPWR_c_159_n 0.00512659f $X=1.475 $Y=1.545 $X2=0 $Y2=0
cc_87 N_Y_c_101_n N_KAPWR_c_159_n 0.00199519f $X=1.615 $Y=1.46 $X2=0 $Y2=0
cc_88 N_Y_M1000_s N_KAPWR_c_160_n 7.38703e-19 $X=0.155 $Y=1.485 $X2=0 $Y2=0
cc_89 N_Y_c_102_n N_KAPWR_c_160_n 0.0247761f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_90 N_Y_c_96_n N_KAPWR_c_160_n 0.0046895f $X=1.045 $Y=1.545 $X2=0 $Y2=0
cc_91 N_Y_c_102_n N_KAPWR_c_165_n 0.00150275f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_92 N_Y_c_96_n N_KAPWR_c_165_n 0.00134299f $X=1.045 $Y=1.545 $X2=0 $Y2=0
cc_93 N_Y_c_111_n N_KAPWR_c_165_n 4.04566e-19 $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_94 N_Y_c_102_n N_KAPWR_c_166_n 0.0261096f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_95 N_Y_c_96_n N_KAPWR_c_166_n 0.0164188f $X=1.045 $Y=1.545 $X2=0 $Y2=0
cc_96 N_Y_c_111_n N_KAPWR_c_166_n 0.0262616f $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_97 N_Y_c_111_n N_KAPWR_c_161_n 0.0262662f $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_98 N_Y_c_98_n N_KAPWR_c_161_n 0.00172789f $X=1.475 $Y=1.545 $X2=0 $Y2=0
cc_99 N_Y_c_101_n N_KAPWR_c_161_n 0.0214627f $X=1.615 $Y=1.46 $X2=0 $Y2=0
cc_100 N_Y_c_92_n N_VGND_c_200_n 0.0027328f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_101 N_Y_c_95_n N_VGND_c_200_n 0.0230152f $X=1.615 $Y=0.895 $X2=0 $Y2=0
cc_102 N_Y_c_91_n N_VGND_c_202_n 0.0117468f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_103 N_Y_c_92_n N_VGND_c_202_n 0.0023442f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_104 N_Y_M1002_d N_VGND_c_204_n 0.00285545f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_105 N_Y_c_91_n N_VGND_c_204_n 0.00845997f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_106 N_Y_c_92_n N_VGND_c_204_n 0.00409036f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_107 N_Y_c_95_n N_VGND_c_204_n 0.00136789f $X=1.615 $Y=0.895 $X2=0 $Y2=0
cc_108 N_Y_c_102_n N_VPWR_c_223_n 0.0125314f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_109 N_Y_c_111_n N_VPWR_c_223_n 0.0104472f $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_110 N_Y_M1000_s N_VPWR_c_222_n 0.00128181f $X=0.155 $Y=1.485 $X2=0 $Y2=0
cc_111 N_Y_M1001_s N_VPWR_c_222_n 0.00151759f $X=1 $Y=1.485 $X2=0 $Y2=0
cc_112 N_Y_c_102_n N_VPWR_c_222_n 0.00207101f $X=0.28 $Y=1.83 $X2=0 $Y2=0
cc_113 N_Y_c_111_n N_VPWR_c_222_n 0.00178601f $X=1.14 $Y=1.83 $X2=0 $Y2=0
cc_114 N_KAPWR_c_159_n N_VPWR_c_223_n 0.00227985f $X=1.44 $Y=2.24 $X2=0 $Y2=0
cc_115 N_KAPWR_c_160_n N_VPWR_c_223_n 0.00147939f $X=0.54 $Y=2.21 $X2=0 $Y2=0
cc_116 N_KAPWR_c_165_n N_VPWR_c_223_n 2.22852e-19 $X=0.83 $Y=2.21 $X2=0 $Y2=0
cc_117 N_KAPWR_c_166_n N_VPWR_c_223_n 0.0189011f $X=0.71 $Y=1.965 $X2=0 $Y2=0
cc_118 N_KAPWR_c_161_n N_VPWR_c_223_n 0.0210176f $X=1.57 $Y=1.965 $X2=0 $Y2=0
cc_119 N_KAPWR_M1000_d N_VPWR_c_222_n 0.00113449f $X=0.57 $Y=1.485 $X2=0 $Y2=0
cc_120 N_KAPWR_M1003_d N_VPWR_c_222_n 0.00109164f $X=1.43 $Y=1.485 $X2=0 $Y2=0
cc_121 N_KAPWR_c_160_n N_VPWR_c_222_n 0.175136f $X=0.54 $Y=2.21 $X2=0 $Y2=0
cc_122 N_KAPWR_c_166_n N_VPWR_c_222_n 0.00295042f $X=0.71 $Y=1.965 $X2=0 $Y2=0
cc_123 N_KAPWR_c_161_n N_VPWR_c_222_n 0.00299364f $X=1.57 $Y=1.965 $X2=0 $Y2=0

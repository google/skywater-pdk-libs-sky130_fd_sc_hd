* File: sky130_fd_sc_hd__dlxtn_1.pxi.spice
* Created: Tue Sep  1 19:06:07 2020
* 
x_PM_SKY130_FD_SC_HD__DLXTN_1%GATE_N N_GATE_N_c_133_n N_GATE_N_c_128_n
+ N_GATE_N_M1016_g N_GATE_N_c_134_n N_GATE_N_M1009_g N_GATE_N_c_129_n
+ N_GATE_N_c_135_n GATE_N GATE_N N_GATE_N_c_131_n N_GATE_N_c_132_n
+ PM_SKY130_FD_SC_HD__DLXTN_1%GATE_N
x_PM_SKY130_FD_SC_HD__DLXTN_1%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1009_s
+ N_A_27_47#_M1010_g N_A_27_47#_M1000_g N_A_27_47#_c_172_n N_A_27_47#_M1015_g
+ N_A_27_47#_c_182_n N_A_27_47#_M1002_g N_A_27_47#_c_326_p N_A_27_47#_c_174_n
+ N_A_27_47#_c_175_n N_A_27_47#_c_184_n N_A_27_47#_c_176_n N_A_27_47#_c_185_n
+ N_A_27_47#_c_177_n N_A_27_47#_c_178_n N_A_27_47#_c_187_n N_A_27_47#_c_188_n
+ N_A_27_47#_c_189_n N_A_27_47#_c_190_n N_A_27_47#_c_191_n N_A_27_47#_c_179_n
+ N_A_27_47#_c_180_n PM_SKY130_FD_SC_HD__DLXTN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLXTN_1%D N_D_c_339_n N_D_c_340_n N_D_M1005_g N_D_c_346_n
+ N_D_M1014_g N_D_c_341_n N_D_c_342_n N_D_c_347_n D N_D_c_343_n N_D_c_344_n
+ PM_SKY130_FD_SC_HD__DLXTN_1%D
x_PM_SKY130_FD_SC_HD__DLXTN_1%A_299_47# N_A_299_47#_M1005_s N_A_299_47#_M1014_s
+ N_A_299_47#_M1007_g N_A_299_47#_c_397_n N_A_299_47#_M1011_g
+ N_A_299_47#_c_405_n N_A_299_47#_c_399_n N_A_299_47#_c_400_n
+ N_A_299_47#_c_401_n N_A_299_47#_c_407_n N_A_299_47#_c_402_n
+ N_A_299_47#_c_403_n PM_SKY130_FD_SC_HD__DLXTN_1%A_299_47#
x_PM_SKY130_FD_SC_HD__DLXTN_1%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1003_g N_A_193_47#_c_490_n N_A_193_47#_M1017_g
+ N_A_193_47#_c_491_n N_A_193_47#_c_492_n N_A_193_47#_c_496_n
+ N_A_193_47#_c_497_n N_A_193_47#_c_498_n N_A_193_47#_c_499_n
+ N_A_193_47#_c_500_n N_A_193_47#_c_501_n N_A_193_47#_c_493_n
+ PM_SKY130_FD_SC_HD__DLXTN_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLXTN_1%A_715_21# N_A_715_21#_M1006_s N_A_715_21#_M1001_s
+ N_A_715_21#_M1012_g N_A_715_21#_M1004_g N_A_715_21#_M1008_g
+ N_A_715_21#_M1013_g N_A_715_21#_c_607_n N_A_715_21#_c_608_n
+ N_A_715_21#_c_619_p N_A_715_21#_c_625_p N_A_715_21#_c_600_n
+ N_A_715_21#_c_609_n N_A_715_21#_c_601_n N_A_715_21#_c_602_n
+ N_A_715_21#_c_621_p N_A_715_21#_c_627_p N_A_715_21#_c_633_p
+ N_A_715_21#_c_603_n PM_SKY130_FD_SC_HD__DLXTN_1%A_715_21#
x_PM_SKY130_FD_SC_HD__DLXTN_1%A_560_47# N_A_560_47#_M1015_d N_A_560_47#_M1003_d
+ N_A_560_47#_c_682_n N_A_560_47#_M1006_g N_A_560_47#_M1001_g
+ N_A_560_47#_c_683_n N_A_560_47#_c_684_n N_A_560_47#_c_694_n
+ N_A_560_47#_c_698_n N_A_560_47#_c_685_n N_A_560_47#_c_691_n
+ N_A_560_47#_c_686_n N_A_560_47#_c_687_n PM_SKY130_FD_SC_HD__DLXTN_1%A_560_47#
x_PM_SKY130_FD_SC_HD__DLXTN_1%VPWR N_VPWR_M1009_d N_VPWR_M1014_d N_VPWR_M1004_d
+ N_VPWR_M1001_d N_VPWR_c_773_n N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n
+ VPWR N_VPWR_c_777_n N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n
+ N_VPWR_c_781_n N_VPWR_c_772_n N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n
+ N_VPWR_c_786_n PM_SKY130_FD_SC_HD__DLXTN_1%VPWR
x_PM_SKY130_FD_SC_HD__DLXTN_1%Q N_Q_M1008_d N_Q_M1013_d Q Q Q Q N_Q_c_872_n
+ PM_SKY130_FD_SC_HD__DLXTN_1%Q
x_PM_SKY130_FD_SC_HD__DLXTN_1%VGND N_VGND_M1016_d N_VGND_M1005_d N_VGND_M1012_d
+ N_VGND_M1006_d N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n
+ N_VGND_c_891_n VGND N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n
+ N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n N_VGND_c_899_n
+ N_VGND_c_900_n PM_SKY130_FD_SC_HD__DLXTN_1%VGND
cc_1 VNB N_GATE_N_c_128_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_N_c_129_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_131_n 0.0212744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_132_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1010_g 0.0406284f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_172_n 0.0306297f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_8 VNB N_A_27_47#_M1015_g 0.0186012f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_9 VNB N_A_27_47#_c_174_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_175_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_176_n 0.00515794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_177_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_178_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_179_n 0.00262586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_180_n 0.0235456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_c_339_n 0.00558205f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.07
cc_17 VNB N_D_c_340_n 0.0171218f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_18 VNB N_D_c_341_n 0.0257161f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_19 VNB N_D_c_342_n 0.0121577f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_20 VNB N_D_c_343_n 0.0131107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_D_c_344_n 0.00647161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_M1007_g 0.0232546f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_23 VNB N_A_299_47#_c_397_n 0.0305912f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_24 VNB N_A_299_47#_M1011_g 0.00427745f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_25 VNB N_A_299_47#_c_399_n 0.00327127f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_26 VNB N_A_299_47#_c_400_n 0.00234194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_299_47#_c_401_n 0.00105735f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_28 VNB N_A_299_47#_c_402_n 0.00177472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_299_47#_c_403_n 0.00192362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_490_n 0.0230889f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_31 VNB N_A_193_47#_c_491_n 0.0200852f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_32 VNB N_A_193_47#_c_492_n 0.0136323f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_493_n 0.0206918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_715_21#_M1012_g 0.047176f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_35 VNB N_A_715_21#_c_600_n 0.0015831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_715_21#_c_601_n 0.00472551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_715_21#_c_602_n 0.0248945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_715_21#_c_603_n 0.0196002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_560_47#_c_682_n 0.0205485f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_40 VNB N_A_560_47#_c_683_n 0.0421338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_560_47#_c_684_n 0.00807219f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_42 VNB N_A_560_47#_c_685_n 0.00230325f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_560_47#_c_686_n 0.00474481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_560_47#_c_687_n 0.00185621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VPWR_c_772_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB Q 0.0130125f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_47 VNB N_Q_c_872_n 0.0247635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_887_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_49 VNB N_VGND_c_888_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_50 VNB N_VGND_c_889_n 0.00919263f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_51 VNB N_VGND_c_890_n 0.0202095f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_52 VNB N_VGND_c_891_n 0.00237086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_892_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_893_n 0.0269775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_894_n 0.0417421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_895_n 0.0165063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_896_n 0.296722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_897_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_898_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_899_n 0.00516539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_900_n 0.00323302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VPB N_GATE_N_c_133_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_63 VPB N_GATE_N_c_134_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_64 VPB N_GATE_N_c_135_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_65 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_66 VPB N_GATE_N_c_131_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_67 VPB N_A_27_47#_M1000_g 0.0397961f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_68 VPB N_A_27_47#_c_182_n 0.0282933f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_69 VPB N_A_27_47#_M1002_g 0.0210872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_184_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_71 VPB N_A_27_47#_c_185_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_177_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_187_n 0.00458212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_188_n 0.0273234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_189_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_190_n 0.0054554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_191_n 0.00123931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_179_n 0.00161824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_180_n 0.011944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_D_c_339_n 0.0196123f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.07
cc_81 VPB N_D_c_346_n 0.0177239f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_82 VPB N_D_c_347_n 0.0207624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_D_c_344_n 0.00156012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_299_47#_M1011_g 0.0388168f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_85 VPB N_A_299_47#_c_405_n 0.00681894f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_86 VPB N_A_299_47#_c_401_n 0.00354472f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_87 VPB N_A_299_47#_c_407_n 0.00734188f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_88 VPB N_A_193_47#_M1003_g 0.0298355f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_89 VPB N_A_193_47#_c_492_n 0.00763939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_193_47#_c_496_n 0.00285357f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_91 VPB N_A_193_47#_c_497_n 0.00425978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_193_47#_c_498_n 0.00237077f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_93 VPB N_A_193_47#_c_499_n 0.00690126f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_94 VPB N_A_193_47#_c_500_n 0.00102715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_193_47#_c_501_n 0.0104024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_193_47#_c_493_n 0.0442437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_715_21#_M1012_g 0.0151334f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_98 VPB N_A_715_21#_M1004_g 0.0258788f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_99 VPB N_A_715_21#_M1013_g 0.0224782f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_100 VPB N_A_715_21#_c_607_n 0.00588124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_715_21#_c_608_n 0.0434235f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_102 VPB N_A_715_21#_c_609_n 0.0023093f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_715_21#_c_601_n 0.00372091f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_715_21#_c_602_n 0.00611128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_560_47#_M1001_g 0.0237898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_560_47#_c_683_n 0.0146909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_560_47#_c_684_n 5.11289e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_108 VPB N_A_560_47#_c_691_n 0.00630581f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_109 VPB N_A_560_47#_c_686_n 0.00205677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_560_47#_c_687_n 0.0011668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_773_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_112 VPB N_VPWR_c_774_n 0.0034306f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_113 VPB N_VPWR_c_775_n 0.00970698f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_114 VPB N_VPWR_c_776_n 0.00197765f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_115 VPB N_VPWR_c_777_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_116 VPB N_VPWR_c_778_n 0.0292999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_779_n 0.0387914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_780_n 0.0176692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_781_n 0.0151046f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_772_n 0.0575776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_783_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_784_n 0.00407272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_785_n 0.00612673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_786_n 0.00421326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB Q 0.00494099f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_126 VPB Q 0.0252202f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_127 VPB N_Q_c_872_n 0.0155144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 N_GATE_N_c_128_n N_A_27_47#_M1010_g 0.0187834f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_129 N_GATE_N_c_132_n N_A_27_47#_M1010_g 0.0041981f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_130 N_GATE_N_c_135_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_131 N_GATE_N_c_131_n N_A_27_47#_M1000_g 0.00527228f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_132 N_GATE_N_c_128_n N_A_27_47#_c_174_n 0.00663556f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_133 N_GATE_N_c_129_n N_A_27_47#_c_174_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_134 N_GATE_N_c_129_n N_A_27_47#_c_175_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_135 GATE_N N_A_27_47#_c_175_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_136 N_GATE_N_c_131_n N_A_27_47#_c_175_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_137 N_GATE_N_c_134_n N_A_27_47#_c_184_n 0.0135489f $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_138 N_GATE_N_c_135_n N_A_27_47#_c_184_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_139 N_GATE_N_c_134_n N_A_27_47#_c_185_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_140 N_GATE_N_c_135_n N_A_27_47#_c_185_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_141 GATE_N N_A_27_47#_c_185_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_142 N_GATE_N_c_131_n N_A_27_47#_c_185_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_143 N_GATE_N_c_131_n N_A_27_47#_c_177_n 0.00319708f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_144 N_GATE_N_c_129_n N_A_27_47#_c_178_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_145 GATE_N N_A_27_47#_c_178_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_146 N_GATE_N_c_132_n N_A_27_47#_c_178_n 0.0015185f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_147 N_GATE_N_c_133_n N_A_27_47#_c_189_n 0.0033897f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_148 N_GATE_N_c_135_n N_A_27_47#_c_189_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_149 GATE_N N_A_27_47#_c_189_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_150 N_GATE_N_c_133_n N_A_27_47#_c_190_n 7.60515e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_151 N_GATE_N_c_135_n N_A_27_47#_c_190_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_152 GATE_N N_A_27_47#_c_180_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_153 N_GATE_N_c_131_n N_A_27_47#_c_180_n 0.0165992f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_154 N_GATE_N_c_134_n N_VPWR_c_773_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_155 N_GATE_N_c_134_n N_VPWR_c_777_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_156 N_GATE_N_c_134_n N_VPWR_c_772_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_157 N_GATE_N_c_128_n N_VGND_c_887_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_158 N_GATE_N_c_128_n N_VGND_c_892_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_159 N_GATE_N_c_129_n N_VGND_c_892_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_160 N_GATE_N_c_128_n N_VGND_c_896_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_188_n N_D_c_339_n 0.00200477f $X=2.89 $Y=1.53 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_180_n N_D_c_339_n 0.00359135f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1010_g N_D_c_341_n 0.00448292f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_188_n N_D_c_341_n 0.00274536f $X=2.89 $Y=1.53 $X2=0 $Y2=0
cc_165 N_A_27_47#_M1000_g N_D_c_347_n 0.00359135f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_180_n N_D_c_343_n 0.00278795f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_188_n N_D_c_344_n 0.00814614f $X=2.89 $Y=1.53 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_172_n N_A_299_47#_M1007_g 0.00907227f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_M1015_g N_A_299_47#_M1007_g 0.0249914f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_176_n N_A_299_47#_M1007_g 5.44921e-19 $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_172_n N_A_299_47#_c_397_n 0.0086961f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_176_n N_A_299_47#_c_397_n 4.5916e-19 $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_188_n N_A_299_47#_c_397_n 5.84142e-19 $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_179_n N_A_299_47#_c_397_n 0.00256866f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_188_n N_A_299_47#_M1011_g 0.00554036f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_179_n N_A_299_47#_M1011_g 6.33457e-19 $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_188_n N_A_299_47#_c_405_n 5.24155e-19 $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_176_n N_A_299_47#_c_399_n 0.00247801f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_172_n N_A_299_47#_c_400_n 3.38968e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_176_n N_A_299_47#_c_400_n 0.0155004f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_179_n N_A_299_47#_c_400_n 0.00571569f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_188_n N_A_299_47#_c_401_n 0.0104974f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_188_n N_A_299_47#_c_407_n 0.0208753f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_188_n N_A_299_47#_c_403_n 0.00655292f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_182_n N_A_193_47#_M1003_g 0.00993622f $X=3.145 $Y=1.88 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_M1002_g N_A_193_47#_M1003_g 0.0190153f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_187_n N_A_193_47#_M1003_g 0.00127697f $X=3.2 $Y=1.745 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_172_n N_A_193_47#_c_490_n 0.00212264f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_M1015_g N_A_193_47#_c_490_n 0.0133872f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_176_n N_A_193_47#_c_490_n 0.00445002f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_172_n N_A_193_47#_c_491_n 0.0152444f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_176_n N_A_193_47#_c_491_n 0.00676112f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_179_n N_A_193_47#_c_491_n 0.00460475f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1010_g N_A_193_47#_c_492_n 0.00507692f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_174_n N_A_193_47#_c_492_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_177_n N_A_193_47#_c_492_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_178_n N_A_193_47#_c_492_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_188_n N_A_193_47#_c_492_n 0.0183655f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_189_n N_A_193_47#_c_492_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_190_n N_A_193_47#_c_492_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_184_n N_A_193_47#_c_496_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_188_n N_A_193_47#_c_496_n 0.00195186f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_180_n N_A_193_47#_c_496_n 0.00507692f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_188_n N_A_193_47#_c_497_n 0.084973f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_M1000_g N_A_193_47#_c_498_n 0.00448406f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_184_n N_A_193_47#_c_498_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_188_n N_A_193_47#_c_498_n 0.0259095f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_190_n N_A_193_47#_c_498_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_M1000_g N_A_193_47#_c_499_n 0.00507692f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_187_n N_A_193_47#_c_500_n 9.27234e-19 $X=3.2 $Y=1.745 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_188_n N_A_193_47#_c_500_n 0.0255946f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_172_n N_A_193_47#_c_501_n 8.34423e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_182_n N_A_193_47#_c_501_n 2.75547e-19 $X=3.145 $Y=1.88 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1002_g N_A_193_47#_c_501_n 3.99123e-19 $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_215 N_A_27_47#_c_176_n N_A_193_47#_c_501_n 0.00917896f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_188_n N_A_193_47#_c_501_n 0.0252542f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_191_n N_A_193_47#_c_501_n 0.00265117f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_179_n N_A_193_47#_c_501_n 0.0400279f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_172_n N_A_193_47#_c_493_n 0.0203374f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_182_n N_A_193_47#_c_493_n 0.0203336f $X=3.145 $Y=1.88 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_176_n N_A_193_47#_c_493_n 0.00304605f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_187_n N_A_193_47#_c_493_n 4.6339e-19 $X=3.2 $Y=1.745 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_188_n N_A_193_47#_c_493_n 0.00536625f $X=2.89 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_191_n N_A_193_47#_c_493_n 0.00304207f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_179_n N_A_193_47#_c_493_n 0.0223835f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_176_n N_A_715_21#_M1012_g 3.00701e-19 $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_179_n N_A_715_21#_M1012_g 0.00107396f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1002_g N_A_715_21#_M1004_g 0.0238373f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_182_n N_A_715_21#_c_608_n 0.0167028f $X=3.145 $Y=1.88 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_187_n N_A_715_21#_c_608_n 5.08354e-19 $X=3.2 $Y=1.745 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_182_n N_A_560_47#_c_694_n 5.15715e-19 $X=3.145 $Y=1.88 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1002_g N_A_560_47#_c_694_n 0.00925302f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_233 N_A_27_47#_c_187_n N_A_560_47#_c_694_n 0.0102887f $X=3.2 $Y=1.745 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_191_n N_A_560_47#_c_694_n 0.0028874f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_172_n N_A_560_47#_c_698_n 5.57351e-19 $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_M1015_g N_A_560_47#_c_698_n 0.00434196f $X=2.725 $Y=0.415
+ $X2=0 $Y2=0
cc_237 N_A_27_47#_c_176_n N_A_560_47#_c_698_n 0.0284217f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_176_n N_A_560_47#_c_685_n 0.0207576f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_182_n N_A_560_47#_c_691_n 0.00435126f $X=3.145 $Y=1.88 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1002_g N_A_560_47#_c_691_n 0.00741258f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_241 N_A_27_47#_c_187_n N_A_560_47#_c_691_n 0.0264085f $X=3.2 $Y=1.745 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_191_n N_A_560_47#_c_691_n 0.00113328f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_179_n N_A_560_47#_c_691_n 0.00733228f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_176_n N_A_560_47#_c_687_n 0.0040221f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_191_n N_A_560_47#_c_687_n 2.15684e-19 $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_179_n N_A_560_47#_c_687_n 0.0334614f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_184_n N_VPWR_M1009_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_248 N_A_27_47#_M1000_g N_VPWR_c_773_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_184_n N_VPWR_c_773_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_185_n N_VPWR_c_773_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_189_n N_VPWR_c_773_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_188_n N_VPWR_c_774_n 9.13039e-19 $X=2.89 $Y=1.53 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_184_n N_VPWR_c_777_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_185_n N_VPWR_c_777_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_255 N_A_27_47#_M1000_g N_VPWR_c_778_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1002_g N_VPWR_c_779_n 0.00366111f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1000_g N_VPWR_c_772_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1002_g N_VPWR_c_772_n 0.00549784f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_184_n N_VPWR_c_772_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_185_n N_VPWR_c_772_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_174_n N_VGND_M1016_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_262 N_A_27_47#_M1010_g N_VGND_c_887_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_174_n N_VGND_c_887_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_177_n N_VGND_c_887_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_180_n N_VGND_c_887_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1015_g N_VGND_c_888_n 0.00183847f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_326_p N_VGND_c_892_n 0.00713694f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_174_n N_VGND_c_892_n 0.00243651f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1010_g N_VGND_c_893_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_172_n N_VGND_c_894_n 0.00125974f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1015_g N_VGND_c_894_n 0.00425347f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_176_n N_VGND_c_894_n 0.00279347f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1016_s N_VGND_c_896_n 0.003754f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_274 N_A_27_47#_M1010_g N_VGND_c_896_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_172_n N_VGND_c_896_n 0.00214803f $X=2.725 $Y=0.73 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1015_g N_VGND_c_896_n 0.00620714f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_326_p N_VGND_c_896_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_174_n N_VGND_c_896_n 0.00549708f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_176_n N_VGND_c_896_n 0.00520594f $X=2.95 $Y=0.887 $X2=0
+ $Y2=0
cc_280 N_D_c_340_n N_A_299_47#_M1007_g 0.0162452f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_281 N_D_c_341_n N_A_299_47#_M1007_g 0.00370069f $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_282 N_D_c_343_n N_A_299_47#_M1007_g 5.33326e-19 $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_283 N_D_c_343_n N_A_299_47#_c_397_n 0.0111849f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_284 N_D_c_344_n N_A_299_47#_c_397_n 7.68839e-19 $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_285 N_D_c_339_n N_A_299_47#_M1011_g 0.00858502f $X=1.66 $Y=1.62 $X2=0 $Y2=0
cc_286 N_D_c_347_n N_A_299_47#_M1011_g 0.0168373f $X=1.83 $Y=1.695 $X2=0 $Y2=0
cc_287 N_D_c_346_n N_A_299_47#_c_405_n 0.00860661f $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_288 N_D_c_347_n N_A_299_47#_c_405_n 0.0097543f $X=1.83 $Y=1.695 $X2=0 $Y2=0
cc_289 N_D_c_340_n N_A_299_47#_c_399_n 0.00669663f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_290 N_D_c_341_n N_A_299_47#_c_399_n 0.00844874f $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_291 N_D_c_344_n N_A_299_47#_c_399_n 0.00439477f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_292 N_D_c_341_n N_A_299_47#_c_400_n 0.00266829f $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_293 N_D_c_343_n N_A_299_47#_c_400_n 0.00226522f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_294 N_D_c_344_n N_A_299_47#_c_400_n 0.0293831f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_295 N_D_c_339_n N_A_299_47#_c_401_n 0.00386135f $X=1.66 $Y=1.62 $X2=0 $Y2=0
cc_296 N_D_c_339_n N_A_299_47#_c_407_n 0.00630992f $X=1.66 $Y=1.62 $X2=0 $Y2=0
cc_297 N_D_c_341_n N_A_299_47#_c_407_n 0.00288327f $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_298 N_D_c_342_n N_A_299_47#_c_407_n 5.67148e-19 $X=1.6 $Y=1.205 $X2=0 $Y2=0
cc_299 N_D_c_347_n N_A_299_47#_c_407_n 0.00758651f $X=1.83 $Y=1.695 $X2=0 $Y2=0
cc_300 N_D_c_344_n N_A_299_47#_c_407_n 0.0218847f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_301 N_D_c_340_n N_A_299_47#_c_402_n 6.93328e-19 $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_302 N_D_c_341_n N_A_299_47#_c_402_n 0.00748673f $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_303 N_D_c_344_n N_A_299_47#_c_402_n 0.0154053f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_304 N_D_c_342_n N_A_299_47#_c_403_n 4.30918e-19 $X=1.6 $Y=1.205 $X2=0 $Y2=0
cc_305 N_D_c_339_n N_A_193_47#_c_492_n 0.00362684f $X=1.66 $Y=1.62 $X2=0 $Y2=0
cc_306 N_D_c_341_n N_A_193_47#_c_492_n 0.00351194f $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_307 N_D_c_343_n N_A_193_47#_c_492_n 8.97548e-19 $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_308 N_D_c_344_n N_A_193_47#_c_492_n 0.0224186f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_309 N_D_c_346_n N_A_193_47#_c_496_n 9.35223e-19 $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_310 N_D_c_347_n N_A_193_47#_c_496_n 2.37785e-19 $X=1.83 $Y=1.695 $X2=0 $Y2=0
cc_311 N_D_c_346_n N_A_193_47#_c_497_n 0.00269203f $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_312 N_D_c_346_n N_VPWR_c_774_n 0.00302106f $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_313 N_D_c_346_n N_VPWR_c_778_n 0.00543342f $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_314 N_D_c_346_n N_VPWR_c_772_n 0.00734866f $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_315 N_D_c_340_n N_VGND_c_888_n 0.0108532f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_316 N_D_c_340_n N_VGND_c_893_n 0.00337001f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_317 N_D_c_341_n N_VGND_c_893_n 4.6442e-19 $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_318 N_D_c_340_n N_VGND_c_896_n 0.0053254f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_319 N_D_c_341_n N_VGND_c_896_n 0.00104331f $X=1.6 $Y=0.88 $X2=0 $Y2=0
cc_320 N_A_299_47#_M1011_g N_A_193_47#_M1003_g 0.0347134f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_321 N_A_299_47#_c_405_n N_A_193_47#_c_492_n 0.00120694f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_322 N_A_299_47#_c_407_n N_A_193_47#_c_492_n 0.00924877f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_323 N_A_299_47#_c_402_n N_A_193_47#_c_492_n 0.0204455f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_324 N_A_299_47#_c_405_n N_A_193_47#_c_496_n 0.0521161f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_325 N_A_299_47#_M1011_g N_A_193_47#_c_497_n 0.00376202f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_326 N_A_299_47#_c_405_n N_A_193_47#_c_497_n 0.0218599f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_327 N_A_299_47#_c_407_n N_A_193_47#_c_497_n 0.00554627f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_328 N_A_299_47#_c_405_n N_A_193_47#_c_498_n 0.00277234f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_329 N_A_299_47#_M1011_g N_A_193_47#_c_500_n 0.00151683f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_330 N_A_299_47#_c_405_n N_A_193_47#_c_500_n 9.6273e-19 $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_331 N_A_299_47#_M1011_g N_A_193_47#_c_501_n 0.00542783f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_332 N_A_299_47#_c_405_n N_A_193_47#_c_501_n 0.0035756f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_333 N_A_299_47#_c_401_n N_A_193_47#_c_501_n 0.00654233f $X=2.03 $Y=1.495
+ $X2=0 $Y2=0
cc_334 N_A_299_47#_c_407_n N_A_193_47#_c_501_n 0.00750275f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_397_n N_A_193_47#_c_493_n 6.92043e-19 $X=2.25 $Y=1.235
+ $X2=0 $Y2=0
cc_336 N_A_299_47#_M1011_g N_A_193_47#_c_493_n 0.0223288f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_337 N_A_299_47#_M1011_g N_A_560_47#_c_694_n 5.23712e-19 $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_338 N_A_299_47#_M1007_g N_A_560_47#_c_698_n 6.71856e-19 $X=2.25 $Y=0.445
+ $X2=0 $Y2=0
cc_339 N_A_299_47#_c_397_n N_VPWR_c_774_n 2.48532e-19 $X=2.25 $Y=1.235 $X2=0
+ $Y2=0
cc_340 N_A_299_47#_M1011_g N_VPWR_c_774_n 0.0192422f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_341 N_A_299_47#_c_405_n N_VPWR_c_774_n 0.0234125f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_342 N_A_299_47#_c_407_n N_VPWR_c_774_n 0.0106739f $X=2.03 $Y=1.58 $X2=0 $Y2=0
cc_343 N_A_299_47#_c_403_n N_VPWR_c_774_n 0.00164085f $X=2.215 $Y=1.07 $X2=0
+ $Y2=0
cc_344 N_A_299_47#_c_405_n N_VPWR_c_778_n 0.0173028f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_345 N_A_299_47#_M1011_g N_VPWR_c_779_n 0.00310428f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_M1014_s N_VPWR_c_772_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_347 N_A_299_47#_M1011_g N_VPWR_c_772_n 0.00335906f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_348 N_A_299_47#_c_405_n N_VPWR_c_772_n 0.00621325f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_349 N_A_299_47#_c_399_n N_VGND_M1005_d 0.00209965f $X=1.945 $Y=0.7 $X2=0
+ $Y2=0
cc_350 N_A_299_47#_M1007_g N_VGND_c_888_n 0.00940518f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_351 N_A_299_47#_c_397_n N_VGND_c_888_n 2.98383e-19 $X=2.25 $Y=1.235 $X2=0
+ $Y2=0
cc_352 N_A_299_47#_c_399_n N_VGND_c_888_n 0.0174457f $X=1.945 $Y=0.7 $X2=0 $Y2=0
cc_353 N_A_299_47#_c_399_n N_VGND_c_893_n 0.00255672f $X=1.945 $Y=0.7 $X2=0
+ $Y2=0
cc_354 N_A_299_47#_c_402_n N_VGND_c_893_n 0.00819232f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_355 N_A_299_47#_M1007_g N_VGND_c_894_n 0.0046653f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_356 N_A_299_47#_M1005_s N_VGND_c_896_n 0.00252595f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_357 N_A_299_47#_M1007_g N_VGND_c_896_n 0.00456069f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_299_47#_c_399_n N_VGND_c_896_n 0.00976593f $X=1.945 $Y=0.7 $X2=0
+ $Y2=0
cc_359 N_A_299_47#_c_402_n N_VGND_c_896_n 0.00698341f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_360 N_A_193_47#_c_490_n N_A_715_21#_M1012_g 0.0499857f $X=3.175 $Y=0.685
+ $X2=0 $Y2=0
cc_361 N_A_193_47#_c_493_n N_A_715_21#_M1012_g 9.80014e-19 $X=2.725 $Y=1.42
+ $X2=0 $Y2=0
cc_362 N_A_193_47#_M1003_g N_A_560_47#_c_694_n 0.00524459f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_363 N_A_193_47#_c_501_n N_A_560_47#_c_694_n 0.00171185f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_364 N_A_193_47#_c_490_n N_A_560_47#_c_698_n 0.00870331f $X=3.175 $Y=0.685
+ $X2=0 $Y2=0
cc_365 N_A_193_47#_c_490_n N_A_560_47#_c_685_n 0.00567426f $X=3.175 $Y=0.685
+ $X2=0 $Y2=0
cc_366 N_A_193_47#_c_501_n N_A_560_47#_c_691_n 0.00249299f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_367 N_A_193_47#_c_491_n N_A_560_47#_c_687_n 0.00288095f $X=3.21 $Y=1.175
+ $X2=0 $Y2=0
cc_368 N_A_193_47#_c_497_n N_VPWR_M1014_d 6.81311e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_193_47#_c_499_n N_VPWR_c_773_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_M1003_g N_VPWR_c_774_n 0.00338485f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_c_497_n N_VPWR_c_774_n 0.0155454f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_372 N_A_193_47#_c_500_n N_VPWR_c_774_n 0.0013453f $X=2.53 $Y=1.87 $X2=0 $Y2=0
cc_373 N_A_193_47#_c_501_n N_VPWR_c_774_n 0.00973315f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_499_n N_VPWR_c_778_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_375 N_A_193_47#_M1003_g N_VPWR_c_779_n 0.00410595f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_376 N_A_193_47#_c_501_n N_VPWR_c_779_n 0.00482885f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_M1003_g N_VPWR_c_772_n 0.00585915f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_378 N_A_193_47#_c_497_n N_VPWR_c_772_n 0.0504141f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_498_n N_VPWR_c_772_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_380 N_A_193_47#_c_499_n N_VPWR_c_772_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_381 N_A_193_47#_c_500_n N_VPWR_c_772_n 0.0151254f $X=2.53 $Y=1.87 $X2=0 $Y2=0
cc_382 N_A_193_47#_c_501_n N_VPWR_c_772_n 0.00454439f $X=2.69 $Y=1.52 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_c_497_n A_465_369# 8.37444e-19 $X=2.385 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_384 N_A_193_47#_c_500_n A_465_369# 0.00120144f $X=2.53 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_385 N_A_193_47#_c_501_n A_465_369# 0.00371441f $X=2.69 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_386 N_A_193_47#_c_492_n N_VGND_c_893_n 0.00732874f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_387 N_A_193_47#_c_490_n N_VGND_c_894_n 0.00378965f $X=3.175 $Y=0.685 $X2=0
+ $Y2=0
cc_388 N_A_193_47#_M1010_d N_VGND_c_896_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_389 N_A_193_47#_c_490_n N_VGND_c_896_n 0.00557387f $X=3.175 $Y=0.685 $X2=0
+ $Y2=0
cc_390 N_A_193_47#_c_492_n N_VGND_c_896_n 0.00616598f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_391 N_A_715_21#_c_619_p N_A_560_47#_c_682_n 0.00397711f $X=4.38 $Y=0.425
+ $X2=0 $Y2=0
cc_392 N_A_715_21#_c_600_n N_A_560_47#_c_682_n 0.00954296f $X=4.455 $Y=0.995
+ $X2=0 $Y2=0
cc_393 N_A_715_21#_c_621_p N_A_560_47#_c_682_n 0.00329065f $X=4.417 $Y=0.72
+ $X2=0 $Y2=0
cc_394 N_A_715_21#_c_603_n N_A_560_47#_c_682_n 0.0189912f $X=5.022 $Y=0.995
+ $X2=0 $Y2=0
cc_395 N_A_715_21#_M1013_g N_A_560_47#_M1001_g 0.0207717f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_396 N_A_715_21#_c_608_n N_A_560_47#_M1001_g 0.00371851f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_397 N_A_715_21#_c_625_p N_A_560_47#_M1001_g 0.00849361f $X=4.38 $Y=2.27 $X2=0
+ $Y2=0
cc_398 N_A_715_21#_c_609_n N_A_560_47#_M1001_g 0.00723855f $X=4.455 $Y=1.535
+ $X2=0 $Y2=0
cc_399 N_A_715_21#_c_627_p N_A_560_47#_M1001_g 0.00421774f $X=4.38 $Y=1.755
+ $X2=0 $Y2=0
cc_400 N_A_715_21#_M1012_g N_A_560_47#_c_683_n 0.0168568f $X=3.65 $Y=0.445 $X2=0
+ $Y2=0
cc_401 N_A_715_21#_c_607_n N_A_560_47#_c_683_n 0.00752066f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_402 N_A_715_21#_c_608_n N_A_560_47#_c_683_n 0.00335173f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_403 N_A_715_21#_c_621_p N_A_560_47#_c_683_n 0.00278344f $X=4.417 $Y=0.72
+ $X2=0 $Y2=0
cc_404 N_A_715_21#_c_627_p N_A_560_47#_c_683_n 0.00319255f $X=4.38 $Y=1.755
+ $X2=0 $Y2=0
cc_405 N_A_715_21#_c_633_p N_A_560_47#_c_683_n 0.0161731f $X=4.455 $Y=1.16 $X2=0
+ $Y2=0
cc_406 N_A_715_21#_c_601_n N_A_560_47#_c_684_n 0.0186811f $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_407 N_A_715_21#_c_602_n N_A_560_47#_c_684_n 0.0215009f $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_408 N_A_715_21#_c_633_p N_A_560_47#_c_684_n 7.76856e-19 $X=4.455 $Y=1.16
+ $X2=0 $Y2=0
cc_409 N_A_715_21#_M1012_g N_A_560_47#_c_698_n 0.00453048f $X=3.65 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_715_21#_M1012_g N_A_560_47#_c_685_n 0.021917f $X=3.65 $Y=0.445 $X2=0
+ $Y2=0
cc_411 N_A_715_21#_M1012_g N_A_560_47#_c_691_n 0.00499902f $X=3.65 $Y=0.445
+ $X2=0 $Y2=0
cc_412 N_A_715_21#_M1004_g N_A_560_47#_c_691_n 0.0192147f $X=3.65 $Y=2.275 $X2=0
+ $Y2=0
cc_413 N_A_715_21#_c_607_n N_A_560_47#_c_691_n 0.0251783f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_414 N_A_715_21#_c_608_n N_A_560_47#_c_691_n 0.00913418f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_415 N_A_715_21#_c_625_p N_A_560_47#_c_691_n 0.00604896f $X=4.38 $Y=2.27 $X2=0
+ $Y2=0
cc_416 N_A_715_21#_M1012_g N_A_560_47#_c_686_n 0.0135129f $X=3.65 $Y=0.445 $X2=0
+ $Y2=0
cc_417 N_A_715_21#_c_607_n N_A_560_47#_c_686_n 0.0257843f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_418 N_A_715_21#_c_608_n N_A_560_47#_c_686_n 0.0073464f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_419 N_A_715_21#_c_633_p N_A_560_47#_c_686_n 0.0277655f $X=4.455 $Y=1.16 $X2=0
+ $Y2=0
cc_420 N_A_715_21#_M1012_g N_A_560_47#_c_687_n 0.0135786f $X=3.65 $Y=0.445 $X2=0
+ $Y2=0
cc_421 N_A_715_21#_M1004_g N_VPWR_c_775_n 0.00456783f $X=3.65 $Y=2.275 $X2=0
+ $Y2=0
cc_422 N_A_715_21#_c_607_n N_VPWR_c_775_n 0.0136604f $X=4.295 $Y=1.7 $X2=0 $Y2=0
cc_423 N_A_715_21#_c_608_n N_VPWR_c_775_n 0.00604449f $X=3.9 $Y=1.7 $X2=0 $Y2=0
cc_424 N_A_715_21#_c_625_p N_VPWR_c_775_n 0.0184545f $X=4.38 $Y=2.27 $X2=0 $Y2=0
cc_425 N_A_715_21#_M1013_g N_VPWR_c_776_n 0.0185361f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_A_715_21#_c_601_n N_VPWR_c_776_n 0.0161993f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A_715_21#_c_602_n N_VPWR_c_776_n 0.00202662f $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_428 N_A_715_21#_M1004_g N_VPWR_c_779_n 0.00498701f $X=3.65 $Y=2.275 $X2=0
+ $Y2=0
cc_429 N_A_715_21#_c_625_p N_VPWR_c_780_n 0.012607f $X=4.38 $Y=2.27 $X2=0 $Y2=0
cc_430 N_A_715_21#_M1013_g N_VPWR_c_781_n 0.0046653f $X=5.05 $Y=1.985 $X2=0
+ $Y2=0
cc_431 N_A_715_21#_M1001_s N_VPWR_c_772_n 0.00238199f $X=4.255 $Y=1.485 $X2=0
+ $Y2=0
cc_432 N_A_715_21#_M1004_g N_VPWR_c_772_n 0.00974648f $X=3.65 $Y=2.275 $X2=0
+ $Y2=0
cc_433 N_A_715_21#_M1013_g N_VPWR_c_772_n 0.008846f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_434 N_A_715_21#_c_607_n N_VPWR_c_772_n 0.00834132f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_435 N_A_715_21#_c_608_n N_VPWR_c_772_n 0.00110429f $X=3.9 $Y=1.7 $X2=0 $Y2=0
cc_436 N_A_715_21#_c_625_p N_VPWR_c_772_n 0.00909897f $X=4.38 $Y=2.27 $X2=0
+ $Y2=0
cc_437 N_A_715_21#_M1013_g N_Q_c_872_n 0.0102086f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_438 N_A_715_21#_c_601_n N_Q_c_872_n 0.02621f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_439 N_A_715_21#_c_602_n N_Q_c_872_n 0.00793017f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_440 N_A_715_21#_c_603_n N_Q_c_872_n 0.00828285f $X=5.022 $Y=0.995 $X2=0 $Y2=0
cc_441 N_A_715_21#_M1012_g N_VGND_c_889_n 0.00451776f $X=3.65 $Y=0.445 $X2=0
+ $Y2=0
cc_442 N_A_715_21#_c_619_p N_VGND_c_889_n 0.0170259f $X=4.38 $Y=0.425 $X2=0
+ $Y2=0
cc_443 N_A_715_21#_c_619_p N_VGND_c_890_n 0.0144146f $X=4.38 $Y=0.425 $X2=0
+ $Y2=0
cc_444 N_A_715_21#_c_619_p N_VGND_c_891_n 0.0279714f $X=4.38 $Y=0.425 $X2=0
+ $Y2=0
cc_445 N_A_715_21#_c_601_n N_VGND_c_891_n 0.011251f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_446 N_A_715_21#_c_602_n N_VGND_c_891_n 0.00196734f $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_447 N_A_715_21#_c_603_n N_VGND_c_891_n 0.0150774f $X=5.022 $Y=0.995 $X2=0
+ $Y2=0
cc_448 N_A_715_21#_M1012_g N_VGND_c_894_n 0.00544232f $X=3.65 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_715_21#_c_603_n N_VGND_c_895_n 0.00564095f $X=5.022 $Y=0.995 $X2=0
+ $Y2=0
cc_450 N_A_715_21#_M1006_s N_VGND_c_896_n 0.00351772f $X=4.255 $Y=0.235 $X2=0
+ $Y2=0
cc_451 N_A_715_21#_M1012_g N_VGND_c_896_n 0.0110078f $X=3.65 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_715_21#_c_619_p N_VGND_c_896_n 0.00912528f $X=4.38 $Y=0.425 $X2=0
+ $Y2=0
cc_453 N_A_715_21#_c_603_n N_VGND_c_896_n 0.0104943f $X=5.022 $Y=0.995 $X2=0
+ $Y2=0
cc_454 N_A_560_47#_c_694_n N_VPWR_c_774_n 0.00549517f $X=3.295 $Y=2.34 $X2=0
+ $Y2=0
cc_455 N_A_560_47#_M1001_g N_VPWR_c_775_n 0.00201034f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_456 N_A_560_47#_M1001_g N_VPWR_c_776_n 0.00248304f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_457 N_A_560_47#_c_694_n N_VPWR_c_779_n 0.023646f $X=3.295 $Y=2.34 $X2=0 $Y2=0
cc_458 N_A_560_47#_c_691_n N_VPWR_c_779_n 0.0160426f $X=3.55 $Y=2.01 $X2=0 $Y2=0
cc_459 N_A_560_47#_M1001_g N_VPWR_c_780_n 0.00549943f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_460 N_A_560_47#_M1003_d N_VPWR_c_772_n 0.00217615f $X=2.8 $Y=2.065 $X2=0
+ $Y2=0
cc_461 N_A_560_47#_M1001_g N_VPWR_c_772_n 0.0112391f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_462 N_A_560_47#_c_694_n N_VPWR_c_772_n 0.0188931f $X=3.295 $Y=2.34 $X2=0
+ $Y2=0
cc_463 N_A_560_47#_c_691_n N_VPWR_c_772_n 0.0124455f $X=3.55 $Y=2.01 $X2=0 $Y2=0
cc_464 N_A_560_47#_c_694_n A_644_413# 3.96979e-19 $X=3.295 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_465 N_A_560_47#_c_691_n A_644_413# 0.00655118f $X=3.55 $Y=2.01 $X2=-0.19
+ $Y2=-0.24
cc_466 N_A_560_47#_c_698_n N_VGND_c_888_n 0.00235802f $X=3.435 $Y=0.45 $X2=0
+ $Y2=0
cc_467 N_A_560_47#_c_682_n N_VGND_c_889_n 0.00246239f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_468 N_A_560_47#_c_683_n N_VGND_c_889_n 0.00123674f $X=4.515 $Y=1.16 $X2=0
+ $Y2=0
cc_469 N_A_560_47#_c_686_n N_VGND_c_889_n 0.011199f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_470 N_A_560_47#_c_682_n N_VGND_c_890_n 0.00549117f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_471 N_A_560_47#_c_682_n N_VGND_c_891_n 0.00512998f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_560_47#_c_698_n N_VGND_c_894_n 0.0277584f $X=3.435 $Y=0.45 $X2=0
+ $Y2=0
cc_473 N_A_560_47#_M1015_d N_VGND_c_896_n 0.00254978f $X=2.8 $Y=0.235 $X2=0
+ $Y2=0
cc_474 N_A_560_47#_c_682_n N_VGND_c_896_n 0.011316f $X=4.59 $Y=0.995 $X2=0 $Y2=0
cc_475 N_A_560_47#_c_698_n N_VGND_c_896_n 0.0283424f $X=3.435 $Y=0.45 $X2=0
+ $Y2=0
cc_476 N_A_560_47#_c_698_n A_650_47# 0.00734648f $X=3.435 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_477 N_A_560_47#_c_685_n A_650_47# 0.00139441f $X=3.52 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_478 N_VPWR_c_772_n A_465_369# 0.00356403f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_479 N_VPWR_c_772_n A_644_413# 0.00288164f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_480 N_VPWR_c_772_n N_Q_M1013_d 0.00383158f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_481 N_VPWR_c_781_n Q 0.0169196f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_482 N_VPWR_c_772_n Q 0.00988906f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_c_776_n N_Q_c_872_n 0.0052414f $X=4.84 $Y=1.735 $X2=0 $Y2=0
cc_484 Q N_VGND_c_895_n 0.00867248f $X=5.23 $Y=0.425 $X2=0 $Y2=0
cc_485 N_Q_M1008_d N_VGND_c_896_n 0.00405593f $X=5.125 $Y=0.235 $X2=0 $Y2=0
cc_486 Q N_VGND_c_896_n 0.00898293f $X=5.23 $Y=0.425 $X2=0 $Y2=0
cc_487 N_VGND_c_896_n A_465_47# 0.0112288f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24
cc_488 N_VGND_c_896_n A_650_47# 0.00276125f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__fahcon_1.pxi.spice
* Created: Thu Aug 27 14:21:38 2020
* 
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_67_199# N_A_67_199#_M1023_d N_A_67_199#_M1015_s
+ N_A_67_199#_M1017_d N_A_67_199#_M1010_d N_A_67_199#_M1019_d
+ N_A_67_199#_M1012_g N_A_67_199#_M1018_g N_A_67_199#_c_209_n
+ N_A_67_199#_c_216_n N_A_67_199#_c_210_n N_A_67_199#_c_231_p
+ N_A_67_199#_c_319_p N_A_67_199#_c_226_p N_A_67_199#_c_227_p
+ N_A_67_199#_c_211_n N_A_67_199#_c_217_n N_A_67_199#_c_218_n
+ N_A_67_199#_c_212_n N_A_67_199#_c_239_p N_A_67_199#_c_220_n
+ N_A_67_199#_c_221_n N_A_67_199#_c_222_n N_A_67_199#_c_223_n
+ N_A_67_199#_c_255_p N_A_67_199#_c_213_n PM_SKY130_FD_SC_HD__FAHCON_1%A_67_199#
x_PM_SKY130_FD_SC_HD__FAHCON_1%A N_A_c_384_n N_A_M1023_g N_A_M1017_g A
+ N_A_c_386_n PM_SKY130_FD_SC_HD__FAHCON_1%A
x_PM_SKY130_FD_SC_HD__FAHCON_1%B N_B_c_428_n N_B_M1009_g N_B_M1028_g N_B_M1019_g
+ N_B_M1031_g N_B_M1000_g N_B_c_429_n N_B_M1027_g N_B_c_430_n N_B_c_431_n
+ N_B_M1005_g N_B_M1001_g N_B_c_432_n N_B_c_433_n N_B_c_434_n N_B_c_435_n
+ N_B_c_436_n N_B_c_437_n N_B_c_438_n B N_B_c_440_n N_B_c_441_n B N_B_c_442_n
+ N_B_c_443_n PM_SKY130_FD_SC_HD__FAHCON_1%B
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_488_21# N_A_488_21#_M1027_s N_A_488_21#_M1000_s
+ N_A_488_21#_c_607_n N_A_488_21#_M1002_g N_A_488_21#_M1010_g
+ N_A_488_21#_c_608_n N_A_488_21#_M1015_g N_A_488_21#_M1014_g
+ N_A_488_21#_c_609_n N_A_488_21#_c_610_n N_A_488_21#_c_611_n
+ N_A_488_21#_c_612_n N_A_488_21#_c_650_n N_A_488_21#_c_618_n
+ N_A_488_21#_c_619_n N_A_488_21#_c_670_p N_A_488_21#_c_620_n
+ N_A_488_21#_c_621_n N_A_488_21#_c_622_n PM_SKY130_FD_SC_HD__FAHCON_1%A_488_21#
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_434_49# N_A_434_49#_M1009_d N_A_434_49#_M1028_d
+ N_A_434_49#_M1025_g N_A_434_49#_c_727_n N_A_434_49#_M1013_g
+ N_A_434_49#_M1008_g N_A_434_49#_M1022_g N_A_434_49#_c_728_n
+ N_A_434_49#_c_750_n N_A_434_49#_c_729_n N_A_434_49#_c_730_n
+ N_A_434_49#_c_731_n N_A_434_49#_c_732_n N_A_434_49#_c_733_n
+ N_A_434_49#_c_734_n N_A_434_49#_c_735_n N_A_434_49#_c_736_n
+ N_A_434_49#_c_737_n PM_SKY130_FD_SC_HD__FAHCON_1%A_434_49#
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_726_47# N_A_726_47#_M1015_d N_A_726_47#_M1014_d
+ N_A_726_47#_M1004_g N_A_726_47#_c_903_n N_A_726_47#_M1029_g
+ N_A_726_47#_c_904_n N_A_726_47#_M1007_g N_A_726_47#_c_912_n
+ N_A_726_47#_M1024_g N_A_726_47#_c_905_n N_A_726_47#_c_906_n
+ N_A_726_47#_c_907_n N_A_726_47#_c_916_n N_A_726_47#_c_917_n
+ N_A_726_47#_c_918_n N_A_726_47#_c_908_n N_A_726_47#_c_932_n
+ N_A_726_47#_c_947_n N_A_726_47#_c_933_n N_A_726_47#_c_952_n
+ N_A_726_47#_c_919_n N_A_726_47#_c_953_n N_A_726_47#_c_920_n
+ N_A_726_47#_c_909_n N_A_726_47#_c_910_n N_A_726_47#_c_923_n
+ PM_SKY130_FD_SC_HD__FAHCON_1%A_726_47#
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_1589_49# N_A_1589_49#_M1007_s
+ N_A_1589_49#_M1003_d N_A_1589_49#_M1022_d N_A_1589_49#_M1016_d
+ N_A_1589_49#_M1020_g N_A_1589_49#_M1030_g N_A_1589_49#_c_1108_n
+ N_A_1589_49#_c_1094_n N_A_1589_49#_c_1095_n N_A_1589_49#_c_1096_n
+ N_A_1589_49#_c_1097_n N_A_1589_49#_c_1173_p N_A_1589_49#_c_1098_n
+ N_A_1589_49#_c_1104_n N_A_1589_49#_c_1105_n N_A_1589_49#_c_1160_p
+ N_A_1589_49#_c_1099_n N_A_1589_49#_c_1100_n N_A_1589_49#_c_1107_n
+ PM_SKY130_FD_SC_HD__FAHCON_1%A_1589_49#
x_PM_SKY130_FD_SC_HD__FAHCON_1%CI N_CI_M1016_g N_CI_c_1242_n N_CI_M1003_g
+ N_CI_c_1243_n N_CI_M1026_g N_CI_M1021_g N_CI_c_1244_n N_CI_c_1245_n
+ N_CI_c_1246_n CI PM_SKY130_FD_SC_HD__FAHCON_1%CI
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_1710_49# N_A_1710_49#_M1007_d
+ N_A_1710_49#_M1024_d N_A_1710_49#_M1011_g N_A_1710_49#_M1006_g
+ N_A_1710_49#_c_1307_n N_A_1710_49#_c_1313_n N_A_1710_49#_c_1329_n
+ N_A_1710_49#_c_1348_n N_A_1710_49#_c_1330_n N_A_1710_49#_c_1314_n
+ N_A_1710_49#_c_1315_n N_A_1710_49#_c_1316_n N_A_1710_49#_c_1308_n
+ N_A_1710_49#_c_1309_n N_A_1710_49#_c_1310_n
+ PM_SKY130_FD_SC_HD__FAHCON_1%A_1710_49#
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_28_47# N_A_28_47#_M1012_s N_A_28_47#_M1002_d
+ N_A_28_47#_M1031_d N_A_28_47#_M1018_s N_A_28_47#_M1028_s N_A_28_47#_M1014_s
+ N_A_28_47#_c_1431_n N_A_28_47#_c_1425_n N_A_28_47#_c_1446_n
+ N_A_28_47#_c_1455_n N_A_28_47#_c_1490_n N_A_28_47#_c_1432_n
+ N_A_28_47#_c_1433_n N_A_28_47#_c_1426_n N_A_28_47#_c_1464_n
+ N_A_28_47#_c_1465_n N_A_28_47#_c_1427_n N_A_28_47#_c_1435_n
+ N_A_28_47#_c_1428_n N_A_28_47#_c_1437_n N_A_28_47#_c_1438_n
+ N_A_28_47#_c_1429_n N_A_28_47#_c_1430_n N_A_28_47#_c_1505_n
+ PM_SKY130_FD_SC_HD__FAHCON_1%A_28_47#
x_PM_SKY130_FD_SC_HD__FAHCON_1%VPWR N_VPWR_M1018_d N_VPWR_M1000_d N_VPWR_M1030_d
+ N_VPWR_M1021_d N_VPWR_c_1578_n N_VPWR_c_1579_n N_VPWR_c_1580_n N_VPWR_c_1581_n
+ N_VPWR_c_1582_n VPWR N_VPWR_c_1583_n N_VPWR_c_1584_n N_VPWR_c_1585_n
+ N_VPWR_c_1586_n N_VPWR_c_1577_n N_VPWR_c_1588_n N_VPWR_c_1589_n
+ N_VPWR_c_1590_n N_VPWR_c_1591_n PM_SKY130_FD_SC_HD__FAHCON_1%VPWR
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_1144_49# N_A_1144_49#_M1005_d
+ N_A_1144_49#_M1029_d N_A_1144_49#_M1001_d N_A_1144_49#_c_1710_n
+ N_A_1144_49#_c_1706_n N_A_1144_49#_c_1724_n N_A_1144_49#_c_1714_n
+ N_A_1144_49#_c_1730_n N_A_1144_49#_c_1707_n N_A_1144_49#_c_1709_n
+ N_A_1144_49#_c_1715_n N_A_1144_49#_c_1716_n
+ PM_SKY130_FD_SC_HD__FAHCON_1%A_1144_49#
x_PM_SKY130_FD_SC_HD__FAHCON_1%COUT_N N_COUT_N_M1013_d N_COUT_N_M1025_d COUT_N
+ COUT_N N_COUT_N_c_1780_n COUT_N PM_SKY130_FD_SC_HD__FAHCON_1%COUT_N
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_1261_49# N_A_1261_49#_M1013_s
+ N_A_1261_49#_M1026_s N_A_1261_49#_M1004_d N_A_1261_49#_M1021_s
+ N_A_1261_49#_c_1807_n N_A_1261_49#_c_1837_n N_A_1261_49#_c_1813_n
+ N_A_1261_49#_c_1814_n N_A_1261_49#_c_1857_n N_A_1261_49#_c_1808_n
+ N_A_1261_49#_c_1815_n N_A_1261_49#_c_1858_n N_A_1261_49#_c_1809_n
+ N_A_1261_49#_c_1810_n N_A_1261_49#_c_1811_n N_A_1261_49#_c_1870_n
+ N_A_1261_49#_c_1812_n PM_SKY130_FD_SC_HD__FAHCON_1%A_1261_49#
x_PM_SKY130_FD_SC_HD__FAHCON_1%A_1634_315# N_A_1634_315#_M1008_d
+ N_A_1634_315#_M1024_s N_A_1634_315#_M1030_s N_A_1634_315#_c_1942_n
+ N_A_1634_315#_c_1939_n N_A_1634_315#_c_1940_n N_A_1634_315#_c_1944_n
+ N_A_1634_315#_c_1961_n N_A_1634_315#_c_1964_n N_A_1634_315#_c_1968_n
+ N_A_1634_315#_c_1938_n PM_SKY130_FD_SC_HD__FAHCON_1%A_1634_315#
x_PM_SKY130_FD_SC_HD__FAHCON_1%SUM N_SUM_M1006_d N_SUM_M1011_d SUM SUM SUM SUM
+ SUM SUM N_SUM_c_1997_n PM_SKY130_FD_SC_HD__FAHCON_1%SUM
x_PM_SKY130_FD_SC_HD__FAHCON_1%VGND N_VGND_M1012_d N_VGND_M1027_d N_VGND_M1020_d
+ N_VGND_M1026_d N_VGND_c_2015_n N_VGND_c_2016_n N_VGND_c_2017_n N_VGND_c_2018_n
+ VGND N_VGND_c_2019_n N_VGND_c_2020_n N_VGND_c_2021_n N_VGND_c_2022_n
+ N_VGND_c_2023_n N_VGND_c_2024_n N_VGND_c_2025_n N_VGND_c_2026_n
+ N_VGND_c_2027_n PM_SKY130_FD_SC_HD__FAHCON_1%VGND
cc_1 VNB N_A_67_199#_c_209_n 0.00625651f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.325
cc_2 VNB N_A_67_199#_c_210_n 0.00333527f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.82
cc_3 VNB N_A_67_199#_c_211_n 0.00591028f $X=-0.19 $Y=-0.24 $X2=3.24 $Y2=0.36
cc_4 VNB N_A_67_199#_c_212_n 0.026083f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_5 VNB N_A_67_199#_c_213_n 0.0205236f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_6 VNB N_A_c_384_n 0.020424f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.235
cc_7 VNB A 0.00179467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_c_386_n 0.0300339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_c_428_n 0.0202452f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.235
cc_10 VNB N_B_c_429_n 0.0197241f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.325
cc_11 VNB N_B_c_430_n 0.0150305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_431_n 0.0199356f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.5
cc_13 VNB N_B_c_432_n 0.0343277f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_14 VNB N_B_c_433_n 0.00893089f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_15 VNB N_B_c_434_n 0.0181943f $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=0.36
cc_16 VNB N_B_c_435_n 0.021911f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.36
cc_17 VNB N_B_c_436_n 0.0481181f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.96
cc_18 VNB N_B_c_437_n 0.005593f $X=-0.19 $Y=-0.24 $X2=2.725 $Y2=1.96
cc_19 VNB N_B_c_438_n 0.0123608f $X=-0.19 $Y=-0.24 $X2=2.725 $Y2=1.96
cc_20 VNB B 0.00422851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B_c_440_n 0.00527227f $X=-0.19 $Y=-0.24 $X2=0.602 $Y2=1.16
cc_22 VNB N_B_c_441_n 0.00284671f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_23 VNB N_B_c_442_n 8.60476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_B_c_443_n 7.51502e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_488_21#_c_607_n 0.0206704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_488_21#_c_608_n 0.0233256f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_488_21#_c_609_n 0.00892974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_488_21#_c_610_n 0.0462984f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.325
cc_29 VNB N_A_488_21#_c_611_n 0.0139107f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.5
cc_30 VNB N_A_488_21#_c_612_n 0.00187979f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.585
cc_31 VNB N_A_434_49#_c_727_n 0.0189404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_434_49#_c_728_n 0.00827173f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_33 VNB N_A_434_49#_c_729_n 0.0035785f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.325
cc_34 VNB N_A_434_49#_c_730_n 0.00285941f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.5
cc_35 VNB N_A_434_49#_c_731_n 0.00626672f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_36 VNB N_A_434_49#_c_732_n 0.00194186f $X=-0.19 $Y=-0.24 $X2=3.24 $Y2=0.36
cc_37 VNB N_A_434_49#_c_733_n 0.0360802f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_38 VNB N_A_434_49#_c_734_n 0.0276015f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_39 VNB N_A_434_49#_c_735_n 0.00324736f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.36
cc_40 VNB N_A_434_49#_c_736_n 0.020976f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.38
cc_41 VNB N_A_434_49#_c_737_n 7.72485e-19 $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.665
cc_42 VNB N_A_726_47#_c_903_n 0.020289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_726_47#_c_904_n 0.0209104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_726_47#_c_905_n 0.0133977f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_45 VNB N_A_726_47#_c_906_n 0.0519294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_726_47#_c_907_n 0.0299111f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.325
cc_47 VNB N_A_726_47#_c_908_n 0.00273809f $X=-0.19 $Y=-0.24 $X2=3.24 $Y2=0.36
cc_48 VNB N_A_726_47#_c_909_n 0.00151294f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.67
cc_49 VNB N_A_726_47#_c_910_n 0.00385168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1589_49#_c_1094_n 0.00827772f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.82
cc_51 VNB N_A_1589_49#_c_1095_n 0.00311702f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_52 VNB N_A_1589_49#_c_1096_n 0.00517348f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.735
cc_53 VNB N_A_1589_49#_c_1097_n 0.00423574f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_54 VNB N_A_1589_49#_c_1098_n 0.00589542f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.96
cc_55 VNB N_A_1589_49#_c_1099_n 0.0224911f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.665
cc_56 VNB N_A_1589_49#_c_1100_n 0.0202796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_CI_c_1242_n 0.0207742f $X=-0.19 $Y=-0.24 $X2=4.16 $Y2=1.61
cc_58 VNB N_CI_c_1243_n 0.0206681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_CI_c_1244_n 0.0116244f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_60 VNB N_CI_c_1245_n 0.0437832f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.555
cc_61 VNB N_CI_c_1246_n 0.0101793f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.555
cc_62 VNB N_A_1710_49#_c_1307_n 0.00258682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1710_49#_c_1308_n 0.0226007f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.36
cc_64 VNB N_A_1710_49#_c_1309_n 0.00585462f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.38
cc_65 VNB N_A_1710_49#_c_1310_n 0.0201404f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.96
cc_66 VNB N_A_28_47#_c_1425_n 0.0188266f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.585
cc_67 VNB N_A_28_47#_c_1426_n 0.00133361f $X=-0.19 $Y=-0.24 $X2=0.602 $Y2=1.16
cc_68 VNB N_A_28_47#_c_1427_n 0.00297172f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.585
cc_69 VNB N_A_28_47#_c_1428_n 0.0227417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_28_47#_c_1429_n 0.00923293f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.87
cc_71 VNB N_A_28_47#_c_1430_n 0.00372175f $X=-0.19 $Y=-0.24 $X2=4.295 $Y2=1.87
cc_72 VNB N_VPWR_c_1577_n 0.516438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1144_49#_c_1706_n 0.00834334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1144_49#_c_1707_n 0.00120965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB COUT_N 0.00193947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_COUT_N_c_1780_n 8.43544e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1261_49#_c_1807_n 0.00556039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1261_49#_c_1808_n 0.0044801f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.465
cc_79 VNB N_A_1261_49#_c_1809_n 0.0198906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1261_49#_c_1810_n 0.00445149f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_81 VNB N_A_1261_49#_c_1811_n 0.0128096f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_82 VNB N_A_1261_49#_c_1812_n 0.00135949f $X=-0.19 $Y=-0.24 $X2=1.365
+ $Y2=1.585
cc_83 VNB N_A_1634_315#_c_1938_n 0.00801383f $X=-0.19 $Y=-0.24 $X2=1.28
+ $Y2=1.585
cc_84 VNB SUM 0.0294705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_SUM_c_1997_n 0.0160045f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.5
cc_86 VNB N_VGND_c_2015_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.555
cc_87 VNB N_VGND_c_2016_n 0.00288723f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_88 VNB N_VGND_c_2017_n 0.00470301f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.82
cc_89 VNB N_VGND_c_2018_n 0.00545133f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.465
cc_90 VNB N_VGND_c_2019_n 0.103626f $X=-0.19 $Y=-0.24 $X2=3.24 $Y2=0.36
cc_91 VNB N_VGND_c_2020_n 0.114166f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_92 VNB N_VGND_c_2021_n 0.0311583f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.665
cc_93 VNB N_VGND_c_2022_n 0.0177767f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.87
cc_94 VNB N_VGND_c_2023_n 0.62285f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.87
cc_95 VNB N_VGND_c_2024_n 0.0220858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_2025_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=4.295 $Y2=1.87
cc_97 VNB N_VGND_c_2026_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_98 VNB N_VGND_c_2027_n 0.00554706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VPB N_A_67_199#_M1018_g 0.023979f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_100 VPB N_A_67_199#_c_209_n 0.00109618f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_101 VPB N_A_67_199#_c_216_n 0.00272323f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.5
cc_102 VPB N_A_67_199#_c_217_n 0.00222197f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.96
cc_103 VPB N_A_67_199#_c_218_n 0.0104579f $X=-0.19 $Y=1.305 $X2=2.725 $Y2=1.96
cc_104 VPB N_A_67_199#_c_212_n 0.00620175f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_105 VPB N_A_67_199#_c_220_n 0.00631565f $X=-0.19 $Y=1.305 $X2=4.15 $Y2=1.87
cc_106 VPB N_A_67_199#_c_221_n 0.00149388f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=1.87
cc_107 VPB N_A_67_199#_c_222_n 5.31139e-19 $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.87
cc_108 VPB N_A_67_199#_c_223_n 0.00346908f $X=-0.19 $Y=1.305 $X2=4.295 $Y2=1.87
cc_109 VPB N_A_M1017_g 0.0270986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_c_386_n 0.00854837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_B_M1028_g 0.0221422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_B_M1019_g 0.0348546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_B_M1000_g 0.0239944f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_114 VPB N_B_c_430_n 0.00654745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_B_M1001_g 0.0226713f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.465
cc_116 VPB N_B_c_432_n 0.0161045f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_117 VPB N_B_c_433_n 5.76186e-19 $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_118 VPB N_B_c_434_n 0.00225379f $X=-0.19 $Y=1.305 $X2=1.325 $Y2=0.36
cc_119 VPB N_B_c_436_n 0.0214716f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.96
cc_120 VPB N_B_c_437_n 3.60839e-19 $X=-0.19 $Y=1.305 $X2=2.725 $Y2=1.96
cc_121 VPB N_B_c_438_n 8.22615e-19 $X=-0.19 $Y=1.305 $X2=2.725 $Y2=1.96
cc_122 VPB B 0.00388628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_B_c_443_n 0.00287175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_488_21#_M1010_g 0.0196215f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_488_21#_M1014_g 0.021858f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_126 VPB N_A_488_21#_c_609_n 5.76112e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_488_21#_c_610_n 0.0247236f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_128 VPB N_A_488_21#_c_611_n 0.00120001f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.5
cc_129 VPB N_A_488_21#_c_618_n 0.0171974f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_130 VPB N_A_488_21#_c_619_n 0.00304619f $X=-0.19 $Y=1.305 $X2=3.24 $Y2=0.36
cc_131 VPB N_A_488_21#_c_620_n 0.00761145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_488_21#_c_621_n 0.00593283f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_133 VPB N_A_488_21#_c_622_n 9.59248e-19 $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.585
cc_134 VPB N_A_434_49#_M1025_g 0.0208531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_434_49#_M1022_g 0.0283351f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_136 VPB N_A_434_49#_c_730_n 4.7406e-19 $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.5
cc_137 VPB N_A_434_49#_c_731_n 8.12858e-19 $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_138 VPB N_A_434_49#_c_733_n 0.0115302f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_139 VPB N_A_434_49#_c_734_n 0.00581379f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_140 VPB N_A_434_49#_c_737_n 0.0062423f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.665
cc_141 VPB N_A_726_47#_M1004_g 0.0216864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_726_47#_c_912_n 0.017473f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_143 VPB N_A_726_47#_c_905_n 0.00248297f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_144 VPB N_A_726_47#_c_906_n 0.0335564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_726_47#_c_907_n 0.0385191f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_146 VPB N_A_726_47#_c_916_n 0.00370412f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.585
cc_147 VPB N_A_726_47#_c_917_n 0.0181555f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.465
cc_148 VPB N_A_726_47#_c_918_n 0.00233537f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.735
cc_149 VPB N_A_726_47#_c_919_n 0.0226589f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_150 VPB N_A_726_47#_c_920_n 0.0184882f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_151 VPB N_A_726_47#_c_909_n 0.00278828f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.67
cc_152 VPB N_A_726_47#_c_910_n 0.00179342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_726_47#_c_923_n 0.00763073f $X=-0.19 $Y=1.305 $X2=4.15 $Y2=1.87
cc_154 VPB N_A_1589_49#_M1030_g 0.0222279f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_155 VPB N_A_1589_49#_c_1094_n 0.00492816f $X=-0.19 $Y=1.305 $X2=0.995
+ $Y2=0.82
cc_156 VPB N_A_1589_49#_c_1097_n 0.00548399f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_157 VPB N_A_1589_49#_c_1104_n 0.00203469f $X=-0.19 $Y=1.305 $X2=2.725
+ $Y2=1.96
cc_158 VPB N_A_1589_49#_c_1105_n 0.00146841f $X=-0.19 $Y=1.305 $X2=2.725
+ $Y2=1.96
cc_159 VPB N_A_1589_49#_c_1099_n 0.0049967f $X=-0.19 $Y=1.305 $X2=1.365
+ $Y2=1.665
cc_160 VPB N_A_1589_49#_c_1107_n 0.00863914f $X=-0.19 $Y=1.305 $X2=3.325
+ $Y2=0.42
cc_161 VPB N_CI_M1016_g 0.0230099f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.485
cc_162 VPB N_CI_M1021_g 0.023149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_CI_c_1244_n 7.09285e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_164 VPB N_CI_c_1245_n 0.0204495f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_165 VPB N_CI_c_1246_n 6.56727e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_166 VPB N_A_1710_49#_M1011_g 0.0220957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_1710_49#_c_1307_n 0.00140835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1710_49#_c_1313_n 0.00387345f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=0.995
cc_169 VPB N_A_1710_49#_c_1314_n 0.022756f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.5
cc_170 VPB N_A_1710_49#_c_1315_n 0.00164955f $X=-0.19 $Y=1.305 $X2=0.995
+ $Y2=0.82
cc_171 VPB N_A_1710_49#_c_1316_n 0.00131607f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_172 VPB N_A_1710_49#_c_1308_n 0.00600825f $X=-0.19 $Y=1.305 $X2=1.885
+ $Y2=0.36
cc_173 VPB N_A_1710_49#_c_1309_n 0.00253093f $X=-0.19 $Y=1.305 $X2=1.885
+ $Y2=0.38
cc_174 VPB N_A_28_47#_c_1431_n 0.0183122f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_175 VPB N_A_28_47#_c_1432_n 0.0114055f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.96
cc_176 VPB N_A_28_47#_c_1433_n 7.77626e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_28_47#_c_1426_n 0.00212054f $X=-0.19 $Y=1.305 $X2=0.602 $Y2=1.16
cc_178 VPB N_A_28_47#_c_1435_n 0.0201963f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.875
cc_179 VPB N_A_28_47#_c_1428_n 0.00898972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_28_47#_c_1437_n 0.0102409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_28_47#_c_1438_n 0.00240158f $X=-0.19 $Y=1.305 $X2=4.15 $Y2=1.87
cc_182 VPB N_VPWR_c_1578_n 0.00465796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1579_n 0.106101f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_184 VPB N_VPWR_c_1580_n 0.00276876f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_185 VPB N_VPWR_c_1581_n 4.89207e-19 $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.82
cc_186 VPB N_VPWR_c_1582_n 0.00231609f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.465
cc_187 VPB N_VPWR_c_1583_n 0.0172154f $X=-0.19 $Y=1.305 $X2=3.24 $Y2=0.36
cc_188 VPB N_VPWR_c_1584_n 0.104283f $X=-0.19 $Y=1.305 $X2=2.725 $Y2=1.96
cc_189 VPB N_VPWR_c_1585_n 0.0289725f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.38
cc_190 VPB N_VPWR_c_1586_n 0.0165146f $X=-0.19 $Y=1.305 $X2=3.325 $Y2=0.42
cc_191 VPB N_VPWR_c_1577_n 0.109739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1588_n 0.00323923f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.87
cc_193 VPB N_VPWR_c_1589_n 0.00506918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1590_n 0.00442675f $X=-0.19 $Y=1.305 $X2=4.295 $Y2=1.87
cc_195 VPB N_VPWR_c_1591_n 0.0036033f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=0.995
cc_196 VPB N_A_1144_49#_c_1706_n 0.00448095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1144_49#_c_1709_n 0.00150393f $X=-0.19 $Y=1.305 $X2=0.695
+ $Y2=1.325
cc_198 VPB COUT_N 0.00104353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1261_49#_c_1813_n 0.00145761f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.325
cc_200 VPB N_A_1261_49#_c_1814_n 0.00851012f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.985
cc_201 VPB N_A_1261_49#_c_1815_n 0.00293746f $X=-0.19 $Y=1.305 $X2=1.325
+ $Y2=0.36
cc_202 VPB N_A_1261_49#_c_1812_n 0.00188532f $X=-0.19 $Y=1.305 $X2=1.365
+ $Y2=1.585
cc_203 VPB N_A_1634_315#_c_1939_n 0.0132669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1634_315#_c_1940_n 0.00185585f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1634_315#_c_1938_n 0.00373506f $X=-0.19 $Y=1.305 $X2=1.28
+ $Y2=1.585
cc_206 VPB SUM 0.0203847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB SUM 0.0283032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 N_A_67_199#_c_209_n N_A_c_384_n 0.0068634f $X=0.695 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_209 N_A_67_199#_c_210_n N_A_c_384_n 0.0105647f $X=0.995 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_210 N_A_67_199#_c_226_p N_A_c_384_n 0.00258977f $X=1.16 $Y=0.465 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_67_199#_c_227_p N_A_c_384_n 0.00439001f $X=1.16 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_212 N_A_67_199#_c_213_n N_A_c_384_n 0.0190131f $X=0.5 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_213 N_A_67_199#_M1018_g N_A_M1017_g 0.0350328f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_67_199#_c_216_n N_A_M1017_g 0.00394699f $X=0.695 $Y=1.5 $X2=0 $Y2=0
cc_215 N_A_67_199#_c_231_p N_A_M1017_g 0.0129341f $X=1.28 $Y=1.585 $X2=0 $Y2=0
cc_216 N_A_67_199#_c_217_n N_A_M1017_g 0.00107008f $X=1.45 $Y=1.96 $X2=0 $Y2=0
cc_217 N_A_67_199#_c_221_n N_A_M1017_g 0.00224374f $X=1.51 $Y=1.87 $X2=0 $Y2=0
cc_218 N_A_67_199#_c_222_n N_A_M1017_g 0.00529642f $X=1.365 $Y=1.87 $X2=0 $Y2=0
cc_219 N_A_67_199#_c_209_n A 0.0161919f $X=0.695 $Y=1.325 $X2=0 $Y2=0
cc_220 N_A_67_199#_c_210_n A 0.0298669f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_221 N_A_67_199#_c_231_p A 0.0166344f $X=1.28 $Y=1.585 $X2=0 $Y2=0
cc_222 N_A_67_199#_c_211_n A 4.10315e-19 $X=3.24 $Y=0.36 $X2=0 $Y2=0
cc_223 N_A_67_199#_c_239_p A 0.00360789f $X=1.365 $Y=1.67 $X2=0 $Y2=0
cc_224 N_A_67_199#_c_221_n A 4.23853e-19 $X=1.51 $Y=1.87 $X2=0 $Y2=0
cc_225 N_A_67_199#_c_210_n N_A_c_386_n 0.00739621f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_226 N_A_67_199#_c_231_p N_A_c_386_n 0.00510798f $X=1.28 $Y=1.585 $X2=0 $Y2=0
cc_227 N_A_67_199#_c_212_n N_A_c_386_n 0.0208492f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_67_199#_c_239_p N_A_c_386_n 7.13664e-19 $X=1.365 $Y=1.67 $X2=0 $Y2=0
cc_229 N_A_67_199#_c_227_p N_B_c_428_n 0.00298527f $X=1.16 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_230 N_A_67_199#_c_211_n N_B_c_428_n 0.00856778f $X=3.24 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_231 N_A_67_199#_c_218_n N_B_M1028_g 0.0114816f $X=2.725 $Y=1.96 $X2=0 $Y2=0
cc_232 N_A_67_199#_c_239_p N_B_M1028_g 0.00103814f $X=1.365 $Y=1.67 $X2=0 $Y2=0
cc_233 N_A_67_199#_c_220_n N_B_M1028_g 0.00280807f $X=4.15 $Y=1.87 $X2=0 $Y2=0
cc_234 N_A_67_199#_c_221_n N_B_M1028_g 8.91012e-19 $X=1.51 $Y=1.87 $X2=0 $Y2=0
cc_235 N_A_67_199#_c_222_n N_B_M1028_g 0.00310207f $X=1.365 $Y=1.87 $X2=0 $Y2=0
cc_236 N_A_67_199#_c_220_n N_B_M1019_g 0.00433663f $X=4.15 $Y=1.87 $X2=0 $Y2=0
cc_237 N_A_67_199#_c_223_n N_B_M1019_g 9.92956e-19 $X=4.295 $Y=1.87 $X2=0 $Y2=0
cc_238 N_A_67_199#_c_223_n N_B_M1000_g 0.00221665f $X=4.295 $Y=1.87 $X2=0 $Y2=0
cc_239 N_A_67_199#_c_255_p N_B_M1000_g 0.00210622f $X=4.295 $Y=1.87 $X2=0 $Y2=0
cc_240 N_A_67_199#_c_211_n N_B_c_432_n 0.00588727f $X=3.24 $Y=0.36 $X2=0 $Y2=0
cc_241 N_A_67_199#_c_218_n N_B_c_432_n 0.00500074f $X=2.725 $Y=1.96 $X2=0 $Y2=0
cc_242 N_A_67_199#_c_220_n N_B_c_432_n 0.00350789f $X=4.15 $Y=1.87 $X2=0 $Y2=0
cc_243 N_A_67_199#_c_255_p N_B_c_434_n 9.81759e-19 $X=4.295 $Y=1.87 $X2=0 $Y2=0
cc_244 N_A_67_199#_M1023_d B 0.00712543f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_245 N_A_67_199#_c_210_n B 0.0110733f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_246 N_A_67_199#_c_227_p B 0.00181773f $X=1.16 $Y=0.72 $X2=0 $Y2=0
cc_247 N_A_67_199#_c_211_n B 0.0131806f $X=3.24 $Y=0.36 $X2=0 $Y2=0
cc_248 N_A_67_199#_c_218_n B 0.00496235f $X=2.725 $Y=1.96 $X2=0 $Y2=0
cc_249 N_A_67_199#_c_220_n B 0.00586246f $X=4.15 $Y=1.87 $X2=0 $Y2=0
cc_250 N_A_67_199#_M1023_d N_B_c_440_n 0.00149043f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_251 N_A_67_199#_c_211_n N_B_c_440_n 0.0138827f $X=3.24 $Y=0.36 $X2=0 $Y2=0
cc_252 N_A_67_199#_M1023_d N_B_c_441_n 0.00163049f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_253 N_A_67_199#_c_210_n N_B_c_441_n 0.00585767f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_254 N_A_67_199#_c_211_n N_B_c_441_n 0.00242222f $X=3.24 $Y=0.36 $X2=0 $Y2=0
cc_255 N_A_67_199#_c_255_p N_B_c_443_n 0.00245985f $X=4.295 $Y=1.87 $X2=0 $Y2=0
cc_256 N_A_67_199#_c_211_n N_A_488_21#_c_607_n 0.0170367f $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_257 N_A_67_199#_c_218_n N_A_488_21#_M1010_g 0.00951573f $X=2.725 $Y=1.96
+ $X2=0 $Y2=0
cc_258 N_A_67_199#_c_220_n N_A_488_21#_M1010_g 0.00258762f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_259 N_A_67_199#_c_220_n N_A_488_21#_M1014_g 0.00637693f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_260 N_A_67_199#_c_211_n N_A_488_21#_c_610_n 5.76737e-19 $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_261 N_A_67_199#_c_218_n N_A_488_21#_c_610_n 7.35213e-19 $X=2.725 $Y=1.96
+ $X2=0 $Y2=0
cc_262 N_A_67_199#_c_220_n N_A_488_21#_c_618_n 0.0779927f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_263 N_A_67_199#_c_223_n N_A_488_21#_c_618_n 0.0267379f $X=4.295 $Y=1.87 $X2=0
+ $Y2=0
cc_264 N_A_67_199#_c_255_p N_A_488_21#_c_618_n 8.7652e-19 $X=4.295 $Y=1.87 $X2=0
+ $Y2=0
cc_265 N_A_67_199#_M1010_d N_A_488_21#_c_619_n 3.52047e-19 $X=2.59 $Y=1.485
+ $X2=0 $Y2=0
cc_266 N_A_67_199#_c_218_n N_A_488_21#_c_619_n 2.41221e-19 $X=2.725 $Y=1.96
+ $X2=0 $Y2=0
cc_267 N_A_67_199#_c_220_n N_A_488_21#_c_619_n 0.0303498f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_268 N_A_67_199#_M1010_d N_A_488_21#_c_621_n 0.00362735f $X=2.59 $Y=1.485
+ $X2=0 $Y2=0
cc_269 N_A_67_199#_c_218_n N_A_488_21#_c_621_n 0.0122649f $X=2.725 $Y=1.96 $X2=0
+ $Y2=0
cc_270 N_A_67_199#_c_220_n N_A_488_21#_c_621_n 0.00408223f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_271 N_A_67_199#_c_211_n N_A_434_49#_M1009_d 0.00305293f $X=3.24 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_272 N_A_67_199#_c_218_n N_A_434_49#_M1028_d 0.00234544f $X=2.725 $Y=1.96
+ $X2=0 $Y2=0
cc_273 N_A_67_199#_c_220_n N_A_434_49#_M1028_d 0.00178317f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_274 N_A_67_199#_c_218_n N_A_434_49#_c_728_n 0.00176169f $X=2.725 $Y=1.96
+ $X2=0 $Y2=0
cc_275 N_A_67_199#_c_220_n N_A_434_49#_c_728_n 0.0271339f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_276 N_A_67_199#_c_218_n N_A_434_49#_c_750_n 4.53831e-19 $X=2.725 $Y=1.96
+ $X2=0 $Y2=0
cc_277 N_A_67_199#_c_220_n N_A_434_49#_c_750_n 0.0134988f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_278 N_A_67_199#_c_211_n N_A_434_49#_c_737_n 0.0235577f $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_279 N_A_67_199#_c_218_n N_A_434_49#_c_737_n 0.0256325f $X=2.725 $Y=1.96 $X2=0
+ $Y2=0
cc_280 N_A_67_199#_c_220_n N_A_434_49#_c_737_n 0.00616255f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_281 N_A_67_199#_c_220_n N_A_726_47#_M1014_d 0.00280973f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_282 N_A_67_199#_c_220_n N_A_726_47#_c_916_n 0.0142723f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_283 N_A_67_199#_c_223_n N_A_726_47#_c_916_n 0.00217224f $X=4.295 $Y=1.87
+ $X2=0 $Y2=0
cc_284 N_A_67_199#_c_255_p N_A_726_47#_c_916_n 0.00858155f $X=4.295 $Y=1.87
+ $X2=0 $Y2=0
cc_285 N_A_67_199#_M1019_d N_A_726_47#_c_917_n 0.00350822f $X=4.16 $Y=1.61 $X2=0
+ $Y2=0
cc_286 N_A_67_199#_c_220_n N_A_726_47#_c_917_n 0.00567245f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_287 N_A_67_199#_c_223_n N_A_726_47#_c_917_n 0.00373424f $X=4.295 $Y=1.87
+ $X2=0 $Y2=0
cc_288 N_A_67_199#_c_255_p N_A_726_47#_c_917_n 0.00926398f $X=4.295 $Y=1.87
+ $X2=0 $Y2=0
cc_289 N_A_67_199#_c_255_p N_A_726_47#_c_932_n 9.91724e-19 $X=4.295 $Y=1.87
+ $X2=0 $Y2=0
cc_290 N_A_67_199#_c_223_n N_A_726_47#_c_933_n 0.00251694f $X=4.295 $Y=1.87
+ $X2=0 $Y2=0
cc_291 N_A_67_199#_c_255_p N_A_726_47#_c_933_n 0.00487705f $X=4.295 $Y=1.87
+ $X2=0 $Y2=0
cc_292 N_A_67_199#_c_211_n N_A_28_47#_M1002_d 0.00723162f $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_293 N_A_67_199#_c_218_n N_A_28_47#_M1028_s 0.00588535f $X=2.725 $Y=1.96 $X2=0
+ $Y2=0
cc_294 N_A_67_199#_c_220_n N_A_28_47#_M1028_s 0.00344091f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_295 N_A_67_199#_c_220_n N_A_28_47#_M1014_s 0.00278187f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_67_199#_M1018_g N_A_28_47#_c_1431_n 0.00625347f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_297 N_A_67_199#_c_227_p N_A_28_47#_c_1425_n 0.00527756f $X=1.16 $Y=0.72 $X2=0
+ $Y2=0
cc_298 N_A_67_199#_c_213_n N_A_28_47#_c_1425_n 0.00700681f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_299 N_A_67_199#_M1017_d N_A_28_47#_c_1446_n 0.00164288f $X=1.05 $Y=1.485
+ $X2=0 $Y2=0
cc_300 N_A_67_199#_M1018_g N_A_28_47#_c_1446_n 0.0101197f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_301 N_A_67_199#_c_209_n N_A_28_47#_c_1446_n 0.00414367f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_302 N_A_67_199#_c_231_p N_A_28_47#_c_1446_n 0.0156825f $X=1.28 $Y=1.585 $X2=0
+ $Y2=0
cc_303 N_A_67_199#_c_319_p N_A_28_47#_c_1446_n 0.0137412f $X=0.78 $Y=1.585 $X2=0
+ $Y2=0
cc_304 N_A_67_199#_c_217_n N_A_28_47#_c_1446_n 0.0100843f $X=1.45 $Y=1.96 $X2=0
+ $Y2=0
cc_305 N_A_67_199#_c_212_n N_A_28_47#_c_1446_n 3.28412e-19 $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_306 N_A_67_199#_c_221_n N_A_28_47#_c_1446_n 0.00524508f $X=1.51 $Y=1.87 $X2=0
+ $Y2=0
cc_307 N_A_67_199#_c_222_n N_A_28_47#_c_1446_n 0.00241061f $X=1.365 $Y=1.87
+ $X2=0 $Y2=0
cc_308 N_A_67_199#_M1017_d N_A_28_47#_c_1455_n 0.00680972f $X=1.05 $Y=1.485
+ $X2=0 $Y2=0
cc_309 N_A_67_199#_M1018_g N_A_28_47#_c_1455_n 5.25648e-19 $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_310 N_A_67_199#_c_217_n N_A_28_47#_c_1455_n 0.00281104f $X=1.45 $Y=1.96 $X2=0
+ $Y2=0
cc_311 N_A_67_199#_M1010_d N_A_28_47#_c_1432_n 0.00255556f $X=2.59 $Y=1.485
+ $X2=0 $Y2=0
cc_312 N_A_67_199#_c_218_n N_A_28_47#_c_1432_n 0.0136635f $X=2.725 $Y=1.96 $X2=0
+ $Y2=0
cc_313 N_A_67_199#_c_220_n N_A_28_47#_c_1432_n 0.0101207f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_314 N_A_67_199#_c_220_n N_A_28_47#_c_1433_n 0.00242718f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_315 N_A_67_199#_c_218_n N_A_28_47#_c_1426_n 0.00733634f $X=2.725 $Y=1.96
+ $X2=0 $Y2=0
cc_316 N_A_67_199#_c_220_n N_A_28_47#_c_1426_n 0.0154617f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_317 N_A_67_199#_c_211_n N_A_28_47#_c_1464_n 0.0111988f $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_318 N_A_67_199#_c_211_n N_A_28_47#_c_1465_n 0.0133617f $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_319 N_A_67_199#_c_209_n N_A_28_47#_c_1427_n 0.00556977f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_320 N_A_67_199#_c_212_n N_A_28_47#_c_1427_n 0.00146618f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_321 N_A_67_199#_c_213_n N_A_28_47#_c_1427_n 0.00216178f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_322 N_A_67_199#_M1018_g N_A_28_47#_c_1435_n 0.00819617f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_323 N_A_67_199#_c_209_n N_A_28_47#_c_1435_n 0.0010813f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_324 N_A_67_199#_c_319_p N_A_28_47#_c_1435_n 0.0141105f $X=0.78 $Y=1.585 $X2=0
+ $Y2=0
cc_325 N_A_67_199#_c_212_n N_A_28_47#_c_1435_n 0.00150157f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_326 N_A_67_199#_M1018_g N_A_28_47#_c_1428_n 0.00270966f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_327 N_A_67_199#_c_209_n N_A_28_47#_c_1428_n 0.0315979f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_328 N_A_67_199#_c_216_n N_A_28_47#_c_1428_n 0.00561378f $X=0.695 $Y=1.5 $X2=0
+ $Y2=0
cc_329 N_A_67_199#_c_212_n N_A_28_47#_c_1428_n 0.00822704f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A_67_199#_c_213_n N_A_28_47#_c_1428_n 0.00268818f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A_67_199#_M1017_d N_A_28_47#_c_1437_n 0.00591258f $X=1.05 $Y=1.485
+ $X2=0 $Y2=0
cc_332 N_A_67_199#_c_231_p N_A_28_47#_c_1437_n 0.00363279f $X=1.28 $Y=1.585
+ $X2=0 $Y2=0
cc_333 N_A_67_199#_c_217_n N_A_28_47#_c_1437_n 0.0123158f $X=1.45 $Y=1.96 $X2=0
+ $Y2=0
cc_334 N_A_67_199#_c_218_n N_A_28_47#_c_1437_n 0.058811f $X=2.725 $Y=1.96 $X2=0
+ $Y2=0
cc_335 N_A_67_199#_c_220_n N_A_28_47#_c_1437_n 0.00358352f $X=4.15 $Y=1.87 $X2=0
+ $Y2=0
cc_336 N_A_67_199#_c_221_n N_A_28_47#_c_1437_n 0.00209461f $X=1.51 $Y=1.87 $X2=0
+ $Y2=0
cc_337 N_A_67_199#_M1015_s N_A_28_47#_c_1429_n 0.00295741f $X=3.2 $Y=0.235 $X2=0
+ $Y2=0
cc_338 N_A_67_199#_c_211_n N_A_28_47#_c_1429_n 0.044404f $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_339 N_A_67_199#_c_216_n N_VPWR_M1018_d 3.11669e-19 $X=0.695 $Y=1.5 $X2=-0.19
+ $Y2=-0.24
cc_340 N_A_67_199#_c_231_p N_VPWR_M1018_d 0.0018145f $X=1.28 $Y=1.585 $X2=-0.19
+ $Y2=-0.24
cc_341 N_A_67_199#_c_319_p N_VPWR_M1018_d 0.00417692f $X=0.78 $Y=1.585 $X2=-0.19
+ $Y2=-0.24
cc_342 N_A_67_199#_M1018_g N_VPWR_c_1578_n 0.00280412f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_67_199#_M1018_g N_VPWR_c_1583_n 0.0042268f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_67_199#_M1017_d N_VPWR_c_1577_n 0.00190284f $X=1.05 $Y=1.485 $X2=0
+ $Y2=0
cc_345 N_A_67_199#_M1018_g N_VPWR_c_1577_n 0.00684251f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_A_67_199#_c_220_n N_VPWR_c_1577_n 0.126171f $X=4.15 $Y=1.87 $X2=0 $Y2=0
cc_347 N_A_67_199#_c_221_n N_VPWR_c_1577_n 0.0163456f $X=1.51 $Y=1.87 $X2=0
+ $Y2=0
cc_348 N_A_67_199#_c_223_n N_VPWR_c_1577_n 0.0151773f $X=4.295 $Y=1.87 $X2=0
+ $Y2=0
cc_349 N_A_67_199#_c_209_n N_VGND_M1012_d 0.00396202f $X=0.695 $Y=1.325
+ $X2=-0.19 $Y2=-0.24
cc_350 N_A_67_199#_c_210_n N_VGND_M1012_d 5.44633e-19 $X=0.995 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_351 N_A_67_199#_c_209_n N_VGND_c_2015_n 0.0117147f $X=0.695 $Y=1.325 $X2=0
+ $Y2=0
cc_352 N_A_67_199#_c_210_n N_VGND_c_2015_n 0.00132365f $X=0.995 $Y=0.82 $X2=0
+ $Y2=0
cc_353 N_A_67_199#_c_226_p N_VGND_c_2015_n 0.0148348f $X=1.16 $Y=0.465 $X2=0
+ $Y2=0
cc_354 N_A_67_199#_c_227_p N_VGND_c_2015_n 0.00527979f $X=1.16 $Y=0.72 $X2=0
+ $Y2=0
cc_355 N_A_67_199#_c_213_n N_VGND_c_2015_n 0.00383303f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_67_199#_c_210_n N_VGND_c_2019_n 0.00224601f $X=0.995 $Y=0.82 $X2=0
+ $Y2=0
cc_357 N_A_67_199#_c_226_p N_VGND_c_2019_n 0.0210601f $X=1.16 $Y=0.465 $X2=0
+ $Y2=0
cc_358 N_A_67_199#_c_211_n N_VGND_c_2019_n 0.127391f $X=3.24 $Y=0.36 $X2=0 $Y2=0
cc_359 N_A_67_199#_M1023_d N_VGND_c_2023_n 0.00438671f $X=1.025 $Y=0.235 $X2=0
+ $Y2=0
cc_360 N_A_67_199#_M1015_s N_VGND_c_2023_n 0.00206736f $X=3.2 $Y=0.235 $X2=0
+ $Y2=0
cc_361 N_A_67_199#_c_209_n N_VGND_c_2023_n 0.00127085f $X=0.695 $Y=1.325 $X2=0
+ $Y2=0
cc_362 N_A_67_199#_c_210_n N_VGND_c_2023_n 0.00458421f $X=0.995 $Y=0.82 $X2=0
+ $Y2=0
cc_363 N_A_67_199#_c_226_p N_VGND_c_2023_n 0.0124843f $X=1.16 $Y=0.465 $X2=0
+ $Y2=0
cc_364 N_A_67_199#_c_211_n N_VGND_c_2023_n 0.0379351f $X=3.24 $Y=0.36 $X2=0
+ $Y2=0
cc_365 N_A_67_199#_c_213_n N_VGND_c_2023_n 0.0106925f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A_67_199#_c_209_n N_VGND_c_2024_n 3.07438e-19 $X=0.695 $Y=1.325 $X2=0
+ $Y2=0
cc_367 N_A_67_199#_c_213_n N_VGND_c_2024_n 0.00541359f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_368 A N_B_c_432_n 6.60282e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_369 N_A_c_386_n N_B_c_432_n 0.0214042f $X=1.175 $Y=1.16 $X2=0 $Y2=0
cc_370 N_A_c_384_n B 0.00222756f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_371 A B 0.0161706f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_372 N_A_c_386_n B 0.00341979f $X=1.175 $Y=1.16 $X2=0 $Y2=0
cc_373 N_A_c_384_n N_B_c_441_n 0.00127453f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A_M1017_g N_A_28_47#_c_1431_n 5.78297e-19 $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_375 N_A_c_384_n N_A_28_47#_c_1425_n 5.98586e-19 $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A_M1017_g N_A_28_47#_c_1446_n 0.0104009f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_377 N_A_M1017_g N_A_28_47#_c_1455_n 0.0075453f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_378 N_A_M1017_g N_A_28_47#_c_1490_n 0.00814033f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A_M1017_g N_A_28_47#_c_1435_n 0.00103455f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A_M1017_g N_VPWR_c_1578_n 0.0059862f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A_M1017_g N_VPWR_c_1579_n 0.00390371f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_382 N_A_M1017_g N_VPWR_c_1577_n 0.00710619f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_383 N_A_c_384_n N_VGND_c_2015_n 0.00384648f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A_c_384_n N_VGND_c_2019_n 0.00422898f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_385 N_A_c_384_n N_VGND_c_2023_n 0.0072906f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_386 N_B_c_428_n N_A_488_21#_c_607_n 0.0268178f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_387 N_B_c_440_n N_A_488_21#_c_607_n 0.00472557f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_388 N_B_M1028_g N_A_488_21#_M1010_g 0.0268178f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_389 N_B_c_435_n N_A_488_21#_c_608_n 0.0137515f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_390 N_B_M1019_g N_A_488_21#_M1014_g 0.028599f $X=4.085 $Y=2.03 $X2=0 $Y2=0
cc_391 N_B_c_433_n N_A_488_21#_c_609_n 0.0268178f $X=2.095 $Y=1.16 $X2=0 $Y2=0
cc_392 N_B_c_440_n N_A_488_21#_c_610_n 0.00609439f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_393 N_B_c_434_n N_A_488_21#_c_611_n 0.0129174f $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_394 N_B_c_429_n N_A_488_21#_c_612_n 0.00477107f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_395 N_B_c_435_n N_A_488_21#_c_612_n 0.00378031f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_396 N_B_c_442_n N_A_488_21#_c_612_n 0.00674342f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_397 N_B_c_443_n N_A_488_21#_c_612_n 0.025901f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_398 N_B_c_436_n N_A_488_21#_c_650_n 0.0114462f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_399 N_B_c_437_n N_A_488_21#_c_650_n 0.0121397f $X=5.145 $Y=1.16 $X2=0 $Y2=0
cc_400 N_B_M1019_g N_A_488_21#_c_618_n 0.00686235f $X=4.085 $Y=2.03 $X2=0 $Y2=0
cc_401 N_B_c_434_n N_A_488_21#_c_618_n 0.00321777f $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_402 N_B_c_443_n N_A_488_21#_c_618_n 0.00546712f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_403 N_B_M1019_g N_A_488_21#_c_620_n 0.0074008f $X=4.085 $Y=2.03 $X2=0 $Y2=0
cc_404 N_B_M1000_g N_A_488_21#_c_620_n 0.0121212f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_405 N_B_c_436_n N_A_488_21#_c_620_n 0.00636812f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_406 N_B_c_440_n N_A_488_21#_c_621_n 0.00272545f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_407 N_B_M1019_g N_A_488_21#_c_622_n 0.00129959f $X=4.085 $Y=2.03 $X2=0 $Y2=0
cc_408 N_B_M1000_g N_A_488_21#_c_622_n 0.00258145f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_409 N_B_M1001_g N_A_488_21#_c_622_n 0.00153733f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_410 N_B_c_436_n N_A_488_21#_c_622_n 0.00860517f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_411 N_B_c_437_n N_A_488_21#_c_622_n 0.00524923f $X=5.145 $Y=1.16 $X2=0 $Y2=0
cc_412 N_B_c_430_n N_A_434_49#_c_728_n 0.0192977f $X=5.57 $Y=1.16 $X2=0 $Y2=0
cc_413 N_B_c_434_n N_A_434_49#_c_728_n 0.00300711f $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_414 N_B_c_436_n N_A_434_49#_c_728_n 0.0130034f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_415 N_B_c_437_n N_A_434_49#_c_728_n 0.00330725f $X=5.145 $Y=1.16 $X2=0 $Y2=0
cc_416 N_B_c_438_n N_A_434_49#_c_728_n 0.0116991f $X=5.645 $Y=1.16 $X2=0 $Y2=0
cc_417 N_B_c_440_n N_A_434_49#_c_728_n 0.158533f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_418 N_B_c_442_n N_A_434_49#_c_728_n 0.0253176f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_419 N_B_c_443_n N_A_434_49#_c_728_n 0.0128229f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_420 N_B_c_432_n N_A_434_49#_c_750_n 0.00241151f $X=2.02 $Y=1.16 $X2=0 $Y2=0
cc_421 B N_A_434_49#_c_750_n 0.00651693f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_422 N_B_c_440_n N_A_434_49#_c_750_n 0.0253204f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_423 N_B_c_431_n N_A_434_49#_c_731_n 0.00149902f $X=5.645 $Y=0.995 $X2=0 $Y2=0
cc_424 N_B_c_438_n N_A_434_49#_c_733_n 0.0069216f $X=5.645 $Y=1.16 $X2=0 $Y2=0
cc_425 N_B_c_428_n N_A_434_49#_c_737_n 0.0138347f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_426 N_B_M1028_g N_A_434_49#_c_737_n 0.014908f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_427 N_B_c_432_n N_A_434_49#_c_737_n 0.00723239f $X=2.02 $Y=1.16 $X2=0 $Y2=0
cc_428 N_B_c_433_n N_A_434_49#_c_737_n 0.00848015f $X=2.095 $Y=1.16 $X2=0 $Y2=0
cc_429 B N_A_434_49#_c_737_n 0.0356367f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_430 N_B_c_440_n N_A_434_49#_c_737_n 0.0270152f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_431 N_B_c_441_n N_A_434_49#_c_737_n 6.92027e-19 $X=1.755 $Y=0.85 $X2=0 $Y2=0
cc_432 N_B_c_440_n N_A_726_47#_M1015_d 0.00187267f $X=4.25 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_433 N_B_c_434_n N_A_726_47#_c_916_n 0.0165126f $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_434 N_B_c_443_n N_A_726_47#_c_916_n 2.05789e-19 $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_435 N_B_M1019_g N_A_726_47#_c_917_n 0.0123794f $X=4.085 $Y=2.03 $X2=0 $Y2=0
cc_436 N_B_M1000_g N_A_726_47#_c_917_n 0.00637456f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_437 N_B_c_434_n N_A_726_47#_c_908_n 0.00599801f $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_438 N_B_c_435_n N_A_726_47#_c_908_n 0.00115759f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_439 N_B_c_440_n N_A_726_47#_c_908_n 0.0108825f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_440 N_B_c_442_n N_A_726_47#_c_908_n 0.00226876f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_441 N_B_c_443_n N_A_726_47#_c_908_n 0.0280077f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_442 N_B_M1000_g N_A_726_47#_c_932_n 0.00815313f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_443 N_B_M1001_g N_A_726_47#_c_932_n 5.55638e-19 $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_444 N_B_M1000_g N_A_726_47#_c_947_n 0.00916731f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_445 N_B_c_430_n N_A_726_47#_c_947_n 0.00451048f $X=5.57 $Y=1.16 $X2=0 $Y2=0
cc_446 N_B_M1001_g N_A_726_47#_c_947_n 0.0156501f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_447 N_B_M1000_g N_A_726_47#_c_933_n 0.00428892f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_448 N_B_c_436_n N_A_726_47#_c_933_n 3.24364e-19 $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_449 N_B_M1001_g N_A_726_47#_c_952_n 0.00743023f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_450 N_B_M1001_g N_A_726_47#_c_953_n 0.00383087f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_451 N_B_c_434_n N_A_726_47#_c_910_n 0.00614786f $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_452 N_B_c_440_n N_A_726_47#_c_910_n 0.00133263f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_453 N_B_c_443_n N_A_726_47#_c_910_n 0.011552f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_454 N_B_c_440_n N_A_28_47#_M1002_d 3.94762e-19 $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_455 N_B_c_442_n N_A_28_47#_M1031_d 0.00174146f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_456 N_B_c_443_n N_A_28_47#_M1031_d 0.00452825f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_457 N_B_c_434_n N_A_28_47#_c_1426_n 2.97394e-19 $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_458 N_B_c_435_n N_A_28_47#_c_1464_n 0.00259971f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_459 N_B_M1028_g N_A_28_47#_c_1437_n 0.0116015f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_460 N_B_M1028_g N_A_28_47#_c_1438_n 0.00184265f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_461 N_B_c_440_n N_A_28_47#_c_1429_n 0.0462428f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_462 N_B_c_429_n N_A_28_47#_c_1430_n 0.00376413f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_463 N_B_c_435_n N_A_28_47#_c_1430_n 0.0019893f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_464 N_B_c_436_n N_A_28_47#_c_1430_n 0.0026102f $X=5.06 $Y=1.16 $X2=0 $Y2=0
cc_465 N_B_c_442_n N_A_28_47#_c_1430_n 0.00164354f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_466 N_B_c_443_n N_A_28_47#_c_1430_n 0.0137147f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_467 N_B_c_434_n N_A_28_47#_c_1505_n 2.48926e-19 $X=4.295 $Y=1.16 $X2=0 $Y2=0
cc_468 N_B_c_435_n N_A_28_47#_c_1505_n 0.00813469f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_469 N_B_c_440_n N_A_28_47#_c_1505_n 0.0082305f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_470 N_B_c_442_n N_A_28_47#_c_1505_n 3.07703e-19 $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_471 N_B_M1028_g N_VPWR_c_1579_n 0.00394444f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_472 N_B_M1019_g N_VPWR_c_1579_n 0.00335164f $X=4.085 $Y=2.03 $X2=0 $Y2=0
cc_473 N_B_M1000_g N_VPWR_c_1579_n 0.00409261f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_474 N_B_M1000_g N_VPWR_c_1580_n 0.00537106f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_475 N_B_M1001_g N_VPWR_c_1580_n 0.00902456f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_476 N_B_M1001_g N_VPWR_c_1584_n 0.00341689f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_477 N_B_M1028_g N_VPWR_c_1577_n 0.00381947f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_478 N_B_M1019_g N_VPWR_c_1577_n 0.00687674f $X=4.085 $Y=2.03 $X2=0 $Y2=0
cc_479 N_B_M1000_g N_VPWR_c_1577_n 0.00725684f $X=5.135 $Y=1.985 $X2=0 $Y2=0
cc_480 N_B_M1001_g N_VPWR_c_1577_n 0.00540327f $X=5.645 $Y=1.985 $X2=0 $Y2=0
cc_481 N_B_c_431_n N_A_1144_49#_c_1710_n 0.00325851f $X=5.645 $Y=0.995 $X2=0
+ $Y2=0
cc_482 N_B_M1000_g N_A_1144_49#_c_1706_n 5.46372e-19 $X=5.135 $Y=1.985 $X2=0
+ $Y2=0
cc_483 N_B_c_431_n N_A_1144_49#_c_1706_n 0.0142331f $X=5.645 $Y=0.995 $X2=0
+ $Y2=0
cc_484 N_B_M1001_g N_A_1144_49#_c_1706_n 0.00573601f $X=5.645 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_B_M1001_g N_A_1144_49#_c_1714_n 0.00281901f $X=5.645 $Y=1.985 $X2=0
+ $Y2=0
cc_486 N_B_c_431_n N_A_1144_49#_c_1715_n 0.00264124f $X=5.645 $Y=0.995 $X2=0
+ $Y2=0
cc_487 N_B_M1001_g N_A_1144_49#_c_1716_n 8.4745e-19 $X=5.645 $Y=1.985 $X2=0
+ $Y2=0
cc_488 N_B_c_431_n N_A_1261_49#_c_1808_n 0.00354077f $X=5.645 $Y=0.995 $X2=0
+ $Y2=0
cc_489 N_B_c_429_n N_VGND_c_2016_n 0.0158626f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_490 N_B_c_430_n N_VGND_c_2016_n 0.00695882f $X=5.57 $Y=1.16 $X2=0 $Y2=0
cc_491 N_B_c_431_n N_VGND_c_2016_n 0.00588266f $X=5.645 $Y=0.995 $X2=0 $Y2=0
cc_492 N_B_c_428_n N_VGND_c_2019_n 0.00357877f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_493 N_B_c_429_n N_VGND_c_2019_n 0.0046653f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_494 N_B_c_435_n N_VGND_c_2019_n 0.00351226f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_495 N_B_c_431_n N_VGND_c_2020_n 0.00549826f $X=5.645 $Y=0.995 $X2=0 $Y2=0
cc_496 N_B_c_428_n N_VGND_c_2023_n 0.00661646f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_497 N_B_c_429_n N_VGND_c_2023_n 0.00934473f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_498 N_B_c_431_n N_VGND_c_2023_n 0.0113103f $X=5.645 $Y=0.995 $X2=0 $Y2=0
cc_499 N_B_c_435_n N_VGND_c_2023_n 0.00686244f $X=4.152 $Y=0.995 $X2=0 $Y2=0
cc_500 N_B_c_440_n N_VGND_c_2023_n 0.11709f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_501 N_B_c_441_n N_VGND_c_2023_n 0.0148637f $X=1.755 $Y=0.85 $X2=0 $Y2=0
cc_502 N_B_c_442_n N_VGND_c_2023_n 0.0148223f $X=4.395 $Y=0.85 $X2=0 $Y2=0
cc_503 N_A_488_21#_c_609_n N_A_434_49#_c_728_n 0.00276606f $X=2.515 $Y=1.16
+ $X2=0 $Y2=0
cc_504 N_A_488_21#_c_610_n N_A_434_49#_c_728_n 0.00359514f $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_505 N_A_488_21#_c_611_n N_A_434_49#_c_728_n 0.00466411f $X=3.582 $Y=1.16
+ $X2=0 $Y2=0
cc_506 N_A_488_21#_c_650_n N_A_434_49#_c_728_n 0.0201244f $X=5.01 $Y=1.165 $X2=0
+ $Y2=0
cc_507 N_A_488_21#_c_618_n N_A_434_49#_c_728_n 0.122617f $X=4.71 $Y=1.53 $X2=0
+ $Y2=0
cc_508 N_A_488_21#_c_619_n N_A_434_49#_c_728_n 0.0276606f $X=3.16 $Y=1.53 $X2=0
+ $Y2=0
cc_509 N_A_488_21#_c_670_p N_A_434_49#_c_728_n 0.0254409f $X=4.855 $Y=1.53 $X2=0
+ $Y2=0
cc_510 N_A_488_21#_c_620_n N_A_434_49#_c_728_n 0.00419315f $X=4.855 $Y=1.53
+ $X2=0 $Y2=0
cc_511 N_A_488_21#_c_621_n N_A_434_49#_c_728_n 0.020679f $X=2.81 $Y=1.16 $X2=0
+ $Y2=0
cc_512 N_A_488_21#_c_622_n N_A_434_49#_c_728_n 0.0181199f $X=4.94 $Y=1.385 $X2=0
+ $Y2=0
cc_513 N_A_488_21#_c_621_n N_A_434_49#_c_750_n 3.81879e-19 $X=2.81 $Y=1.16 $X2=0
+ $Y2=0
cc_514 N_A_488_21#_c_607_n N_A_434_49#_c_737_n 0.00829859f $X=2.515 $Y=0.995
+ $X2=0 $Y2=0
cc_515 N_A_488_21#_M1010_g N_A_434_49#_c_737_n 0.00873699f $X=2.515 $Y=1.905
+ $X2=0 $Y2=0
cc_516 N_A_488_21#_c_609_n N_A_434_49#_c_737_n 0.0113589f $X=2.515 $Y=1.16 $X2=0
+ $Y2=0
cc_517 N_A_488_21#_c_619_n N_A_434_49#_c_737_n 0.00215433f $X=3.16 $Y=1.53 $X2=0
+ $Y2=0
cc_518 N_A_488_21#_c_621_n N_A_434_49#_c_737_n 0.0353631f $X=2.81 $Y=1.16 $X2=0
+ $Y2=0
cc_519 N_A_488_21#_c_618_n N_A_726_47#_M1014_d 8.0571e-19 $X=4.71 $Y=1.53 $X2=0
+ $Y2=0
cc_520 N_A_488_21#_M1014_g N_A_726_47#_c_916_n 0.0039967f $X=3.6 $Y=1.905 $X2=0
+ $Y2=0
cc_521 N_A_488_21#_c_618_n N_A_726_47#_c_916_n 0.0133874f $X=4.71 $Y=1.53 $X2=0
+ $Y2=0
cc_522 N_A_488_21#_M1000_s N_A_726_47#_c_917_n 0.00410738f $X=4.8 $Y=1.485 $X2=0
+ $Y2=0
cc_523 N_A_488_21#_c_620_n N_A_726_47#_c_917_n 0.00578738f $X=4.855 $Y=1.53
+ $X2=0 $Y2=0
cc_524 N_A_488_21#_M1014_g N_A_726_47#_c_918_n 0.00133802f $X=3.6 $Y=1.905 $X2=0
+ $Y2=0
cc_525 N_A_488_21#_c_608_n N_A_726_47#_c_908_n 0.00202271f $X=3.555 $Y=0.995
+ $X2=0 $Y2=0
cc_526 N_A_488_21#_c_611_n N_A_726_47#_c_908_n 0.00140297f $X=3.582 $Y=1.16
+ $X2=0 $Y2=0
cc_527 N_A_488_21#_M1000_s N_A_726_47#_c_932_n 0.00843142f $X=4.8 $Y=1.485 $X2=0
+ $Y2=0
cc_528 N_A_488_21#_c_620_n N_A_726_47#_c_947_n 0.0059838f $X=4.855 $Y=1.53 $X2=0
+ $Y2=0
cc_529 N_A_488_21#_M1000_s N_A_726_47#_c_933_n 0.00432451f $X=4.8 $Y=1.485 $X2=0
+ $Y2=0
cc_530 N_A_488_21#_c_670_p N_A_726_47#_c_933_n 8.54896e-19 $X=4.855 $Y=1.53
+ $X2=0 $Y2=0
cc_531 N_A_488_21#_c_620_n N_A_726_47#_c_933_n 0.0138423f $X=4.855 $Y=1.53 $X2=0
+ $Y2=0
cc_532 N_A_488_21#_c_611_n N_A_726_47#_c_910_n 0.00177791f $X=3.582 $Y=1.16
+ $X2=0 $Y2=0
cc_533 N_A_488_21#_c_618_n N_A_726_47#_c_910_n 0.00523631f $X=4.71 $Y=1.53 $X2=0
+ $Y2=0
cc_534 N_A_488_21#_c_618_n N_A_28_47#_M1014_s 0.00150278f $X=4.71 $Y=1.53 $X2=0
+ $Y2=0
cc_535 N_A_488_21#_M1010_g N_A_28_47#_c_1432_n 0.005828f $X=2.515 $Y=1.905 $X2=0
+ $Y2=0
cc_536 N_A_488_21#_M1014_g N_A_28_47#_c_1433_n 0.00593769f $X=3.6 $Y=1.905 $X2=0
+ $Y2=0
cc_537 N_A_488_21#_c_607_n N_A_28_47#_c_1426_n 0.00159539f $X=2.515 $Y=0.995
+ $X2=0 $Y2=0
cc_538 N_A_488_21#_M1010_g N_A_28_47#_c_1426_n 0.00817981f $X=2.515 $Y=1.905
+ $X2=0 $Y2=0
cc_539 N_A_488_21#_c_608_n N_A_28_47#_c_1426_n 5.11963e-19 $X=3.555 $Y=0.995
+ $X2=0 $Y2=0
cc_540 N_A_488_21#_M1014_g N_A_28_47#_c_1426_n 0.0141056f $X=3.6 $Y=1.905 $X2=0
+ $Y2=0
cc_541 N_A_488_21#_c_610_n N_A_28_47#_c_1426_n 0.0226016f $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_542 N_A_488_21#_c_618_n N_A_28_47#_c_1426_n 0.0112473f $X=4.71 $Y=1.53 $X2=0
+ $Y2=0
cc_543 N_A_488_21#_c_619_n N_A_28_47#_c_1426_n 0.0034311f $X=3.16 $Y=1.53 $X2=0
+ $Y2=0
cc_544 N_A_488_21#_c_621_n N_A_28_47#_c_1426_n 0.0361586f $X=2.81 $Y=1.16 $X2=0
+ $Y2=0
cc_545 N_A_488_21#_c_608_n N_A_28_47#_c_1464_n 0.0106545f $X=3.555 $Y=0.995
+ $X2=0 $Y2=0
cc_546 N_A_488_21#_c_608_n N_A_28_47#_c_1465_n 0.00557927f $X=3.555 $Y=0.995
+ $X2=0 $Y2=0
cc_547 N_A_488_21#_M1010_g N_A_28_47#_c_1438_n 0.0109534f $X=2.515 $Y=1.905
+ $X2=0 $Y2=0
cc_548 N_A_488_21#_c_607_n N_A_28_47#_c_1429_n 0.00495001f $X=2.515 $Y=0.995
+ $X2=0 $Y2=0
cc_549 N_A_488_21#_c_608_n N_A_28_47#_c_1429_n 0.0152145f $X=3.555 $Y=0.995
+ $X2=0 $Y2=0
cc_550 N_A_488_21#_c_610_n N_A_28_47#_c_1429_n 0.0175468f $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_551 N_A_488_21#_c_611_n N_A_28_47#_c_1429_n 0.00289939f $X=3.582 $Y=1.16
+ $X2=0 $Y2=0
cc_552 N_A_488_21#_c_621_n N_A_28_47#_c_1429_n 0.0288026f $X=2.81 $Y=1.16 $X2=0
+ $Y2=0
cc_553 N_A_488_21#_M1010_g N_VPWR_c_1579_n 9.63786e-19 $X=2.515 $Y=1.905 $X2=0
+ $Y2=0
cc_554 N_A_488_21#_M1014_g N_VPWR_c_1579_n 0.00513163f $X=3.6 $Y=1.905 $X2=0
+ $Y2=0
cc_555 N_A_488_21#_M1000_s N_VPWR_c_1577_n 0.00210129f $X=4.8 $Y=1.485 $X2=0
+ $Y2=0
cc_556 N_A_488_21#_M1014_g N_VPWR_c_1577_n 0.00343753f $X=3.6 $Y=1.905 $X2=0
+ $Y2=0
cc_557 N_A_488_21#_c_650_n N_A_1144_49#_c_1706_n 0.0120043f $X=5.01 $Y=1.165
+ $X2=0 $Y2=0
cc_558 N_A_488_21#_c_620_n N_A_1144_49#_c_1706_n 0.00614439f $X=4.855 $Y=1.53
+ $X2=0 $Y2=0
cc_559 N_A_488_21#_c_607_n N_VGND_c_2019_n 0.00357877f $X=2.515 $Y=0.995 $X2=0
+ $Y2=0
cc_560 N_A_488_21#_c_608_n N_VGND_c_2019_n 0.00413718f $X=3.555 $Y=0.995 $X2=0
+ $Y2=0
cc_561 N_A_488_21#_c_612_n N_VGND_c_2019_n 0.00481203f $X=4.945 $Y=0.73 $X2=0
+ $Y2=0
cc_562 N_A_488_21#_M1027_s N_VGND_c_2023_n 0.00475007f $X=4.82 $Y=0.605 $X2=0
+ $Y2=0
cc_563 N_A_488_21#_c_607_n N_VGND_c_2023_n 0.00661646f $X=2.515 $Y=0.995 $X2=0
+ $Y2=0
cc_564 N_A_488_21#_c_608_n N_VGND_c_2023_n 0.00745794f $X=3.555 $Y=0.995 $X2=0
+ $Y2=0
cc_565 N_A_488_21#_c_612_n N_VGND_c_2023_n 0.00619044f $X=4.945 $Y=0.73 $X2=0
+ $Y2=0
cc_566 N_A_434_49#_M1025_g N_A_726_47#_M1004_g 0.0371801f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_567 N_A_434_49#_c_727_n N_A_726_47#_c_903_n 0.0260017f $X=6.64 $Y=0.995 $X2=0
+ $Y2=0
cc_568 N_A_434_49#_c_736_n N_A_726_47#_c_904_n 0.021801f $X=8.96 $Y=0.995 $X2=0
+ $Y2=0
cc_569 N_A_434_49#_c_729_n N_A_726_47#_c_905_n 0.0101614f $X=8.85 $Y=1.19 $X2=0
+ $Y2=0
cc_570 N_A_434_49#_c_733_n N_A_726_47#_c_905_n 0.0214585f $X=6.64 $Y=1.16 $X2=0
+ $Y2=0
cc_571 N_A_434_49#_c_729_n N_A_726_47#_c_906_n 0.0153043f $X=8.85 $Y=1.19 $X2=0
+ $Y2=0
cc_572 N_A_434_49#_M1022_g N_A_726_47#_c_907_n 0.0263406f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_573 N_A_434_49#_c_729_n N_A_726_47#_c_907_n 0.0127568f $X=8.85 $Y=1.19 $X2=0
+ $Y2=0
cc_574 N_A_434_49#_c_734_n N_A_726_47#_c_907_n 0.0163799f $X=8.945 $Y=1.16 $X2=0
+ $Y2=0
cc_575 N_A_434_49#_c_735_n N_A_726_47#_c_907_n 7.30793e-19 $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_576 N_A_434_49#_c_728_n N_A_726_47#_c_916_n 2.63373e-19 $X=6.09 $Y=1.19 $X2=0
+ $Y2=0
cc_577 N_A_434_49#_c_728_n N_A_726_47#_c_908_n 0.00412821f $X=6.09 $Y=1.19 $X2=0
+ $Y2=0
cc_578 N_A_434_49#_M1025_g N_A_726_47#_c_952_n 0.00350227f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_579 N_A_434_49#_M1025_g N_A_726_47#_c_919_n 0.0119433f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_580 N_A_434_49#_c_729_n N_A_726_47#_c_909_n 0.0166904f $X=8.85 $Y=1.19 $X2=0
+ $Y2=0
cc_581 N_A_434_49#_c_728_n N_A_726_47#_c_910_n 0.0135249f $X=6.09 $Y=1.19 $X2=0
+ $Y2=0
cc_582 N_A_434_49#_c_729_n N_A_726_47#_c_923_n 0.00362829f $X=8.85 $Y=1.19 $X2=0
+ $Y2=0
cc_583 N_A_434_49#_c_734_n N_A_1589_49#_c_1108_n 0.00187737f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_584 N_A_434_49#_c_735_n N_A_1589_49#_c_1108_n 0.00202234f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_585 N_A_434_49#_c_736_n N_A_1589_49#_c_1108_n 0.0124748f $X=8.96 $Y=0.995
+ $X2=0 $Y2=0
cc_586 N_A_434_49#_M1022_g N_A_1589_49#_c_1094_n 0.0039232f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_587 N_A_434_49#_c_732_n N_A_1589_49#_c_1094_n 0.00768453f $X=8.995 $Y=1.19
+ $X2=0 $Y2=0
cc_588 N_A_434_49#_c_734_n N_A_1589_49#_c_1094_n 0.00317608f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_589 N_A_434_49#_c_735_n N_A_1589_49#_c_1094_n 0.0185336f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_590 N_A_434_49#_c_736_n N_A_1589_49#_c_1094_n 0.0122115f $X=8.96 $Y=0.995
+ $X2=0 $Y2=0
cc_591 N_A_434_49#_c_729_n N_A_1589_49#_c_1098_n 0.0012513f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_592 N_A_434_49#_M1022_g N_A_1589_49#_c_1107_n 0.0114385f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_593 N_A_434_49#_c_732_n N_A_1589_49#_c_1107_n 2.98178e-19 $X=8.995 $Y=1.19
+ $X2=0 $Y2=0
cc_594 N_A_434_49#_c_734_n N_A_1589_49#_c_1107_n 8.86285e-19 $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_595 N_A_434_49#_c_735_n N_A_1589_49#_c_1107_n 0.00182047f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_596 N_A_434_49#_M1022_g N_A_1710_49#_c_1307_n 0.00100967f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_597 N_A_434_49#_c_729_n N_A_1710_49#_c_1307_n 0.0114746f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_598 N_A_434_49#_c_732_n N_A_1710_49#_c_1307_n 0.00125349f $X=8.995 $Y=1.19
+ $X2=0 $Y2=0
cc_599 N_A_434_49#_c_734_n N_A_1710_49#_c_1307_n 0.0012474f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_600 N_A_434_49#_c_735_n N_A_1710_49#_c_1307_n 0.020673f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_601 N_A_434_49#_c_736_n N_A_1710_49#_c_1307_n 0.00157684f $X=8.96 $Y=0.995
+ $X2=0 $Y2=0
cc_602 N_A_434_49#_M1022_g N_A_1710_49#_c_1313_n 0.00225168f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_603 N_A_434_49#_c_729_n N_A_1710_49#_c_1313_n 0.00276081f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_604 N_A_434_49#_c_734_n N_A_1710_49#_c_1313_n 0.00144337f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_605 N_A_434_49#_c_735_n N_A_1710_49#_c_1313_n 0.00524068f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_606 N_A_434_49#_M1022_g N_A_1710_49#_c_1329_n 0.0059407f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_607 N_A_434_49#_c_735_n N_A_1710_49#_c_1330_n 0.00352613f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_608 N_A_434_49#_c_736_n N_A_1710_49#_c_1330_n 0.00478173f $X=8.96 $Y=0.995
+ $X2=0 $Y2=0
cc_609 N_A_434_49#_M1022_g N_A_1710_49#_c_1314_n 0.00845332f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_610 N_A_434_49#_c_729_n N_A_1710_49#_c_1314_n 0.0134523f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_611 N_A_434_49#_c_732_n N_A_1710_49#_c_1314_n 0.0274167f $X=8.995 $Y=1.19
+ $X2=0 $Y2=0
cc_612 N_A_434_49#_c_734_n N_A_1710_49#_c_1314_n 0.00240935f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_613 N_A_434_49#_c_735_n N_A_1710_49#_c_1314_n 0.00348359f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_614 N_A_434_49#_M1022_g N_A_1710_49#_c_1315_n 4.4878e-19 $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_615 N_A_434_49#_c_729_n N_A_1710_49#_c_1315_n 0.0260853f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_616 N_A_434_49#_c_728_n N_A_28_47#_c_1426_n 0.0115149f $X=6.09 $Y=1.19 $X2=0
+ $Y2=0
cc_617 N_A_434_49#_M1028_d N_A_28_47#_c_1437_n 0.00146558f $X=2.17 $Y=1.485
+ $X2=0 $Y2=0
cc_618 N_A_434_49#_c_728_n N_A_28_47#_c_1429_n 0.0130352f $X=6.09 $Y=1.19 $X2=0
+ $Y2=0
cc_619 N_A_434_49#_c_737_n N_A_28_47#_c_1429_n 0.0122149f $X=2.305 $Y=0.72 $X2=0
+ $Y2=0
cc_620 N_A_434_49#_M1025_g N_VPWR_c_1584_n 9.44495e-19 $X=6.585 $Y=1.905 $X2=0
+ $Y2=0
cc_621 N_A_434_49#_M1022_g N_VPWR_c_1584_n 0.00313972f $X=8.945 $Y=1.995 $X2=0
+ $Y2=0
cc_622 N_A_434_49#_M1022_g N_VPWR_c_1577_n 0.00519382f $X=8.945 $Y=1.995 $X2=0
+ $Y2=0
cc_623 N_A_434_49#_c_727_n N_A_1144_49#_c_1710_n 0.00310651f $X=6.64 $Y=0.995
+ $X2=0 $Y2=0
cc_624 N_A_434_49#_M1025_g N_A_1144_49#_c_1706_n 0.00356489f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_625 N_A_434_49#_c_728_n N_A_1144_49#_c_1706_n 0.0307657f $X=6.09 $Y=1.19
+ $X2=0 $Y2=0
cc_626 N_A_434_49#_c_730_n N_A_1144_49#_c_1706_n 0.00275249f $X=6.38 $Y=1.19
+ $X2=0 $Y2=0
cc_627 N_A_434_49#_c_733_n N_A_1144_49#_c_1706_n 9.64063e-19 $X=6.64 $Y=1.16
+ $X2=0 $Y2=0
cc_628 N_A_434_49#_M1025_g N_A_1144_49#_c_1724_n 0.00382305f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_629 N_A_434_49#_c_728_n N_A_1144_49#_c_1724_n 0.00437461f $X=6.09 $Y=1.19
+ $X2=0 $Y2=0
cc_630 N_A_434_49#_c_730_n N_A_1144_49#_c_1724_n 0.00433012f $X=6.38 $Y=1.19
+ $X2=0 $Y2=0
cc_631 N_A_434_49#_c_731_n N_A_1144_49#_c_1724_n 0.013108f $X=6.235 $Y=1.19
+ $X2=0 $Y2=0
cc_632 N_A_434_49#_c_733_n N_A_1144_49#_c_1724_n 0.00363059f $X=6.64 $Y=1.16
+ $X2=0 $Y2=0
cc_633 N_A_434_49#_M1025_g N_A_1144_49#_c_1714_n 0.00215498f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_634 N_A_434_49#_M1025_g N_A_1144_49#_c_1730_n 0.00931505f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_635 N_A_434_49#_c_729_n N_A_1144_49#_c_1707_n 0.0201739f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_636 N_A_434_49#_M1025_g N_A_1144_49#_c_1709_n 6.70022e-19 $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_637 N_A_434_49#_c_729_n N_A_1144_49#_c_1709_n 0.0101391f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_638 N_A_434_49#_c_728_n N_A_1144_49#_c_1715_n 0.00464233f $X=6.09 $Y=1.19
+ $X2=0 $Y2=0
cc_639 N_A_434_49#_c_731_n N_A_1144_49#_c_1715_n 0.0441479f $X=6.235 $Y=1.19
+ $X2=0 $Y2=0
cc_640 N_A_434_49#_M1025_g N_A_1144_49#_c_1716_n 0.00321587f $X=6.585 $Y=1.905
+ $X2=0 $Y2=0
cc_641 N_A_434_49#_c_731_n N_A_1144_49#_c_1716_n 0.00169815f $X=6.235 $Y=1.19
+ $X2=0 $Y2=0
cc_642 N_A_434_49#_c_733_n N_A_1144_49#_c_1716_n 0.00214523f $X=6.64 $Y=1.16
+ $X2=0 $Y2=0
cc_643 N_A_434_49#_M1025_g COUT_N 0.00635668f $X=6.585 $Y=1.905 $X2=0 $Y2=0
cc_644 N_A_434_49#_c_727_n COUT_N 0.00161643f $X=6.64 $Y=0.995 $X2=0 $Y2=0
cc_645 N_A_434_49#_c_729_n COUT_N 0.0330527f $X=8.85 $Y=1.19 $X2=0 $Y2=0
cc_646 N_A_434_49#_c_730_n COUT_N 5.6439e-19 $X=6.38 $Y=1.19 $X2=0 $Y2=0
cc_647 N_A_434_49#_c_731_n COUT_N 0.0271315f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_648 N_A_434_49#_c_733_n COUT_N 0.0101219f $X=6.64 $Y=1.16 $X2=0 $Y2=0
cc_649 N_A_434_49#_M1025_g COUT_N 0.00293392f $X=6.585 $Y=1.905 $X2=0 $Y2=0
cc_650 N_A_434_49#_c_727_n N_COUT_N_c_1780_n 0.00522673f $X=6.64 $Y=0.995 $X2=0
+ $Y2=0
cc_651 N_A_434_49#_c_729_n N_COUT_N_c_1780_n 0.002594f $X=8.85 $Y=1.19 $X2=0
+ $Y2=0
cc_652 N_A_434_49#_c_731_n N_COUT_N_c_1780_n 0.0129305f $X=6.235 $Y=1.19 $X2=0
+ $Y2=0
cc_653 N_A_434_49#_c_731_n N_A_1261_49#_M1013_s 0.00314604f $X=6.235 $Y=1.19
+ $X2=-0.19 $Y2=-0.24
cc_654 N_A_434_49#_c_727_n N_A_1261_49#_c_1807_n 0.00808644f $X=6.64 $Y=0.995
+ $X2=0 $Y2=0
cc_655 N_A_434_49#_c_727_n N_A_1261_49#_c_1808_n 0.00530807f $X=6.64 $Y=0.995
+ $X2=0 $Y2=0
cc_656 N_A_434_49#_c_729_n N_A_1261_49#_c_1808_n 0.00490782f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_657 N_A_434_49#_c_730_n N_A_1261_49#_c_1808_n 4.57094e-19 $X=6.38 $Y=1.19
+ $X2=0 $Y2=0
cc_658 N_A_434_49#_c_731_n N_A_1261_49#_c_1808_n 0.0133397f $X=6.235 $Y=1.19
+ $X2=0 $Y2=0
cc_659 N_A_434_49#_c_733_n N_A_1261_49#_c_1808_n 0.00400012f $X=6.64 $Y=1.16
+ $X2=0 $Y2=0
cc_660 N_A_434_49#_c_729_n N_A_1261_49#_c_1815_n 0.0253117f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_661 N_A_434_49#_c_729_n N_A_1261_49#_c_1809_n 0.0874609f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_662 N_A_434_49#_c_732_n N_A_1261_49#_c_1809_n 0.0263368f $X=8.995 $Y=1.19
+ $X2=0 $Y2=0
cc_663 N_A_434_49#_c_734_n N_A_1261_49#_c_1809_n 0.00250551f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_664 N_A_434_49#_c_735_n N_A_1261_49#_c_1809_n 0.00354077f $X=8.945 $Y=1.16
+ $X2=0 $Y2=0
cc_665 N_A_434_49#_c_736_n N_A_1261_49#_c_1809_n 0.00574413f $X=8.96 $Y=0.995
+ $X2=0 $Y2=0
cc_666 N_A_434_49#_c_729_n N_A_1261_49#_c_1810_n 0.0258329f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_667 N_A_434_49#_c_729_n N_A_1634_315#_c_1942_n 0.00544491f $X=8.85 $Y=1.19
+ $X2=0 $Y2=0
cc_668 N_A_434_49#_M1022_g N_A_1634_315#_c_1939_n 0.0170018f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_669 N_A_434_49#_c_736_n N_A_1634_315#_c_1944_n 0.00114584f $X=8.96 $Y=0.995
+ $X2=0 $Y2=0
cc_670 N_A_434_49#_M1022_g N_A_1634_315#_c_1938_n 0.00288021f $X=8.945 $Y=1.995
+ $X2=0 $Y2=0
cc_671 N_A_434_49#_c_728_n N_VGND_c_2016_n 0.0136256f $X=6.09 $Y=1.19 $X2=0
+ $Y2=0
cc_672 N_A_434_49#_c_727_n N_VGND_c_2020_n 0.00352679f $X=6.64 $Y=0.995 $X2=0
+ $Y2=0
cc_673 N_A_434_49#_c_731_n N_VGND_c_2020_n 0.00189339f $X=6.235 $Y=1.19 $X2=0
+ $Y2=0
cc_674 N_A_434_49#_c_736_n N_VGND_c_2020_n 0.00357877f $X=8.96 $Y=0.995 $X2=0
+ $Y2=0
cc_675 N_A_434_49#_c_727_n N_VGND_c_2023_n 0.00646238f $X=6.64 $Y=0.995 $X2=0
+ $Y2=0
cc_676 N_A_434_49#_c_731_n N_VGND_c_2023_n 0.00355378f $X=6.235 $Y=1.19 $X2=0
+ $Y2=0
cc_677 N_A_434_49#_c_736_n N_VGND_c_2023_n 0.00676309f $X=8.96 $Y=0.995 $X2=0
+ $Y2=0
cc_678 N_A_726_47#_c_904_n N_A_1589_49#_c_1108_n 0.0116053f $X=8.475 $Y=0.995
+ $X2=0 $Y2=0
cc_679 N_A_726_47#_c_907_n N_A_1589_49#_c_1108_n 0.00103372f $X=8.475 $Y=1.247
+ $X2=0 $Y2=0
cc_680 N_A_726_47#_c_904_n N_A_1589_49#_c_1098_n 0.011097f $X=8.475 $Y=0.995
+ $X2=0 $Y2=0
cc_681 N_A_726_47#_c_906_n N_A_1589_49#_c_1098_n 7.35476e-19 $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_682 N_A_726_47#_c_907_n N_A_1589_49#_c_1098_n 0.00859402f $X=8.475 $Y=1.247
+ $X2=0 $Y2=0
cc_683 N_A_726_47#_c_909_n N_A_1589_49#_c_1098_n 0.00742174f $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_684 N_A_726_47#_c_904_n N_A_1710_49#_c_1307_n 0.00750834f $X=8.475 $Y=0.995
+ $X2=0 $Y2=0
cc_685 N_A_726_47#_c_907_n N_A_1710_49#_c_1307_n 0.0168582f $X=8.475 $Y=1.247
+ $X2=0 $Y2=0
cc_686 N_A_726_47#_c_909_n N_A_1710_49#_c_1307_n 0.0134898f $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_687 N_A_726_47#_c_912_n N_A_1710_49#_c_1313_n 0.00675957f $X=8.525 $Y=1.5
+ $X2=0 $Y2=0
cc_688 N_A_726_47#_c_907_n N_A_1710_49#_c_1313_n 0.0022202f $X=8.475 $Y=1.247
+ $X2=0 $Y2=0
cc_689 N_A_726_47#_c_909_n N_A_1710_49#_c_1313_n 0.00416498f $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_690 N_A_726_47#_c_912_n N_A_1710_49#_c_1329_n 0.00740019f $X=8.525 $Y=1.5
+ $X2=0 $Y2=0
cc_691 N_A_726_47#_c_920_n N_A_1710_49#_c_1329_n 0.00183499f $X=7.875 $Y=2.295
+ $X2=0 $Y2=0
cc_692 N_A_726_47#_c_923_n N_A_1710_49#_c_1329_n 0.0029706f $X=7.917 $Y=1.72
+ $X2=0 $Y2=0
cc_693 N_A_726_47#_c_904_n N_A_1710_49#_c_1348_n 0.00431321f $X=8.475 $Y=0.995
+ $X2=0 $Y2=0
cc_694 N_A_726_47#_c_912_n N_A_1710_49#_c_1315_n 0.0054666f $X=8.525 $Y=1.5
+ $X2=0 $Y2=0
cc_695 N_A_726_47#_c_907_n N_A_1710_49#_c_1315_n 0.00190534f $X=8.475 $Y=1.247
+ $X2=0 $Y2=0
cc_696 N_A_726_47#_c_909_n N_A_1710_49#_c_1315_n 0.00623789f $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_697 N_A_726_47#_c_918_n N_A_28_47#_c_1433_n 0.0128907f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_698 N_A_726_47#_c_916_n N_A_28_47#_c_1426_n 0.0285419f $X=3.81 $Y=1.7 $X2=0
+ $Y2=0
cc_699 N_A_726_47#_c_908_n N_A_28_47#_c_1426_n 0.00539181f $X=4.01 $Y=0.76 $X2=0
+ $Y2=0
cc_700 N_A_726_47#_c_910_n N_A_28_47#_c_1426_n 0.00742461f $X=4.01 $Y=1.235
+ $X2=0 $Y2=0
cc_701 N_A_726_47#_M1015_d N_A_28_47#_c_1464_n 0.00381449f $X=3.63 $Y=0.235
+ $X2=0 $Y2=0
cc_702 N_A_726_47#_c_908_n N_A_28_47#_c_1464_n 0.0112862f $X=4.01 $Y=0.76 $X2=0
+ $Y2=0
cc_703 N_A_726_47#_M1015_d N_A_28_47#_c_1465_n 6.15829e-19 $X=3.63 $Y=0.235
+ $X2=0 $Y2=0
cc_704 N_A_726_47#_M1015_d N_A_28_47#_c_1429_n 6.97451e-19 $X=3.63 $Y=0.235
+ $X2=0 $Y2=0
cc_705 N_A_726_47#_c_908_n N_A_28_47#_c_1429_n 0.0119356f $X=4.01 $Y=0.76 $X2=0
+ $Y2=0
cc_706 N_A_726_47#_c_910_n N_A_28_47#_c_1429_n 0.00136905f $X=4.01 $Y=1.235
+ $X2=0 $Y2=0
cc_707 N_A_726_47#_M1015_d N_A_28_47#_c_1505_n 0.00895089f $X=3.63 $Y=0.235
+ $X2=0 $Y2=0
cc_708 N_A_726_47#_c_908_n N_A_28_47#_c_1505_n 0.0114751f $X=4.01 $Y=0.76 $X2=0
+ $Y2=0
cc_709 N_A_726_47#_c_947_n N_VPWR_M1000_d 0.00794628f $X=5.835 $Y=1.98 $X2=0
+ $Y2=0
cc_710 N_A_726_47#_c_917_n N_VPWR_c_1579_n 0.0761665f $X=4.875 $Y=2.38 $X2=0
+ $Y2=0
cc_711 N_A_726_47#_c_918_n N_VPWR_c_1579_n 0.0121882f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_712 N_A_726_47#_c_947_n N_VPWR_c_1579_n 0.00228295f $X=5.835 $Y=1.98 $X2=0
+ $Y2=0
cc_713 N_A_726_47#_c_917_n N_VPWR_c_1580_n 0.0140085f $X=4.875 $Y=2.38 $X2=0
+ $Y2=0
cc_714 N_A_726_47#_c_932_n N_VPWR_c_1580_n 0.0044937f $X=4.987 $Y=2.295 $X2=0
+ $Y2=0
cc_715 N_A_726_47#_c_947_n N_VPWR_c_1580_n 0.0206205f $X=5.835 $Y=1.98 $X2=0
+ $Y2=0
cc_716 N_A_726_47#_c_952_n N_VPWR_c_1580_n 0.003425f $X=5.92 $Y=2.295 $X2=0
+ $Y2=0
cc_717 N_A_726_47#_c_953_n N_VPWR_c_1580_n 0.0109407f $X=6.005 $Y=2.38 $X2=0
+ $Y2=0
cc_718 N_A_726_47#_M1004_g N_VPWR_c_1584_n 9.44495e-19 $X=7.005 $Y=1.905 $X2=0
+ $Y2=0
cc_719 N_A_726_47#_c_912_n N_VPWR_c_1584_n 0.00313972f $X=8.525 $Y=1.5 $X2=0
+ $Y2=0
cc_720 N_A_726_47#_c_947_n N_VPWR_c_1584_n 0.00335963f $X=5.835 $Y=1.98 $X2=0
+ $Y2=0
cc_721 N_A_726_47#_c_919_n N_VPWR_c_1584_n 0.126769f $X=7.79 $Y=2.38 $X2=0 $Y2=0
cc_722 N_A_726_47#_c_953_n N_VPWR_c_1584_n 0.0118015f $X=6.005 $Y=2.38 $X2=0
+ $Y2=0
cc_723 N_A_726_47#_c_912_n N_VPWR_c_1577_n 0.00519382f $X=8.525 $Y=1.5 $X2=0
+ $Y2=0
cc_724 N_A_726_47#_c_917_n N_VPWR_c_1577_n 0.0333818f $X=4.875 $Y=2.38 $X2=0
+ $Y2=0
cc_725 N_A_726_47#_c_918_n N_VPWR_c_1577_n 0.00311866f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_726 N_A_726_47#_c_947_n N_VPWR_c_1577_n 0.0116076f $X=5.835 $Y=1.98 $X2=0
+ $Y2=0
cc_727 N_A_726_47#_c_919_n N_VPWR_c_1577_n 0.0730221f $X=7.79 $Y=2.38 $X2=0
+ $Y2=0
cc_728 N_A_726_47#_c_953_n N_VPWR_c_1577_n 0.00651702f $X=6.005 $Y=2.38 $X2=0
+ $Y2=0
cc_729 N_A_726_47#_c_947_n N_A_1144_49#_M1001_d 0.00626813f $X=5.835 $Y=1.98
+ $X2=0 $Y2=0
cc_730 N_A_726_47#_c_952_n N_A_1144_49#_M1001_d 0.00716186f $X=5.92 $Y=2.295
+ $X2=0 $Y2=0
cc_731 N_A_726_47#_c_919_n N_A_1144_49#_M1001_d 0.0128212f $X=7.79 $Y=2.38 $X2=0
+ $Y2=0
cc_732 N_A_726_47#_c_953_n N_A_1144_49#_M1001_d 0.00490995f $X=6.005 $Y=2.38
+ $X2=0 $Y2=0
cc_733 N_A_726_47#_c_947_n N_A_1144_49#_c_1706_n 0.0223447f $X=5.835 $Y=1.98
+ $X2=0 $Y2=0
cc_734 N_A_726_47#_c_947_n N_A_1144_49#_c_1724_n 0.0019685f $X=5.835 $Y=1.98
+ $X2=0 $Y2=0
cc_735 N_A_726_47#_c_919_n N_A_1144_49#_c_1724_n 0.00601442f $X=7.79 $Y=2.38
+ $X2=0 $Y2=0
cc_736 N_A_726_47#_M1004_g N_A_1144_49#_c_1730_n 0.01446f $X=7.005 $Y=1.905
+ $X2=0 $Y2=0
cc_737 N_A_726_47#_c_919_n N_A_1144_49#_c_1730_n 0.0083871f $X=7.79 $Y=2.38
+ $X2=0 $Y2=0
cc_738 N_A_726_47#_c_903_n N_A_1144_49#_c_1707_n 0.00664727f $X=7.065 $Y=0.995
+ $X2=0 $Y2=0
cc_739 N_A_726_47#_c_905_n N_A_1144_49#_c_1707_n 0.00505614f $X=7.035 $Y=1.16
+ $X2=0 $Y2=0
cc_740 N_A_726_47#_c_906_n N_A_1144_49#_c_1707_n 0.0117706f $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_741 N_A_726_47#_M1004_g N_A_1144_49#_c_1709_n 0.0187858f $X=7.005 $Y=1.905
+ $X2=0 $Y2=0
cc_742 N_A_726_47#_c_905_n N_A_1144_49#_c_1709_n 0.00292034f $X=7.035 $Y=1.16
+ $X2=0 $Y2=0
cc_743 N_A_726_47#_c_906_n N_A_1144_49#_c_1709_n 0.00398638f $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_744 N_A_726_47#_c_947_n N_A_1144_49#_c_1716_n 0.0130086f $X=5.835 $Y=1.98
+ $X2=0 $Y2=0
cc_745 N_A_726_47#_c_952_n N_A_1144_49#_c_1716_n 0.00414373f $X=5.92 $Y=2.295
+ $X2=0 $Y2=0
cc_746 N_A_726_47#_c_919_n N_A_1144_49#_c_1716_n 0.0448489f $X=7.79 $Y=2.38
+ $X2=0 $Y2=0
cc_747 N_A_726_47#_c_919_n N_COUT_N_M1025_d 0.00166235f $X=7.79 $Y=2.38 $X2=0
+ $Y2=0
cc_748 N_A_726_47#_c_903_n COUT_N 5.04756e-19 $X=7.065 $Y=0.995 $X2=0 $Y2=0
cc_749 N_A_726_47#_c_905_n COUT_N 0.00356487f $X=7.035 $Y=1.16 $X2=0 $Y2=0
cc_750 N_A_726_47#_c_903_n N_COUT_N_c_1780_n 2.94306e-19 $X=7.065 $Y=0.995 $X2=0
+ $Y2=0
cc_751 N_A_726_47#_c_905_n N_COUT_N_c_1780_n 2.47785e-19 $X=7.035 $Y=1.16 $X2=0
+ $Y2=0
cc_752 N_A_726_47#_c_919_n N_A_1261_49#_M1004_d 0.0120493f $X=7.79 $Y=2.38 $X2=0
+ $Y2=0
cc_753 N_A_726_47#_c_903_n N_A_1261_49#_c_1807_n 0.0141726f $X=7.065 $Y=0.995
+ $X2=0 $Y2=0
cc_754 N_A_726_47#_c_904_n N_A_1261_49#_c_1807_n 5.53798e-19 $X=8.475 $Y=0.995
+ $X2=0 $Y2=0
cc_755 N_A_726_47#_c_905_n N_A_1261_49#_c_1807_n 8.79554e-19 $X=7.035 $Y=1.16
+ $X2=0 $Y2=0
cc_756 N_A_726_47#_c_906_n N_A_1261_49#_c_1807_n 0.00443758f $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_757 N_A_726_47#_M1004_g N_A_1261_49#_c_1837_n 0.00301685f $X=7.005 $Y=1.905
+ $X2=0 $Y2=0
cc_758 N_A_726_47#_c_919_n N_A_1261_49#_c_1837_n 0.0128008f $X=7.79 $Y=2.38
+ $X2=0 $Y2=0
cc_759 N_A_726_47#_c_909_n N_A_1261_49#_c_1837_n 9.05164e-19 $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_760 N_A_726_47#_c_923_n N_A_1261_49#_c_1837_n 0.034532f $X=7.917 $Y=1.72
+ $X2=0 $Y2=0
cc_761 N_A_726_47#_c_903_n N_A_1261_49#_c_1808_n 7.8676e-19 $X=7.065 $Y=0.995
+ $X2=0 $Y2=0
cc_762 N_A_726_47#_M1004_g N_A_1261_49#_c_1815_n 0.00105176f $X=7.005 $Y=1.905
+ $X2=0 $Y2=0
cc_763 N_A_726_47#_c_906_n N_A_1261_49#_c_1815_n 0.0217605f $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_764 N_A_726_47#_c_907_n N_A_1261_49#_c_1815_n 8.81477e-19 $X=8.475 $Y=1.247
+ $X2=0 $Y2=0
cc_765 N_A_726_47#_c_909_n N_A_1261_49#_c_1815_n 0.0255141f $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_766 N_A_726_47#_c_904_n N_A_1261_49#_c_1809_n 0.0031077f $X=8.475 $Y=0.995
+ $X2=0 $Y2=0
cc_767 N_A_726_47#_c_906_n N_A_1261_49#_c_1809_n 0.00673126f $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_768 N_A_726_47#_c_909_n N_A_1261_49#_c_1809_n 0.00285468f $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_769 N_A_726_47#_c_904_n N_A_1261_49#_c_1810_n 8.14764e-19 $X=8.475 $Y=0.995
+ $X2=0 $Y2=0
cc_770 N_A_726_47#_c_906_n N_A_1261_49#_c_1810_n 0.0020237f $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_771 N_A_726_47#_c_903_n N_A_1261_49#_c_1811_n 0.0050088f $X=7.065 $Y=0.995
+ $X2=0 $Y2=0
cc_772 N_A_726_47#_c_906_n N_A_1261_49#_c_1811_n 0.00920242f $X=8.005 $Y=1.16
+ $X2=0 $Y2=0
cc_773 N_A_726_47#_c_909_n N_A_1261_49#_c_1811_n 0.00725132f $X=7.96 $Y=1.16
+ $X2=0 $Y2=0
cc_774 N_A_726_47#_c_907_n N_A_1634_315#_c_1942_n 0.00681059f $X=8.475 $Y=1.247
+ $X2=0 $Y2=0
cc_775 N_A_726_47#_c_920_n N_A_1634_315#_c_1942_n 0.0270432f $X=7.875 $Y=2.295
+ $X2=0 $Y2=0
cc_776 N_A_726_47#_c_912_n N_A_1634_315#_c_1939_n 0.0118974f $X=8.525 $Y=1.5
+ $X2=0 $Y2=0
cc_777 N_A_726_47#_c_919_n N_A_1634_315#_c_1940_n 0.0112831f $X=7.79 $Y=2.38
+ $X2=0 $Y2=0
cc_778 N_A_726_47#_c_903_n N_VGND_c_2020_n 0.00351226f $X=7.065 $Y=0.995 $X2=0
+ $Y2=0
cc_779 N_A_726_47#_c_904_n N_VGND_c_2020_n 0.00351226f $X=8.475 $Y=0.995 $X2=0
+ $Y2=0
cc_780 N_A_726_47#_M1015_d N_VGND_c_2023_n 0.00240414f $X=3.63 $Y=0.235 $X2=0
+ $Y2=0
cc_781 N_A_726_47#_c_903_n N_VGND_c_2023_n 0.00647149f $X=7.065 $Y=0.995 $X2=0
+ $Y2=0
cc_782 N_A_726_47#_c_904_n N_VGND_c_2023_n 0.00645346f $X=8.475 $Y=0.995 $X2=0
+ $Y2=0
cc_783 N_A_1589_49#_M1030_g N_CI_M1016_g 0.043969f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_784 N_A_1589_49#_c_1097_n N_CI_M1016_g 0.0206783f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_785 N_A_1589_49#_c_1095_n N_CI_c_1242_n 0.00898136f $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_786 N_A_1589_49#_c_1096_n N_CI_c_1242_n 0.00724166f $X=10.73 $Y=0.4 $X2=0
+ $Y2=0
cc_787 N_A_1589_49#_c_1097_n N_CI_c_1242_n 9.635e-19 $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_788 N_A_1589_49#_c_1100_n N_CI_c_1242_n 0.0193004f $X=10.075 $Y=0.995 $X2=0
+ $Y2=0
cc_789 N_A_1589_49#_c_1095_n N_CI_c_1243_n 6.87385e-19 $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_790 N_A_1589_49#_c_1097_n N_CI_M1021_g 0.00117726f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_791 N_A_1589_49#_c_1095_n N_CI_c_1244_n 8.06394e-19 $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_792 N_A_1589_49#_c_1097_n N_CI_c_1244_n 0.00715055f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_793 N_A_1589_49#_c_1099_n N_CI_c_1244_n 0.0215662f $X=10.075 $Y=1.16 $X2=0
+ $Y2=0
cc_794 N_A_1589_49#_c_1095_n N_CI_c_1245_n 0.00578114f $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_795 N_A_1589_49#_c_1097_n N_CI_c_1245_n 0.0044129f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_796 N_A_1589_49#_c_1095_n CI 0.0250787f $X=10.54 $Y=0.82 $X2=0 $Y2=0
cc_797 N_A_1589_49#_c_1097_n CI 0.0368559f $X=10.73 $Y=2.045 $X2=0 $Y2=0
cc_798 N_A_1589_49#_c_1108_n N_A_1710_49#_M1007_d 0.00338156f $X=9.28 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_799 N_A_1589_49#_c_1094_n N_A_1710_49#_c_1307_n 0.0081729f $X=9.365 $Y=1.53
+ $X2=0 $Y2=0
cc_800 N_A_1589_49#_c_1098_n N_A_1710_49#_c_1307_n 0.00410672f $X=8.105 $Y=0.38
+ $X2=0 $Y2=0
cc_801 N_A_1589_49#_c_1094_n N_A_1710_49#_c_1313_n 0.00184268f $X=9.365 $Y=1.53
+ $X2=0 $Y2=0
cc_802 N_A_1589_49#_c_1107_n N_A_1710_49#_c_1313_n 0.00500592f $X=9.235 $Y=1.7
+ $X2=0 $Y2=0
cc_803 N_A_1589_49#_c_1105_n N_A_1710_49#_c_1329_n 0.00121486f $X=9.51 $Y=1.87
+ $X2=0 $Y2=0
cc_804 N_A_1589_49#_c_1108_n N_A_1710_49#_c_1348_n 0.00759547f $X=9.28 $Y=0.34
+ $X2=0 $Y2=0
cc_805 N_A_1589_49#_c_1098_n N_A_1710_49#_c_1348_n 0.0136154f $X=8.105 $Y=0.38
+ $X2=0 $Y2=0
cc_806 N_A_1589_49#_c_1108_n N_A_1710_49#_c_1330_n 0.0146389f $X=9.28 $Y=0.34
+ $X2=0 $Y2=0
cc_807 N_A_1589_49#_c_1094_n N_A_1710_49#_c_1330_n 0.00686482f $X=9.365 $Y=1.53
+ $X2=0 $Y2=0
cc_808 N_A_1589_49#_M1022_d N_A_1710_49#_c_1314_n 0.00186371f $X=9.02 $Y=1.575
+ $X2=0 $Y2=0
cc_809 N_A_1589_49#_M1016_d N_A_1710_49#_c_1314_n 7.60699e-19 $X=10.57 $Y=1.485
+ $X2=0 $Y2=0
cc_810 N_A_1589_49#_M1030_g N_A_1710_49#_c_1314_n 0.00614805f $X=10.075 $Y=1.985
+ $X2=0 $Y2=0
cc_811 N_A_1589_49#_c_1094_n N_A_1710_49#_c_1314_n 0.00844026f $X=9.365 $Y=1.53
+ $X2=0 $Y2=0
cc_812 N_A_1589_49#_c_1095_n N_A_1710_49#_c_1314_n 3.15721e-19 $X=10.54 $Y=0.82
+ $X2=0 $Y2=0
cc_813 N_A_1589_49#_c_1097_n N_A_1710_49#_c_1314_n 0.0570187f $X=10.73 $Y=2.045
+ $X2=0 $Y2=0
cc_814 N_A_1589_49#_c_1104_n N_A_1710_49#_c_1314_n 0.0481824f $X=10.13 $Y=1.87
+ $X2=0 $Y2=0
cc_815 N_A_1589_49#_c_1105_n N_A_1710_49#_c_1314_n 0.0277343f $X=9.51 $Y=1.87
+ $X2=0 $Y2=0
cc_816 N_A_1589_49#_c_1160_p N_A_1710_49#_c_1314_n 0.0253896f $X=10.275 $Y=1.87
+ $X2=0 $Y2=0
cc_817 N_A_1589_49#_c_1099_n N_A_1710_49#_c_1314_n 9.6356e-19 $X=10.075 $Y=1.16
+ $X2=0 $Y2=0
cc_818 N_A_1589_49#_c_1107_n N_A_1710_49#_c_1314_n 0.0181695f $X=9.235 $Y=1.7
+ $X2=0 $Y2=0
cc_819 N_A_1589_49#_c_1094_n N_A_1710_49#_c_1315_n 7.45832e-19 $X=9.365 $Y=1.53
+ $X2=0 $Y2=0
cc_820 N_A_1589_49#_c_1107_n N_A_1710_49#_c_1315_n 2.18508e-19 $X=9.235 $Y=1.7
+ $X2=0 $Y2=0
cc_821 N_A_1589_49#_c_1097_n N_VPWR_M1030_d 0.00285197f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_822 N_A_1589_49#_c_1160_p N_VPWR_M1030_d 5.16085e-19 $X=10.275 $Y=1.87 $X2=0
+ $Y2=0
cc_823 N_A_1589_49#_M1030_g N_VPWR_c_1581_n 0.00826262f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_824 N_A_1589_49#_c_1097_n N_VPWR_c_1581_n 0.0108182f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_825 N_A_1589_49#_c_1104_n N_VPWR_c_1581_n 2.2332e-19 $X=10.13 $Y=1.87 $X2=0
+ $Y2=0
cc_826 N_A_1589_49#_c_1160_p N_VPWR_c_1581_n 0.00287523f $X=10.275 $Y=1.87 $X2=0
+ $Y2=0
cc_827 N_A_1589_49#_M1030_g N_VPWR_c_1584_n 0.0046653f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_828 N_A_1589_49#_c_1097_n N_VPWR_c_1585_n 0.00234007f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_829 N_A_1589_49#_c_1173_p N_VPWR_c_1585_n 0.0145919f $X=10.71 $Y=2.3 $X2=0
+ $Y2=0
cc_830 N_A_1589_49#_M1016_d N_VPWR_c_1577_n 0.00324681f $X=10.57 $Y=1.485 $X2=0
+ $Y2=0
cc_831 N_A_1589_49#_M1030_g N_VPWR_c_1577_n 0.00581646f $X=10.075 $Y=1.985 $X2=0
+ $Y2=0
cc_832 N_A_1589_49#_c_1097_n N_VPWR_c_1577_n 0.00535399f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_833 N_A_1589_49#_c_1173_p N_VPWR_c_1577_n 0.00800522f $X=10.71 $Y=2.3 $X2=0
+ $Y2=0
cc_834 N_A_1589_49#_c_1104_n N_VPWR_c_1577_n 0.0297559f $X=10.13 $Y=1.87 $X2=0
+ $Y2=0
cc_835 N_A_1589_49#_c_1105_n N_VPWR_c_1577_n 0.0162998f $X=9.51 $Y=1.87 $X2=0
+ $Y2=0
cc_836 N_A_1589_49#_c_1160_p N_VPWR_c_1577_n 0.0134077f $X=10.275 $Y=1.87 $X2=0
+ $Y2=0
cc_837 N_A_1589_49#_c_1098_n N_A_1261_49#_c_1807_n 0.0126753f $X=8.105 $Y=0.38
+ $X2=0 $Y2=0
cc_838 N_A_1589_49#_c_1097_n N_A_1261_49#_c_1813_n 0.0362355f $X=10.73 $Y=2.045
+ $X2=0 $Y2=0
cc_839 N_A_1589_49#_c_1173_p N_A_1261_49#_c_1814_n 0.0251865f $X=10.71 $Y=2.3
+ $X2=0 $Y2=0
cc_840 N_A_1589_49#_c_1096_n N_A_1261_49#_c_1857_n 0.0273464f $X=10.73 $Y=0.4
+ $X2=0 $Y2=0
cc_841 N_A_1589_49#_c_1095_n N_A_1261_49#_c_1858_n 0.00872264f $X=10.54 $Y=0.82
+ $X2=0 $Y2=0
cc_842 N_A_1589_49#_M1007_s N_A_1261_49#_c_1809_n 0.00108682f $X=7.945 $Y=0.245
+ $X2=0 $Y2=0
cc_843 N_A_1589_49#_c_1108_n N_A_1261_49#_c_1809_n 0.0115577f $X=9.28 $Y=0.34
+ $X2=0 $Y2=0
cc_844 N_A_1589_49#_c_1094_n N_A_1261_49#_c_1809_n 0.0172142f $X=9.365 $Y=1.53
+ $X2=0 $Y2=0
cc_845 N_A_1589_49#_c_1095_n N_A_1261_49#_c_1809_n 0.0253331f $X=10.54 $Y=0.82
+ $X2=0 $Y2=0
cc_846 N_A_1589_49#_c_1097_n N_A_1261_49#_c_1809_n 0.0209561f $X=10.73 $Y=2.045
+ $X2=0 $Y2=0
cc_847 N_A_1589_49#_c_1098_n N_A_1261_49#_c_1809_n 0.0176953f $X=8.105 $Y=0.38
+ $X2=0 $Y2=0
cc_848 N_A_1589_49#_c_1099_n N_A_1261_49#_c_1809_n 5.57837e-19 $X=10.075 $Y=1.16
+ $X2=0 $Y2=0
cc_849 N_A_1589_49#_c_1100_n N_A_1261_49#_c_1809_n 0.00459474f $X=10.075
+ $Y=0.995 $X2=0 $Y2=0
cc_850 N_A_1589_49#_c_1107_n N_A_1261_49#_c_1809_n 8.1166e-19 $X=9.235 $Y=1.7
+ $X2=0 $Y2=0
cc_851 N_A_1589_49#_c_1098_n N_A_1261_49#_c_1810_n 0.00135069f $X=8.105 $Y=0.38
+ $X2=0 $Y2=0
cc_852 N_A_1589_49#_c_1098_n N_A_1261_49#_c_1811_n 0.0241124f $X=8.105 $Y=0.38
+ $X2=0 $Y2=0
cc_853 N_A_1589_49#_c_1095_n N_A_1261_49#_c_1870_n 3.70194e-19 $X=10.54 $Y=0.82
+ $X2=0 $Y2=0
cc_854 N_A_1589_49#_c_1108_n N_A_1634_315#_M1008_d 0.0118782f $X=9.28 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_855 N_A_1589_49#_c_1094_n N_A_1634_315#_M1008_d 0.0142652f $X=9.365 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_856 N_A_1589_49#_c_1104_n N_A_1634_315#_M1030_s 0.00104271f $X=10.13 $Y=1.87
+ $X2=0 $Y2=0
cc_857 N_A_1589_49#_M1022_d N_A_1634_315#_c_1939_n 0.00429707f $X=9.02 $Y=1.575
+ $X2=0 $Y2=0
cc_858 N_A_1589_49#_c_1104_n N_A_1634_315#_c_1939_n 0.00358285f $X=10.13 $Y=1.87
+ $X2=0 $Y2=0
cc_859 N_A_1589_49#_c_1105_n N_A_1634_315#_c_1939_n 0.00241459f $X=9.51 $Y=1.87
+ $X2=0 $Y2=0
cc_860 N_A_1589_49#_c_1107_n N_A_1634_315#_c_1939_n 0.0264883f $X=9.235 $Y=1.7
+ $X2=0 $Y2=0
cc_861 N_A_1589_49#_c_1108_n N_A_1634_315#_c_1944_n 0.0129306f $X=9.28 $Y=0.34
+ $X2=0 $Y2=0
cc_862 N_A_1589_49#_c_1094_n N_A_1634_315#_c_1944_n 0.0721013f $X=9.365 $Y=1.53
+ $X2=0 $Y2=0
cc_863 N_A_1589_49#_c_1096_n N_A_1634_315#_c_1944_n 0.00518308f $X=10.73 $Y=0.4
+ $X2=0 $Y2=0
cc_864 N_A_1589_49#_c_1100_n N_A_1634_315#_c_1944_n 0.00557231f $X=10.075
+ $Y=0.995 $X2=0 $Y2=0
cc_865 N_A_1589_49#_M1030_g N_A_1634_315#_c_1961_n 0.00577249f $X=10.075
+ $Y=1.985 $X2=0 $Y2=0
cc_866 N_A_1589_49#_c_1097_n N_A_1634_315#_c_1961_n 0.00652238f $X=10.73
+ $Y=2.045 $X2=0 $Y2=0
cc_867 N_A_1589_49#_c_1099_n N_A_1634_315#_c_1961_n 2.65954e-19 $X=10.075
+ $Y=1.16 $X2=0 $Y2=0
cc_868 N_A_1589_49#_c_1104_n N_A_1634_315#_c_1964_n 0.0212408f $X=10.13 $Y=1.87
+ $X2=0 $Y2=0
cc_869 N_A_1589_49#_c_1105_n N_A_1634_315#_c_1964_n 0.00278291f $X=9.51 $Y=1.87
+ $X2=0 $Y2=0
cc_870 N_A_1589_49#_c_1160_p N_A_1634_315#_c_1964_n 0.00233426f $X=10.275
+ $Y=1.87 $X2=0 $Y2=0
cc_871 N_A_1589_49#_c_1107_n N_A_1634_315#_c_1964_n 0.00526993f $X=9.235 $Y=1.7
+ $X2=0 $Y2=0
cc_872 N_A_1589_49#_c_1097_n N_A_1634_315#_c_1968_n 0.00865173f $X=10.73
+ $Y=2.045 $X2=0 $Y2=0
cc_873 N_A_1589_49#_c_1099_n N_A_1634_315#_c_1968_n 8.53648e-19 $X=10.075
+ $Y=1.16 $X2=0 $Y2=0
cc_874 N_A_1589_49#_c_1100_n N_A_1634_315#_c_1968_n 0.00337697f $X=10.075
+ $Y=0.995 $X2=0 $Y2=0
cc_875 N_A_1589_49#_M1030_g N_A_1634_315#_c_1938_n 0.00323567f $X=10.075
+ $Y=1.985 $X2=0 $Y2=0
cc_876 N_A_1589_49#_c_1097_n N_A_1634_315#_c_1938_n 0.0370987f $X=10.73 $Y=2.045
+ $X2=0 $Y2=0
cc_877 N_A_1589_49#_c_1099_n N_A_1634_315#_c_1938_n 0.00752814f $X=10.075
+ $Y=1.16 $X2=0 $Y2=0
cc_878 N_A_1589_49#_c_1100_n N_A_1634_315#_c_1938_n 0.00227138f $X=10.075
+ $Y=0.995 $X2=0 $Y2=0
cc_879 N_A_1589_49#_c_1107_n N_A_1634_315#_c_1938_n 0.0335608f $X=9.235 $Y=1.7
+ $X2=0 $Y2=0
cc_880 N_A_1589_49#_c_1095_n N_VGND_M1020_d 4.32033e-19 $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_881 N_A_1589_49#_c_1097_n N_VGND_M1020_d 0.00375843f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_882 N_A_1589_49#_c_1095_n N_VGND_c_2017_n 6.03982e-19 $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_883 N_A_1589_49#_c_1096_n N_VGND_c_2017_n 0.0209035f $X=10.73 $Y=0.4 $X2=0
+ $Y2=0
cc_884 N_A_1589_49#_c_1097_n N_VGND_c_2017_n 0.0125847f $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_885 N_A_1589_49#_c_1100_n N_VGND_c_2017_n 0.00365114f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_886 N_A_1589_49#_c_1108_n N_VGND_c_2020_n 0.0689497f $X=9.28 $Y=0.34 $X2=0
+ $Y2=0
cc_887 N_A_1589_49#_c_1098_n N_VGND_c_2020_n 0.023271f $X=8.105 $Y=0.38 $X2=0
+ $Y2=0
cc_888 N_A_1589_49#_c_1100_n N_VGND_c_2020_n 0.00501942f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_889 N_A_1589_49#_c_1095_n N_VGND_c_2021_n 0.00191836f $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_890 N_A_1589_49#_c_1096_n N_VGND_c_2021_n 0.0204614f $X=10.73 $Y=0.4 $X2=0
+ $Y2=0
cc_891 N_A_1589_49#_M1003_d N_VGND_c_2023_n 0.0017338f $X=10.595 $Y=0.235 $X2=0
+ $Y2=0
cc_892 N_A_1589_49#_c_1108_n N_VGND_c_2023_n 0.0197304f $X=9.28 $Y=0.34 $X2=0
+ $Y2=0
cc_893 N_A_1589_49#_c_1095_n N_VGND_c_2023_n 0.0017193f $X=10.54 $Y=0.82 $X2=0
+ $Y2=0
cc_894 N_A_1589_49#_c_1096_n N_VGND_c_2023_n 0.00664209f $X=10.73 $Y=0.4 $X2=0
+ $Y2=0
cc_895 N_A_1589_49#_c_1097_n N_VGND_c_2023_n 5.90557e-19 $X=10.73 $Y=2.045 $X2=0
+ $Y2=0
cc_896 N_A_1589_49#_c_1098_n N_VGND_c_2023_n 0.00608687f $X=8.105 $Y=0.38 $X2=0
+ $Y2=0
cc_897 N_A_1589_49#_c_1100_n N_VGND_c_2023_n 0.00730937f $X=10.075 $Y=0.995
+ $X2=0 $Y2=0
cc_898 N_CI_M1021_g N_A_1710_49#_M1011_g 0.0261027f $X=11.46 $Y=1.985 $X2=0
+ $Y2=0
cc_899 N_CI_M1021_g N_A_1710_49#_c_1314_n 0.00976642f $X=11.46 $Y=1.985 $X2=0
+ $Y2=0
cc_900 N_CI_c_1245_n N_A_1710_49#_c_1314_n 0.00446966f $X=11.385 $Y=1.16 $X2=0
+ $Y2=0
cc_901 CI N_A_1710_49#_c_1314_n 0.00508423f $X=10.75 $Y=1.105 $X2=0 $Y2=0
cc_902 N_CI_M1021_g N_A_1710_49#_c_1316_n 0.00144107f $X=11.46 $Y=1.985 $X2=0
+ $Y2=0
cc_903 N_CI_c_1246_n N_A_1710_49#_c_1308_n 0.0216941f $X=11.46 $Y=1.16 $X2=0
+ $Y2=0
cc_904 N_CI_c_1246_n N_A_1710_49#_c_1309_n 0.00446904f $X=11.46 $Y=1.16 $X2=0
+ $Y2=0
cc_905 N_CI_c_1243_n N_A_1710_49#_c_1310_n 0.0196241f $X=11.46 $Y=0.995 $X2=0
+ $Y2=0
cc_906 N_CI_M1016_g N_VPWR_c_1581_n 0.00846058f $X=10.495 $Y=1.985 $X2=0 $Y2=0
cc_907 N_CI_M1021_g N_VPWR_c_1582_n 0.00280208f $X=11.46 $Y=1.985 $X2=0 $Y2=0
cc_908 N_CI_M1016_g N_VPWR_c_1585_n 0.00329498f $X=10.495 $Y=1.985 $X2=0 $Y2=0
cc_909 N_CI_M1021_g N_VPWR_c_1585_n 0.00541359f $X=11.46 $Y=1.985 $X2=0 $Y2=0
cc_910 N_CI_M1016_g N_VPWR_c_1577_n 0.00520039f $X=10.495 $Y=1.985 $X2=0 $Y2=0
cc_911 N_CI_M1021_g N_VPWR_c_1577_n 0.0108548f $X=11.46 $Y=1.985 $X2=0 $Y2=0
cc_912 N_CI_M1016_g N_A_1261_49#_c_1813_n 0.00109032f $X=10.495 $Y=1.985 $X2=0
+ $Y2=0
cc_913 N_CI_M1021_g N_A_1261_49#_c_1813_n 0.00203012f $X=11.46 $Y=1.985 $X2=0
+ $Y2=0
cc_914 N_CI_c_1245_n N_A_1261_49#_c_1813_n 0.00366648f $X=11.385 $Y=1.16 $X2=0
+ $Y2=0
cc_915 N_CI_M1021_g N_A_1261_49#_c_1814_n 0.0101256f $X=11.46 $Y=1.985 $X2=0
+ $Y2=0
cc_916 N_CI_c_1242_n N_A_1261_49#_c_1857_n 9.04978e-19 $X=10.52 $Y=0.995 $X2=0
+ $Y2=0
cc_917 N_CI_c_1243_n N_A_1261_49#_c_1858_n 0.00382698f $X=11.46 $Y=0.995 $X2=0
+ $Y2=0
cc_918 N_CI_c_1242_n N_A_1261_49#_c_1809_n 0.00198631f $X=10.52 $Y=0.995 $X2=0
+ $Y2=0
cc_919 N_CI_c_1244_n N_A_1261_49#_c_1809_n 5.63257e-19 $X=10.507 $Y=1.16 $X2=0
+ $Y2=0
cc_920 N_CI_c_1245_n N_A_1261_49#_c_1809_n 0.00894399f $X=11.385 $Y=1.16 $X2=0
+ $Y2=0
cc_921 CI N_A_1261_49#_c_1809_n 0.00558207f $X=10.75 $Y=1.105 $X2=0 $Y2=0
cc_922 N_CI_c_1243_n N_A_1261_49#_c_1870_n 0.00514817f $X=11.46 $Y=0.995 $X2=0
+ $Y2=0
cc_923 N_CI_M1016_g N_A_1261_49#_c_1812_n 0.00297411f $X=10.495 $Y=1.985 $X2=0
+ $Y2=0
cc_924 N_CI_c_1242_n N_A_1261_49#_c_1812_n 0.00196745f $X=10.52 $Y=0.995 $X2=0
+ $Y2=0
cc_925 N_CI_c_1243_n N_A_1261_49#_c_1812_n 0.00740992f $X=11.46 $Y=0.995 $X2=0
+ $Y2=0
cc_926 N_CI_M1021_g N_A_1261_49#_c_1812_n 0.00393605f $X=11.46 $Y=1.985 $X2=0
+ $Y2=0
cc_927 N_CI_c_1245_n N_A_1261_49#_c_1812_n 0.0220421f $X=11.385 $Y=1.16 $X2=0
+ $Y2=0
cc_928 N_CI_c_1246_n N_A_1261_49#_c_1812_n 0.00395206f $X=11.46 $Y=1.16 $X2=0
+ $Y2=0
cc_929 CI N_A_1261_49#_c_1812_n 0.0136896f $X=10.75 $Y=1.105 $X2=0 $Y2=0
cc_930 N_CI_c_1242_n N_A_1634_315#_c_1944_n 5.47812e-19 $X=10.52 $Y=0.995 $X2=0
+ $Y2=0
cc_931 N_CI_c_1243_n N_SUM_c_1997_n 8.2064e-19 $X=11.46 $Y=0.995 $X2=0 $Y2=0
cc_932 N_CI_c_1242_n N_VGND_c_2017_n 0.00441669f $X=10.52 $Y=0.995 $X2=0 $Y2=0
cc_933 N_CI_c_1243_n N_VGND_c_2018_n 0.00317394f $X=11.46 $Y=0.995 $X2=0 $Y2=0
cc_934 N_CI_c_1242_n N_VGND_c_2021_n 0.00413062f $X=10.52 $Y=0.995 $X2=0 $Y2=0
cc_935 N_CI_c_1243_n N_VGND_c_2021_n 0.00543994f $X=11.46 $Y=0.995 $X2=0 $Y2=0
cc_936 N_CI_c_1242_n N_VGND_c_2023_n 0.00696852f $X=10.52 $Y=0.995 $X2=0 $Y2=0
cc_937 N_CI_c_1243_n N_VGND_c_2023_n 0.00949627f $X=11.46 $Y=0.995 $X2=0 $Y2=0
cc_938 N_A_1710_49#_c_1314_n N_VPWR_M1030_d 3.23615e-19 $X=11.63 $Y=1.53 $X2=0
+ $Y2=0
cc_939 N_A_1710_49#_c_1314_n N_VPWR_M1021_d 0.00228444f $X=11.63 $Y=1.53 $X2=0
+ $Y2=0
cc_940 N_A_1710_49#_c_1316_n N_VPWR_M1021_d 0.00180492f $X=11.775 $Y=1.53 $X2=0
+ $Y2=0
cc_941 N_A_1710_49#_c_1309_n N_VPWR_M1021_d 0.00128737f $X=11.88 $Y=1.16 $X2=0
+ $Y2=0
cc_942 N_A_1710_49#_M1011_g N_VPWR_c_1582_n 0.0135622f $X=11.88 $Y=1.985 $X2=0
+ $Y2=0
cc_943 N_A_1710_49#_c_1314_n N_VPWR_c_1582_n 0.00226154f $X=11.63 $Y=1.53 $X2=0
+ $Y2=0
cc_944 N_A_1710_49#_c_1316_n N_VPWR_c_1582_n 0.00669312f $X=11.775 $Y=1.53 $X2=0
+ $Y2=0
cc_945 N_A_1710_49#_c_1309_n N_VPWR_c_1582_n 0.00992907f $X=11.88 $Y=1.16 $X2=0
+ $Y2=0
cc_946 N_A_1710_49#_M1011_g N_VPWR_c_1586_n 0.00447018f $X=11.88 $Y=1.985 $X2=0
+ $Y2=0
cc_947 N_A_1710_49#_M1011_g N_VPWR_c_1577_n 0.00859957f $X=11.88 $Y=1.985 $X2=0
+ $Y2=0
cc_948 N_A_1710_49#_M1011_g N_A_1261_49#_c_1813_n 7.52739e-19 $X=11.88 $Y=1.985
+ $X2=0 $Y2=0
cc_949 N_A_1710_49#_c_1314_n N_A_1261_49#_c_1813_n 0.0343003f $X=11.63 $Y=1.53
+ $X2=0 $Y2=0
cc_950 N_A_1710_49#_c_1316_n N_A_1261_49#_c_1813_n 0.00177524f $X=11.775 $Y=1.53
+ $X2=0 $Y2=0
cc_951 N_A_1710_49#_c_1310_n N_A_1261_49#_c_1858_n 0.00178776f $X=11.88 $Y=0.995
+ $X2=0 $Y2=0
cc_952 N_A_1710_49#_M1007_d N_A_1261_49#_c_1809_n 0.00149273f $X=8.55 $Y=0.245
+ $X2=0 $Y2=0
cc_953 N_A_1710_49#_c_1307_n N_A_1261_49#_c_1809_n 0.0148048f $X=8.525 $Y=1.445
+ $X2=0 $Y2=0
cc_954 N_A_1710_49#_c_1330_n N_A_1261_49#_c_1809_n 0.00803645f $X=8.705 $Y=0.68
+ $X2=0 $Y2=0
cc_955 N_A_1710_49#_c_1314_n N_A_1261_49#_c_1809_n 0.0895979f $X=11.63 $Y=1.53
+ $X2=0 $Y2=0
cc_956 N_A_1710_49#_c_1314_n N_A_1261_49#_c_1870_n 0.0126255f $X=11.63 $Y=1.53
+ $X2=0 $Y2=0
cc_957 N_A_1710_49#_c_1310_n N_A_1261_49#_c_1870_n 0.00112497f $X=11.88 $Y=0.995
+ $X2=0 $Y2=0
cc_958 N_A_1710_49#_M1011_g N_A_1261_49#_c_1812_n 3.23024e-19 $X=11.88 $Y=1.985
+ $X2=0 $Y2=0
cc_959 N_A_1710_49#_c_1316_n N_A_1261_49#_c_1812_n 0.00125324f $X=11.775 $Y=1.53
+ $X2=0 $Y2=0
cc_960 N_A_1710_49#_c_1308_n N_A_1261_49#_c_1812_n 2.99878e-19 $X=11.88 $Y=1.16
+ $X2=0 $Y2=0
cc_961 N_A_1710_49#_c_1309_n N_A_1261_49#_c_1812_n 0.0342796f $X=11.88 $Y=1.16
+ $X2=0 $Y2=0
cc_962 N_A_1710_49#_c_1315_n N_A_1634_315#_M1024_s 0.0028544f $X=8.68 $Y=1.53
+ $X2=0 $Y2=0
cc_963 N_A_1710_49#_c_1314_n N_A_1634_315#_M1030_s 4.43593e-19 $X=11.63 $Y=1.53
+ $X2=0 $Y2=0
cc_964 N_A_1710_49#_c_1315_n N_A_1634_315#_c_1942_n 5.098e-19 $X=8.68 $Y=1.53
+ $X2=0 $Y2=0
cc_965 N_A_1710_49#_M1024_d N_A_1634_315#_c_1939_n 0.00165831f $X=8.6 $Y=1.575
+ $X2=0 $Y2=0
cc_966 N_A_1710_49#_c_1329_n N_A_1634_315#_c_1939_n 0.0158712f $X=8.735 $Y=1.7
+ $X2=0 $Y2=0
cc_967 N_A_1710_49#_c_1314_n N_A_1634_315#_c_1961_n 0.0110907f $X=11.63 $Y=1.53
+ $X2=0 $Y2=0
cc_968 N_A_1710_49#_c_1314_n N_A_1634_315#_c_1938_n 0.00740659f $X=11.63 $Y=1.53
+ $X2=0 $Y2=0
cc_969 N_A_1710_49#_M1011_g SUM 0.0061778f $X=11.88 $Y=1.985 $X2=0 $Y2=0
cc_970 N_A_1710_49#_c_1316_n SUM 0.00262669f $X=11.775 $Y=1.53 $X2=0 $Y2=0
cc_971 N_A_1710_49#_c_1308_n SUM 0.00756306f $X=11.88 $Y=1.16 $X2=0 $Y2=0
cc_972 N_A_1710_49#_c_1309_n SUM 0.0412654f $X=11.88 $Y=1.16 $X2=0 $Y2=0
cc_973 N_A_1710_49#_c_1310_n SUM 0.00784594f $X=11.88 $Y=0.995 $X2=0 $Y2=0
cc_974 N_A_1710_49#_c_1310_n N_SUM_c_1997_n 0.00484081f $X=11.88 $Y=0.995 $X2=0
+ $Y2=0
cc_975 N_A_1710_49#_c_1308_n N_VGND_c_2018_n 4.46335e-19 $X=11.88 $Y=1.16 $X2=0
+ $Y2=0
cc_976 N_A_1710_49#_c_1309_n N_VGND_c_2018_n 0.00687847f $X=11.88 $Y=1.16 $X2=0
+ $Y2=0
cc_977 N_A_1710_49#_c_1310_n N_VGND_c_2018_n 0.00313438f $X=11.88 $Y=0.995 $X2=0
+ $Y2=0
cc_978 N_A_1710_49#_c_1310_n N_VGND_c_2022_n 0.00564131f $X=11.88 $Y=0.995 $X2=0
+ $Y2=0
cc_979 N_A_1710_49#_c_1310_n N_VGND_c_2023_n 0.0112336f $X=11.88 $Y=0.995 $X2=0
+ $Y2=0
cc_980 N_A_28_47#_c_1446_n N_VPWR_M1018_d 0.00541207f $X=0.94 $Y=1.925 $X2=-0.19
+ $Y2=-0.24
cc_981 N_A_28_47#_c_1446_n N_VPWR_c_1578_n 0.0126308f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_982 N_A_28_47#_c_1455_n N_VPWR_c_1578_n 0.00242328f $X=1.025 $Y=2.215 $X2=0
+ $Y2=0
cc_983 N_A_28_47#_c_1490_n N_VPWR_c_1578_n 0.0133618f $X=1.11 $Y=2.3 $X2=0 $Y2=0
cc_984 N_A_28_47#_c_1446_n N_VPWR_c_1579_n 0.00208831f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_985 N_A_28_47#_c_1490_n N_VPWR_c_1579_n 0.00633644f $X=1.11 $Y=2.3 $X2=0
+ $Y2=0
cc_986 N_A_28_47#_c_1433_n N_VPWR_c_1579_n 0.018373f $X=3.355 $Y=2.295 $X2=0
+ $Y2=0
cc_987 N_A_28_47#_c_1437_n N_VPWR_c_1579_n 0.0534473f $X=2.375 $Y=2.34 $X2=0
+ $Y2=0
cc_988 N_A_28_47#_c_1438_n N_VPWR_c_1579_n 0.05782f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_989 N_A_28_47#_c_1431_n N_VPWR_c_1583_n 0.0221136f $X=0.265 $Y=2.31 $X2=0
+ $Y2=0
cc_990 N_A_28_47#_c_1446_n N_VPWR_c_1583_n 0.00191602f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_991 N_A_28_47#_M1018_s N_VPWR_c_1577_n 0.00209319f $X=0.14 $Y=1.485 $X2=0
+ $Y2=0
cc_992 N_A_28_47#_M1014_s N_VPWR_c_1577_n 0.00202962f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_993 N_A_28_47#_c_1431_n N_VPWR_c_1577_n 0.0130045f $X=0.265 $Y=2.31 $X2=0
+ $Y2=0
cc_994 N_A_28_47#_c_1446_n N_VPWR_c_1577_n 0.00872069f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_995 N_A_28_47#_c_1490_n N_VPWR_c_1577_n 0.00570549f $X=1.11 $Y=2.3 $X2=0
+ $Y2=0
cc_996 N_A_28_47#_c_1433_n N_VPWR_c_1577_n 0.00481919f $X=3.355 $Y=2.295 $X2=0
+ $Y2=0
cc_997 N_A_28_47#_c_1435_n N_VPWR_c_1577_n 2.06696e-19 $X=0.265 $Y=1.63 $X2=0
+ $Y2=0
cc_998 N_A_28_47#_c_1437_n N_VPWR_c_1577_n 0.0215915f $X=2.375 $Y=2.34 $X2=0
+ $Y2=0
cc_999 N_A_28_47#_c_1438_n N_VPWR_c_1577_n 0.0153395f $X=2.545 $Y=2.34 $X2=0
+ $Y2=0
cc_1000 N_A_28_47#_c_1425_n N_VGND_c_2015_n 0.0188898f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_1001 N_A_28_47#_c_1430_n N_VGND_c_2016_n 0.00695297f $X=4.43 $Y=0.39 $X2=0
+ $Y2=0
cc_1002 N_A_28_47#_c_1465_n N_VGND_c_2019_n 0.00985313f $X=3.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1003 N_A_28_47#_c_1429_n N_VGND_c_2019_n 0.00189661f $X=3.355 $Y=0.79 $X2=0
+ $Y2=0
cc_1004 N_A_28_47#_c_1505_n N_VGND_c_2019_n 0.0503423f $X=4.265 $Y=0.365 $X2=0
+ $Y2=0
cc_1005 N_A_28_47#_M1012_s N_VGND_c_2023_n 0.00209319f $X=0.14 $Y=0.235 $X2=0
+ $Y2=0
cc_1006 N_A_28_47#_c_1425_n N_VGND_c_2023_n 0.0123905f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_1007 N_A_28_47#_c_1465_n N_VGND_c_2023_n 0.00300815f $X=3.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1008 N_A_28_47#_c_1427_n N_VGND_c_2023_n 3.91258e-19 $X=0.257 $Y=0.805 $X2=0
+ $Y2=0
cc_1009 N_A_28_47#_c_1429_n N_VGND_c_2023_n 0.00226166f $X=3.355 $Y=0.79 $X2=0
+ $Y2=0
cc_1010 N_A_28_47#_c_1505_n N_VGND_c_2023_n 0.0150372f $X=4.265 $Y=0.365 $X2=0
+ $Y2=0
cc_1011 N_A_28_47#_c_1425_n N_VGND_c_2024_n 0.0209141f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_1012 N_A_28_47#_c_1427_n N_VGND_c_2024_n 2.33971e-19 $X=0.257 $Y=0.805 $X2=0
+ $Y2=0
cc_1013 N_VPWR_c_1577_n N_A_1144_49#_M1001_d 0.00562065f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1577_n N_A_1261_49#_M1021_s 0.00209319f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1015 N_VPWR_c_1585_n N_A_1261_49#_c_1814_n 0.0210382f $X=11.585 $Y=2.72 $X2=0
+ $Y2=0
cc_1016 N_VPWR_c_1577_n N_A_1261_49#_c_1814_n 0.0124268f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1017 N_VPWR_c_1577_n N_A_1634_315#_M1030_s 0.00272942f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1584_n N_A_1634_315#_c_1939_n 0.100484f $X=10.12 $Y=2.72 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1577_n N_A_1634_315#_c_1939_n 0.0412509f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1584_n N_A_1634_315#_c_1940_n 0.0121882f $X=10.12 $Y=2.72 $X2=0
+ $Y2=0
cc_1021 N_VPWR_c_1577_n N_A_1634_315#_c_1940_n 0.006547f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1577_n N_SUM_M1011_d 0.0042075f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1023 N_VPWR_c_1586_n SUM 0.0228079f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1024 N_VPWR_c_1577_n SUM 0.0124341f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1025 N_A_1144_49#_c_1730_n N_COUT_N_M1025_d 0.00324451f $X=7.05 $Y=2.04 $X2=0
+ $Y2=0
cc_1026 N_A_1144_49#_c_1706_n COUT_N 0.00590902f $X=5.895 $Y=1.555 $X2=0 $Y2=0
cc_1027 N_A_1144_49#_c_1707_n COUT_N 0.0199735f $X=7.135 $Y=1.23 $X2=0 $Y2=0
cc_1028 N_A_1144_49#_c_1709_n COUT_N 0.0205108f $X=7.135 $Y=1.955 $X2=0 $Y2=0
cc_1029 N_A_1144_49#_c_1706_n COUT_N 4.18687e-19 $X=5.895 $Y=1.555 $X2=0 $Y2=0
cc_1030 N_A_1144_49#_c_1724_n COUT_N 0.00777354f $X=6.21 $Y=1.64 $X2=0 $Y2=0
cc_1031 N_A_1144_49#_c_1730_n COUT_N 0.015187f $X=7.05 $Y=2.04 $X2=0 $Y2=0
cc_1032 N_A_1144_49#_c_1707_n N_COUT_N_c_1780_n 0.013211f $X=7.135 $Y=1.23 $X2=0
+ $Y2=0
cc_1033 N_A_1144_49#_c_1730_n N_A_1261_49#_M1004_d 0.0027538f $X=7.05 $Y=2.04
+ $X2=0 $Y2=0
cc_1034 N_A_1144_49#_c_1709_n N_A_1261_49#_M1004_d 0.00499655f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_1035 N_A_1144_49#_M1029_d N_A_1261_49#_c_1807_n 0.00648656f $X=7.14 $Y=0.245
+ $X2=0 $Y2=0
cc_1036 N_A_1144_49#_c_1707_n N_A_1261_49#_c_1807_n 0.0156983f $X=7.135 $Y=1.23
+ $X2=0 $Y2=0
cc_1037 N_A_1144_49#_c_1730_n N_A_1261_49#_c_1837_n 0.0138309f $X=7.05 $Y=2.04
+ $X2=0 $Y2=0
cc_1038 N_A_1144_49#_c_1709_n N_A_1261_49#_c_1837_n 0.0307964f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_1039 N_A_1144_49#_c_1710_n N_A_1261_49#_c_1808_n 0.0106106f $X=5.855 $Y=0.58
+ $X2=0 $Y2=0
cc_1040 N_A_1144_49#_c_1707_n N_A_1261_49#_c_1815_n 0.00833805f $X=7.135 $Y=1.23
+ $X2=0 $Y2=0
cc_1041 N_A_1144_49#_c_1709_n N_A_1261_49#_c_1815_n 0.0200829f $X=7.135 $Y=1.955
+ $X2=0 $Y2=0
cc_1042 N_A_1144_49#_c_1707_n N_A_1261_49#_c_1810_n 0.00772608f $X=7.135 $Y=1.23
+ $X2=0 $Y2=0
cc_1043 N_A_1144_49#_c_1707_n N_A_1261_49#_c_1811_n 0.0323518f $X=7.135 $Y=1.23
+ $X2=0 $Y2=0
cc_1044 N_A_1144_49#_c_1710_n N_VGND_c_2020_n 0.0096389f $X=5.855 $Y=0.58 $X2=0
+ $Y2=0
cc_1045 N_A_1144_49#_c_1710_n N_VGND_c_2023_n 0.00983468f $X=5.855 $Y=0.58 $X2=0
+ $Y2=0
cc_1046 N_COUT_N_M1013_d N_A_1261_49#_c_1807_n 0.0031917f $X=6.715 $Y=0.245
+ $X2=0 $Y2=0
cc_1047 N_COUT_N_c_1780_n N_A_1261_49#_c_1807_n 0.0160879f $X=6.745 $Y=0.925
+ $X2=0 $Y2=0
cc_1048 N_A_1261_49#_c_1809_n N_A_1634_315#_M1008_d 0.00533046f $X=11.17 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1049 N_A_1261_49#_c_1809_n N_A_1634_315#_c_1961_n 7.07302e-19 $X=11.17
+ $Y=0.85 $X2=0 $Y2=0
cc_1050 N_A_1261_49#_c_1809_n N_A_1634_315#_c_1968_n 0.0170165f $X=11.17 $Y=0.85
+ $X2=0 $Y2=0
cc_1051 N_A_1261_49#_c_1809_n N_A_1634_315#_c_1938_n 0.00841278f $X=11.17
+ $Y=0.85 $X2=0 $Y2=0
cc_1052 N_A_1261_49#_c_1858_n SUM 0.00267588f $X=11.29 $Y=0.805 $X2=0 $Y2=0
cc_1053 N_A_1261_49#_c_1870_n SUM 0.00182668f $X=11.315 $Y=0.85 $X2=0 $Y2=0
cc_1054 N_A_1261_49#_c_1809_n N_VGND_M1020_d 9.93578e-19 $X=11.17 $Y=0.85 $X2=0
+ $Y2=0
cc_1055 N_A_1261_49#_c_1809_n N_VGND_c_2017_n 8.17573e-19 $X=11.17 $Y=0.85 $X2=0
+ $Y2=0
cc_1056 N_A_1261_49#_c_1807_n N_VGND_c_2020_n 0.0662031f $X=7.53 $Y=0.34 $X2=0
+ $Y2=0
cc_1057 N_A_1261_49#_c_1808_n N_VGND_c_2020_n 0.0200489f $X=6.43 $Y=0.34 $X2=0
+ $Y2=0
cc_1058 N_A_1261_49#_c_1857_n N_VGND_c_2021_n 0.0105862f $X=11.25 $Y=0.55 $X2=0
+ $Y2=0
cc_1059 N_A_1261_49#_c_1858_n N_VGND_c_2021_n 8.99889e-19 $X=11.29 $Y=0.805
+ $X2=0 $Y2=0
cc_1060 N_A_1261_49#_c_1807_n N_VGND_c_2023_n 0.0353042f $X=7.53 $Y=0.34 $X2=0
+ $Y2=0
cc_1061 N_A_1261_49#_c_1857_n N_VGND_c_2023_n 0.00292257f $X=11.25 $Y=0.55 $X2=0
+ $Y2=0
cc_1062 N_A_1261_49#_c_1808_n N_VGND_c_2023_n 0.0122613f $X=6.43 $Y=0.34 $X2=0
+ $Y2=0
cc_1063 N_A_1261_49#_c_1858_n N_VGND_c_2023_n 9.51601e-19 $X=11.29 $Y=0.805
+ $X2=0 $Y2=0
cc_1064 N_A_1261_49#_c_1809_n N_VGND_c_2023_n 0.164575f $X=11.17 $Y=0.85 $X2=0
+ $Y2=0
cc_1065 N_A_1261_49#_c_1810_n N_VGND_c_2023_n 0.0155056f $X=7.76 $Y=0.85 $X2=0
+ $Y2=0
cc_1066 N_A_1261_49#_c_1870_n N_VGND_c_2023_n 0.0149084f $X=11.315 $Y=0.85 $X2=0
+ $Y2=0
cc_1067 N_A_1634_315#_c_1944_n N_VGND_c_2017_n 0.0220959f $X=9.825 $Y=0.4 $X2=0
+ $Y2=0
cc_1068 N_A_1634_315#_c_1944_n N_VGND_c_2020_n 0.0236293f $X=9.825 $Y=0.4 $X2=0
+ $Y2=0
cc_1069 N_A_1634_315#_c_1944_n N_VGND_c_2023_n 0.00660066f $X=9.825 $Y=0.4 $X2=0
+ $Y2=0
cc_1070 N_SUM_c_1997_n N_VGND_c_2022_n 0.0217148f $X=12.16 $Y=0.39 $X2=0 $Y2=0
cc_1071 N_SUM_M1006_d N_VGND_c_2023_n 0.00221616f $X=12.01 $Y=0.235 $X2=0 $Y2=0
cc_1072 N_SUM_c_1997_n N_VGND_c_2023_n 0.0128564f $X=12.16 $Y=0.39 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__sdfstp_1.spice
* Created: Thu Aug 27 14:46:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdfstp_1.spice.pex"
.subckt sky130_fd_sc_hd__sdfstp_1  VNB VPB SCD SCE D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1035 A_109_47# N_SCD_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_181_47#_M1011_d N_SCE_M1011_g A_109_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1018 A_265_47# N_D_M1018_g N_A_181_47#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_A_319_21#_M1027_g A_265_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1218 AS=0.0567 PD=1.42 PS=0.69 NRD=7.14 NRS=22.848 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SCE_M1012_g N_A_319_21#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_CLK_M1000_g N_A_643_369#_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_809_369#_M1033_d N_A_643_369#_M1033_g N_VGND_M1000_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_997_413#_M1019_d N_A_643_369#_M1019_g N_A_181_47#_M1019_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1020 A_1087_47# N_A_809_369#_M1020_g N_A_997_413#_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_1129_21#_M1021_g A_1087_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_1347_47# N_A_997_413#_M1007_g N_A_1129_21#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_SET_B_M1037_g A_1347_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0758774 AS=0.0441 PD=0.764717 PS=0.63 NRD=1.428 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1013 A_1514_47# N_A_997_413#_M1013_g N_VGND_M1037_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2384 AS=0.115623 PD=1.385 PS=1.16528 NRD=59.52 NRS=7.488 M=1 R=4.26667
+ SA=75000.7 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1038 N_A_1597_329#_M1038_d N_A_809_369#_M1038_g A_1514_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.149857 AS=0.2384 PD=1.3283 PS=1.385 NRD=4.68 NRS=59.52 M=1
+ R=4.26667 SA=75001.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1028 A_1815_47# N_A_643_369#_M1028_g N_A_1597_329#_M1038_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0983434 PD=0.63 PS=0.871698 NRD=14.28 NRS=44.28 M=1
+ R=2.8 SA=75002.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1030 A_1887_47# N_A_1781_295#_M1030_g A_1815_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0441 PD=0.75 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8 SA=75002.9
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_SET_B_M1036_g A_1887_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0693 PD=0.84 PS=0.75 NRD=41.424 NRS=31.428 M=1 R=2.8 SA=75003.4
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1009 N_A_1781_295#_M1009_d N_A_1597_329#_M1009_g N_VGND_M1036_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1596 AS=0.0882 PD=1.6 PS=0.84 NRD=32.856 NRS=0 M=1 R=2.8
+ SA=75003.9 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_1597_329#_M1008_g N_A_2227_47#_M1008_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0769738 AS=0.1092 PD=0.769346 PS=1.36 NRD=15.708 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1014 N_Q_M1014_d N_A_2227_47#_M1014_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.119126 PD=1.82 PS=1.19065 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1017 N_VPWR_M1017_d N_SCD_M1017_g N_A_27_369#_M1017_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 A_193_369# N_SCE_M1002_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1003 N_A_181_47#_M1003_d N_D_M1003_g A_193_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_27_369#_M1001_d N_A_319_21#_M1001_g N_A_181_47#_M1003_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_VPWR_M1024_d N_SCE_M1024_g N_A_319_21#_M1024_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.1664 PD=1.8 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1031 N_VPWR_M1031_d N_CLK_M1031_g N_A_643_369#_M1031_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1025 N_A_809_369#_M1025_d N_A_643_369#_M1025_g N_VPWR_M1031_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_997_413#_M1006_d N_A_809_369#_M1006_g N_A_181_47#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1032 A_1081_413# N_A_643_369#_M1032_g N_A_997_413#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0756 AS=0.0567 PD=0.78 PS=0.69 NRD=58.6272 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1034 N_VPWR_M1034_d N_A_1129_21#_M1034_g A_1081_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1029 AS=0.0756 PD=0.91 PS=0.78 NRD=25.7873 NRS=58.6272 M=1 R=2.8
+ SA=75001.1 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_1129_21#_M1004_d N_A_997_413#_M1004_g N_VPWR_M1034_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0714 AS=0.1029 PD=0.76 PS=0.91 NRD=9.3772 NRS=72.693 M=1
+ R=2.8 SA=75001.8 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1026 N_VPWR_M1026_d N_SET_B_M1026_g N_A_1129_21#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0952 AS=0.0714 PD=0.846667 PS=0.76 NRD=18.7544 NRS=18.7544 M=1
+ R=2.8 SA=75002.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1010 A_1525_329# N_A_997_413#_M1010_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.0882 AS=0.1904 PD=1.05 PS=1.69333 NRD=11.7215 NRS=25.7873 M=1 R=5.6
+ SA=75001.5 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1016 N_A_1597_329#_M1016_d N_A_643_369#_M1016_g A_1525_329# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2044 AS=0.0882 PD=1.76 PS=1.05 NRD=34.0022 NRS=11.7215 M=1 R=5.6
+ SA=75001.9 SB=75001 A=0.126 P=1.98 MULT=1
MM1029 A_1723_413# N_A_809_369#_M1029_g N_A_1597_329#_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0609 AS=0.1022 PD=0.71 PS=0.88 NRD=42.1974 NRS=25.7873 M=1 R=2.8
+ SA=75003.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_1781_295#_M1005_g A_1723_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0966 AS=0.0609 PD=0.88 PS=0.71 NRD=60.9715 NRS=42.1974 M=1 R=2.8
+ SA=75004.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1022 N_A_1597_329#_M1022_d N_SET_B_M1022_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0966 PD=1.36 PS=0.88 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75004.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_1781_295#_M1015_d N_A_1597_329#_M1015_g N_VPWR_M1015_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_1597_329#_M1023_g N_A_2227_47#_M1023_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.117541 AS=0.1664 PD=1.03805 PS=1.8 NRD=16.9223 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1039 N_Q_M1039_d N_A_2227_47#_M1039_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.183659 PD=2.52 PS=1.62195 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=20.544 P=28.81
c_124 VNB 0 1.07953e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__sdfstp_1.spice.SKY130_FD_SC_HD__SDFSTP_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a21o_2.pex.spice
* Created: Tue Sep  1 18:52:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21O_2%A_80_199# 1 2 9 11 13 16 18 20 22 25 26 27 31
+ 34 36 45
r72 35 45 2.02521 $w=2.38e-07 $l=1e-08 $layer=POLY_cond $X=1.085 $Y=1.235
+ $X2=1.075 $Y2=1.235
r73 34 36 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=1.16
+ $X2=1.125 $Y2=0.995
r74 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.16 $X2=1.085 $Y2=1.16
r75 29 31 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.77 $Y=0.655
+ $X2=1.77 $Y2=0.42
r76 25 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.675 $Y=0.74
+ $X2=1.77 $Y2=0.655
r77 25 26 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.675 $Y=0.74
+ $X2=1.295 $Y2=0.74
r78 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=0.825
+ $X2=1.295 $Y2=0.74
r79 23 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.21 $Y=0.825
+ $X2=1.21 $Y2=0.995
r80 22 27 25.4039 $w=2.28e-07 $l=5.07e-07 $layer=LI1_cond $X=1.125 $Y=1.805
+ $X2=1.632 $Y2=1.805
r81 21 34 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=1.125 $Y=1.165
+ $X2=1.125 $Y2=1.16
r82 21 22 17.7951 $w=3.38e-07 $l=5.25e-07 $layer=LI1_cond $X=1.125 $Y=1.165
+ $X2=1.125 $Y2=1.69
r83 18 45 13.5836 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.075 $Y=0.995
+ $X2=1.075 $Y2=1.235
r84 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.075 $Y=0.995
+ $X2=1.075 $Y2=0.56
r85 14 45 34.4286 $w=2.38e-07 $l=1.7e-07 $layer=POLY_cond $X=0.905 $Y=1.235
+ $X2=1.075 $Y2=1.235
r86 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r87 11 14 52.6555 $w=2.38e-07 $l=3.60555e-07 $layer=POLY_cond $X=0.645 $Y=0.995
+ $X2=0.905 $Y2=1.235
r88 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.645 $Y=0.995
+ $X2=0.645 $Y2=0.56
r89 7 11 34.4286 $w=2.38e-07 $l=2.33238e-07 $layer=POLY_cond $X=0.475 $Y=1.145
+ $X2=0.645 $Y2=0.995
r90 7 9 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=1.145
+ $X2=0.475 $Y2=1.985
r91 2 27 300 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=1.485 $X2=1.64 $Y2=1.88
r92 1 31 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.235 $X2=1.78 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_2%B1 1 3 6 8 15
r35 13 15 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.655 $Y=1.16
+ $X2=1.855 $Y2=1.16
r36 10 13 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.565 $Y=1.16
+ $X2=1.655 $Y2=1.16
r37 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.16 $X2=1.655 $Y2=1.16
r38 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.325
+ $X2=1.855 $Y2=1.16
r39 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.855 $Y=1.325
+ $X2=1.855 $Y2=1.985
r40 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=0.995
+ $X2=1.565 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.565 $Y=0.995
+ $X2=1.565 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_2%A1 3 6 8 9 13 15
c39 15 0 1.66259e-19 $X=2.3 $Y=0.995
r40 13 16 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.16 $X2=2.3
+ $Y2=1.325
r41 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.16 $X2=2.3
+ $Y2=0.995
r42 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=1.16 $X2=2.325 $Y2=1.16
r43 9 14 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=2.43 $Y=0.85 $X2=2.43
+ $Y2=1.16
r44 8 9 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=2.43 $Y=0.51 $X2=2.43
+ $Y2=0.85
r45 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.285 $Y=1.985
+ $X2=2.285 $Y2=1.325
r46 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.215 $Y=0.56
+ $X2=2.215 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_2%A2 1 3 6 8 11 18
c28 8 0 1.66259e-19 $X=2.91 $Y=1.105
r29 14 18 1.97613 $w=5.73e-07 $l=9.5e-08 $layer=LI1_cond $X=2.895 $Y=1.037
+ $X2=2.99 $Y2=1.037
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.895
+ $Y=1.16 $X2=2.895 $Y2=1.16
r31 11 13 24.0172 $w=2.91e-07 $l=1.45e-07 $layer=POLY_cond $X=2.75 $Y=1.155
+ $X2=2.895 $Y2=1.155
r32 10 11 0.828179 $w=2.91e-07 $l=5e-09 $layer=POLY_cond $X=2.745 $Y=1.155
+ $X2=2.75 $Y2=1.155
r33 8 18 0.104007 $w=5.73e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=1.037
+ $X2=2.99 $Y2=1.037
r34 4 11 18.2534 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.75 $Y=1.305
+ $X2=2.75 $Y2=1.155
r35 4 6 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.75 $Y=1.305 $X2=2.75
+ $Y2=1.985
r36 1 10 18.2534 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.745 $Y=1.005
+ $X2=2.745 $Y2=1.155
r37 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.745 $Y=1.005
+ $X2=2.745 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_2%VPWR 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r46 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=2.72
+ $X2=2.52 $Y2=2.72
r51 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.685 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r53 33 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.12 $Y2=2.72
r56 30 32 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.52 $Y2=2.72
r58 29 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 25 40 4.40339 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r62 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=1.12 $Y2=2.72
r64 24 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 22 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.635
+ $X2=2.52 $Y2=2.72
r68 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.52 $Y=2.635
+ $X2=2.52 $Y2=2.34
r69 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r70 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.34
r71 10 40 3.03446 $w=2.9e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.192 $Y2=2.72
r72 10 12 31.3941 $w=2.88e-07 $l=7.9e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=1.845
r73 3 20 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.485 $X2=2.52 $Y2=2.34
r74 2 16 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=2.34
r75 1 12 300 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_2%X 1 2 9 14 16 19
r19 16 19 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.67 $Y=2.21
+ $X2=0.67 $Y2=1.825
r20 12 19 50.1062 $w=2.28e-07 $l=1e-06 $layer=LI1_cond $X=0.67 $Y=0.825 $X2=0.67
+ $Y2=1.825
r21 12 14 11.0909 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.67 $Y=0.73
+ $X2=0.86 $Y2=0.73
r22 7 14 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.86 $Y=0.635
+ $X2=0.86 $Y2=0.73
r23 7 9 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=0.86 $Y=0.635
+ $X2=0.86 $Y2=0.42
r24 2 19 300 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.825
r25 1 9 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.72
+ $Y=0.235 $X2=0.86 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_2%A_386_297# 1 2 7 9 11 13 15
r17 13 20 3.77276 $w=2.2e-07 $l=1.33e-07 $layer=LI1_cond $X=2.965 $Y=1.935
+ $X2=2.965 $Y2=1.802
r18 13 15 19.1201 $w=2.18e-07 $l=3.65e-07 $layer=LI1_cond $X=2.965 $Y=1.935
+ $X2=2.965 $Y2=2.3
r19 12 18 3.15837 $w=2.65e-07 $l=1.13e-07 $layer=LI1_cond $X=2.185 $Y=1.802
+ $X2=2.072 $Y2=1.802
r20 11 20 3.12033 $w=2.65e-07 $l=1.1e-07 $layer=LI1_cond $X=2.855 $Y=1.802
+ $X2=2.965 $Y2=1.802
r21 11 12 29.1372 $w=2.63e-07 $l=6.7e-07 $layer=LI1_cond $X=2.855 $Y=1.802
+ $X2=2.185 $Y2=1.802
r22 7 18 3.71737 $w=2.25e-07 $l=1.33e-07 $layer=LI1_cond $X=2.072 $Y=1.935
+ $X2=2.072 $Y2=1.802
r23 7 9 18.6952 $w=2.23e-07 $l=3.65e-07 $layer=LI1_cond $X=2.072 $Y=1.935
+ $X2=2.072 $Y2=2.3
r24 2 20 600 $w=1.7e-07 $l=4.272e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.85
r25 2 15 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=2.3
r26 1 18 600 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.485 $X2=2.07 $Y2=1.85
r27 1 9 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.485 $X2=2.07 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A21O_2%VGND 1 2 3 10 12 14 18 20 22 24 26 38 42
r52 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r53 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r55 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r56 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r57 30 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r58 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r59 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r60 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.29
+ $Y2=0
r61 27 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.61
+ $Y2=0
r62 26 41 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=3.012
+ $Y2=0
r63 26 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.53
+ $Y2=0
r64 24 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r65 24 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 20 41 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=3.012 $Y2=0
r67 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0.38
r68 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=0.085
+ $X2=1.29 $Y2=0
r69 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.29 $Y=0.085
+ $X2=1.29 $Y2=0.36
r70 15 35 4.48512 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.297
+ $Y2=0
r71 14 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.29
+ $Y2=0
r72 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.595
+ $Y2=0
r73 10 35 3.28106 $w=3.3e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.43 $Y=0.085
+ $X2=0.297 $Y2=0
r74 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.43 $Y=0.085
+ $X2=0.43 $Y2=0.38
r75 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.235 $X2=2.96 $Y2=0.38
r76 2 18 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.15
+ $Y=0.235 $X2=1.29 $Y2=0.36
r77 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.305
+ $Y=0.235 $X2=0.43 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a311oi_4.pex.spice
* Created: Tue Sep  1 18:54:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A311OI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 47
r70 45 47 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.73 $Y2=1.16
r71 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.395
+ $Y=1.16 $X2=1.395 $Y2=1.16
r72 43 45 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.395 $Y2=1.16
r73 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r74 41 42 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r75 38 41 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.285 $Y=1.16
+ $X2=0.47 $Y2=1.16
r76 32 46 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=1.395 $Y2=1.16
r77 31 46 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=1.395 $Y2=1.16
r78 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=1.155 $Y2=1.16
r79 29 30 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.16
+ $X2=0.695 $Y2=1.16
r80 29 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=1.16 $X2=0.285 $Y2=1.16
r81 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r82 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r83 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r84 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r85 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r86 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r87 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r88 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r89 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r90 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r91 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r92 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r93 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r94 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r95 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r96 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 47
r71 45 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.32 $Y=1.16 $X2=3.41
+ $Y2=1.16
r72 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.32
+ $Y=1.16 $X2=3.32 $Y2=1.16
r73 43 45 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.32 $Y2=1.16
r74 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r75 40 42 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.21 $Y=1.16
+ $X2=2.57 $Y2=1.16
r76 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.21
+ $Y=1.16 $X2=2.21 $Y2=1.16
r77 37 40 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.15 $Y=1.16 $X2=2.21
+ $Y2=1.16
r78 32 46 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.455 $Y=1.16
+ $X2=3.32 $Y2=1.16
r79 31 46 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=3.32 $Y2=1.16
r80 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.16
+ $X2=2.995 $Y2=1.16
r81 30 41 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.535 $Y=1.16
+ $X2=2.21 $Y2=1.16
r82 29 41 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.075 $Y=1.16
+ $X2=2.21 $Y2=1.16
r83 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r85 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r87 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r89 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r91 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r93 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r95 4 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
r97 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995 $X2=2.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%A1 3 7 9 11 14 16 18 21 23 25 26 28 29 30
+ 31 32 49
c68 32 0 1.99742e-19 $X=5.295 $Y=1.19
r69 49 50 58.8488 $w=3.44e-07 $l=4.2e-07 $layer=POLY_cond $X=5.19 $Y=1.17
+ $X2=5.61 $Y2=1.17
r70 48 49 14.0116 $w=3.44e-07 $l=1e-07 $layer=POLY_cond $X=5.09 $Y=1.17 $X2=5.19
+ $Y2=1.17
r71 46 48 12.6105 $w=3.44e-07 $l=9e-08 $layer=POLY_cond $X=5 $Y=1.17 $X2=5.09
+ $Y2=1.17
r72 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5 $Y=1.16
+ $X2=5 $Y2=1.16
r73 44 46 32.2267 $w=3.44e-07 $l=2.3e-07 $layer=POLY_cond $X=4.77 $Y=1.17 $X2=5
+ $Y2=1.17
r74 43 44 14.0116 $w=3.44e-07 $l=1e-07 $layer=POLY_cond $X=4.67 $Y=1.17 $X2=4.77
+ $Y2=1.17
r75 42 43 44.8372 $w=3.44e-07 $l=3.2e-07 $layer=POLY_cond $X=4.35 $Y=1.17
+ $X2=4.67 $Y2=1.17
r76 41 42 14.0116 $w=3.44e-07 $l=1e-07 $layer=POLY_cond $X=4.25 $Y=1.17 $X2=4.35
+ $Y2=1.17
r77 39 41 50.4419 $w=3.44e-07 $l=3.6e-07 $layer=POLY_cond $X=3.89 $Y=1.17
+ $X2=4.25 $Y2=1.17
r78 37 39 8.40698 $w=3.44e-07 $l=6e-08 $layer=POLY_cond $X=3.83 $Y=1.17 $X2=3.89
+ $Y2=1.17
r79 32 47 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.295 $Y=1.16 $X2=5
+ $Y2=1.16
r80 31 47 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=1.16 $X2=5
+ $Y2=1.16
r81 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.375 $Y=1.16
+ $X2=4.835 $Y2=1.16
r82 29 30 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.89 $Y=1.16
+ $X2=4.375 $Y2=1.16
r83 29 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.89
+ $Y=1.16 $X2=3.89 $Y2=1.16
r84 26 50 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.17
r85 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r86 23 49 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.17
r87 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r88 19 48 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.09 $Y=1.345
+ $X2=5.09 $Y2=1.17
r89 19 21 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.09 $Y=1.345
+ $X2=5.09 $Y2=1.985
r90 16 44 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.17
r91 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r92 12 43 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.67 $Y=1.345
+ $X2=4.67 $Y2=1.17
r93 12 14 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.67 $Y=1.345
+ $X2=4.67 $Y2=1.985
r94 9 42 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.17
r95 9 11 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
r96 5 41 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.25 $Y=1.345
+ $X2=4.25 $Y2=1.17
r97 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.25 $Y=1.345 $X2=4.25
+ $Y2=1.985
r98 1 37 22.2144 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.83 $Y=1.345
+ $X2=3.83 $Y2=1.17
r99 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.83 $Y=1.345 $X2=3.83
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 31 33
+ 48 50
c70 50 0 1.99742e-19 $X=7.29 $Y=1.16
r71 49 50 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.87 $Y=1.16
+ $X2=7.29 $Y2=1.16
r72 47 49 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.77 $Y=1.16 $X2=6.87
+ $Y2=1.16
r73 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.16 $X2=6.77 $Y2=1.16
r74 45 47 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=6.45 $Y=1.16
+ $X2=6.77 $Y2=1.16
r75 43 45 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.03 $Y=1.16
+ $X2=6.45 $Y2=1.16
r76 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.03
+ $Y=1.16 $X2=6.03 $Y2=1.16
r77 33 48 1.41269 $w=6.33e-07 $l=7.5e-08 $layer=LI1_cond $X=6.695 $Y=1.312
+ $X2=6.77 $Y2=1.312
r78 31 33 8.66451 $w=6.33e-07 $l=4.6e-07 $layer=LI1_cond $X=6.235 $Y=1.312
+ $X2=6.695 $Y2=1.312
r79 31 44 3.86136 $w=6.33e-07 $l=2.05e-07 $layer=LI1_cond $X=6.235 $Y=1.312
+ $X2=6.03 $Y2=1.312
r80 29 44 4.80315 $w=6.33e-07 $l=2.55e-07 $layer=LI1_cond $X=5.775 $Y=1.312
+ $X2=6.03 $Y2=1.312
r81 25 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.16
r82 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.985
r83 22 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=1.16
r84 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=0.56
r85 18 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.16
r86 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.985
r87 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=1.16
r88 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=0.56
r89 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r90 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r91 8 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r92 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r93 4 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r94 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325 $X2=6.03
+ $Y2=1.985
r95 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r96 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995 $X2=6.03
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%C1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 46
c74 20 0 7.42849e-20 $X=8.77 $Y=1.985
r75 44 46 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=9.19 $Y=1.16
+ $X2=9.415 $Y2=1.16
r76 43 44 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.77 $Y=1.16
+ $X2=9.19 $Y2=1.16
r77 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.35 $Y=1.16
+ $X2=8.77 $Y2=1.16
r78 40 42 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=8.305 $Y=1.16
+ $X2=8.35 $Y2=1.16
r79 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.305
+ $Y=1.16 $X2=8.305 $Y2=1.16
r80 37 40 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=7.93 $Y=1.16
+ $X2=8.305 $Y2=1.16
r81 32 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.415
+ $Y=1.16 $X2=9.415 $Y2=1.16
r82 31 32 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.965 $Y=1.16
+ $X2=9.415 $Y2=1.16
r83 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=8.505 $Y=1.16
+ $X2=8.965 $Y2=1.16
r84 30 41 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=8.505 $Y=1.16 $X2=8.305
+ $Y2=1.16
r85 29 41 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=8.045 $Y=1.16
+ $X2=8.305 $Y2=1.16
r86 25 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.19 $Y=1.325
+ $X2=9.19 $Y2=1.16
r87 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.19 $Y=1.325
+ $X2=9.19 $Y2=1.985
r88 22 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.19 $Y=0.995
+ $X2=9.19 $Y2=1.16
r89 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.19 $Y=0.995
+ $X2=9.19 $Y2=0.56
r90 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.77 $Y=1.325
+ $X2=8.77 $Y2=1.16
r91 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.77 $Y=1.325
+ $X2=8.77 $Y2=1.985
r92 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.77 $Y=0.995
+ $X2=8.77 $Y2=1.16
r93 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.77 $Y=0.995
+ $X2=8.77 $Y2=0.56
r94 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.35 $Y=1.325
+ $X2=8.35 $Y2=1.16
r95 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.35 $Y=1.325
+ $X2=8.35 $Y2=1.985
r96 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.35 $Y=0.995
+ $X2=8.35 $Y2=1.16
r97 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.35 $Y=0.995
+ $X2=8.35 $Y2=0.56
r98 4 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.93 $Y=1.325
+ $X2=7.93 $Y2=1.16
r99 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.93 $Y=1.325 $X2=7.93
+ $Y2=1.985
r100 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.93 $Y=0.995
+ $X2=7.93 $Y2=1.16
r101 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.93 $Y=0.995
+ $X2=7.93 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 44 48
+ 52 55 56 58 59 60 61 62 64 79 89 90 96 99 102
r137 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r138 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r139 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 89 90 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r141 87 90 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=9.43 $Y2=2.72
r142 87 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r143 86 89 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=9.43 $Y2=2.72
r144 86 87 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r145 84 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.3 $Y2=2.72
r146 84 86 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.75 $Y2=2.72
r147 83 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r148 83 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r149 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r150 80 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.46 $Y2=2.72
r151 80 82 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.83 $Y2=2.72
r152 79 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=5.3 $Y2=2.72
r153 79 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=4.83 $Y2=2.72
r154 78 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r155 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r156 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r157 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r158 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r159 72 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r160 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r161 69 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.1 $Y2=2.72
r162 69 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.61 $Y2=2.72
r163 68 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r164 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r165 65 93 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r166 65 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r167 64 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.1 $Y2=2.72
r168 64 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r169 62 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r170 62 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r171 60 77 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.45 $Y2=2.72
r172 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.62 $Y2=2.72
r173 58 74 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.53 $Y2=2.72
r174 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.78 $Y2=2.72
r175 57 77 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.45 $Y2=2.72
r176 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.78 $Y2=2.72
r177 55 71 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.61 $Y2=2.72
r178 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.94 $Y2=2.72
r179 54 74 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.53 $Y2=2.72
r180 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=1.94 $Y2=2.72
r181 50 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.72
r182 50 52 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.34
r183 46 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2.72
r184 46 48 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2
r185 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.62 $Y2=2.72
r186 44 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=4.46 $Y2=2.72
r187 44 45 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=3.785 $Y2=2.72
r188 40 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r189 40 42 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2
r190 36 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r191 36 38 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r192 32 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r193 32 34 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r194 28 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r195 28 30 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r196 24 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r197 22 93 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r198 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r199 7 52 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=2.34
r200 6 48 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=2
r201 5 42 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2
r202 4 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r203 3 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r204 2 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r205 1 27 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r206 1 24 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%A_109_297# 1 2 3 4 5 6 7 8 27 29 30 33 35
+ 39 41 45 47 51 53 59 65 67 68 69 70
r82 63 65 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.24 $Y=2 $X2=7.08
+ $Y2=2
r83 61 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=2 $X2=4.88
+ $Y2=2
r84 61 63 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=4.965 $Y=2
+ $X2=6.24 $Y2=2
r85 57 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=2.085
+ $X2=4.88 $Y2=2
r86 57 59 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.88 $Y=2.085
+ $X2=4.88 $Y2=2.3
r87 56 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=1.915
+ $X2=4.88 $Y2=2
r88 55 56 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.88 $Y=1.665
+ $X2=4.88 $Y2=1.915
r89 54 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=1.58
+ $X2=4.04 $Y2=1.58
r90 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.795 $Y=1.58
+ $X2=4.88 $Y2=1.665
r91 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.795 $Y=1.58
+ $X2=4.125 $Y2=1.58
r92 49 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=1.58
r93 49 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=1.96
r94 48 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=1.58 $X2=3.2
+ $Y2=1.58
r95 47 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=1.58
+ $X2=4.04 $Y2=1.58
r96 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.955 $Y=1.58
+ $X2=3.285 $Y2=1.58
r97 43 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=1.665 $X2=3.2
+ $Y2=1.58
r98 43 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.2 $Y=1.665 $X2=3.2
+ $Y2=1.96
r99 42 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=2.36 $Y2=1.58
r100 41 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=1.58
+ $X2=3.2 $Y2=1.58
r101 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.115 $Y=1.58
+ $X2=2.445 $Y2=1.58
r102 37 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=1.58
r103 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=1.96
r104 36 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.58
+ $X2=1.52 $Y2=1.58
r105 35 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=1.58
+ $X2=2.36 $Y2=1.58
r106 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.275 $Y=1.58
+ $X2=1.605 $Y2=1.58
r107 31 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.58
r108 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.96
r109 29 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=1.58
+ $X2=1.52 $Y2=1.58
r110 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=1.58
+ $X2=0.765 $Y2=1.58
r111 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.765 $Y2=1.58
r112 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.96
r113 8 65 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=2
r114 7 63 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=2
r115 6 72 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=1.96
r116 6 59 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=2.3
r117 5 51 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=1.96
r118 4 45 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.96
r119 3 39 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.96
r120 2 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r121 1 27 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%A_1139_297# 1 2 3 4 5 16 26 28
r41 26 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.44 $Y=2.255
+ $X2=9.44 $Y2=2.34
r42 26 28 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=9.44 $Y=2.255
+ $X2=9.44 $Y2=2
r43 23 25 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=7.5 $Y=2.34
+ $X2=8.56 $Y2=2.34
r44 21 23 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.66 $Y=2.34 $X2=7.5
+ $Y2=2.34
r45 18 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.82 $Y=2.34
+ $X2=6.66 $Y2=2.34
r46 16 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.315 $Y=2.34
+ $X2=9.44 $Y2=2.34
r47 16 25 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.315 $Y=2.34
+ $X2=8.56 $Y2=2.34
r48 5 31 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.485 $X2=9.4 $Y2=2.34
r49 5 28 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.485 $X2=9.4 $Y2=2
r50 4 25 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.425
+ $Y=1.485 $X2=8.56 $Y2=2.34
r51 3 23 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=2.34
r52 2 21 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=2.34
r53 1 18 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.485 $X2=5.82 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%Y 1 2 3 4 5 6 7 8 9 28 38 40 44 46 48 52 56
+ 58 64 66 68 69 71 72 73 74 75 85 91
c110 68 0 7.42849e-20 $X=8.14 $Y=1.63
r111 83 91 0.540208 $w=3.18e-07 $l=1.5e-08 $layer=LI1_cond $X=7.575 $Y=1.545
+ $X2=7.575 $Y2=1.53
r112 82 85 1.62062 $w=3.18e-07 $l=4.5e-08 $layer=LI1_cond $X=7.575 $Y=0.805
+ $X2=7.575 $Y2=0.85
r113 75 94 8.64332 $w=3.18e-07 $l=2.4e-07 $layer=LI1_cond $X=7.575 $Y=1.87
+ $X2=7.575 $Y2=1.63
r114 74 94 1.80069 $w=3.18e-07 $l=5e-08 $layer=LI1_cond $X=7.575 $Y=1.58
+ $X2=7.575 $Y2=1.63
r115 74 83 1.26048 $w=3.18e-07 $l=3.5e-08 $layer=LI1_cond $X=7.575 $Y=1.58
+ $X2=7.575 $Y2=1.545
r116 74 91 1.26048 $w=3.18e-07 $l=3.5e-08 $layer=LI1_cond $X=7.575 $Y=1.495
+ $X2=7.575 $Y2=1.53
r117 73 74 10.9842 $w=3.18e-07 $l=3.05e-07 $layer=LI1_cond $X=7.575 $Y=1.19
+ $X2=7.575 $Y2=1.495
r118 72 82 2.01537 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.575 $Y=0.72
+ $X2=7.575 $Y2=0.805
r119 72 73 11.5244 $w=3.18e-07 $l=3.2e-07 $layer=LI1_cond $X=7.575 $Y=0.87
+ $X2=7.575 $Y2=1.19
r120 72 85 0.720277 $w=3.18e-07 $l=2e-08 $layer=LI1_cond $X=7.575 $Y=0.87
+ $X2=7.575 $Y2=0.85
r121 62 64 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.4 $Y=0.635
+ $X2=9.4 $Y2=0.42
r122 59 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.645 $Y=0.72
+ $X2=8.56 $Y2=0.72
r123 58 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.315 $Y=0.72
+ $X2=9.4 $Y2=0.635
r124 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.315 $Y=0.72
+ $X2=8.645 $Y2=0.72
r125 54 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.56 $Y=0.635
+ $X2=8.56 $Y2=0.72
r126 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.56 $Y=0.635
+ $X2=8.56 $Y2=0.42
r127 53 68 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=8.305 $Y=1.63
+ $X2=8.14 $Y2=1.622
r128 52 71 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.815 $Y=1.63
+ $X2=8.98 $Y2=1.63
r129 52 53 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.815 $Y=1.63
+ $X2=8.305 $Y2=1.63
r130 49 94 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.735 $Y=1.63
+ $X2=7.575 $Y2=1.63
r131 48 68 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=7.975 $Y=1.63
+ $X2=8.14 $Y2=1.622
r132 48 49 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.975 $Y=1.63
+ $X2=7.735 $Y2=1.63
r133 47 72 4.23144 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.735 $Y=0.72
+ $X2=7.575 $Y2=0.72
r134 46 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.475 $Y=0.72
+ $X2=8.56 $Y2=0.72
r135 46 47 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=8.475 $Y=0.72
+ $X2=7.735 $Y2=0.72
r136 42 72 2.01537 $w=1.7e-07 $l=1.16619e-07 $layer=LI1_cond $X=7.5 $Y=0.635
+ $X2=7.575 $Y2=0.72
r137 42 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.5 $Y=0.635
+ $X2=7.5 $Y2=0.42
r138 41 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0.72
+ $X2=6.66 $Y2=0.72
r139 40 72 4.23144 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.415 $Y=0.72
+ $X2=7.575 $Y2=0.72
r140 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.415 $Y=0.72
+ $X2=6.745 $Y2=0.72
r141 36 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0.635
+ $X2=6.66 $Y2=0.72
r142 36 38 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.66 $Y=0.635
+ $X2=6.66 $Y2=0.42
r143 33 35 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.98 $Y=0.72
+ $X2=5.82 $Y2=0.72
r144 30 33 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.72
+ $X2=4.98 $Y2=0.72
r145 28 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0.72
+ $X2=6.66 $Y2=0.72
r146 28 35 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.575 $Y=0.72
+ $X2=5.82 $Y2=0.72
r147 9 71 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.845
+ $Y=1.485 $X2=8.98 $Y2=1.63
r148 8 68 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.005
+ $Y=1.485 $X2=8.14 $Y2=1.63
r149 7 64 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.265
+ $Y=0.235 $X2=9.4 $Y2=0.42
r150 6 56 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.425
+ $Y=0.235 $X2=8.56 $Y2=0.42
r151 5 44 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.5 $Y2=0.42
r152 4 38 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.42
r153 3 35 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.72
r154 2 33 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.72
r155 1 30 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 30 36 38
+ 39
r50 34 36 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=0.72
+ $X2=3.62 $Y2=0.72
r51 32 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.72
+ $X2=1.94 $Y2=0.72
r52 32 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.72
+ $X2=2.78 $Y2=0.72
r53 28 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.635
+ $X2=1.94 $Y2=0.72
r54 28 30 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.94 $Y=0.635
+ $X2=1.94 $Y2=0.42
r55 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.72 $X2=1.1
+ $Y2=0.72
r56 26 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0.72
+ $X2=1.94 $Y2=0.72
r57 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=0.72
+ $X2=1.185 $Y2=0.72
r58 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.635 $X2=1.1
+ $Y2=0.72
r59 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.1 $Y=0.635
+ $X2=1.1 $Y2=0.42
r60 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.72 $X2=1.1
+ $Y2=0.72
r61 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.72
+ $X2=0.345 $Y2=0.72
r62 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r63 16 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.42
r64 5 36 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.72
r65 4 34 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.72
r66 3 30 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.42
r67 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.42
r68 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%VGND 1 2 3 4 5 6 21 25 29 33 35 39 43 45 47
+ 52 57 62 67 74 75 78 81 84 87 90 93
r150 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r151 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r152 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r153 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r154 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r155 81 82 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r156 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r157 75 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=8.97
+ $Y2=0
r158 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r159 72 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=0 $X2=8.98
+ $Y2=0
r160 72 74 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.145 $Y=0
+ $X2=9.43 $Y2=0
r161 71 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.97
+ $Y2=0
r162 71 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.05
+ $Y2=0
r163 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r164 68 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.305 $Y=0 $X2=8.14
+ $Y2=0
r165 68 70 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.305 $Y=0
+ $X2=8.51 $Y2=0
r166 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.815 $Y=0 $X2=8.98
+ $Y2=0
r167 67 70 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.815 $Y=0
+ $X2=8.51 $Y2=0
r168 66 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r169 66 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r170 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r171 63 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=0 $X2=6.24
+ $Y2=0
r172 63 65 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.405 $Y=0
+ $X2=6.67 $Y2=0
r173 62 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=7.08
+ $Y2=0
r174 62 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.67
+ $Y2=0
r175 61 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r176 61 82 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=1.61
+ $Y2=0
r177 60 61 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r178 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.52
+ $Y2=0
r179 58 60 265.203 $w=1.68e-07 $l=4.065e-06 $layer=LI1_cond $X=1.685 $Y=0
+ $X2=5.75 $Y2=0
r180 57 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0 $X2=6.24
+ $Y2=0
r181 57 60 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=5.75 $Y2=0
r182 56 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r183 56 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r184 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r185 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r186 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r187 52 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.52
+ $Y2=0
r188 52 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.15 $Y2=0
r189 47 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r190 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r191 45 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r192 45 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r193 41 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=8.98 $Y2=0
r194 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=8.98 $Y2=0.38
r195 37 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.14 $Y=0.085
+ $X2=8.14 $Y2=0
r196 37 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.14 $Y=0.085
+ $X2=8.14 $Y2=0.38
r197 36 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=0 $X2=7.08
+ $Y2=0
r198 35 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=8.14
+ $Y2=0
r199 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.975 $Y=0
+ $X2=7.245 $Y2=0
r200 31 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0
r201 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0.38
r202 27 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=0.085
+ $X2=6.24 $Y2=0
r203 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.24 $Y=0.085
+ $X2=6.24 $Y2=0.38
r204 23 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r205 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.38
r206 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r207 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r208 6 43 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.845
+ $Y=0.235 $X2=8.98 $Y2=0.38
r209 5 39 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.005
+ $Y=0.235 $X2=8.14 $Y2=0.38
r210 4 33 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.38
r211 3 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.38
r212 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r213 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_4%A_445_47# 1 2 3 4 21
r29 19 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=0.38 $X2=5.4
+ $Y2=0.38
r30 17 19 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.2 $Y=0.38
+ $X2=4.56 $Y2=0.38
r31 14 17 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.38 $X2=3.2
+ $Y2=0.38
r32 4 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.38
r33 3 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.38
r34 2 17 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.38
r35 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.38
.ends


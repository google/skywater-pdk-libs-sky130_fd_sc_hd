* File: sky130_fd_sc_hd__sdlclkp_1.pxi.spice
* Created: Tue Sep  1 19:31:36 2020
* 
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%SCE N_SCE_M1020_g N_SCE_M1010_g SCE SCE
+ N_SCE_c_138_n PM_SKY130_FD_SC_HD__SDLCLKP_1%SCE
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%GATE N_GATE_M1005_g N_GATE_M1008_g GATE GATE
+ N_GATE_c_167_n PM_SKY130_FD_SC_HD__SDLCLKP_1%GATE
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%A_256_147# N_A_256_147#_M1014_d
+ N_A_256_147#_M1006_d N_A_256_147#_M1019_g N_A_256_147#_M1007_g
+ N_A_256_147#_M1011_g N_A_256_147#_M1015_g N_A_256_147#_c_208_n
+ N_A_256_147#_c_209_n N_A_256_147#_c_210_n N_A_256_147#_c_211_n
+ N_A_256_147#_c_218_n N_A_256_147#_c_212_n N_A_256_147#_c_213_n
+ N_A_256_147#_c_214_n N_A_256_147#_c_215_n N_A_256_147#_c_220_n
+ N_A_256_147#_c_232_n N_A_256_147#_c_221_n N_A_256_147#_c_222_n
+ N_A_256_147#_c_223_n N_A_256_147#_c_224_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_1%A_256_147#
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%A_256_243# N_A_256_243#_M1011_s
+ N_A_256_243#_M1015_s N_A_256_243#_M1021_g N_A_256_243#_c_377_n
+ N_A_256_243#_c_378_n N_A_256_243#_M1000_g N_A_256_243#_c_379_n
+ N_A_256_243#_c_380_n N_A_256_243#_c_381_n N_A_256_243#_c_393_n
+ N_A_256_243#_c_382_n N_A_256_243#_c_383_n N_A_256_243#_c_384_n
+ N_A_256_243#_c_385_n N_A_256_243#_c_386_n N_A_256_243#_c_387_n
+ N_A_256_243#_c_388_n PM_SKY130_FD_SC_HD__SDLCLKP_1%A_256_243#
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%A_464_315# N_A_464_315#_M1003_d
+ N_A_464_315#_M1001_d N_A_464_315#_M1017_g N_A_464_315#_M1018_g
+ N_A_464_315#_M1002_g N_A_464_315#_M1016_g N_A_464_315#_c_499_n
+ N_A_464_315#_c_494_n N_A_464_315#_c_513_n N_A_464_315#_c_501_n
+ N_A_464_315#_c_502_n N_A_464_315#_c_503_n N_A_464_315#_c_525_n
+ N_A_464_315#_c_526_n N_A_464_315#_c_504_n N_A_464_315#_c_505_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_1%A_464_315#
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%A_286_413# N_A_286_413#_M1019_d
+ N_A_286_413#_M1021_d N_A_286_413#_c_624_n N_A_286_413#_M1003_g
+ N_A_286_413#_M1001_g N_A_286_413#_c_635_n N_A_286_413#_c_639_n
+ N_A_286_413#_c_630_n N_A_286_413#_c_625_n N_A_286_413#_c_626_n
+ N_A_286_413#_c_627_n N_A_286_413#_c_628_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_1%A_286_413#
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%CLK N_CLK_M1014_g N_CLK_c_724_n N_CLK_M1006_g
+ N_CLK_M1004_g N_CLK_M1012_g N_CLK_c_727_n N_CLK_c_728_n N_CLK_c_729_n
+ N_CLK_c_730_n CLK N_CLK_c_731_n N_CLK_c_735_n N_CLK_c_732_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_1%CLK
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%A_1012_47# N_A_1012_47#_M1002_s
+ N_A_1012_47#_M1016_d N_A_1012_47#_M1013_g N_A_1012_47#_M1009_g
+ N_A_1012_47#_c_798_n N_A_1012_47#_c_799_n N_A_1012_47#_c_800_n
+ N_A_1012_47#_c_801_n N_A_1012_47#_c_802_n N_A_1012_47#_c_803_n
+ N_A_1012_47#_c_804_n PM_SKY130_FD_SC_HD__SDLCLKP_1%A_1012_47#
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%VPWR N_VPWR_M1010_s N_VPWR_M1017_d
+ N_VPWR_M1015_d N_VPWR_M1016_s N_VPWR_M1012_d N_VPWR_c_857_n N_VPWR_c_858_n
+ N_VPWR_c_859_n N_VPWR_c_860_n N_VPWR_c_861_n VPWR N_VPWR_c_862_n
+ N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_856_n N_VPWR_c_866_n N_VPWR_c_867_n
+ N_VPWR_c_868_n N_VPWR_c_869_n PM_SKY130_FD_SC_HD__SDLCLKP_1%VPWR
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%A_27_47# N_A_27_47#_M1020_s N_A_27_47#_M1008_d
+ N_A_27_47#_M1005_d N_A_27_47#_c_948_n N_A_27_47#_c_952_n N_A_27_47#_c_949_n
+ N_A_27_47#_c_950_n N_A_27_47#_c_959_n N_A_27_47#_c_969_n N_A_27_47#_c_979_n
+ N_A_27_47#_c_951_n N_A_27_47#_c_954_n PM_SKY130_FD_SC_HD__SDLCLKP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%GCLK N_GCLK_M1013_d N_GCLK_M1009_d
+ N_GCLK_c_1004_n N_GCLK_c_1007_n N_GCLK_c_1005_n GCLK GCLK GCLK N_GCLK_c_1006_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_1%GCLK
x_PM_SKY130_FD_SC_HD__SDLCLKP_1%VGND N_VGND_M1020_d N_VGND_M1018_d
+ N_VGND_M1011_d N_VGND_M1004_d N_VGND_c_1021_n N_VGND_c_1022_n N_VGND_c_1023_n
+ VGND N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n
+ N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n
+ N_VGND_c_1032_n N_VGND_c_1033_n PM_SKY130_FD_SC_HD__SDLCLKP_1%VGND
cc_1 VNB N_SCE_M1020_g 0.0353283f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB SCE 0.0152489f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_SCE_c_138_n 0.0345609f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_GATE_M1008_g 0.0275832f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_5 VNB GATE 0.00454478f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_6 VNB N_GATE_c_167_n 0.027114f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_7 VNB N_A_256_147#_M1019_g 0.019494f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_256_147#_M1011_g 0.0381097f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_9 VNB N_A_256_147#_c_208_n 0.00683226f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_256_147#_c_209_n 0.0268988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_256_147#_c_210_n 7.88187e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_256_147#_c_211_n 0.00847412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_256_147#_c_212_n 0.00234051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_256_147#_c_213_n 0.00341068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_256_147#_c_214_n 0.00214682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_256_147#_c_215_n 0.0238041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_256_243#_c_377_n 0.0152184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_256_243#_c_378_n 0.00503804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_256_243#_c_379_n 0.0111999f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_20 VNB N_A_256_243#_c_380_n 0.00769152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_256_243#_c_381_n 0.00732811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_256_243#_c_382_n 0.00867647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_256_243#_c_383_n 0.00127255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_256_243#_c_384_n 0.00212966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_256_243#_c_385_n 0.00436356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_256_243#_c_386_n 0.0269987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_256_243#_c_387_n 0.00250527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_256_243#_c_388_n 0.0189173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_464_315#_M1018_g 0.0445515f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_30 VNB N_A_464_315#_M1002_g 0.0483469f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_31 VNB N_A_464_315#_c_494_n 0.00912014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_286_413#_c_624_n 0.0210526f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_33 VNB N_A_286_413#_c_625_n 0.0018369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_286_413#_c_626_n 0.00624625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_286_413#_c_627_n 0.00187427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_286_413#_c_628_n 0.0292618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_CLK_c_724_n 0.0200497f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_38 VNB N_CLK_M1004_g 0.0246477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_CLK_M1012_g 0.00619163f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_40 VNB N_CLK_c_727_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_41 VNB N_CLK_c_728_n 0.0303536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_CLK_c_729_n 0.0183112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_CLK_c_730_n 0.0282361f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.53
cc_44 VNB N_CLK_c_731_n 0.0152659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_CLK_c_732_n 4.78612e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1012_47#_c_798_n 0.00361747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1012_47#_c_799_n 0.00459884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1012_47#_c_800_n 0.00424431f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_49 VNB N_A_1012_47#_c_801_n 0.00205783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1012_47#_c_802_n 9.07783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1012_47#_c_803_n 0.0227875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1012_47#_c_804_n 0.019243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VPWR_c_856_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_27_47#_c_948_n 0.0141546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_27_47#_c_949_n 0.00553702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_27_47#_c_950_n 0.0102032f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_57 VNB N_A_27_47#_c_951_n 0.00399709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_GCLK_c_1004_n 0.00545527f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_59 VNB N_GCLK_c_1005_n 0.0221381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_GCLK_c_1006_n 0.016761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1021_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_62 VNB N_VGND_c_1022_n 0.00566341f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_63 VNB N_VGND_c_1023_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1024_n 0.0142589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1025_n 0.0433008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1026_n 0.0278025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1027_n 0.0156121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1028_n 0.34215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1029_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1030_n 0.00663229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1031_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1032_n 0.027081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1033_n 0.0157552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VPB N_SCE_M1010_g 0.0419269f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_75 VPB SCE 0.0188038f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_76 VPB N_SCE_c_138_n 0.0111553f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_77 VPB N_GATE_M1005_g 0.0361864f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_78 VPB GATE 0.00752588f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_79 VPB N_GATE_c_167_n 0.00591646f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_80 VPB N_A_256_147#_M1007_g 0.0211245f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_81 VPB N_A_256_147#_c_210_n 0.00334009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_256_147#_c_218_n 0.00519656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_256_147#_c_215_n 0.00658814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_256_147#_c_220_n 0.0169889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_256_147#_c_221_n 0.00400932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_256_147#_c_222_n 7.50236e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_256_147#_c_223_n 0.0266048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_256_147#_c_224_n 0.0455041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_256_243#_M1021_g 0.0504347f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_90 VPB N_A_256_243#_c_377_n 0.0163673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_256_243#_c_378_n 0.00221325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_256_243#_c_381_n 0.0046398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_256_243#_c_393_n 0.00292655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_464_315#_M1017_g 0.022326f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_95 VPB N_A_464_315#_M1018_g 0.0170562f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_96 VPB N_A_464_315#_M1002_g 0.00537539f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_97 VPB N_A_464_315#_M1016_g 0.0229485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_464_315#_c_499_n 0.0033307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_464_315#_c_494_n 0.00397244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_464_315#_c_501_n 0.0151177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_464_315#_c_502_n 0.00526649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_464_315#_c_503_n 0.0310341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_464_315#_c_504_n 0.00417089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_464_315#_c_505_n 0.0297319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_286_413#_M1001_g 0.0243607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_286_413#_c_630_n 0.0134653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_286_413#_c_626_n 0.00269176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_286_413#_c_627_n 0.00386605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_286_413#_c_628_n 0.0083407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_CLK_M1012_g 0.0363646f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_111 VPB N_CLK_c_731_n 0.00852177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_CLK_c_735_n 0.0475815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_CLK_c_732_n 2.27341e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_1012_47#_M1009_g 0.0227544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_1012_47#_c_801_n 0.00858661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_1012_47#_c_803_n 0.00478448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_857_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_858_n 0.0319263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_859_n 0.00225253f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.53
cc_120 VPB N_VPWR_c_860_n 0.0131233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_861_n 0.01418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_862_n 0.0332005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_863_n 0.0135884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_864_n 0.015618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_856_n 0.0452937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_866_n 0.0488492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_867_n 0.0138042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_868_n 0.00455555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_869_n 0.00521963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_952_n 5.07672e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_131 VPB N_A_27_47#_c_951_n 9.33202e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_954_n 0.00214923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_GCLK_c_1007_n 0.00545527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_GCLK_c_1005_n 0.00890457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB GCLK 0.032128f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_136 N_SCE_M1010_g N_GATE_M1005_g 0.0494929f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_137 N_SCE_M1020_g N_GATE_M1008_g 0.0256158f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_138 N_SCE_M1020_g GATE 3.1151e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_139 N_SCE_M1010_g GATE 4.94095e-19 $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_140 N_SCE_c_138_n N_GATE_c_167_n 0.0494929f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_141 N_SCE_M1010_g N_VPWR_c_858_n 0.00473096f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_142 SCE N_VPWR_c_858_n 0.0237825f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_143 N_SCE_c_138_n N_VPWR_c_858_n 0.00105941f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_144 N_SCE_M1010_g N_VPWR_c_856_n 0.0112477f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_145 N_SCE_M1010_g N_VPWR_c_866_n 0.00577794f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_146 N_SCE_M1010_g N_A_27_47#_c_952_n 0.00815687f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_147 N_SCE_M1020_g N_A_27_47#_c_950_n 0.0157772f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_148 SCE N_A_27_47#_c_950_n 0.0214425f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_149 N_SCE_c_138_n N_A_27_47#_c_950_n 0.00349016f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_150 N_SCE_M1010_g N_A_27_47#_c_959_n 0.00646992f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_151 N_SCE_M1020_g N_A_27_47#_c_951_n 0.00897123f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_152 N_SCE_M1010_g N_A_27_47#_c_951_n 0.00221953f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_153 SCE N_A_27_47#_c_951_n 0.0512439f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_154 N_SCE_c_138_n N_A_27_47#_c_951_n 0.00730885f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_155 N_SCE_M1010_g N_A_27_47#_c_954_n 0.00938762f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_156 N_SCE_M1020_g N_VGND_c_1021_n 0.00809304f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_157 N_SCE_M1020_g N_VGND_c_1024_n 0.00337001f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_158 N_SCE_M1020_g N_VGND_c_1028_n 0.00485988f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_159 N_GATE_M1008_g N_A_256_147#_M1019_g 0.00956705f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_160 N_GATE_M1008_g N_A_256_147#_c_208_n 9.85224e-19 $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_161 GATE N_A_256_147#_c_208_n 0.030663f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_162 N_GATE_c_167_n N_A_256_147#_c_208_n 0.00116492f $X=0.935 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_GATE_M1008_g N_A_256_147#_c_209_n 0.00976894f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_164 GATE N_A_256_147#_c_209_n 3.958e-19 $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_165 N_GATE_c_167_n N_A_256_147#_c_209_n 6.18775e-19 $X=0.935 $Y=1.16 $X2=0
+ $Y2=0
cc_166 GATE N_A_256_147#_c_232_n 0.00153887f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_167 N_GATE_M1005_g N_A_256_147#_c_221_n 4.35899e-19 $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_168 GATE N_A_256_147#_c_221_n 0.0482195f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_169 GATE N_A_256_243#_M1021_g 0.0045356f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_170 N_GATE_M1005_g N_A_256_243#_c_378_n 0.0263234f $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_171 GATE N_A_256_243#_c_378_n 0.00193079f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_172 N_GATE_c_167_n N_A_256_243#_c_378_n 0.00718876f $X=0.935 $Y=1.16 $X2=0
+ $Y2=0
cc_173 N_GATE_M1005_g N_VPWR_c_856_n 0.00535424f $X=0.83 $Y=2.165 $X2=0 $Y2=0
cc_174 N_GATE_M1005_g N_VPWR_c_866_n 0.00357877f $X=0.83 $Y=2.165 $X2=0 $Y2=0
cc_175 GATE N_A_27_47#_M1005_d 0.00337146f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_176 N_GATE_M1008_g N_A_27_47#_c_949_n 0.0121516f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_177 GATE N_A_27_47#_c_949_n 0.0289312f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_178 N_GATE_c_167_n N_A_27_47#_c_949_n 0.00307889f $X=0.935 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_GATE_M1005_g N_A_27_47#_c_969_n 0.0153806f $X=0.83 $Y=2.165 $X2=0 $Y2=0
cc_180 GATE N_A_27_47#_c_969_n 0.0238941f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_181 N_GATE_M1008_g N_A_27_47#_c_951_n 0.0038793f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_182 GATE N_A_27_47#_c_951_n 0.0368851f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_183 N_GATE_c_167_n N_A_27_47#_c_951_n 0.00292348f $X=0.935 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_GATE_M1005_g N_A_27_47#_c_954_n 0.00332185f $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_185 GATE N_A_27_47#_c_954_n 0.0336367f $X=1.065 $Y=1.785 $X2=0 $Y2=0
cc_186 N_GATE_M1008_g N_VGND_c_1021_n 0.00763107f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_187 N_GATE_M1008_g N_VGND_c_1025_n 0.00337001f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_188 N_GATE_M1008_g N_VGND_c_1028_n 0.00407348f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_256_147#_M1007_g N_A_256_243#_M1021_g 0.0138034f $X=1.835 $Y=2.275
+ $X2=0 $Y2=0
cc_190 N_A_256_147#_c_221_n N_A_256_243#_M1021_g 0.0149056f $X=1.61 $Y=1.53
+ $X2=0 $Y2=0
cc_191 N_A_256_147#_c_223_n N_A_256_243#_M1021_g 0.021304f $X=1.775 $Y=1.74
+ $X2=0 $Y2=0
cc_192 N_A_256_147#_c_214_n N_A_256_243#_c_377_n 0.0105586f $X=1.61 $Y=1.325
+ $X2=0 $Y2=0
cc_193 N_A_256_147#_c_220_n N_A_256_243#_c_377_n 0.00213361f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_194 N_A_256_147#_c_221_n N_A_256_243#_c_377_n 0.00868281f $X=1.61 $Y=1.53
+ $X2=0 $Y2=0
cc_195 N_A_256_147#_c_223_n N_A_256_243#_c_377_n 0.0180583f $X=1.775 $Y=1.74
+ $X2=0 $Y2=0
cc_196 N_A_256_147#_c_209_n N_A_256_243#_c_378_n 0.0227923f $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_197 N_A_256_147#_c_214_n N_A_256_243#_c_378_n 0.00433366f $X=1.61 $Y=1.325
+ $X2=0 $Y2=0
cc_198 N_A_256_147#_c_221_n N_A_256_243#_c_378_n 4.44282e-19 $X=1.61 $Y=1.53
+ $X2=0 $Y2=0
cc_199 N_A_256_147#_c_214_n N_A_256_243#_c_379_n 0.00150324f $X=1.61 $Y=1.325
+ $X2=0 $Y2=0
cc_200 N_A_256_147#_M1011_g N_A_256_243#_c_380_n 0.00282429f $X=4.035 $Y=0.445
+ $X2=0 $Y2=0
cc_201 N_A_256_147#_c_212_n N_A_256_243#_c_380_n 0.00771195f $X=4.705 $Y=0.615
+ $X2=0 $Y2=0
cc_202 N_A_256_147#_M1011_g N_A_256_243#_c_381_n 0.00236246f $X=4.035 $Y=0.445
+ $X2=0 $Y2=0
cc_203 N_A_256_147#_c_210_n N_A_256_243#_c_381_n 0.0101973f $X=4.312 $Y=1.495
+ $X2=0 $Y2=0
cc_204 N_A_256_147#_c_211_n N_A_256_243#_c_381_n 0.0193569f $X=4.32 $Y=1.105
+ $X2=0 $Y2=0
cc_205 N_A_256_147#_c_215_n N_A_256_243#_c_381_n 0.00376938f $X=4.085 $Y=1.19
+ $X2=0 $Y2=0
cc_206 N_A_256_147#_c_220_n N_A_256_243#_c_381_n 0.0103533f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_207 N_A_256_147#_c_222_n N_A_256_243#_c_381_n 2.68226e-19 $X=4.38 $Y=1.53
+ $X2=0 $Y2=0
cc_208 N_A_256_147#_c_224_n N_A_256_243#_c_381_n 0.00385034f $X=4.085 $Y=1.325
+ $X2=0 $Y2=0
cc_209 N_A_256_147#_c_210_n N_A_256_243#_c_393_n 0.00660951f $X=4.312 $Y=1.495
+ $X2=0 $Y2=0
cc_210 N_A_256_147#_c_211_n N_A_256_243#_c_393_n 0.00185537f $X=4.32 $Y=1.105
+ $X2=0 $Y2=0
cc_211 N_A_256_147#_c_215_n N_A_256_243#_c_393_n 7.57315e-19 $X=4.085 $Y=1.19
+ $X2=0 $Y2=0
cc_212 N_A_256_147#_c_220_n N_A_256_243#_c_393_n 0.00987276f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_213 N_A_256_147#_c_222_n N_A_256_243#_c_393_n 2.78941e-19 $X=4.38 $Y=1.53
+ $X2=0 $Y2=0
cc_214 N_A_256_147#_c_224_n N_A_256_243#_c_393_n 0.00246207f $X=4.085 $Y=1.325
+ $X2=0 $Y2=0
cc_215 N_A_256_147#_c_220_n N_A_256_243#_c_382_n 0.0689878f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_216 N_A_256_147#_c_208_n N_A_256_243#_c_383_n 0.00155066f $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_217 N_A_256_147#_c_220_n N_A_256_243#_c_383_n 0.0132091f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_218 N_A_256_147#_M1011_g N_A_256_243#_c_384_n 0.00504445f $X=4.035 $Y=0.445
+ $X2=0 $Y2=0
cc_219 N_A_256_147#_c_211_n N_A_256_243#_c_384_n 0.00817201f $X=4.32 $Y=1.105
+ $X2=0 $Y2=0
cc_220 N_A_256_147#_c_212_n N_A_256_243#_c_384_n 0.00144026f $X=4.705 $Y=0.615
+ $X2=0 $Y2=0
cc_221 N_A_256_147#_c_215_n N_A_256_243#_c_384_n 7.14969e-19 $X=4.085 $Y=1.19
+ $X2=0 $Y2=0
cc_222 N_A_256_147#_c_220_n N_A_256_243#_c_384_n 0.0150763f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_223 N_A_256_147#_M1011_g N_A_256_243#_c_385_n 0.00636449f $X=4.035 $Y=0.445
+ $X2=0 $Y2=0
cc_224 N_A_256_147#_c_211_n N_A_256_243#_c_385_n 0.0148946f $X=4.32 $Y=1.105
+ $X2=0 $Y2=0
cc_225 N_A_256_147#_c_212_n N_A_256_243#_c_385_n 0.00132326f $X=4.705 $Y=0.615
+ $X2=0 $Y2=0
cc_226 N_A_256_147#_c_215_n N_A_256_243#_c_385_n 8.95761e-19 $X=4.085 $Y=1.19
+ $X2=0 $Y2=0
cc_227 N_A_256_147#_c_220_n N_A_256_243#_c_385_n 9.85771e-19 $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_228 N_A_256_147#_c_208_n N_A_256_243#_c_386_n 0.00708004f $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_229 N_A_256_147#_c_209_n N_A_256_243#_c_386_n 0.0165261f $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_230 N_A_256_147#_c_220_n N_A_256_243#_c_386_n 8.52878e-19 $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_231 N_A_256_147#_c_208_n N_A_256_243#_c_387_n 0.0242697f $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_232 N_A_256_147#_c_209_n N_A_256_243#_c_387_n 2.60953e-19 $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_233 N_A_256_147#_c_220_n N_A_256_243#_c_387_n 0.00446365f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_234 N_A_256_147#_M1019_g N_A_256_243#_c_388_n 0.0107241f $X=1.37 $Y=0.415
+ $X2=0 $Y2=0
cc_235 N_A_256_147#_c_220_n N_A_464_315#_M1001_d 2.81924e-19 $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_236 N_A_256_147#_M1007_g N_A_464_315#_M1017_g 0.0155568f $X=1.835 $Y=2.275
+ $X2=0 $Y2=0
cc_237 N_A_256_147#_c_220_n N_A_464_315#_M1018_g 0.00428067f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_238 N_A_256_147#_c_212_n N_A_464_315#_M1002_g 4.14369e-19 $X=4.705 $Y=0.615
+ $X2=0 $Y2=0
cc_239 N_A_256_147#_c_220_n N_A_464_315#_c_499_n 0.0228159f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_240 N_A_256_147#_M1011_g N_A_464_315#_c_494_n 4.90665e-19 $X=4.035 $Y=0.445
+ $X2=0 $Y2=0
cc_241 N_A_256_147#_c_220_n N_A_464_315#_c_494_n 0.027217f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_242 N_A_256_147#_c_224_n N_A_464_315#_c_513_n 0.00469714f $X=4.085 $Y=1.325
+ $X2=0 $Y2=0
cc_243 N_A_256_147#_M1006_d N_A_464_315#_c_501_n 0.00479771f $X=4.66 $Y=1.515
+ $X2=0 $Y2=0
cc_244 N_A_256_147#_c_210_n N_A_464_315#_c_501_n 0.0210881f $X=4.312 $Y=1.495
+ $X2=0 $Y2=0
cc_245 N_A_256_147#_c_211_n N_A_464_315#_c_501_n 0.00128309f $X=4.32 $Y=1.105
+ $X2=0 $Y2=0
cc_246 N_A_256_147#_c_218_n N_A_464_315#_c_501_n 0.0286514f $X=4.795 $Y=1.66
+ $X2=0 $Y2=0
cc_247 N_A_256_147#_c_215_n N_A_464_315#_c_501_n 2.59847e-19 $X=4.085 $Y=1.19
+ $X2=0 $Y2=0
cc_248 N_A_256_147#_c_220_n N_A_464_315#_c_501_n 0.0136002f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_249 N_A_256_147#_c_222_n N_A_464_315#_c_501_n 0.00169866f $X=4.38 $Y=1.53
+ $X2=0 $Y2=0
cc_250 N_A_256_147#_c_224_n N_A_464_315#_c_501_n 0.0145602f $X=4.085 $Y=1.325
+ $X2=0 $Y2=0
cc_251 N_A_256_147#_c_218_n N_A_464_315#_c_502_n 0.0116692f $X=4.795 $Y=1.66
+ $X2=0 $Y2=0
cc_252 N_A_256_147#_c_220_n N_A_464_315#_c_503_n 0.0039188f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_253 N_A_256_147#_c_223_n N_A_464_315#_c_503_n 0.00753208f $X=1.775 $Y=1.74
+ $X2=0 $Y2=0
cc_254 N_A_256_147#_c_220_n N_A_464_315#_c_525_n 0.00517255f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_255 N_A_256_147#_c_224_n N_A_464_315#_c_526_n 0.00339261f $X=4.085 $Y=1.325
+ $X2=0 $Y2=0
cc_256 N_A_256_147#_c_210_n N_A_464_315#_c_504_n 9.55812e-19 $X=4.312 $Y=1.495
+ $X2=0 $Y2=0
cc_257 N_A_256_147#_c_218_n N_A_464_315#_c_504_n 0.00920802f $X=4.795 $Y=1.66
+ $X2=0 $Y2=0
cc_258 N_A_256_147#_c_222_n N_A_464_315#_c_504_n 0.00163332f $X=4.38 $Y=1.53
+ $X2=0 $Y2=0
cc_259 N_A_256_147#_c_218_n N_A_464_315#_c_505_n 5.57199e-19 $X=4.795 $Y=1.66
+ $X2=0 $Y2=0
cc_260 N_A_256_147#_c_220_n N_A_286_413#_M1001_g 0.0074801f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_261 N_A_256_147#_M1019_g N_A_286_413#_c_635_n 0.00581223f $X=1.37 $Y=0.415
+ $X2=0 $Y2=0
cc_262 N_A_256_147#_c_208_n N_A_286_413#_c_635_n 0.0249382f $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_263 N_A_256_147#_c_209_n N_A_286_413#_c_635_n 9.8177e-19 $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_264 N_A_256_147#_c_214_n N_A_286_413#_c_635_n 0.00398233f $X=1.61 $Y=1.325
+ $X2=0 $Y2=0
cc_265 N_A_256_147#_M1007_g N_A_286_413#_c_639_n 0.0131252f $X=1.835 $Y=2.275
+ $X2=0 $Y2=0
cc_266 N_A_256_147#_c_220_n N_A_286_413#_c_639_n 0.00594058f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_267 N_A_256_147#_c_232_n N_A_286_413#_c_639_n 0.00121651f $X=1.755 $Y=1.53
+ $X2=0 $Y2=0
cc_268 N_A_256_147#_c_221_n N_A_286_413#_c_639_n 0.0302261f $X=1.61 $Y=1.53
+ $X2=0 $Y2=0
cc_269 N_A_256_147#_c_223_n N_A_286_413#_c_639_n 6.45937e-19 $X=1.775 $Y=1.74
+ $X2=0 $Y2=0
cc_270 N_A_256_147#_c_220_n N_A_286_413#_c_630_n 0.0205826f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_271 N_A_256_147#_c_232_n N_A_286_413#_c_630_n 5.20192e-19 $X=1.755 $Y=1.53
+ $X2=0 $Y2=0
cc_272 N_A_256_147#_c_221_n N_A_286_413#_c_630_n 0.0436285f $X=1.61 $Y=1.53
+ $X2=0 $Y2=0
cc_273 N_A_256_147#_c_223_n N_A_286_413#_c_630_n 0.00709868f $X=1.775 $Y=1.74
+ $X2=0 $Y2=0
cc_274 N_A_256_147#_c_208_n N_A_286_413#_c_626_n 0.00602675f $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_275 N_A_256_147#_c_214_n N_A_286_413#_c_626_n 0.0146898f $X=1.61 $Y=1.325
+ $X2=0 $Y2=0
cc_276 N_A_256_147#_c_220_n N_A_286_413#_c_626_n 0.00783084f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_277 N_A_256_147#_c_220_n N_A_286_413#_c_627_n 0.00746407f $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_278 N_A_256_147#_c_220_n N_A_286_413#_c_628_n 3.93021e-19 $X=4.235 $Y=1.53
+ $X2=0 $Y2=0
cc_279 N_A_256_147#_M1011_g N_CLK_c_724_n 0.00386856f $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_280 N_A_256_147#_c_211_n N_CLK_c_724_n 0.00562288f $X=4.32 $Y=1.105 $X2=0
+ $Y2=0
cc_281 N_A_256_147#_c_215_n N_CLK_c_724_n 0.012847f $X=4.085 $Y=1.19 $X2=0 $Y2=0
cc_282 N_A_256_147#_M1011_g N_CLK_c_727_n 0.0199171f $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_283 N_A_256_147#_c_212_n N_CLK_c_727_n 0.00705718f $X=4.705 $Y=0.615 $X2=0
+ $Y2=0
cc_284 N_A_256_147#_c_211_n N_CLK_c_728_n 0.00792429f $X=4.32 $Y=1.105 $X2=0
+ $Y2=0
cc_285 N_A_256_147#_c_218_n N_CLK_c_728_n 9.73222e-19 $X=4.795 $Y=1.66 $X2=0
+ $Y2=0
cc_286 N_A_256_147#_c_212_n N_CLK_c_728_n 0.0204503f $X=4.705 $Y=0.615 $X2=0
+ $Y2=0
cc_287 N_A_256_147#_c_213_n N_CLK_c_728_n 0.00148768f $X=4.665 $Y=0.465 $X2=0
+ $Y2=0
cc_288 N_A_256_147#_c_222_n N_CLK_c_728_n 0.00109922f $X=4.38 $Y=1.53 $X2=0
+ $Y2=0
cc_289 N_A_256_147#_c_218_n N_CLK_c_729_n 0.00193807f $X=4.795 $Y=1.66 $X2=0
+ $Y2=0
cc_290 N_A_256_147#_c_210_n N_CLK_c_731_n 0.00433288f $X=4.312 $Y=1.495 $X2=0
+ $Y2=0
cc_291 N_A_256_147#_c_218_n N_CLK_c_731_n 0.00772226f $X=4.795 $Y=1.66 $X2=0
+ $Y2=0
cc_292 N_A_256_147#_c_218_n N_CLK_c_735_n 0.0158328f $X=4.795 $Y=1.66 $X2=0
+ $Y2=0
cc_293 N_A_256_147#_c_222_n N_CLK_c_735_n 0.00279615f $X=4.38 $Y=1.53 $X2=0
+ $Y2=0
cc_294 N_A_256_147#_c_224_n N_CLK_c_735_n 0.0381082f $X=4.085 $Y=1.325 $X2=0
+ $Y2=0
cc_295 N_A_256_147#_c_210_n N_CLK_c_732_n 0.00286067f $X=4.312 $Y=1.495 $X2=0
+ $Y2=0
cc_296 N_A_256_147#_c_211_n N_CLK_c_732_n 0.0204944f $X=4.32 $Y=1.105 $X2=0
+ $Y2=0
cc_297 N_A_256_147#_c_218_n N_CLK_c_732_n 0.0171796f $X=4.795 $Y=1.66 $X2=0
+ $Y2=0
cc_298 N_A_256_147#_c_212_n N_CLK_c_732_n 0.00864905f $X=4.705 $Y=0.615 $X2=0
+ $Y2=0
cc_299 N_A_256_147#_c_213_n N_A_1012_47#_c_798_n 0.0276513f $X=4.665 $Y=0.465
+ $X2=0 $Y2=0
cc_300 N_A_256_147#_c_212_n N_A_1012_47#_c_800_n 0.0148221f $X=4.705 $Y=0.615
+ $X2=0 $Y2=0
cc_301 N_A_256_147#_c_220_n N_VPWR_M1017_d 0.0020643f $X=4.235 $Y=1.53 $X2=0
+ $Y2=0
cc_302 N_A_256_147#_c_210_n N_VPWR_M1015_d 0.00511429f $X=4.312 $Y=1.495 $X2=0
+ $Y2=0
cc_303 N_A_256_147#_c_220_n N_VPWR_M1015_d 4.60476e-19 $X=4.235 $Y=1.53 $X2=0
+ $Y2=0
cc_304 N_A_256_147#_c_224_n N_VPWR_c_862_n 0.0230773f $X=4.085 $Y=1.325 $X2=0
+ $Y2=0
cc_305 N_A_256_147#_M1007_g N_VPWR_c_856_n 0.00579685f $X=1.835 $Y=2.275 $X2=0
+ $Y2=0
cc_306 N_A_256_147#_c_221_n N_VPWR_c_856_n 0.00150144f $X=1.61 $Y=1.53 $X2=0
+ $Y2=0
cc_307 N_A_256_147#_M1007_g N_VPWR_c_866_n 0.00357877f $X=1.835 $Y=2.275 $X2=0
+ $Y2=0
cc_308 N_A_256_147#_M1007_g N_VPWR_c_867_n 0.00145256f $X=1.835 $Y=2.275 $X2=0
+ $Y2=0
cc_309 N_A_256_147#_c_220_n N_VPWR_c_867_n 7.31718e-19 $X=4.235 $Y=1.53 $X2=0
+ $Y2=0
cc_310 N_A_256_147#_M1019_g N_A_27_47#_c_949_n 0.00296433f $X=1.37 $Y=0.415
+ $X2=0 $Y2=0
cc_311 N_A_256_147#_c_208_n N_A_27_47#_c_949_n 0.0067219f $X=1.445 $Y=0.87 $X2=0
+ $Y2=0
cc_312 N_A_256_147#_c_209_n N_A_27_47#_c_949_n 4.39845e-19 $X=1.445 $Y=0.87
+ $X2=0 $Y2=0
cc_313 N_A_256_147#_M1019_g N_A_27_47#_c_979_n 0.00230184f $X=1.37 $Y=0.415
+ $X2=0 $Y2=0
cc_314 N_A_256_147#_c_212_n N_VGND_M1011_d 0.00192931f $X=4.705 $Y=0.615 $X2=0
+ $Y2=0
cc_315 N_A_256_147#_M1019_g N_VGND_c_1021_n 0.0010609f $X=1.37 $Y=0.415 $X2=0
+ $Y2=0
cc_316 N_A_256_147#_M1011_g N_VGND_c_1023_n 0.00853729f $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_317 N_A_256_147#_c_211_n N_VGND_c_1023_n 0.00151747f $X=4.32 $Y=1.105 $X2=0
+ $Y2=0
cc_318 N_A_256_147#_c_212_n N_VGND_c_1023_n 0.0132365f $X=4.705 $Y=0.615 $X2=0
+ $Y2=0
cc_319 N_A_256_147#_c_215_n N_VGND_c_1023_n 8.45001e-19 $X=4.085 $Y=1.19 $X2=0
+ $Y2=0
cc_320 N_A_256_147#_M1019_g N_VGND_c_1025_n 0.00456464f $X=1.37 $Y=0.415 $X2=0
+ $Y2=0
cc_321 N_A_256_147#_c_209_n N_VGND_c_1025_n 2.64403e-19 $X=1.445 $Y=0.87 $X2=0
+ $Y2=0
cc_322 N_A_256_147#_M1011_g N_VGND_c_1026_n 0.0046653f $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_323 N_A_256_147#_M1014_d N_VGND_c_1028_n 0.00227267f $X=4.53 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_A_256_147#_M1019_g N_VGND_c_1028_n 0.0079756f $X=1.37 $Y=0.415 $X2=0
+ $Y2=0
cc_325 N_A_256_147#_M1011_g N_VGND_c_1028_n 0.0060162f $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_326 N_A_256_147#_c_209_n N_VGND_c_1028_n 3.36535e-19 $X=1.445 $Y=0.87 $X2=0
+ $Y2=0
cc_327 N_A_256_147#_c_212_n N_VGND_c_1028_n 0.00544468f $X=4.705 $Y=0.615 $X2=0
+ $Y2=0
cc_328 N_A_256_147#_c_213_n N_VGND_c_1028_n 0.00940011f $X=4.665 $Y=0.465 $X2=0
+ $Y2=0
cc_329 N_A_256_147#_c_212_n N_VGND_c_1032_n 0.00258611f $X=4.705 $Y=0.615 $X2=0
+ $Y2=0
cc_330 N_A_256_147#_c_213_n N_VGND_c_1032_n 0.0165187f $X=4.665 $Y=0.465 $X2=0
+ $Y2=0
cc_331 N_A_256_243#_c_382_n N_A_464_315#_M1003_d 5.67759e-19 $X=3.775 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_332 N_A_256_243#_c_379_n N_A_464_315#_M1018_g 0.00692236f $X=1.895 $Y=1.215
+ $X2=0 $Y2=0
cc_333 N_A_256_243#_c_382_n N_A_464_315#_M1018_g 0.00340334f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_334 N_A_256_243#_c_386_n N_A_464_315#_M1018_g 0.0115616f $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_335 N_A_256_243#_c_387_n N_A_464_315#_M1018_g 7.79891e-19 $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_336 N_A_256_243#_c_388_n N_A_464_315#_M1018_g 0.0139526f $X=1.955 $Y=0.705
+ $X2=0 $Y2=0
cc_337 N_A_256_243#_c_380_n N_A_464_315#_c_494_n 0.0964478f $X=3.825 $Y=0.465
+ $X2=0 $Y2=0
cc_338 N_A_256_243#_c_393_n N_A_464_315#_c_494_n 0.00430195f $X=3.825 $Y=1.66
+ $X2=0 $Y2=0
cc_339 N_A_256_243#_c_382_n N_A_464_315#_c_494_n 0.0209151f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_340 N_A_256_243#_c_384_n N_A_464_315#_c_494_n 2.93344e-19 $X=3.92 $Y=0.85
+ $X2=0 $Y2=0
cc_341 N_A_256_243#_M1015_s N_A_464_315#_c_501_n 0.00457358f $X=3.7 $Y=1.515
+ $X2=0 $Y2=0
cc_342 N_A_256_243#_c_393_n N_A_464_315#_c_501_n 0.0240592f $X=3.825 $Y=1.66
+ $X2=0 $Y2=0
cc_343 N_A_256_243#_c_393_n N_A_464_315#_c_526_n 0.00924997f $X=3.825 $Y=1.66
+ $X2=0 $Y2=0
cc_344 N_A_256_243#_c_382_n N_A_286_413#_c_624_n 0.00842195f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_345 N_A_256_243#_c_393_n N_A_286_413#_M1001_g 4.99393e-19 $X=3.825 $Y=1.66
+ $X2=0 $Y2=0
cc_346 N_A_256_243#_c_377_n N_A_286_413#_c_635_n 7.07243e-19 $X=1.82 $Y=1.29
+ $X2=0 $Y2=0
cc_347 N_A_256_243#_c_382_n N_A_286_413#_c_635_n 0.00173863f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_348 N_A_256_243#_c_383_n N_A_286_413#_c_635_n 0.0020338f $X=2.215 $Y=0.85
+ $X2=0 $Y2=0
cc_349 N_A_256_243#_c_386_n N_A_286_413#_c_635_n 0.00258224f $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_350 N_A_256_243#_c_387_n N_A_286_413#_c_635_n 0.0175669f $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_351 N_A_256_243#_c_388_n N_A_286_413#_c_635_n 0.0128508f $X=1.955 $Y=0.705
+ $X2=0 $Y2=0
cc_352 N_A_256_243#_M1021_g N_A_286_413#_c_639_n 0.00300731f $X=1.355 $Y=2.275
+ $X2=0 $Y2=0
cc_353 N_A_256_243#_M1021_g N_A_286_413#_c_630_n 6.3244e-19 $X=1.355 $Y=2.275
+ $X2=0 $Y2=0
cc_354 N_A_256_243#_c_382_n N_A_286_413#_c_625_n 0.0162752f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_355 N_A_256_243#_c_383_n N_A_286_413#_c_625_n 0.00275249f $X=2.215 $Y=0.85
+ $X2=0 $Y2=0
cc_356 N_A_256_243#_c_386_n N_A_286_413#_c_625_n 7.44567e-19 $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_357 N_A_256_243#_c_387_n N_A_286_413#_c_625_n 0.0205672f $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_358 N_A_256_243#_c_388_n N_A_286_413#_c_625_n 0.00302624f $X=1.955 $Y=0.705
+ $X2=0 $Y2=0
cc_359 N_A_256_243#_c_379_n N_A_286_413#_c_626_n 0.00377955f $X=1.895 $Y=1.215
+ $X2=0 $Y2=0
cc_360 N_A_256_243#_c_382_n N_A_286_413#_c_626_n 0.00154998f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_361 N_A_256_243#_c_383_n N_A_286_413#_c_626_n 0.00160742f $X=2.215 $Y=0.85
+ $X2=0 $Y2=0
cc_362 N_A_256_243#_c_386_n N_A_286_413#_c_626_n 0.00153556f $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_363 N_A_256_243#_c_387_n N_A_286_413#_c_626_n 0.0128543f $X=1.955 $Y=0.87
+ $X2=0 $Y2=0
cc_364 N_A_256_243#_c_382_n N_A_286_413#_c_627_n 0.0106635f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_365 N_A_256_243#_c_382_n N_A_286_413#_c_628_n 0.00450205f $X=3.775 $Y=0.85
+ $X2=0 $Y2=0
cc_366 N_A_256_243#_M1021_g N_VPWR_c_856_n 0.0103224f $X=1.355 $Y=2.275 $X2=0
+ $Y2=0
cc_367 N_A_256_243#_M1021_g N_VPWR_c_866_n 0.00577801f $X=1.355 $Y=2.275 $X2=0
+ $Y2=0
cc_368 N_A_256_243#_c_382_n N_VGND_M1018_d 2.83879e-19 $X=3.775 $Y=0.85 $X2=0
+ $Y2=0
cc_369 N_A_256_243#_c_382_n N_VGND_c_1022_n 0.0140539f $X=3.775 $Y=0.85 $X2=0
+ $Y2=0
cc_370 N_A_256_243#_c_388_n N_VGND_c_1025_n 0.00357877f $X=1.955 $Y=0.705 $X2=0
+ $Y2=0
cc_371 N_A_256_243#_c_380_n N_VGND_c_1026_n 0.0230197f $X=3.825 $Y=0.465 $X2=0
+ $Y2=0
cc_372 N_A_256_243#_M1011_s N_VGND_c_1028_n 0.0018314f $X=3.7 $Y=0.235 $X2=0
+ $Y2=0
cc_373 N_A_256_243#_c_380_n N_VGND_c_1028_n 0.00590194f $X=3.825 $Y=0.465 $X2=0
+ $Y2=0
cc_374 N_A_256_243#_c_382_n N_VGND_c_1028_n 0.0729689f $X=3.775 $Y=0.85 $X2=0
+ $Y2=0
cc_375 N_A_256_243#_c_383_n N_VGND_c_1028_n 0.014828f $X=2.215 $Y=0.85 $X2=0
+ $Y2=0
cc_376 N_A_256_243#_c_384_n N_VGND_c_1028_n 0.0153387f $X=3.92 $Y=0.85 $X2=0
+ $Y2=0
cc_377 N_A_256_243#_c_385_n N_VGND_c_1028_n 8.78282e-19 $X=3.92 $Y=0.85 $X2=0
+ $Y2=0
cc_378 N_A_256_243#_c_388_n N_VGND_c_1028_n 0.00589934f $X=1.955 $Y=0.705 $X2=0
+ $Y2=0
cc_379 N_A_464_315#_M1018_g N_A_286_413#_c_624_n 0.0194843f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_380 N_A_464_315#_c_494_n N_A_286_413#_c_624_n 0.0102198f $X=3.305 $Y=0.42
+ $X2=0 $Y2=0
cc_381 N_A_464_315#_M1017_g N_A_286_413#_M1001_g 0.0129074f $X=2.425 $Y=2.275
+ $X2=0 $Y2=0
cc_382 N_A_464_315#_M1018_g N_A_286_413#_M1001_g 0.00670688f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_383 N_A_464_315#_c_499_n N_A_286_413#_M1001_g 0.014088f $X=3.18 $Y=1.77 $X2=0
+ $Y2=0
cc_384 N_A_464_315#_c_503_n N_A_286_413#_M1001_g 0.00808806f $X=2.455 $Y=1.74
+ $X2=0 $Y2=0
cc_385 N_A_464_315#_c_525_n N_A_286_413#_M1001_g 2.06052e-19 $X=2.54 $Y=1.74
+ $X2=0 $Y2=0
cc_386 N_A_464_315#_c_526_n N_A_286_413#_M1001_g 0.0131723f $X=3.29 $Y=1.86
+ $X2=0 $Y2=0
cc_387 N_A_464_315#_M1018_g N_A_286_413#_c_635_n 0.00892805f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_388 N_A_464_315#_M1017_g N_A_286_413#_c_639_n 0.00282173f $X=2.425 $Y=2.275
+ $X2=0 $Y2=0
cc_389 N_A_464_315#_M1017_g N_A_286_413#_c_630_n 0.00426352f $X=2.425 $Y=2.275
+ $X2=0 $Y2=0
cc_390 N_A_464_315#_M1018_g N_A_286_413#_c_630_n 0.00550388f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_391 N_A_464_315#_c_503_n N_A_286_413#_c_630_n 0.00271662f $X=2.455 $Y=1.74
+ $X2=0 $Y2=0
cc_392 N_A_464_315#_c_525_n N_A_286_413#_c_630_n 0.0255746f $X=2.54 $Y=1.74
+ $X2=0 $Y2=0
cc_393 N_A_464_315#_M1018_g N_A_286_413#_c_625_n 0.0114266f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_394 N_A_464_315#_M1018_g N_A_286_413#_c_626_n 0.00791638f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_395 N_A_464_315#_c_503_n N_A_286_413#_c_626_n 0.00300149f $X=2.455 $Y=1.74
+ $X2=0 $Y2=0
cc_396 N_A_464_315#_c_525_n N_A_286_413#_c_626_n 0.00700208f $X=2.54 $Y=1.74
+ $X2=0 $Y2=0
cc_397 N_A_464_315#_M1018_g N_A_286_413#_c_627_n 0.00928658f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_398 N_A_464_315#_c_499_n N_A_286_413#_c_627_n 0.0171291f $X=3.18 $Y=1.77
+ $X2=0 $Y2=0
cc_399 N_A_464_315#_c_494_n N_A_286_413#_c_627_n 0.0310043f $X=3.305 $Y=0.42
+ $X2=0 $Y2=0
cc_400 N_A_464_315#_c_525_n N_A_286_413#_c_627_n 0.00230595f $X=2.54 $Y=1.74
+ $X2=0 $Y2=0
cc_401 N_A_464_315#_M1018_g N_A_286_413#_c_628_n 0.0213485f $X=2.505 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_464_315#_c_499_n N_A_286_413#_c_628_n 0.00123339f $X=3.18 $Y=1.77
+ $X2=0 $Y2=0
cc_403 N_A_464_315#_c_494_n N_A_286_413#_c_628_n 0.0189458f $X=3.305 $Y=0.42
+ $X2=0 $Y2=0
cc_404 N_A_464_315#_M1002_g N_CLK_M1004_g 0.0232879f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_405 N_A_464_315#_M1002_g N_CLK_M1012_g 0.00642463f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_406 N_A_464_315#_c_505_n N_CLK_M1012_g 0.0375236f $X=5.535 $Y=1.52 $X2=0
+ $Y2=0
cc_407 N_A_464_315#_M1002_g N_CLK_c_728_n 0.019113f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_408 N_A_464_315#_M1002_g N_CLK_c_729_n 0.016478f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_409 N_A_464_315#_c_501_n N_CLK_c_729_n 0.00555749f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_410 N_A_464_315#_c_504_n N_CLK_c_729_n 0.0352231f $X=5.445 $Y=1.52 $X2=0
+ $Y2=0
cc_411 N_A_464_315#_c_505_n N_CLK_c_729_n 0.00488951f $X=5.535 $Y=1.52 $X2=0
+ $Y2=0
cc_412 N_A_464_315#_M1002_g N_CLK_c_730_n 0.0176924f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_464_315#_M1002_g N_CLK_c_735_n 0.00135629f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_414 N_A_464_315#_c_501_n N_CLK_c_735_n 0.0130686f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_415 N_A_464_315#_c_502_n N_CLK_c_735_n 0.00317597f $X=5.295 $Y=1.915 $X2=0
+ $Y2=0
cc_416 N_A_464_315#_c_504_n N_CLK_c_735_n 7.48866e-19 $X=5.445 $Y=1.52 $X2=0
+ $Y2=0
cc_417 N_A_464_315#_c_505_n N_CLK_c_735_n 0.00324658f $X=5.535 $Y=1.52 $X2=0
+ $Y2=0
cc_418 N_A_464_315#_M1002_g N_CLK_c_732_n 3.43508e-19 $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_464_315#_M1002_g N_A_1012_47#_c_799_n 0.0125526f $X=5.395 $Y=0.445
+ $X2=0 $Y2=0
cc_420 N_A_464_315#_M1016_g N_A_1012_47#_c_801_n 9.63993e-19 $X=5.535 $Y=2.165
+ $X2=0 $Y2=0
cc_421 N_A_464_315#_c_502_n N_A_1012_47#_c_801_n 0.0143305f $X=5.295 $Y=1.915
+ $X2=0 $Y2=0
cc_422 N_A_464_315#_c_504_n N_A_1012_47#_c_801_n 0.0144034f $X=5.445 $Y=1.52
+ $X2=0 $Y2=0
cc_423 N_A_464_315#_c_505_n N_A_1012_47#_c_801_n 0.002146f $X=5.535 $Y=1.52
+ $X2=0 $Y2=0
cc_424 N_A_464_315#_c_499_n N_VPWR_M1017_d 0.00488989f $X=3.18 $Y=1.77 $X2=0
+ $Y2=0
cc_425 N_A_464_315#_c_501_n N_VPWR_M1015_d 0.00607953f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_426 N_A_464_315#_c_501_n N_VPWR_M1016_s 0.00399258f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_427 N_A_464_315#_c_502_n N_VPWR_M1016_s 7.75292e-19 $X=5.295 $Y=1.915 $X2=0
+ $Y2=0
cc_428 N_A_464_315#_c_513_n N_VPWR_c_860_n 0.0169548f $X=3.315 $Y=2.3 $X2=0
+ $Y2=0
cc_429 N_A_464_315#_c_501_n N_VPWR_c_860_n 0.110903f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_430 N_A_464_315#_c_513_n N_VPWR_c_861_n 0.0133789f $X=3.315 $Y=2.3 $X2=0
+ $Y2=0
cc_431 N_A_464_315#_c_501_n N_VPWR_c_861_n 0.00234498f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_432 N_A_464_315#_c_501_n N_VPWR_c_862_n 0.0216591f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_433 N_A_464_315#_M1016_g N_VPWR_c_863_n 0.0046653f $X=5.535 $Y=2.165 $X2=0
+ $Y2=0
cc_434 N_A_464_315#_M1001_d N_VPWR_c_856_n 0.00223109f $X=3.18 $Y=1.485 $X2=0
+ $Y2=0
cc_435 N_A_464_315#_M1017_g N_VPWR_c_856_n 0.002381f $X=2.425 $Y=2.275 $X2=0
+ $Y2=0
cc_436 N_A_464_315#_M1016_g N_VPWR_c_856_n 0.00794739f $X=5.535 $Y=2.165 $X2=0
+ $Y2=0
cc_437 N_A_464_315#_c_499_n N_VPWR_c_856_n 0.00506605f $X=3.18 $Y=1.77 $X2=0
+ $Y2=0
cc_438 N_A_464_315#_c_513_n N_VPWR_c_856_n 0.00839556f $X=3.315 $Y=2.3 $X2=0
+ $Y2=0
cc_439 N_A_464_315#_c_501_n N_VPWR_c_856_n 0.0140823f $X=5.14 $Y=2 $X2=0 $Y2=0
cc_440 N_A_464_315#_c_503_n N_VPWR_c_856_n 6.86139e-19 $X=2.455 $Y=1.74 $X2=0
+ $Y2=0
cc_441 N_A_464_315#_c_525_n N_VPWR_c_856_n 0.00214472f $X=2.54 $Y=1.74 $X2=0
+ $Y2=0
cc_442 N_A_464_315#_M1017_g N_VPWR_c_866_n 7.6274e-19 $X=2.425 $Y=2.275 $X2=0
+ $Y2=0
cc_443 N_A_464_315#_M1017_g N_VPWR_c_867_n 0.0247949f $X=2.425 $Y=2.275 $X2=0
+ $Y2=0
cc_444 N_A_464_315#_c_503_n N_VPWR_c_867_n 0.0022365f $X=2.455 $Y=1.74 $X2=0
+ $Y2=0
cc_445 N_A_464_315#_c_525_n N_VPWR_c_867_n 0.044273f $X=2.54 $Y=1.74 $X2=0 $Y2=0
cc_446 N_A_464_315#_M1016_g N_VPWR_c_868_n 0.00882421f $X=5.535 $Y=2.165 $X2=0
+ $Y2=0
cc_447 N_A_464_315#_c_504_n N_VPWR_c_868_n 8.53981e-19 $X=5.445 $Y=1.52 $X2=0
+ $Y2=0
cc_448 N_A_464_315#_c_505_n N_VPWR_c_868_n 4.82886e-19 $X=5.535 $Y=1.52 $X2=0
+ $Y2=0
cc_449 N_A_464_315#_M1018_g N_VGND_c_1022_n 0.00841619f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_450 N_A_464_315#_c_494_n N_VGND_c_1022_n 0.00161158f $X=3.305 $Y=0.42 $X2=0
+ $Y2=0
cc_451 N_A_464_315#_M1018_g N_VGND_c_1025_n 0.00486707f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_464_315#_c_494_n N_VGND_c_1026_n 0.0137273f $X=3.305 $Y=0.42 $X2=0
+ $Y2=0
cc_453 N_A_464_315#_M1003_d N_VGND_c_1028_n 0.00204319f $X=3.17 $Y=0.235 $X2=0
+ $Y2=0
cc_454 N_A_464_315#_M1018_g N_VGND_c_1028_n 0.00671579f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_455 N_A_464_315#_M1002_g N_VGND_c_1028_n 0.0073887f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_456 N_A_464_315#_c_494_n N_VGND_c_1028_n 0.00399922f $X=3.305 $Y=0.42 $X2=0
+ $Y2=0
cc_457 N_A_464_315#_M1002_g N_VGND_c_1032_n 0.00422112f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_464_315#_M1002_g N_VGND_c_1033_n 0.00469598f $X=5.395 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_A_286_413#_M1001_g N_VPWR_c_860_n 0.00214227f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_460 N_A_286_413#_M1001_g N_VPWR_c_861_n 0.00468308f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_461 N_A_286_413#_M1021_d N_VPWR_c_856_n 0.00263412f $X=1.43 $Y=2.065 $X2=0
+ $Y2=0
cc_462 N_A_286_413#_M1001_g N_VPWR_c_856_n 0.00796283f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_463 N_A_286_413#_c_639_n N_VPWR_c_856_n 0.0285676f $X=2.03 $Y=2.295 $X2=0
+ $Y2=0
cc_464 N_A_286_413#_c_639_n N_VPWR_c_866_n 0.0463617f $X=2.03 $Y=2.295 $X2=0
+ $Y2=0
cc_465 N_A_286_413#_M1001_g N_VPWR_c_867_n 0.0051638f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_466 N_A_286_413#_c_639_n N_VPWR_c_867_n 0.0295853f $X=2.03 $Y=2.295 $X2=0
+ $Y2=0
cc_467 N_A_286_413#_c_630_n N_VPWR_c_867_n 0.00379592f $X=2.115 $Y=2.125 $X2=0
+ $Y2=0
cc_468 N_A_286_413#_c_635_n N_A_27_47#_c_979_n 0.0218946f $X=2.325 $Y=0.395
+ $X2=0 $Y2=0
cc_469 N_A_286_413#_c_639_n A_382_413# 0.00832946f $X=2.03 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_470 N_A_286_413#_c_630_n A_382_413# 0.00151526f $X=2.115 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_471 N_A_286_413#_c_624_n N_VGND_c_1022_n 0.00741046f $X=3.095 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_286_413#_c_635_n N_VGND_c_1022_n 0.0231479f $X=2.325 $Y=0.395 $X2=0
+ $Y2=0
cc_473 N_A_286_413#_c_625_n N_VGND_c_1022_n 0.0210362f $X=2.41 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_286_413#_c_627_n N_VGND_c_1022_n 0.0221749f $X=2.925 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_A_286_413#_c_628_n N_VGND_c_1022_n 0.00483796f $X=3.105 $Y=1.16 $X2=0
+ $Y2=0
cc_476 N_A_286_413#_c_635_n N_VGND_c_1025_n 0.0673769f $X=2.325 $Y=0.395 $X2=0
+ $Y2=0
cc_477 N_A_286_413#_c_624_n N_VGND_c_1026_n 0.00585385f $X=3.095 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_286_413#_M1019_d N_VGND_c_1028_n 0.00299551f $X=1.445 $Y=0.235 $X2=0
+ $Y2=0
cc_479 N_A_286_413#_c_624_n N_VGND_c_1028_n 0.00789762f $X=3.095 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_A_286_413#_c_635_n N_VGND_c_1028_n 0.0299006f $X=2.325 $Y=0.395 $X2=0
+ $Y2=0
cc_481 N_A_286_413#_c_635_n A_394_47# 0.00874765f $X=2.325 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_482 N_A_286_413#_c_625_n A_394_47# 0.00160798f $X=2.41 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_483 N_CLK_M1012_g N_A_1012_47#_M1009_g 0.035715f $X=5.955 $Y=2.165 $X2=0
+ $Y2=0
cc_484 N_CLK_M1004_g N_A_1012_47#_c_799_n 0.0115624f $X=5.955 $Y=0.445 $X2=0
+ $Y2=0
cc_485 N_CLK_c_729_n N_A_1012_47#_c_799_n 0.0553291f $X=5.845 $Y=1.05 $X2=0
+ $Y2=0
cc_486 N_CLK_c_730_n N_A_1012_47#_c_799_n 0.00451117f $X=5.845 $Y=1.05 $X2=0
+ $Y2=0
cc_487 N_CLK_c_727_n N_A_1012_47#_c_800_n 3.83662e-19 $X=4.655 $Y=0.73 $X2=0
+ $Y2=0
cc_488 N_CLK_c_728_n N_A_1012_47#_c_800_n 6.28557e-19 $X=4.655 $Y=0.88 $X2=0
+ $Y2=0
cc_489 N_CLK_c_729_n N_A_1012_47#_c_800_n 0.022455f $X=5.845 $Y=1.05 $X2=0 $Y2=0
cc_490 N_CLK_M1012_g N_A_1012_47#_c_801_n 0.0269046f $X=5.955 $Y=2.165 $X2=0
+ $Y2=0
cc_491 N_CLK_c_729_n N_A_1012_47#_c_801_n 0.045368f $X=5.845 $Y=1.05 $X2=0 $Y2=0
cc_492 N_CLK_c_730_n N_A_1012_47#_c_801_n 0.00645493f $X=5.845 $Y=1.05 $X2=0
+ $Y2=0
cc_493 N_CLK_M1004_g N_A_1012_47#_c_802_n 0.00394742f $X=5.955 $Y=0.445 $X2=0
+ $Y2=0
cc_494 N_CLK_c_729_n N_A_1012_47#_c_802_n 0.00294772f $X=5.845 $Y=1.05 $X2=0
+ $Y2=0
cc_495 N_CLK_c_729_n N_A_1012_47#_c_803_n 2.92443e-19 $X=5.845 $Y=1.05 $X2=0
+ $Y2=0
cc_496 N_CLK_c_730_n N_A_1012_47#_c_803_n 0.0201268f $X=5.845 $Y=1.05 $X2=0
+ $Y2=0
cc_497 N_CLK_M1004_g N_A_1012_47#_c_804_n 0.0205784f $X=5.955 $Y=0.445 $X2=0
+ $Y2=0
cc_498 N_CLK_M1012_g N_VPWR_c_859_n 0.00166155f $X=5.955 $Y=2.165 $X2=0 $Y2=0
cc_499 N_CLK_c_735_n N_VPWR_c_862_n 0.0240974f $X=4.72 $Y=1.325 $X2=0 $Y2=0
cc_500 N_CLK_M1012_g N_VPWR_c_863_n 0.00424239f $X=5.955 $Y=2.165 $X2=0 $Y2=0
cc_501 N_CLK_M1012_g N_VPWR_c_856_n 0.00576116f $X=5.955 $Y=2.165 $X2=0 $Y2=0
cc_502 N_CLK_M1012_g N_VPWR_c_868_n 5.79077e-19 $X=5.955 $Y=2.165 $X2=0 $Y2=0
cc_503 N_CLK_c_727_n N_VGND_c_1023_n 0.00809304f $X=4.655 $Y=0.73 $X2=0 $Y2=0
cc_504 N_CLK_c_727_n N_VGND_c_1028_n 0.0053254f $X=4.655 $Y=0.73 $X2=0 $Y2=0
cc_505 N_CLK_c_728_n N_VGND_c_1028_n 0.00262886f $X=4.655 $Y=0.88 $X2=0 $Y2=0
cc_506 N_CLK_c_727_n N_VGND_c_1032_n 0.00337001f $X=4.655 $Y=0.73 $X2=0 $Y2=0
cc_507 N_CLK_c_728_n N_VGND_c_1032_n 0.00230382f $X=4.655 $Y=0.88 $X2=0 $Y2=0
cc_508 N_CLK_M1004_g N_VGND_c_1033_n 0.0161364f $X=5.955 $Y=0.445 $X2=0 $Y2=0
cc_509 N_A_1012_47#_c_801_n N_VPWR_M1012_d 0.00224468f $X=5.745 $Y=2.085 $X2=0
+ $Y2=0
cc_510 N_A_1012_47#_M1009_g N_VPWR_c_859_n 0.00679186f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_A_1012_47#_c_801_n N_VPWR_c_859_n 0.0180293f $X=5.745 $Y=2.085 $X2=0
+ $Y2=0
cc_512 N_A_1012_47#_c_801_n N_VPWR_c_863_n 0.0145632f $X=5.745 $Y=2.085 $X2=0
+ $Y2=0
cc_513 N_A_1012_47#_M1009_g N_VPWR_c_864_n 0.00564095f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_514 N_A_1012_47#_M1016_d N_VPWR_c_856_n 0.00411223f $X=5.61 $Y=1.845 $X2=0
+ $Y2=0
cc_515 N_A_1012_47#_M1009_g N_VPWR_c_856_n 0.0104943f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_516 N_A_1012_47#_c_801_n N_VPWR_c_856_n 0.013348f $X=5.745 $Y=2.085 $X2=0
+ $Y2=0
cc_517 N_A_1012_47#_M1009_g N_GCLK_c_1005_n 0.00252176f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_518 N_A_1012_47#_c_801_n N_GCLK_c_1005_n 0.0289114f $X=5.745 $Y=2.085 $X2=0
+ $Y2=0
cc_519 N_A_1012_47#_c_802_n N_GCLK_c_1005_n 0.00580475f $X=6.275 $Y=0.995 $X2=0
+ $Y2=0
cc_520 N_A_1012_47#_c_803_n N_GCLK_c_1005_n 0.00745796f $X=6.375 $Y=1.16 $X2=0
+ $Y2=0
cc_521 N_A_1012_47#_c_804_n N_GCLK_c_1005_n 0.00252314f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_522 N_A_1012_47#_c_799_n N_VGND_M1004_d 0.00383986f $X=6.19 $Y=0.7 $X2=0
+ $Y2=0
cc_523 N_A_1012_47#_c_802_n N_VGND_M1004_d 0.00114081f $X=6.275 $Y=0.995 $X2=0
+ $Y2=0
cc_524 N_A_1012_47#_c_804_n N_VGND_c_1027_n 0.00564095f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_525 N_A_1012_47#_M1002_s N_VGND_c_1028_n 0.00226128f $X=5.06 $Y=0.235 $X2=0
+ $Y2=0
cc_526 N_A_1012_47#_c_798_n N_VGND_c_1028_n 0.00987224f $X=5.185 $Y=0.46 $X2=0
+ $Y2=0
cc_527 N_A_1012_47#_c_799_n N_VGND_c_1028_n 0.00996785f $X=6.19 $Y=0.7 $X2=0
+ $Y2=0
cc_528 N_A_1012_47#_c_804_n N_VGND_c_1028_n 0.0103332f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_529 N_A_1012_47#_c_798_n N_VGND_c_1032_n 0.0176791f $X=5.185 $Y=0.46 $X2=0
+ $Y2=0
cc_530 N_A_1012_47#_c_799_n N_VGND_c_1032_n 0.00343228f $X=6.19 $Y=0.7 $X2=0
+ $Y2=0
cc_531 N_A_1012_47#_c_799_n N_VGND_c_1033_n 0.0499364f $X=6.19 $Y=0.7 $X2=0
+ $Y2=0
cc_532 N_A_1012_47#_c_803_n N_VGND_c_1033_n 3.22676e-19 $X=6.375 $Y=1.16 $X2=0
+ $Y2=0
cc_533 N_A_1012_47#_c_804_n N_VGND_c_1033_n 0.00694329f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_534 N_A_1012_47#_c_799_n A_1094_47# 0.00313031f $X=6.19 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_535 N_VPWR_c_856_n A_109_369# 0.00168632f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_536 N_VPWR_c_856_n N_A_27_47#_M1005_d 0.00382866f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_537 N_VPWR_c_858_n N_A_27_47#_c_952_n 0.00910312f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_538 N_VPWR_c_856_n N_A_27_47#_c_959_n 0.00651891f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_c_866_n N_A_27_47#_c_959_n 0.00953989f $X=2.37 $Y=2.44 $X2=0 $Y2=0
cc_540 N_VPWR_c_856_n N_A_27_47#_c_969_n 0.0198554f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_541 N_VPWR_c_866_n N_A_27_47#_c_969_n 0.0317135f $X=2.37 $Y=2.44 $X2=0 $Y2=0
cc_542 N_VPWR_c_856_n A_382_413# 0.00809303f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_543 N_VPWR_c_856_n N_GCLK_M1009_d 0.00300383f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_544 N_VPWR_c_864_n GCLK 0.0188881f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_545 N_VPWR_c_856_n GCLK 0.0108988f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_546 A_109_369# N_A_27_47#_c_959_n 9.38831e-19 $X=0.545 $Y=1.845 $X2=6.195
+ $Y2=2.635
cc_547 N_A_27_47#_c_949_n N_VGND_M1020_d 7.84403e-19 $X=1.015 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_548 N_A_27_47#_c_950_n N_VGND_M1020_d 7.9459e-19 $X=0.68 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_549 N_A_27_47#_c_950_n N_VGND_c_1021_n 0.0158273f $X=0.68 $Y=0.7 $X2=0 $Y2=0
cc_550 N_A_27_47#_c_948_n N_VGND_c_1024_n 0.0172026f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_551 N_A_27_47#_c_950_n N_VGND_c_1024_n 0.00258611f $X=0.68 $Y=0.7 $X2=0 $Y2=0
cc_552 N_A_27_47#_c_949_n N_VGND_c_1025_n 0.00256355f $X=1.015 $Y=0.7 $X2=0
+ $Y2=0
cc_553 N_A_27_47#_c_979_n N_VGND_c_1025_n 0.0117453f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_554 N_A_27_47#_M1020_s N_VGND_c_1028_n 0.00226128f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_555 N_A_27_47#_M1008_d N_VGND_c_1028_n 0.00611112f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_556 N_A_27_47#_c_948_n N_VGND_c_1028_n 0.00977915f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_557 N_A_27_47#_c_949_n N_VGND_c_1028_n 0.00427891f $X=1.015 $Y=0.7 $X2=0
+ $Y2=0
cc_558 N_A_27_47#_c_950_n N_VGND_c_1028_n 0.00582244f $X=0.68 $Y=0.7 $X2=0 $Y2=0
cc_559 N_A_27_47#_c_979_n N_VGND_c_1028_n 0.00661975f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_560 N_GCLK_c_1006_n N_VGND_c_1027_n 0.0188134f $X=6.64 $Y=0.42 $X2=0 $Y2=0
cc_561 N_GCLK_M1013_d N_VGND_c_1028_n 0.00296108f $X=6.505 $Y=0.235 $X2=0 $Y2=0
cc_562 N_GCLK_c_1006_n N_VGND_c_1028_n 0.0108787f $X=6.64 $Y=0.42 $X2=0 $Y2=0
cc_563 N_VGND_c_1028_n A_394_47# 0.00299863f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_564 N_VGND_c_1028_n A_1094_47# 3.8732e-19 $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_565 N_VGND_c_1033_n A_1094_47# 0.00502403f $X=6.36 $Y=0.18 $X2=-0.19
+ $Y2=-0.24

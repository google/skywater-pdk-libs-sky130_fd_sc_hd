* File: sky130_fd_sc_hd__o41a_1.pex.spice
* Created: Tue Sep  1 19:26:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O41A_1%A_103_21# 1 2 7 9 12 15 18 22 26 27 33
c53 27 0 1.07318e-19 $X=0.975 $Y=1
c54 26 0 1.56343e-19 $X=0.69 $Y=1.16
c55 15 0 1.81202e-19 $X=0.975 $Y=1.455
r56 31 33 1.58958 $w=2.88e-07 $l=4e-08 $layer=LI1_cond $X=1.47 $Y=1.6 $X2=1.51
+ $Y2=1.6
r57 29 31 19.671 $w=2.88e-07 $l=4.95e-07 $layer=LI1_cond $X=0.975 $Y=1.6
+ $X2=1.47 $Y2=1.6
r58 26 37 16.3642 $w=3.24e-07 $l=1.1e-07 $layer=POLY_cond $X=0.69 $Y=1.16
+ $X2=0.8 $Y2=1.16
r59 26 35 14.8765 $w=3.24e-07 $l=1e-07 $layer=POLY_cond $X=0.69 $Y=1.16 $X2=0.59
+ $Y2=1.16
r60 25 27 10.2265 $w=3.4e-07 $l=3.56125e-07 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.975 $Y2=1
r61 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.16 $X2=0.69 $Y2=1.16
r62 20 31 1.60663 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=1.47 $Y=1.745
+ $X2=1.47 $Y2=1.6
r63 20 22 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.47 $Y=1.745
+ $X2=1.47 $Y2=1.96
r64 16 27 12.3794 $w=3.4e-07 $l=4.66208e-07 $layer=LI1_cond $X=1.32 $Y=0.715
+ $X2=0.975 $Y2=1
r65 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.32 $Y=0.715
+ $X2=1.32 $Y2=0.38
r66 15 29 1.37394 $w=2.6e-07 $l=1.45e-07 $layer=LI1_cond $X=0.975 $Y=1.455
+ $X2=0.975 $Y2=1.6
r67 14 27 2.31059 $w=2.6e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=1.285
+ $X2=0.975 $Y2=1
r68 14 15 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.975 $Y=1.285
+ $X2=0.975 $Y2=1.455
r69 10 37 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.8 $Y=1.325
+ $X2=0.8 $Y2=1.16
r70 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.8 $Y=1.325 $X2=0.8
+ $Y2=1.985
r71 7 35 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=0.995
+ $X2=0.59 $Y2=1.16
r72 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.59 $Y=0.995 $X2=0.59
+ $Y2=0.56
r73 2 33 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=1.295
+ $Y=1.485 $X2=1.51 $Y2=1.62
r74 2 22 300 $w=1.7e-07 $l=5.72495e-07 $layer=licon1_PDIFF $count=2 $X=1.295
+ $Y=1.485 $X2=1.51 $Y2=1.96
r75 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.195
+ $Y=0.235 $X2=1.32 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%B1 3 5 7 8 12
c30 8 0 1.56343e-19 $X=1.61 $Y=1.19
r31 12 14 14.6554 $w=2.96e-07 $l=9e-08 $layer=POLY_cond $X=1.44 $Y=1.16 $X2=1.53
+ $Y2=1.16
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.44
+ $Y=1.16 $X2=1.44 $Y2=1.16
r33 10 12 35.8243 $w=2.96e-07 $l=2.2e-07 $layer=POLY_cond $X=1.22 $Y=1.16
+ $X2=1.44 $Y2=1.16
r34 8 13 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=1.61 $Y=1.18 $X2=1.44
+ $Y2=1.18
r35 5 14 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=1.16
r36 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.53 $Y=0.995 $X2=1.53
+ $Y2=0.56
r37 1 10 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.325
+ $X2=1.22 $Y2=1.16
r38 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.22 $Y=1.325 $X2=1.22
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%A4 1 3 5 7 8 9 10 16
c38 5 0 1.07318e-19 $X=1.95 $Y=0.995
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.16 $X2=2.03 $Y2=1.16
r40 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.03 $Y=1.87 $X2=2.03
+ $Y2=2.21
r41 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.03 $Y=1.53 $X2=2.03
+ $Y2=1.87
r42 8 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.03 $Y=1.53 $X2=2.03
+ $Y2=1.16
r43 5 15 38.9379 $w=3.62e-07 $l=1.90526e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=2.005 $Y2=1.16
r44 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995 $X2=1.95
+ $Y2=0.56
r45 1 15 38.9379 $w=3.62e-07 $l=2.14942e-07 $layer=POLY_cond $X=1.89 $Y=1.325
+ $X2=2.005 $Y2=1.16
r46 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.89 $Y=1.325 $X2=1.89
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%A3 3 6 8 9 10 15 16 17
r34 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.57 $Y2=1.325
r35 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.57 $Y2=0.995
r36 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.16 $X2=2.57 $Y2=1.16
r37 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.57 $Y=1.87 $X2=2.57
+ $Y2=2.21
r38 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.57 $Y=1.53 $X2=2.57
+ $Y2=1.87
r39 8 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.57 $Y=1.53 $X2=2.57
+ $Y2=1.16
r40 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.48 $Y=1.985
+ $X2=2.48 $Y2=1.325
r41 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.48 $Y=0.56 $X2=2.48
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%A2 3 6 8 9 10 15 16 17
r35 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.16
+ $X2=3.11 $Y2=1.325
r36 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.16
+ $X2=3.11 $Y2=0.995
r37 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.16 $X2=3.11 $Y2=1.16
r38 9 10 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.09 $Y=1.87 $X2=3.09
+ $Y2=2.21
r39 8 9 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.09 $Y=1.53 $X2=3.09
+ $Y2=1.87
r40 8 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=1.53 $X2=3.09
+ $Y2=1.16
r41 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.02 $Y=1.985
+ $X2=3.02 $Y2=1.325
r42 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.02 $Y=0.56 $X2=3.02
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%A1 3 6 8 11 13
r25 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.16
+ $X2=3.65 $Y2=1.325
r26 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.16
+ $X2=3.65 $Y2=0.995
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.65
+ $Y=1.16 $X2=3.65 $Y2=1.16
r28 8 12 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=3.91 $Y=1.2 $X2=3.65
+ $Y2=1.2
r29 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.56 $Y=1.985
+ $X2=3.56 $Y2=1.325
r30 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.56 $Y=0.56 $X2=3.56
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%X 1 2 7 8 9 10 11 12 23 43 46
r21 46 47 4.52128 $w=5.23e-07 $l=7.5e-08 $layer=LI1_cond $X=0.347 $Y=1.53
+ $X2=0.347 $Y2=1.455
r22 43 44 1.7075 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=0.255 $Y=0.85
+ $X2=0.255 $Y2=0.885
r23 33 50 1.98207 $w=5.23e-07 $l=8.7e-08 $layer=LI1_cond $X=0.347 $Y=1.717
+ $X2=0.347 $Y2=1.63
r24 12 39 2.27824 $w=5.23e-07 $l=1e-07 $layer=LI1_cond $X=0.347 $Y=2.21
+ $X2=0.347 $Y2=2.31
r25 11 12 7.74603 $w=5.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.347 $Y=1.87
+ $X2=0.347 $Y2=2.21
r26 11 33 3.48571 $w=5.23e-07 $l=1.53e-07 $layer=LI1_cond $X=0.347 $Y=1.87
+ $X2=0.347 $Y2=1.717
r27 10 50 2.16433 $w=5.23e-07 $l=9.5e-08 $layer=LI1_cond $X=0.347 $Y=1.535
+ $X2=0.347 $Y2=1.63
r28 10 46 0.113912 $w=5.23e-07 $l=5e-09 $layer=LI1_cond $X=0.347 $Y=1.535
+ $X2=0.347 $Y2=1.53
r29 10 47 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=0.22 $Y=1.45 $X2=0.22
+ $Y2=1.455
r30 9 10 11.0976 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.22 $Y=1.19 $X2=0.22
+ $Y2=1.45
r31 8 43 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=0.255 $Y=0.825
+ $X2=0.255 $Y2=0.85
r32 8 21 3.72849 $w=3.38e-07 $l=1.1e-07 $layer=LI1_cond $X=0.255 $Y=0.825
+ $X2=0.255 $Y2=0.715
r33 8 9 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.22 $Y=0.91 $X2=0.22
+ $Y2=1.19
r34 8 44 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.22 $Y=0.91 $X2=0.22
+ $Y2=0.885
r35 7 21 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.255 $Y=0.51
+ $X2=0.255 $Y2=0.715
r36 7 23 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=0.51
+ $X2=0.255 $Y2=0.38
r37 2 50 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.445 $Y2=1.63
r38 2 39 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.445 $Y2=2.31
r39 1 23 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%VPWR 1 2 9 11 13 17 19 24 30 34
r46 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r47 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r49 28 31 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 25 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=2.72
+ $X2=1.01 $Y2=2.72
r52 25 27 148.422 $w=1.68e-07 $l=2.275e-06 $layer=LI1_cond $X=1.175 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 24 33 4.56733 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=3.605 $Y=2.72
+ $X2=3.872 $Y2=2.72
r54 24 27 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.605 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 22 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.01 $Y2=2.72
r58 19 21 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 17 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 13 16 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.77 $Y=1.66
+ $X2=3.77 $Y2=2.34
r61 11 33 3.19884 $w=3.3e-07 $l=1.38109e-07 $layer=LI1_cond $X=3.77 $Y=2.635
+ $X2=3.872 $Y2=2.72
r62 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.77 $Y=2.635
+ $X2=3.77 $Y2=2.34
r63 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.01 $Y=2.635 $X2=1.01
+ $Y2=2.72
r64 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.01 $Y=2.635
+ $X2=1.01 $Y2=2
r65 2 16 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.485 $X2=3.77 $Y2=2.34
r66 2 13 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.485 $X2=3.77 $Y2=1.66
r67 1 9 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.875
+ $Y=1.485 $X2=1.01 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%VGND 1 2 3 12 16 20 23 24 26 27 28 34 43 44
+ 47
r60 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r61 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r62 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r63 41 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r64 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r65 38 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.215
+ $Y2=0
r66 38 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.99
+ $Y2=0
r67 37 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r68 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.215
+ $Y2=0
r70 34 36 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=1.15
+ $Y2=0
r71 32 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r72 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r73 28 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r74 26 40 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=2.99
+ $Y2=0
r75 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.29
+ $Y2=0
r76 25 43 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.91
+ $Y2=0
r77 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.29
+ $Y2=0
r78 23 31 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.69
+ $Y2=0
r79 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.8
+ $Y2=0
r80 22 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.15
+ $Y2=0
r81 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.8
+ $Y2=0
r82 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0
r83 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.29 $Y=0.085
+ $X2=3.29 $Y2=0.38
r84 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0
r85 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0.38
r86 10 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r87 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0.38
r88 3 20 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.235 $X2=3.29 $Y2=0.38
r89 2 16 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.215 $Y2=0.38
r90 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.665
+ $Y=0.235 $X2=0.8 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_1%A_321_47# 1 2 3 12 14 15 18 20 24 26
r44 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.79 $Y=0.735
+ $X2=3.79 $Y2=0.4
r45 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=0.82
+ $X2=2.745 $Y2=0.82
r46 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.625 $Y=0.82
+ $X2=3.79 $Y2=0.735
r47 20 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.625 $Y=0.82
+ $X2=2.91 $Y2=0.82
r48 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=0.735
+ $X2=2.745 $Y2=0.82
r49 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.745 $Y=0.735
+ $X2=2.745 $Y2=0.4
r50 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0.82
+ $X2=2.745 $Y2=0.82
r51 14 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.58 $Y=0.82
+ $X2=1.825 $Y2=0.82
r52 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.74 $Y=0.735
+ $X2=1.825 $Y2=0.82
r53 10 12 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.74 $Y=0.735
+ $X2=1.74 $Y2=0.58
r54 3 24 91 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=2 $X=3.635
+ $Y=0.235 $X2=3.79 $Y2=0.4
r55 2 18 91 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=2 $X=2.555
+ $Y=0.235 $X2=2.745 $Y2=0.4
r56 1 12 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.235 $X2=1.74 $Y2=0.58
.ends


* File: sky130_fd_sc_hd__a211o_4.pxi.spice
* Created: Tue Sep  1 18:50:58 2020
* 
x_PM_SKY130_FD_SC_HD__A211O_4%A_79_204# N_A_79_204#_M1014_d N_A_79_204#_M1007_d
+ N_A_79_204#_M1018_s N_A_79_204#_M1008_s N_A_79_204#_M1000_g
+ N_A_79_204#_M1003_g N_A_79_204#_M1004_g N_A_79_204#_M1011_g
+ N_A_79_204#_M1012_g N_A_79_204#_M1013_g N_A_79_204#_M1015_g
+ N_A_79_204#_M1022_g N_A_79_204#_c_172_p N_A_79_204#_c_106_n
+ N_A_79_204#_c_113_n N_A_79_204#_c_120_p N_A_79_204#_c_201_p
+ N_A_79_204#_c_114_n N_A_79_204#_c_122_p N_A_79_204#_c_242_p
+ N_A_79_204#_c_147_p N_A_79_204#_c_140_p N_A_79_204#_c_153_p
+ N_A_79_204#_c_107_n N_A_79_204#_c_115_n N_A_79_204#_c_116_n
+ N_A_79_204#_c_133_p N_A_79_204#_c_139_p N_A_79_204#_c_108_n
+ PM_SKY130_FD_SC_HD__A211O_4%A_79_204#
x_PM_SKY130_FD_SC_HD__A211O_4%B1 N_B1_M1014_g N_B1_M1023_g N_B1_M1010_g
+ N_B1_M1017_g N_B1_c_266_n N_B1_c_267_n B1 N_B1_c_268_n N_B1_c_269_n
+ N_B1_c_270_n N_B1_c_278_n PM_SKY130_FD_SC_HD__A211O_4%B1
x_PM_SKY130_FD_SC_HD__A211O_4%C1 N_C1_c_359_n N_C1_M1002_g N_C1_M1008_g
+ N_C1_c_360_n N_C1_M1007_g N_C1_M1020_g C1 PM_SKY130_FD_SC_HD__A211O_4%C1
x_PM_SKY130_FD_SC_HD__A211O_4%A2 N_A2_M1001_g N_A2_M1005_g N_A2_M1006_g
+ N_A2_M1009_g N_A2_c_403_n N_A2_c_404_n N_A2_c_433_p N_A2_c_428_n N_A2_c_405_n
+ N_A2_c_406_n A2 N_A2_c_414_n N_A2_c_407_n N_A2_c_453_p
+ PM_SKY130_FD_SC_HD__A211O_4%A2
x_PM_SKY130_FD_SC_HD__A211O_4%A1 N_A1_M1018_g N_A1_M1016_g N_A1_M1019_g
+ N_A1_M1021_g A1 N_A1_c_486_n PM_SKY130_FD_SC_HD__A211O_4%A1
x_PM_SKY130_FD_SC_HD__A211O_4%VPWR N_VPWR_M1000_d N_VPWR_M1004_d N_VPWR_M1015_d
+ N_VPWR_M1001_d N_VPWR_M1021_s N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n
+ VPWR N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n
+ N_VPWR_c_532_n N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_c_548_n
+ PM_SKY130_FD_SC_HD__A211O_4%VPWR
x_PM_SKY130_FD_SC_HD__A211O_4%X N_X_M1003_d N_X_M1013_d N_X_M1000_s N_X_M1012_s
+ N_X_c_638_n N_X_c_646_n N_X_c_641_n N_X_c_671_n N_X_c_648_n N_X_c_683_p
+ N_X_c_652_n N_X_c_675_n N_X_c_681_p N_X_c_659_n N_X_c_661_n X N_X_c_640_n
+ PM_SKY130_FD_SC_HD__A211O_4%X
x_PM_SKY130_FD_SC_HD__A211O_4%A_473_297# N_A_473_297#_M1023_d
+ N_A_473_297#_M1010_d N_A_473_297#_M1016_d N_A_473_297#_M1009_s
+ N_A_473_297#_c_696_n N_A_473_297#_c_716_n N_A_473_297#_c_720_n
+ N_A_473_297#_c_721_n N_A_473_297#_c_697_n N_A_473_297#_c_698_n
+ N_A_473_297#_c_712_n N_A_473_297#_c_728_n N_A_473_297#_c_699_n
+ PM_SKY130_FD_SC_HD__A211O_4%A_473_297#
x_PM_SKY130_FD_SC_HD__A211O_4%VGND N_VGND_M1003_s N_VGND_M1011_s N_VGND_M1022_s
+ N_VGND_M1002_s N_VGND_M1017_s N_VGND_M1006_d N_VGND_c_771_n N_VGND_c_772_n
+ N_VGND_c_773_n N_VGND_c_774_n N_VGND_c_775_n N_VGND_c_776_n N_VGND_c_777_n
+ N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n
+ VGND N_VGND_c_783_n N_VGND_c_784_n N_VGND_c_785_n N_VGND_c_786_n
+ N_VGND_c_787_n N_VGND_c_788_n PM_SKY130_FD_SC_HD__A211O_4%VGND
cc_1 VNB N_A_79_204#_M1003_g 0.0205675f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.56
cc_2 VNB N_A_79_204#_M1011_g 0.0172777f $X=-0.19 $Y=-0.24 $X2=1.295 $Y2=0.56
cc_3 VNB N_A_79_204#_M1013_g 0.0174281f $X=-0.19 $Y=-0.24 $X2=1.725 $Y2=0.56
cc_4 VNB N_A_79_204#_M1022_g 0.0169336f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.56
cc_5 VNB N_A_79_204#_c_106_n 0.00129982f $X=-0.19 $Y=-0.24 $X2=2.282 $Y2=1.045
cc_6 VNB N_A_79_204#_c_107_n 0.00154767f $X=-0.19 $Y=-0.24 $X2=2.277 $Y2=1.185
cc_7 VNB N_A_79_204#_c_108_n 0.083674f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.185
cc_8 VNB N_B1_M1014_g 0.0179991f $X=-0.19 $Y=-0.24 $X2=5.185 $Y2=0.235
cc_9 VNB N_B1_c_266_n 0.00327371f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.02
cc_10 VNB N_B1_c_267_n 0.0225317f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.56
cc_11 VNB N_B1_c_268_n 0.0283686f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.35
cc_12 VNB N_B1_c_269_n 0.00170273f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_13 VNB N_B1_c_270_n 0.018232f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_14 VNB N_C1_c_359_n 0.0167819f $X=-0.19 $Y=-0.24 $X2=2.68 $Y2=0.235
cc_15 VNB N_C1_c_360_n 0.0500746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB C1 0.00763388f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_17 VNB N_A2_M1005_g 0.0194047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_403_n 0.00181812f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.02
cc_19 VNB N_A2_c_404_n 0.0257502f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.56
cc_20 VNB N_A2_c_405_n 0.0236892f $X=-0.19 $Y=-0.24 $X2=1.295 $Y2=0.56
cc_21 VNB N_A2_c_406_n 0.0274483f $X=-0.19 $Y=-0.24 $X2=1.295 $Y2=0.56
cc_22 VNB N_A2_c_407_n 0.0226581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A1_M1018_g 0.0177577f $X=-0.19 $Y=-0.24 $X2=5.185 $Y2=0.235
cc_24 VNB N_A1_M1019_g 0.0177577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB A1 0.00187742f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.02
cc_26 VNB N_A1_c_486_n 0.0284649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_532_n 0.269736f $X=-0.19 $Y=-0.24 $X2=2.847 $Y2=0.615
cc_28 VNB N_X_c_638_n 0.00564768f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.35
cc_29 VNB X 0.0231545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_640_n 0.0154224f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.56
cc_31 VNB N_VGND_c_771_n 0.0118295f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.35
cc_32 VNB N_VGND_c_772_n 3.11777e-19 $X=-0.19 $Y=-0.24 $X2=1.295 $Y2=1.02
cc_33 VNB N_VGND_c_773_n 3.2118e-19 $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.35
cc_34 VNB N_VGND_c_774_n 0.00283357f $X=-0.19 $Y=-0.24 $X2=1.725 $Y2=1.02
cc_35 VNB N_VGND_c_775_n 0.0103361f $X=-0.19 $Y=-0.24 $X2=1.725 $Y2=0.56
cc_36 VNB N_VGND_c_776_n 0.02635f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.35
cc_37 VNB N_VGND_c_777_n 0.011382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_778_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.02
cc_39 VNB N_VGND_c_779_n 0.0126059f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.56
cc_40 VNB N_VGND_c_780_n 0.00442675f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_781_n 0.0125844f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=1.185
cc_42 VNB N_VGND_c_782_n 0.00518879f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=1.16
cc_43 VNB N_VGND_c_783_n 0.015802f $X=-0.19 $Y=-0.24 $X2=1.76 $Y2=1.185
cc_44 VNB N_VGND_c_784_n 0.0177311f $X=-0.19 $Y=-0.24 $X2=2.847 $Y2=0.615
cc_45 VNB N_VGND_c_785_n 0.0394683f $X=-0.19 $Y=-0.24 $X2=3.64 $Y2=0.71
cc_46 VNB N_VGND_c_786_n 0.00510127f $X=-0.19 $Y=-0.24 $X2=2.32 $Y2=1.505
cc_47 VNB N_VGND_c_787_n 0.0129739f $X=-0.19 $Y=-0.24 $X2=3.835 $Y2=0.38
cc_48 VNB N_VGND_c_788_n 0.317454f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.185
cc_49 VPB N_A_79_204#_M1000_g 0.0197402f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_50 VPB N_A_79_204#_M1004_g 0.017272f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_51 VPB N_A_79_204#_M1012_g 0.0172777f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_52 VPB N_A_79_204#_M1015_g 0.0203042f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.985
cc_53 VPB N_A_79_204#_c_113_n 0.00268425f $X=-0.19 $Y=1.305 $X2=2.367 $Y2=1.87
cc_54 VPB N_A_79_204#_c_114_n 0.00279781f $X=-0.19 $Y=1.305 $X2=2.455 $Y2=1.955
cc_55 VPB N_A_79_204#_c_115_n 0.00285344f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=1.505
cc_56 VPB N_A_79_204#_c_116_n 0.00652825f $X=-0.19 $Y=1.305 $X2=2.32 $Y2=1.675
cc_57 VPB N_A_79_204#_c_108_n 0.0334604f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.185
cc_58 VPB N_B1_M1023_g 0.0210125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B1_M1010_g 0.0178502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_B1_c_266_n 0.00285595f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=1.02
cc_61 VPB N_B1_c_267_n 0.00858112f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.56
cc_62 VPB B1 3.31243e-19 $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.35
cc_63 VPB N_B1_c_268_n 0.00835654f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.35
cc_64 VPB N_B1_c_269_n 0.00177664f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_65 VPB N_B1_c_278_n 0.00894491f $X=-0.19 $Y=1.305 $X2=1.725 $Y2=1.02
cc_66 VPB N_C1_M1008_g 0.0170078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_C1_c_360_n 0.00882467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_C1_M1020_g 0.0173901f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.35
cc_69 VPB N_A2_M1009_g 0.0240847f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.35
cc_70 VPB N_A2_c_403_n 9.11121e-19 $X=-0.19 $Y=1.305 $X2=0.865 $Y2=1.02
cc_71 VPB N_A2_c_404_n 0.0121347f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.56
cc_72 VPB N_A2_c_405_n 0.00208175f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.56
cc_73 VPB N_A2_c_406_n 0.00872176f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.56
cc_74 VPB A2 0.00364793f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.35
cc_75 VPB N_A2_c_414_n 0.0161941f $X=-0.19 $Y=1.305 $X2=1.725 $Y2=0.56
cc_76 VPB N_A1_M1016_g 0.0184144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A1_M1021_g 0.0174653f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_78 VPB N_A1_c_486_n 0.00663166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_533_n 0.0101444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_534_n 0.0268137f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.56
cc_81 VPB N_VPWR_c_535_n 3.08203e-19 $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_82 VPB N_VPWR_c_536_n 0.00231076f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.56
cc_83 VPB N_VPWR_c_537_n 0.00227979f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_84 VPB N_VPWR_c_538_n 4.16958e-19 $X=-0.19 $Y=1.305 $X2=1.725 $Y2=0.56
cc_85 VPB N_VPWR_c_539_n 0.0129398f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.35
cc_86 VPB N_VPWR_c_540_n 0.00356964f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.985
cc_87 VPB N_VPWR_c_541_n 0.0128277f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.02
cc_88 VPB N_VPWR_c_542_n 0.0588538f $X=-0.19 $Y=1.305 $X2=1.76 $Y2=1.185
cc_89 VPB N_VPWR_c_543_n 0.0149278f $X=-0.19 $Y=1.305 $X2=2.367 $Y2=1.675
cc_90 VPB N_VPWR_c_544_n 0.014469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_532_n 0.0524445f $X=-0.19 $Y=1.305 $X2=2.847 $Y2=0.615
cc_92 VPB N_VPWR_c_546_n 0.00436868f $X=-0.19 $Y=1.305 $X2=5.16 $Y2=0.71
cc_93 VPB N_VPWR_c_547_n 0.00510002f $X=-0.19 $Y=1.305 $X2=5.325 $Y2=0.36
cc_94 VPB N_VPWR_c_548_n 0.00436029f $X=-0.19 $Y=1.305 $X2=2.277 $Y2=1.185
cc_95 VPB N_X_c_641_n 0.00955713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB X 0.00939098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_473_297#_c_696_n 0.00328414f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.35
cc_98 VPB N_A_473_297#_c_697_n 0.014905f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=0.56
cc_99 VPB N_A_473_297#_c_698_n 0.013765f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_100 VPB N_A_473_297#_c_699_n 0.00949656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 N_A_79_204#_M1022_g N_B1_M1014_g 0.0250239f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_102 N_A_79_204#_c_106_n N_B1_M1014_g 0.00397747f $X=2.282 $Y=1.045 $X2=0
+ $Y2=0
cc_103 N_A_79_204#_c_120_p N_B1_M1014_g 0.0119808f $X=2.725 $Y=0.71 $X2=0 $Y2=0
cc_104 N_A_79_204#_c_113_n N_B1_M1023_g 0.00582257f $X=2.367 $Y=1.87 $X2=0 $Y2=0
cc_105 N_A_79_204#_c_122_p N_B1_M1023_g 0.0119077f $X=3.345 $Y=1.955 $X2=0 $Y2=0
cc_106 N_A_79_204#_c_115_n N_B1_M1023_g 0.00101667f $X=2.32 $Y=1.505 $X2=0 $Y2=0
cc_107 N_A_79_204#_c_116_n N_B1_M1023_g 0.00143344f $X=2.32 $Y=1.675 $X2=0 $Y2=0
cc_108 N_A_79_204#_c_122_p N_B1_M1010_g 5.29143e-19 $X=3.345 $Y=1.955 $X2=0
+ $Y2=0
cc_109 N_A_79_204#_M1022_g N_B1_c_266_n 3.00175e-19 $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A_79_204#_c_106_n N_B1_c_266_n 0.00439264f $X=2.282 $Y=1.045 $X2=0
+ $Y2=0
cc_111 N_A_79_204#_c_120_p N_B1_c_266_n 0.0119685f $X=2.725 $Y=0.71 $X2=0 $Y2=0
cc_112 N_A_79_204#_c_122_p N_B1_c_266_n 0.0131379f $X=3.345 $Y=1.955 $X2=0 $Y2=0
cc_113 N_A_79_204#_c_107_n N_B1_c_266_n 0.0233774f $X=2.277 $Y=1.185 $X2=0 $Y2=0
cc_114 N_A_79_204#_c_115_n N_B1_c_266_n 0.00988314f $X=2.32 $Y=1.505 $X2=0 $Y2=0
cc_115 N_A_79_204#_c_116_n N_B1_c_266_n 0.0157389f $X=2.32 $Y=1.675 $X2=0 $Y2=0
cc_116 N_A_79_204#_c_133_p N_B1_c_266_n 0.00647074f $X=2.847 $Y=0.71 $X2=0 $Y2=0
cc_117 N_A_79_204#_c_120_p N_B1_c_267_n 0.00156926f $X=2.725 $Y=0.71 $X2=0 $Y2=0
cc_118 N_A_79_204#_c_122_p N_B1_c_267_n 0.00362731f $X=3.345 $Y=1.955 $X2=0
+ $Y2=0
cc_119 N_A_79_204#_c_107_n N_B1_c_267_n 0.00203629f $X=2.277 $Y=1.185 $X2=0
+ $Y2=0
cc_120 N_A_79_204#_c_133_p N_B1_c_267_n 4.17163e-19 $X=2.847 $Y=0.71 $X2=0 $Y2=0
cc_121 N_A_79_204#_c_108_n N_B1_c_267_n 0.0199074f $X=2.17 $Y=1.185 $X2=0 $Y2=0
cc_122 N_A_79_204#_c_139_p N_B1_c_268_n 0.00116933f $X=3.835 $Y=0.38 $X2=0 $Y2=0
cc_123 N_A_79_204#_c_140_p N_B1_c_269_n 0.0111378f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_124 N_A_79_204#_c_139_p N_B1_c_269_n 0.0121488f $X=3.835 $Y=0.38 $X2=0 $Y2=0
cc_125 N_A_79_204#_c_140_p N_B1_c_270_n 0.0110655f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_126 N_A_79_204#_M1008_s N_B1_c_278_n 0.00179116f $X=3.205 $Y=1.485 $X2=0
+ $Y2=0
cc_127 N_A_79_204#_c_122_p N_B1_c_278_n 0.0370441f $X=3.345 $Y=1.955 $X2=0 $Y2=0
cc_128 N_A_79_204#_c_133_p N_B1_c_278_n 0.00482114f $X=2.847 $Y=0.71 $X2=0 $Y2=0
cc_129 N_A_79_204#_c_139_p N_B1_c_278_n 0.00561844f $X=3.835 $Y=0.38 $X2=0 $Y2=0
cc_130 N_A_79_204#_c_147_p N_C1_c_359_n 0.0121401f $X=3.64 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_79_204#_c_122_p N_C1_M1008_g 0.00837887f $X=3.345 $Y=1.955 $X2=0
+ $Y2=0
cc_132 N_A_79_204#_c_147_p N_C1_c_360_n 0.0127867f $X=3.64 $Y=0.71 $X2=0 $Y2=0
cc_133 N_A_79_204#_c_122_p N_C1_M1020_g 0.00385536f $X=3.345 $Y=1.955 $X2=0
+ $Y2=0
cc_134 N_A_79_204#_c_147_p C1 0.0425562f $X=3.64 $Y=0.71 $X2=0 $Y2=0
cc_135 N_A_79_204#_c_140_p N_A2_M1005_g 0.0135371f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_136 N_A_79_204#_c_153_p N_A2_M1005_g 0.00134108f $X=5.325 $Y=0.36 $X2=0 $Y2=0
cc_137 N_A_79_204#_c_140_p N_A2_c_403_n 0.0177345f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_138 N_A_79_204#_c_140_p N_A2_c_404_n 9.05102e-19 $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_139 N_A_79_204#_c_140_p N_A2_c_407_n 5.56146e-19 $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_140 N_A_79_204#_c_153_p N_A2_c_407_n 9.9802e-19 $X=5.325 $Y=0.36 $X2=0 $Y2=0
cc_141 N_A_79_204#_c_140_p N_A1_M1018_g 0.00988501f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_142 N_A_79_204#_c_153_p N_A1_M1018_g 0.00645865f $X=5.325 $Y=0.36 $X2=0 $Y2=0
cc_143 N_A_79_204#_c_140_p N_A1_M1019_g 0.00446953f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_144 N_A_79_204#_c_153_p N_A1_M1019_g 0.0061047f $X=5.325 $Y=0.36 $X2=0 $Y2=0
cc_145 N_A_79_204#_c_140_p A1 0.0200141f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_146 N_A_79_204#_c_140_p N_A1_c_486_n 0.00225214f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_147 N_A_79_204#_M1000_g N_VPWR_c_534_n 0.0117695f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_79_204#_M1004_g N_VPWR_c_534_n 6.17801e-19 $X=0.9 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_79_204#_M1000_g N_VPWR_c_535_n 6.09718e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_79_204#_M1004_g N_VPWR_c_535_n 0.0102886f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_79_204#_M1012_g N_VPWR_c_535_n 0.0103003f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_79_204#_M1015_g N_VPWR_c_535_n 6.11735e-19 $X=1.76 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_79_204#_M1012_g N_VPWR_c_536_n 6.18318e-19 $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_79_204#_M1015_g N_VPWR_c_536_n 0.0118732f $X=1.76 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_79_204#_c_172_p N_VPWR_c_536_n 0.00741008f $X=2.185 $Y=1.185 $X2=0
+ $Y2=0
cc_156 N_A_79_204#_c_113_n N_VPWR_c_536_n 0.00218651f $X=2.367 $Y=1.87 $X2=0
+ $Y2=0
cc_157 N_A_79_204#_c_114_n N_VPWR_c_536_n 0.0120391f $X=2.455 $Y=1.955 $X2=0
+ $Y2=0
cc_158 N_A_79_204#_c_108_n N_VPWR_c_536_n 0.00433518f $X=2.17 $Y=1.185 $X2=0
+ $Y2=0
cc_159 N_A_79_204#_M1012_g N_VPWR_c_539_n 0.00486043f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_79_204#_M1015_g N_VPWR_c_539_n 0.00486043f $X=1.76 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_79_204#_M1000_g N_VPWR_c_541_n 0.0046653f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_79_204#_M1004_g N_VPWR_c_541_n 0.00486043f $X=0.9 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_79_204#_c_114_n N_VPWR_c_542_n 7.41891e-19 $X=2.455 $Y=1.955 $X2=0
+ $Y2=0
cc_164 N_A_79_204#_M1008_s N_VPWR_c_532_n 0.00224864f $X=3.205 $Y=1.485 $X2=0
+ $Y2=0
cc_165 N_A_79_204#_M1000_g N_VPWR_c_532_n 0.00791817f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_79_204#_M1004_g N_VPWR_c_532_n 0.00822531f $X=0.9 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_79_204#_M1012_g N_VPWR_c_532_n 0.00822531f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_79_204#_M1015_g N_VPWR_c_532_n 0.00822531f $X=1.76 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_79_204#_c_114_n N_VPWR_c_532_n 0.0014742f $X=2.455 $Y=1.955 $X2=0
+ $Y2=0
cc_170 N_A_79_204#_M1003_g N_X_c_638_n 0.017146f $X=0.865 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A_79_204#_c_172_p N_X_c_638_n 0.0301455f $X=2.185 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A_79_204#_c_108_n N_X_c_638_n 0.0109112f $X=2.17 $Y=1.185 $X2=0 $Y2=0
cc_173 N_A_79_204#_M1000_g N_X_c_646_n 0.0184451f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_79_204#_c_172_p N_X_c_646_n 0.00326148f $X=2.185 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A_79_204#_M1004_g N_X_c_648_n 0.0153878f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_79_204#_M1012_g N_X_c_648_n 0.0150066f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_79_204#_c_172_p N_X_c_648_n 0.0556757f $X=2.185 $Y=1.185 $X2=0 $Y2=0
cc_178 N_A_79_204#_c_108_n N_X_c_648_n 0.00500468f $X=2.17 $Y=1.185 $X2=0 $Y2=0
cc_179 N_A_79_204#_M1011_g N_X_c_652_n 0.0148918f $X=1.295 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A_79_204#_M1013_g N_X_c_652_n 0.0143581f $X=1.725 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_79_204#_M1022_g N_X_c_652_n 0.00208147f $X=2.17 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_79_204#_c_172_p N_X_c_652_n 0.0558478f $X=2.185 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A_79_204#_c_106_n N_X_c_652_n 0.00550154f $X=2.282 $Y=1.045 $X2=0 $Y2=0
cc_184 N_A_79_204#_c_201_p N_X_c_652_n 0.0166066f $X=2.37 $Y=0.71 $X2=0 $Y2=0
cc_185 N_A_79_204#_c_108_n N_X_c_652_n 0.00522281f $X=2.17 $Y=1.185 $X2=0 $Y2=0
cc_186 N_A_79_204#_c_172_p N_X_c_659_n 0.0142514f $X=2.185 $Y=1.185 $X2=0 $Y2=0
cc_187 N_A_79_204#_c_108_n N_X_c_659_n 0.00240082f $X=2.17 $Y=1.185 $X2=0 $Y2=0
cc_188 N_A_79_204#_c_172_p N_X_c_661_n 0.0143339f $X=2.185 $Y=1.185 $X2=0 $Y2=0
cc_189 N_A_79_204#_c_108_n N_X_c_661_n 0.00253191f $X=2.17 $Y=1.185 $X2=0 $Y2=0
cc_190 N_A_79_204#_M1003_g X 0.0038525f $X=0.865 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_79_204#_c_172_p X 0.021458f $X=2.185 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A_79_204#_c_108_n X 0.0167247f $X=2.17 $Y=1.185 $X2=0 $Y2=0
cc_193 N_A_79_204#_c_113_n N_A_473_297#_M1023_d 0.00301386f $X=2.367 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_194 N_A_79_204#_c_114_n N_A_473_297#_M1023_d 0.00164948f $X=2.455 $Y=1.955
+ $X2=-0.19 $Y2=-0.24
cc_195 N_A_79_204#_c_122_p N_A_473_297#_M1023_d 0.00285768f $X=3.345 $Y=1.955
+ $X2=-0.19 $Y2=-0.24
cc_196 N_A_79_204#_c_116_n N_A_473_297#_M1023_d 0.00579173f $X=2.32 $Y=1.675
+ $X2=-0.19 $Y2=-0.24
cc_197 N_A_79_204#_M1008_s N_A_473_297#_c_696_n 0.00336985f $X=3.205 $Y=1.485
+ $X2=0 $Y2=0
cc_198 N_A_79_204#_c_114_n N_A_473_297#_c_696_n 0.0107845f $X=2.455 $Y=1.955
+ $X2=0 $Y2=0
cc_199 N_A_79_204#_c_122_p N_A_473_297#_c_696_n 0.0535599f $X=3.345 $Y=1.955
+ $X2=0 $Y2=0
cc_200 N_A_79_204#_c_122_p A_555_297# 0.00348375f $X=3.345 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_201 N_A_79_204#_c_106_n N_VGND_M1022_s 9.13545e-19 $X=2.282 $Y=1.045 $X2=0
+ $Y2=0
cc_202 N_A_79_204#_c_120_p N_VGND_M1022_s 0.00464239f $X=2.725 $Y=0.71 $X2=0
+ $Y2=0
cc_203 N_A_79_204#_c_201_p N_VGND_M1022_s 7.2107e-19 $X=2.37 $Y=0.71 $X2=0 $Y2=0
cc_204 N_A_79_204#_c_147_p N_VGND_M1002_s 0.00431889f $X=3.64 $Y=0.71 $X2=0
+ $Y2=0
cc_205 N_A_79_204#_c_140_p N_VGND_M1017_s 0.0146538f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_206 N_A_79_204#_M1003_g N_VGND_c_771_n 0.00752096f $X=0.865 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_79_204#_M1011_g N_VGND_c_771_n 5.0423e-19 $X=1.295 $Y=0.56 $X2=0
+ $Y2=0
cc_208 N_A_79_204#_M1003_g N_VGND_c_772_n 4.98572e-19 $X=0.865 $Y=0.56 $X2=0
+ $Y2=0
cc_209 N_A_79_204#_M1011_g N_VGND_c_772_n 0.00625485f $X=1.295 $Y=0.56 $X2=0
+ $Y2=0
cc_210 N_A_79_204#_M1013_g N_VGND_c_772_n 0.00629587f $X=1.725 $Y=0.56 $X2=0
+ $Y2=0
cc_211 N_A_79_204#_M1022_g N_VGND_c_772_n 4.94948e-19 $X=2.17 $Y=0.56 $X2=0
+ $Y2=0
cc_212 N_A_79_204#_M1013_g N_VGND_c_773_n 5.023e-19 $X=1.725 $Y=0.56 $X2=0 $Y2=0
cc_213 N_A_79_204#_M1022_g N_VGND_c_773_n 0.00639155f $X=2.17 $Y=0.56 $X2=0
+ $Y2=0
cc_214 N_A_79_204#_c_120_p N_VGND_c_773_n 0.00950629f $X=2.725 $Y=0.71 $X2=0
+ $Y2=0
cc_215 N_A_79_204#_c_201_p N_VGND_c_773_n 0.00753832f $X=2.37 $Y=0.71 $X2=0
+ $Y2=0
cc_216 N_A_79_204#_c_147_p N_VGND_c_774_n 0.0174773f $X=3.64 $Y=0.71 $X2=0 $Y2=0
cc_217 N_A_79_204#_c_140_p N_VGND_c_776_n 0.00600822f $X=5.16 $Y=0.71 $X2=0
+ $Y2=0
cc_218 N_A_79_204#_c_153_p N_VGND_c_776_n 0.0101237f $X=5.325 $Y=0.36 $X2=0
+ $Y2=0
cc_219 N_A_79_204#_M1003_g N_VGND_c_777_n 0.00353537f $X=0.865 $Y=0.56 $X2=0
+ $Y2=0
cc_220 N_A_79_204#_M1011_g N_VGND_c_777_n 0.00351072f $X=1.295 $Y=0.56 $X2=0
+ $Y2=0
cc_221 N_A_79_204#_M1013_g N_VGND_c_779_n 0.00351072f $X=1.725 $Y=0.56 $X2=0
+ $Y2=0
cc_222 N_A_79_204#_M1022_g N_VGND_c_779_n 0.00459896f $X=2.17 $Y=0.56 $X2=0
+ $Y2=0
cc_223 N_A_79_204#_c_201_p N_VGND_c_779_n 4.60047e-19 $X=2.37 $Y=0.71 $X2=0
+ $Y2=0
cc_224 N_A_79_204#_c_120_p N_VGND_c_781_n 0.00260553f $X=2.725 $Y=0.71 $X2=0
+ $Y2=0
cc_225 N_A_79_204#_c_242_p N_VGND_c_781_n 0.0155765f $X=2.82 $Y=0.485 $X2=0
+ $Y2=0
cc_226 N_A_79_204#_c_147_p N_VGND_c_781_n 0.00270984f $X=3.64 $Y=0.71 $X2=0
+ $Y2=0
cc_227 N_A_79_204#_c_147_p N_VGND_c_784_n 0.00278633f $X=3.64 $Y=0.71 $X2=0
+ $Y2=0
cc_228 N_A_79_204#_c_140_p N_VGND_c_784_n 0.00278969f $X=5.16 $Y=0.71 $X2=0
+ $Y2=0
cc_229 N_A_79_204#_c_139_p N_VGND_c_784_n 0.0227297f $X=3.835 $Y=0.38 $X2=0
+ $Y2=0
cc_230 N_A_79_204#_c_140_p N_VGND_c_785_n 0.00944283f $X=5.16 $Y=0.71 $X2=0
+ $Y2=0
cc_231 N_A_79_204#_c_153_p N_VGND_c_785_n 0.0165645f $X=5.325 $Y=0.36 $X2=0
+ $Y2=0
cc_232 N_A_79_204#_c_140_p N_VGND_c_787_n 0.0241284f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_233 N_A_79_204#_M1014_d N_VGND_c_788_n 0.00280564f $X=2.68 $Y=0.235 $X2=0
+ $Y2=0
cc_234 N_A_79_204#_M1007_d N_VGND_c_788_n 0.00309226f $X=3.635 $Y=0.235 $X2=0
+ $Y2=0
cc_235 N_A_79_204#_M1018_s N_VGND_c_788_n 0.00224096f $X=5.185 $Y=0.235 $X2=0
+ $Y2=0
cc_236 N_A_79_204#_M1003_g N_VGND_c_788_n 0.00411309f $X=0.865 $Y=0.56 $X2=0
+ $Y2=0
cc_237 N_A_79_204#_M1011_g N_VGND_c_788_n 0.0040731f $X=1.295 $Y=0.56 $X2=0
+ $Y2=0
cc_238 N_A_79_204#_M1013_g N_VGND_c_788_n 0.00411174f $X=1.725 $Y=0.56 $X2=0
+ $Y2=0
cc_239 N_A_79_204#_M1022_g N_VGND_c_788_n 0.00739987f $X=2.17 $Y=0.56 $X2=0
+ $Y2=0
cc_240 N_A_79_204#_c_120_p N_VGND_c_788_n 0.00515062f $X=2.725 $Y=0.71 $X2=0
+ $Y2=0
cc_241 N_A_79_204#_c_201_p N_VGND_c_788_n 0.00144425f $X=2.37 $Y=0.71 $X2=0
+ $Y2=0
cc_242 N_A_79_204#_c_242_p N_VGND_c_788_n 0.00930702f $X=2.82 $Y=0.485 $X2=0
+ $Y2=0
cc_243 N_A_79_204#_c_147_p N_VGND_c_788_n 0.00986322f $X=3.64 $Y=0.71 $X2=0
+ $Y2=0
cc_244 N_A_79_204#_c_140_p N_VGND_c_788_n 0.0217274f $X=5.16 $Y=0.71 $X2=0 $Y2=0
cc_245 N_A_79_204#_c_153_p N_VGND_c_788_n 0.01206f $X=5.325 $Y=0.36 $X2=0 $Y2=0
cc_246 N_A_79_204#_c_139_p N_VGND_c_788_n 0.0144776f $X=3.835 $Y=0.38 $X2=0
+ $Y2=0
cc_247 N_A_79_204#_c_140_p A_951_47# 0.00890637f $X=5.16 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_248 N_B1_M1014_g N_C1_c_359_n 0.0208517f $X=2.605 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_249 N_B1_c_266_n N_C1_c_359_n 8.60781e-19 $X=2.625 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_250 N_B1_M1023_g N_C1_M1008_g 0.058562f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B1_c_266_n N_C1_M1008_g 0.00171189f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B1_c_278_n N_C1_M1008_g 0.0137268f $X=3.845 $Y=1.572 $X2=0 $Y2=0
cc_253 N_B1_M1023_g N_C1_c_360_n 2.71034e-19 $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_254 N_B1_M1010_g N_C1_c_360_n 0.0495622f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B1_c_266_n N_C1_c_360_n 0.00174844f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_c_267_n N_C1_c_360_n 0.0215453f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B1_c_268_n N_C1_c_360_n 0.0235655f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B1_c_269_n N_C1_c_360_n 0.00308208f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B1_c_270_n N_C1_c_360_n 0.0165826f $X=4.01 $Y=0.985 $X2=0 $Y2=0
cc_260 N_B1_c_278_n N_C1_c_360_n 0.00414722f $X=3.845 $Y=1.572 $X2=0 $Y2=0
cc_261 N_B1_c_278_n N_C1_M1020_g 0.0155119f $X=3.845 $Y=1.572 $X2=0 $Y2=0
cc_262 N_B1_c_266_n C1 0.0251634f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B1_c_267_n C1 9.12379e-19 $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B1_c_268_n C1 0.0017833f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_265 N_B1_c_269_n C1 0.0214727f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_266 N_B1_c_278_n C1 0.0504207f $X=3.845 $Y=1.572 $X2=0 $Y2=0
cc_267 N_B1_c_270_n N_A2_M1005_g 0.0210266f $X=4.01 $Y=0.985 $X2=0 $Y2=0
cc_268 B1 N_A2_c_403_n 0.00335513f $X=3.83 $Y=1.445 $X2=0 $Y2=0
cc_269 N_B1_c_268_n N_A2_c_403_n 0.00133301f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B1_c_269_n N_A2_c_403_n 0.0195747f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B1_M1010_g N_A2_c_404_n 0.0270294f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B1_c_268_n N_A2_c_404_n 0.0119984f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B1_c_269_n N_A2_c_404_n 0.00200466f $X=4.01 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B1_M1010_g N_A2_c_428_n 2.19015e-19 $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_275 B1 N_A2_c_428_n 0.0101827f $X=3.83 $Y=1.445 $X2=0 $Y2=0
cc_276 B1 N_A2_c_414_n 0.00140553f $X=3.83 $Y=1.445 $X2=0 $Y2=0
cc_277 N_B1_M1023_g N_VPWR_c_536_n 0.00603533f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B1_M1010_g N_VPWR_c_537_n 9.23139e-19 $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B1_M1023_g N_VPWR_c_542_n 0.00357877f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B1_M1010_g N_VPWR_c_542_n 0.00357877f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B1_M1023_g N_VPWR_c_532_n 0.00660494f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_282 N_B1_M1010_g N_VPWR_c_532_n 0.00567005f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_283 B1 N_A_473_297#_M1010_d 0.00272324f $X=3.83 $Y=1.445 $X2=0 $Y2=0
cc_284 N_B1_M1023_g N_A_473_297#_c_696_n 0.00986058f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_285 N_B1_M1010_g N_A_473_297#_c_696_n 0.0119193f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_286 B1 N_A_473_297#_c_696_n 0.00674978f $X=3.83 $Y=1.445 $X2=0 $Y2=0
cc_287 N_B1_c_278_n N_A_473_297#_c_696_n 0.00889077f $X=3.845 $Y=1.572 $X2=0
+ $Y2=0
cc_288 B1 N_A_473_297#_c_712_n 0.00111423f $X=3.83 $Y=1.445 $X2=0 $Y2=0
cc_289 N_B1_c_278_n A_555_297# 0.00179116f $X=3.845 $Y=1.572 $X2=-0.19 $Y2=-0.24
cc_290 B1 A_727_297# 9.96181e-19 $X=3.83 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_291 N_B1_c_278_n A_727_297# 0.00281364f $X=3.845 $Y=1.572 $X2=-0.19 $Y2=-0.24
cc_292 N_B1_M1014_g N_VGND_c_773_n 0.0063832f $X=2.605 $Y=0.56 $X2=0 $Y2=0
cc_293 N_B1_M1014_g N_VGND_c_774_n 5.16106e-19 $X=2.605 $Y=0.56 $X2=0 $Y2=0
cc_294 N_B1_M1014_g N_VGND_c_781_n 0.00351072f $X=2.605 $Y=0.56 $X2=0 $Y2=0
cc_295 N_B1_c_270_n N_VGND_c_784_n 0.00422112f $X=4.01 $Y=0.985 $X2=0 $Y2=0
cc_296 N_B1_c_270_n N_VGND_c_787_n 0.00336173f $X=4.01 $Y=0.985 $X2=0 $Y2=0
cc_297 N_B1_M1014_g N_VGND_c_788_n 0.00424039f $X=2.605 $Y=0.56 $X2=0 $Y2=0
cc_298 N_B1_c_270_n N_VGND_c_788_n 0.00619761f $X=4.01 $Y=0.985 $X2=0 $Y2=0
cc_299 N_C1_M1008_g N_VPWR_c_542_n 0.00357877f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_300 N_C1_M1020_g N_VPWR_c_542_n 0.00357877f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_301 N_C1_M1008_g N_VPWR_c_532_n 0.00534514f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_302 N_C1_M1020_g N_VPWR_c_532_n 0.00544245f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_303 N_C1_M1008_g N_A_473_297#_c_696_n 0.0129288f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_304 N_C1_M1020_g N_A_473_297#_c_696_n 0.0147139f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_305 N_C1_c_359_n N_VGND_c_773_n 5.35333e-19 $X=3.075 $Y=0.99 $X2=0 $Y2=0
cc_306 N_C1_c_359_n N_VGND_c_774_n 0.0055489f $X=3.075 $Y=0.99 $X2=0 $Y2=0
cc_307 N_C1_c_360_n N_VGND_c_774_n 0.0031831f $X=3.56 $Y=0.99 $X2=0 $Y2=0
cc_308 N_C1_c_359_n N_VGND_c_781_n 0.00393283f $X=3.075 $Y=0.99 $X2=0 $Y2=0
cc_309 N_C1_c_360_n N_VGND_c_784_n 0.00422112f $X=3.56 $Y=0.99 $X2=0 $Y2=0
cc_310 N_C1_c_359_n N_VGND_c_788_n 0.00466354f $X=3.075 $Y=0.99 $X2=0 $Y2=0
cc_311 N_C1_c_360_n N_VGND_c_788_n 0.00604366f $X=3.56 $Y=0.99 $X2=0 $Y2=0
cc_312 N_A2_M1005_g N_A1_M1018_g 0.042588f $X=4.68 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A2_c_403_n N_A1_M1016_g 0.00256389f $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A2_c_433_p N_A1_M1016_g 0.011925f $X=5.635 $Y=1.605 $X2=0 $Y2=0
cc_315 N_A2_c_414_n N_A1_M1016_g 0.0311662f $X=4.66 $Y=1.4 $X2=0 $Y2=0
cc_316 N_A2_c_407_n N_A1_M1019_g 0.0316679f $X=6.06 $Y=1.01 $X2=0 $Y2=0
cc_317 N_A2_M1009_g N_A1_M1021_g 0.0316679f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A2_c_433_p N_A1_M1021_g 0.0154705f $X=5.635 $Y=1.605 $X2=0 $Y2=0
cc_319 N_A2_c_403_n A1 0.0196691f $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A2_c_404_n A1 0.00107409f $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A2_c_433_p A1 0.0220708f $X=5.635 $Y=1.605 $X2=0 $Y2=0
cc_322 N_A2_c_405_n A1 0.018457f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A2_c_406_n A1 2.00143e-19 $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_324 A2 A1 5.10986e-19 $X=5.67 $Y=1.445 $X2=0 $Y2=0
cc_325 N_A2_c_403_n N_A1_c_486_n 8.75327e-19 $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A2_c_404_n N_A1_c_486_n 0.0241698f $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A2_c_433_p N_A1_c_486_n 0.0022867f $X=5.635 $Y=1.605 $X2=0 $Y2=0
cc_328 N_A2_c_405_n N_A1_c_486_n 0.00354268f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A2_c_406_n N_A1_c_486_n 0.0316679f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_330 A2 N_A1_c_486_n 0.00427033f $X=5.67 $Y=1.445 $X2=0 $Y2=0
cc_331 N_A2_c_403_n N_VPWR_M1001_d 3.10304e-19 $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A2_c_433_p N_VPWR_M1001_d 0.00773396f $X=5.635 $Y=1.605 $X2=0 $Y2=0
cc_333 N_A2_c_428_n N_VPWR_M1001_d 0.00138647f $X=4.825 $Y=1.605 $X2=0 $Y2=0
cc_334 N_A2_c_453_p N_VPWR_M1021_s 0.00228437f $X=5.74 $Y=1.51 $X2=0 $Y2=0
cc_335 N_A2_c_414_n N_VPWR_c_537_n 0.007566f $X=4.66 $Y=1.4 $X2=0 $Y2=0
cc_336 N_A2_M1009_g N_VPWR_c_538_n 0.00785369f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A2_c_414_n N_VPWR_c_542_n 0.00351072f $X=4.66 $Y=1.4 $X2=0 $Y2=0
cc_338 N_A2_M1009_g N_VPWR_c_544_n 0.00351042f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A2_M1009_g N_VPWR_c_532_n 0.00500047f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_340 N_A2_c_414_n N_VPWR_c_532_n 0.00439456f $X=4.66 $Y=1.4 $X2=0 $Y2=0
cc_341 N_A2_c_433_p N_A_473_297#_M1016_d 0.00416797f $X=5.635 $Y=1.605 $X2=0
+ $Y2=0
cc_342 N_A2_c_404_n N_A_473_297#_c_716_n 5.85636e-19 $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A2_c_433_p N_A_473_297#_c_716_n 0.0192404f $X=5.635 $Y=1.605 $X2=0
+ $Y2=0
cc_344 N_A2_c_428_n N_A_473_297#_c_716_n 0.0207817f $X=4.825 $Y=1.605 $X2=0
+ $Y2=0
cc_345 N_A2_c_414_n N_A_473_297#_c_716_n 0.0132115f $X=4.66 $Y=1.4 $X2=0 $Y2=0
cc_346 N_A2_c_414_n N_A_473_297#_c_720_n 5.22362e-19 $X=4.66 $Y=1.4 $X2=0 $Y2=0
cc_347 N_A2_M1009_g N_A_473_297#_c_721_n 0.0106958f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A2_c_433_p N_A_473_297#_c_721_n 0.0100092f $X=5.635 $Y=1.605 $X2=0
+ $Y2=0
cc_349 N_A2_c_405_n N_A_473_297#_c_721_n 0.0041785f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_350 N_A2_c_453_p N_A_473_297#_c_721_n 0.0125989f $X=5.74 $Y=1.51 $X2=0 $Y2=0
cc_351 N_A2_M1009_g N_A_473_297#_c_697_n 0.00659641f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A2_c_405_n N_A_473_297#_c_697_n 0.0120152f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A2_c_406_n N_A_473_297#_c_697_n 0.00406248f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A2_c_433_p N_A_473_297#_c_728_n 0.0146911f $X=5.635 $Y=1.605 $X2=0
+ $Y2=0
cc_355 N_A2_M1009_g N_A_473_297#_c_699_n 0.00578728f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A2_c_405_n N_VGND_c_776_n 0.0120411f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_357 N_A2_c_406_n N_VGND_c_776_n 0.00396828f $X=6.06 $Y=1.16 $X2=0 $Y2=0
cc_358 N_A2_c_407_n N_VGND_c_776_n 0.0165734f $X=6.06 $Y=1.01 $X2=0 $Y2=0
cc_359 N_A2_M1005_g N_VGND_c_785_n 0.00422112f $X=4.68 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A2_c_407_n N_VGND_c_785_n 0.0046653f $X=6.06 $Y=1.01 $X2=0 $Y2=0
cc_361 N_A2_M1005_g N_VGND_c_787_n 0.0044652f $X=4.68 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A2_M1005_g N_VGND_c_788_n 0.00613204f $X=4.68 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A2_c_407_n N_VGND_c_788_n 0.00802136f $X=6.06 $Y=1.01 $X2=0 $Y2=0
cc_364 N_A1_M1016_g N_VPWR_c_537_n 0.00350443f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_365 N_A1_M1016_g N_VPWR_c_538_n 4.87602e-19 $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A1_M1021_g N_VPWR_c_538_n 0.00646256f $X=5.54 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A1_M1016_g N_VPWR_c_543_n 0.0041289f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A1_M1021_g N_VPWR_c_543_n 0.00351072f $X=5.54 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A1_M1016_g N_VPWR_c_532_n 0.00598322f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_370 N_A1_M1021_g N_VPWR_c_532_n 0.0040731f $X=5.54 $Y=1.985 $X2=0 $Y2=0
cc_371 N_A1_M1016_g N_A_473_297#_c_716_n 0.0104909f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_372 N_A1_M1016_g N_A_473_297#_c_720_n 0.00561143f $X=5.11 $Y=1.985 $X2=0
+ $Y2=0
cc_373 N_A1_M1021_g N_A_473_297#_c_721_n 0.0136689f $X=5.54 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A1_M1021_g N_A_473_297#_c_697_n 0.00100796f $X=5.54 $Y=1.985 $X2=0
+ $Y2=0
cc_375 N_A1_M1016_g N_A_473_297#_c_728_n 0.00357313f $X=5.11 $Y=1.985 $X2=0
+ $Y2=0
cc_376 N_A1_M1019_g N_VGND_c_776_n 0.0027958f $X=5.54 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A1_M1018_g N_VGND_c_785_n 0.00413555f $X=5.11 $Y=0.56 $X2=0 $Y2=0
cc_378 N_A1_M1019_g N_VGND_c_785_n 0.00549615f $X=5.54 $Y=0.56 $X2=0 $Y2=0
cc_379 N_A1_M1018_g N_VGND_c_788_n 0.00576772f $X=5.11 $Y=0.56 $X2=0 $Y2=0
cc_380 N_A1_M1019_g N_VGND_c_788_n 0.00996598f $X=5.54 $Y=0.56 $X2=0 $Y2=0
cc_381 N_VPWR_c_532_n N_X_M1000_s 0.0055303f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_532_n N_X_M1012_s 0.00535672f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_534_n N_X_c_646_n 0.00219958f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_384 N_VPWR_M1000_d N_X_c_641_n 0.00317633f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_385 N_VPWR_c_534_n N_X_c_641_n 0.0224255f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_386 N_VPWR_c_541_n N_X_c_671_n 0.0122764f $X=0.95 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_532_n N_X_c_671_n 0.00704765f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_M1004_d N_X_c_648_n 0.00331972f $X=0.975 $Y=1.485 $X2=0 $Y2=0
cc_389 N_VPWR_c_535_n N_X_c_648_n 0.0173266f $X=1.115 $Y=1.96 $X2=0 $Y2=0
cc_390 N_VPWR_c_539_n N_X_c_675_n 0.0124538f $X=1.81 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_c_532_n N_X_c_675_n 0.00724021f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_c_532_n N_A_473_297#_M1023_d 0.00209344f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_393 N_VPWR_c_532_n N_A_473_297#_M1010_d 0.00325886f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_532_n N_A_473_297#_M1016_d 0.0023722f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_532_n N_A_473_297#_M1009_s 0.00223246f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_536_n N_A_473_297#_c_696_n 0.0159069f $X=1.97 $Y=2 $X2=0 $Y2=0
cc_397 N_VPWR_c_542_n N_A_473_297#_c_696_n 0.103728f $X=4.62 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_c_532_n N_A_473_297#_c_696_n 0.0647613f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_399 N_VPWR_M1001_d N_A_473_297#_c_716_n 0.00625586f $X=4.645 $Y=1.485 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_537_n N_A_473_297#_c_716_n 0.0207638f $X=4.785 $Y=2.36 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_542_n N_A_473_297#_c_716_n 0.00262823f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_543_n N_A_473_297#_c_716_n 0.00327411f $X=5.59 $Y=2.72 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_532_n N_A_473_297#_c_716_n 0.0114067f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_537_n N_A_473_297#_c_720_n 0.0123205f $X=4.785 $Y=2.36 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_543_n N_A_473_297#_c_720_n 0.0155449f $X=5.59 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_532_n N_A_473_297#_c_720_n 0.00971527f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_M1021_s N_A_473_297#_c_721_n 0.00352893f $X=5.615 $Y=1.485 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_538_n N_A_473_297#_c_721_n 0.0162045f $X=5.755 $Y=2.36 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_543_n N_A_473_297#_c_721_n 0.00263536f $X=5.59 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_544_n N_A_473_297#_c_721_n 0.00164049f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_532_n N_A_473_297#_c_721_n 0.00815182f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_544_n N_A_473_297#_c_698_n 0.0174615f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_532_n N_A_473_297#_c_698_n 0.00974347f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_542_n N_A_473_297#_c_712_n 0.0210413f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_532_n N_A_473_297#_c_712_n 0.0125824f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_544_n N_A_473_297#_c_699_n 0.00100665f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_532_n N_A_473_297#_c_699_n 0.00205685f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_532_n A_555_297# 0.00224864f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_419 N_VPWR_c_532_n A_727_297# 0.00256987f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_420 N_X_c_638_n N_VGND_M1003_s 0.00497736f $X=0.985 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_421 N_X_c_652_n N_VGND_M1011_s 0.00326709f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_422 N_X_c_638_n N_VGND_c_771_n 0.0211043f $X=0.985 $Y=0.755 $X2=0 $Y2=0
cc_423 N_X_c_652_n N_VGND_c_772_n 0.0163619f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_424 N_X_c_681_p N_VGND_c_773_n 0.0126877f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_425 N_X_c_638_n N_VGND_c_777_n 0.00252074f $X=0.985 $Y=0.755 $X2=0 $Y2=0
cc_426 N_X_c_683_p N_VGND_c_777_n 0.0123751f $X=1.08 $Y=0.42 $X2=0 $Y2=0
cc_427 N_X_c_652_n N_VGND_c_777_n 0.00265538f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_428 N_X_c_652_n N_VGND_c_779_n 0.00265538f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_429 N_X_c_681_p N_VGND_c_779_n 0.0120547f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_430 N_X_c_638_n N_VGND_c_783_n 0.00269748f $X=0.985 $Y=0.755 $X2=0 $Y2=0
cc_431 N_X_c_640_n N_VGND_c_783_n 0.00517761f $X=0.212 $Y=0.875 $X2=0 $Y2=0
cc_432 N_X_M1003_d N_VGND_c_788_n 0.00252469f $X=0.94 $Y=0.235 $X2=0 $Y2=0
cc_433 N_X_M1013_d N_VGND_c_788_n 0.00492275f $X=1.8 $Y=0.235 $X2=0 $Y2=0
cc_434 N_X_c_638_n N_VGND_c_788_n 0.00993411f $X=0.985 $Y=0.755 $X2=0 $Y2=0
cc_435 N_X_c_683_p N_VGND_c_788_n 0.00722272f $X=1.08 $Y=0.42 $X2=0 $Y2=0
cc_436 N_X_c_652_n N_VGND_c_788_n 0.0102135f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_437 N_X_c_681_p N_VGND_c_788_n 0.00683853f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_438 N_X_c_640_n N_VGND_c_788_n 0.00767249f $X=0.212 $Y=0.875 $X2=0 $Y2=0
cc_439 N_A_473_297#_c_696_n A_555_297# 0.00336985f $X=4.12 $Y=2.337 $X2=-0.19
+ $Y2=1.305
cc_440 N_A_473_297#_c_696_n A_727_297# 0.0057713f $X=4.12 $Y=2.337 $X2=-0.19
+ $Y2=1.305
cc_441 N_VGND_c_788_n A_951_47# 0.00318969f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_442 N_VGND_c_788_n A_1123_47# 0.0119688f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24

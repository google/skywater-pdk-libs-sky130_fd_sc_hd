* File: sky130_fd_sc_hd__o41a_1.spice
* Created: Tue Sep  1 19:26:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o41a_1.pex.spice"
.subckt sky130_fd_sc_hd__o41a_1  VNB VPB B1 A4 A3 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_103_21#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.247 PD=1.82 PS=2.06 NRD=0 NRS=21.228 M=1 R=4.33333 SA=75000.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_321_47#_M1004_d N_B1_M1004_g N_A_103_21#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A4_M1007_g N_A_321_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.08775 PD=1.03 PS=0.92 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_321_47#_M1005_d N_A3_M1005_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.1235 PD=1.04 PS=1.03 NRD=9.228 NRS=9.228 M=1 R=4.33333
+ SA=75001.1 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_321_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.12675 PD=1.04 PS=1.04 NRD=10.152 NRS=11.076 M=1 R=4.33333
+ SA=75001.7 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1003 N_A_321_47#_M1003_d N_A1_M1003_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.195 AS=0.12675 PD=1.9 PS=1.04 NRD=2.76 NRS=10.152 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_103_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.425 PD=1.27 PS=2.85 NRD=0 NRS=27.5603 M=1 R=6.66667 SA=75000.3
+ SB=75003 A=0.15 P=2.3 MULT=1
MM1000 N_A_103_21#_M1000_d N_B1_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=1.52 PS=1.27 NRD=14.775 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1008 A_393_297# N_A4_M1008_g N_A_103_21#_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.22 AS=0.26 PD=1.44 PS=1.52 NRD=32.4853 NRS=32.4853 M=1 R=6.66667
+ SA=75001.4 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1001 A_511_297# N_A3_M1001_g A_393_297# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.22 PD=1.39 PS=1.44 NRD=27.5603 NRS=32.4853 M=1 R=6.66667 SA=75002
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1006 A_619_297# N_A2_M1006_g A_511_297# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.195 PD=1.39 PS=1.39 NRD=27.5603 NRS=27.5603 M=1 R=6.66667 SA=75002.6
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_619_297# VPB PHIGHVT L=0.15 W=1 AD=0.28
+ AS=0.195 PD=2.56 PS=1.39 NRD=0 NRS=27.5603 M=1 R=6.66667 SA=75003.1 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_37 VNB 0 1.81202e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__o41a_1.pxi.spice"
*
.ends
*
*

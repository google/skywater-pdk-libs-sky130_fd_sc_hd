* File: sky130_fd_sc_hd__clkdlybuf4s50_1.spice
* Created: Thu Aug 27 14:12:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkdlybuf4s50_1.pex.spice"
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819196 AS=0.1134 PD=0.792897 PS=1.38 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_A_283_47#_M1001_d N_A_27_47#_M1001_g N_VGND_M1002_d VNB NSHORT L=0.5
+ W=0.65 AD=0.169 AS=0.12678 PD=1.82 PS=1.2271 NRD=0 NRS=4.608 M=1 R=1.3
+ SA=250000 SB=250000 A=0.325 P=2.3 MULT=1
MM1006 N_VGND_M1006_d N_A_283_47#_M1006_g N_A_390_47#_M1006_s VNB NSHORT L=0.5
+ W=0.65 AD=0.11785 AS=0.17225 PD=1.18458 PS=1.83 NRD=0 NRS=0 M=1 R=1.3
+ SA=250000 SB=250000 A=0.325 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_390_47#_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1491 AS=0.0761495 PD=1.55 PS=0.765421 NRD=4.284 NRS=12.852 M=1 R=2.8
+ SA=75001 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_47#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.186923 AS=0.27 PD=1.49451 PS=2.54 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1005 N_A_283_47#_M1005_d N_A_27_47#_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.5
+ W=0.82 AD=0.2173 AS=0.153277 PD=2.17 PS=1.22549 NRD=0 NRS=2.3837 M=1 R=1.64
+ SA=250001 SB=250000 A=0.41 P=2.64 MULT=1
MM1004 N_VPWR_M1004_d N_A_283_47#_M1004_g N_A_390_47#_M1004_s VPB PHIGHVT L=0.5
+ W=0.82 AD=0.140346 AS=0.2173 PD=1.19396 PS=2.17 NRD=0 NRS=0 M=1 R=1.64
+ SA=250000 SB=250001 A=0.41 P=2.64 MULT=1
MM1007 N_X_M1007_d N_A_390_47#_M1007_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.355 AS=0.171154 PD=2.71 PS=1.45604 NRD=2.9353 NRS=8.8453 M=1 R=6.66667
+ SA=75000.9 SB=75000.3 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_58 VPB 0 7.48979e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__clkdlybuf4s50_1.pxi.spice"
*
.ends
*
*

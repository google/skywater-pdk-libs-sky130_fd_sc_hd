* File: sky130_fd_sc_hd__dfrbp_2.pex.spice
* Created: Tue Sep  1 19:02:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFRBP_2%CLK 1 2 3 5 6 8 11 13 14
c40 6 0 9.23148e-20 $X=0.47 $Y=1.74
c41 1 0 2.71124e-20 $X=0.305 $Y=1.325
r42 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=1.16
+ $X2=0.265 $Y2=1.53
r43 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r44 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r47 3 18 88.7086 $w=2.58e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r50 1 18 39.2009 $w=2.58e-07 $l=1.75656e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.327 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_27_47# 1 2 9 13 17 20 21 22 25 27 29 33 37
+ 41 42 43 46 49 50 51 52 55 61 68 71 72 77
c236 77 0 4.56546e-20 $X=6.07 $Y=1.11
c237 61 0 1.76704e-20 $X=6.11 $Y=1.19
c238 51 0 1.58851e-19 $X=5.965 $Y=1.19
c239 29 0 4.11863e-20 $X=5.845 $Y=2.275
c240 22 0 1.90473e-19 $X=2.72 $Y=1.32
r241 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=1.11 $X2=6.07 $Y2=1.11
r242 71 74 47.4498 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=1.095
r243 71 73 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=0.765
r244 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=0.93 $X2=2.585 $Y2=0.93
r245 65 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r246 61 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.19
+ $X2=6.11 $Y2=1.19
r247 59 72 8.56101 $w=3.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.56 $Y=1.19
+ $X2=2.56 $Y2=0.93
r248 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r249 55 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r250 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.19
+ $X2=0.695 $Y2=1.19
r251 52 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.19
+ $X2=2.53 $Y2=1.19
r252 51 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=6.11 $Y2=1.19
r253 51 52 4.07177 $w=1.4e-07 $l=3.29e-06 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=2.675 $Y2=1.19
r254 50 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.19
+ $X2=0.695 $Y2=1.19
r255 49 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r256 49 50 1.91213 $w=1.4e-07 $l=1.545e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.84 $Y2=1.19
r257 48 55 30.3143 $w=2.28e-07 $l=6.05e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.19
r258 47 55 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.19
r259 44 46 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r260 43 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.795
r261 43 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r262 41 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r263 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r264 35 42 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.345 $Y2=0.72
r265 35 37 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.51
r266 31 76 38.5991 $w=2.92e-07 $l=1.76125e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=5.987 $Y2=1.11
r267 31 33 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=6.01 $Y2=0.415
r268 27 76 58.4073 $w=2.92e-07 $l=3.48848e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.987 $Y2=1.11
r269 27 29 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.845 $Y2=2.275
r270 23 25 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.18 $Y=1.395
+ $X2=3.18 $Y2=2.275
r271 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=3.18 $Y2=1.395
r272 21 22 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=2.72 $Y2=1.32
r273 20 22 26.9401 $w=1.5e-07 $l=1.09243e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.72 $Y2=1.32
r274 20 74 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.642 $Y2=1.095
r275 17 73 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.64 $Y=0.415
+ $X2=2.64 $Y2=0.765
r276 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r277 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r278 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r279 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r280 2 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r281 1 37 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%D 3 7 9 10 15 19
c53 10 0 1.85993e-19 $X=2.09 $Y=1.3
c54 7 0 1.77283e-19 $X=2.225 $Y=2.275
r55 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.465 $X2=1.79 $Y2=1.465
r56 15 19 1.96287 $w=4.04e-07 $l=6.5e-08 $layer=LI1_cond $X=1.615 $Y=1.53
+ $X2=1.615 $Y2=1.465
r57 9 18 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.09 $Y=1.465 $X2=1.79
+ $Y2=1.465
r58 9 10 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.465
+ $X2=2.09 $Y2=1.3
r59 5 10 37.0704 $w=1.5e-07 $l=3.91727e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.09 $Y2=1.3
r60 5 7 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.225 $Y2=2.275
r61 1 10 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.165 $Y=1.3 $X2=2.09
+ $Y2=1.3
r62 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.165 $Y=1.3
+ $X2=2.165 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_193_47# 1 2 9 13 15 17 20 23 26 27 29 30
+ 34 35 37 38 39 40 47 49 53 65 66 70
c212 66 0 3.94709e-20 $X=6.265 $Y=1.74
c213 47 0 1.77283e-19 $X=2.99 $Y=1.87
c214 39 0 1.36782e-20 $X=5.965 $Y=1.87
c215 38 0 9.23148e-20 $X=1.245 $Y=1.87
c216 37 0 1.20979e-19 $X=2.845 $Y=1.87
c217 35 0 1.61046e-19 $X=3.095 $Y=0.9
c218 29 0 1.76704e-20 $X=5.97 $Y=1.58
c219 26 0 1.28114e-19 $X=5.59 $Y=0.87
r220 65 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.74
+ $X2=6.265 $Y2=1.905
r221 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.265
+ $Y=1.74 $X2=6.265 $Y2=1.74
r222 53 56 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.695 $Y=1.74
+ $X2=2.695 $Y2=1.875
r223 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.74 $X2=2.695 $Y2=1.74
r224 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.87
+ $X2=6.11 $Y2=1.87
r225 47 54 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=1.77
+ $X2=2.695 $Y2=1.77
r226 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.87
+ $X2=2.99 $Y2=1.87
r227 43 70 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.1 $Y=1.87
+ $X2=1.1 $Y2=0.51
r228 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=1.87 $X2=1.1
+ $Y2=1.87
r229 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.87
+ $X2=2.99 $Y2=1.87
r230 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=6.11 $Y2=1.87
r231 39 40 3.50247 $w=1.4e-07 $l=2.83e-06 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=3.135 $Y2=1.87
r232 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=1.87
+ $X2=1.1 $Y2=1.87
r233 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=2.99 $Y2=1.87
r234 37 38 1.98019 $w=1.4e-07 $l=1.6e-06 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=1.245 $Y2=1.87
r235 35 58 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.095 $Y=0.9
+ $X2=3.095 $Y2=0.765
r236 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=0.9 $X2=3.095 $Y2=0.9
r237 31 34 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.875
+ $X2=3.095 $Y2=0.875
r238 29 66 5.43733 $w=3.59e-07 $l=2.995e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=6.2 $Y2=1.74
r239 29 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=5.675 $Y2=1.58
r240 27 60 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.59 $Y=0.87
+ $X2=5.465 $Y2=0.87
r241 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=0.87 $X2=5.59 $Y2=0.87
r242 24 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.675 $Y2=1.58
r243 24 26 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.57 $Y2=0.87
r244 23 47 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.99 $Y=1.575
+ $X2=2.99 $Y2=1.77
r245 22 31 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=0.875
r246 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=1.575
r247 20 68 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.275 $Y=2.275
+ $X2=6.275 $Y2=1.905
r248 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.87
r249 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.415
r250 13 58 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.12 $Y=0.415
+ $X2=3.12 $Y2=0.765
r251 9 56 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.685 $Y=2.275
+ $X2=2.685 $Y2=1.875
r252 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r253 1 70 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_761_289# 1 2 9 13 15 18 21 23 25 26 27 30
+ 33 36 37
c109 36 0 1.00332e-19 $X=5.145 $Y=0.835
c110 23 0 4.11863e-20 $X=5.19 $Y=1.525
r111 33 35 3.58511 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.36
+ $X2=5.19 $Y2=0.445
r112 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.58 $Y=2.005
+ $X2=5.58 $Y2=2.3
r113 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.58 $Y2=2.005
r114 26 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.275 $Y2=1.92
r115 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.19 $Y=1.835
+ $X2=5.275 $Y2=1.92
r116 24 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.61
r117 24 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.835
r118 23 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=1.61
r119 23 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=0.835
r120 21 36 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.835
r121 21 35 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.445
r122 18 40 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.775
r123 18 39 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.445
r124 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.61 $X2=3.94 $Y2=1.61
r125 15 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=5.19 $Y2=1.61
r126 15 17 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=3.94 $Y2=1.61
r127 13 39 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.95 $Y=0.445
+ $X2=3.95 $Y2=1.445
r128 9 40 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.88 $Y=2.275 $X2=3.88
+ $Y2=1.775
r129 2 30 600 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.645 $X2=5.58 $Y2=2.3
r130 1 33 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.2 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%RESET_B 3 6 10 14 16 17 20 23 25 26 27 29 37
+ 39 42 57
c153 37 0 1.00332e-19 $X=4.37 $Y=0.93
c154 29 0 4.83118e-21 $X=7.19 $Y=1.165
c155 23 0 6.10372e-20 $X=4.25 $Y=0.85
c156 14 0 1.03533e-19 $X=7.235 $Y=2.275
c157 10 0 4.70414e-20 $X=7.235 $Y=0.445
r158 49 57 3.2703 $w=2.4e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=1.035
+ $X2=7.525 $Y2=1.22
r159 42 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=1.285
r160 42 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=0.955
r161 37 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=1.095
r162 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=0.765
r163 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.27
+ $Y=1.12 $X2=7.27 $Y2=1.12
r164 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.19 $Y=1.165
+ $X2=7.19 $Y2=1.165
r165 27 34 0.181159 $w=2.07e-07 $l=3e-07 $layer=MET1_cond $X=7.19 $Y=0.85
+ $X2=7.49 $Y2=0.85
r166 27 29 0.0979621 $w=2.9e-07 $l=2e-07 $layer=MET1_cond $X=7.19 $Y=0.965
+ $X2=7.19 $Y2=1.165
r167 25 27 0.10072 $w=2.07e-07 $l=1.45e-07 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=7.19 $Y2=0.85
r168 25 26 3.2797 $w=1.4e-07 $l=2.65e-06 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=4.395 $Y2=0.85
r169 23 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=0.93 $X2=4.37 $Y2=0.93
r170 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.25 $Y=0.85
+ $X2=4.25 $Y2=0.85
r171 20 26 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.395 $Y2=0.85
r172 20 22 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.25 $Y2=0.85
r173 17 57 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.49 $Y=1.22
+ $X2=7.525 $Y2=1.22
r174 17 30 9.34413 $w=3.68e-07 $l=3e-07 $layer=LI1_cond $X=7.49 $Y=1.22 $X2=7.19
+ $Y2=1.22
r175 16 49 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=0.85
+ $X2=7.525 $Y2=1.035
r176 16 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.49 $Y=0.85
+ $X2=7.49 $Y2=0.85
r177 14 45 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=7.235 $Y=2.275
+ $X2=7.235 $Y2=1.285
r178 10 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.235 $Y=0.445
+ $X2=7.235 $Y2=0.955
r179 6 40 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=4.365 $Y=2.275
+ $X2=4.365 $Y2=1.095
r180 3 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.31 $Y=0.445
+ $X2=4.31 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_543_47# 1 2 9 11 13 15 16 20 25 27 28 29
+ 34 35
c126 35 0 6.10372e-20 $X=4.85 $Y=1.17
c127 29 0 1.61046e-19 $X=3.6 $Y=1.27
c128 11 0 1.36782e-20 $X=5.275 $Y=1.495
c129 9 0 1.28114e-19 $X=4.97 $Y=0.555
r130 34 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.85 $Y=1.17 $X2=4.85
+ $Y2=1.27
r131 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.17 $X2=4.85 $Y2=1.17
r132 30 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.33 $Y=1.27
+ $X2=3.515 $Y2=1.27
r133 29 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.27
+ $X2=3.515 $Y2=1.27
r134 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=4.85 $Y2=1.27
r135 28 29 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=3.6 $Y2=1.27
r136 27 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=1.185
+ $X2=3.515 $Y2=1.27
r137 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.515 $Y=0.475
+ $X2=3.515 $Y2=1.185
r138 24 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=1.27
r139 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=2.135
r140 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=3.515 $Y2=0.475
r141 20 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=2.91 $Y2=0.39
r142 16 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=3.33 $Y2=2.135
r143 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=2.9 $Y2=2.3
r144 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.35 $Y=1.57
+ $X2=5.35 $Y2=2.065
r145 12 35 61.4314 $w=2.55e-07 $l=3.99061e-07 $layer=POLY_cond $X=5.045 $Y=1.495
+ $X2=4.88 $Y2=1.17
r146 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.35 $Y2=1.57
r147 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.045 $Y2=1.495
r148 7 35 39.2931 $w=2.55e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.88 $Y2=1.17
r149 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.97 $Y2=0.555
r150 2 18 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.065 $X2=2.9 $Y2=2.33
r151 1 22 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.91 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_1283_21# 1 2 9 13 17 21 23 24 25 27 30 32
+ 34 37 40 44 48 49 50 53 55 56 57 58 60 61 63 68 75
c200 75 0 6.15427e-20 $X=6.695 $Y=0.98
c201 68 0 1.94811e-19 $X=7.15 $Y=0.78
c202 40 0 6.54241e-20 $X=9.575 $Y=1.16
c203 13 0 2.35828e-20 $X=6.695 $Y=2.275
r204 72 73 6.79936 $w=3.14e-07 $l=1.75e-07 $layer=LI1_cond $X=7.9 $Y=1.16
+ $X2=8.075 $Y2=1.16
r205 64 79 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=8.485 $Y=1.16
+ $X2=8.63 $Y2=1.16
r206 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.485
+ $Y=1.16 $X2=8.485 $Y2=1.16
r207 61 73 3.84416 $w=3.14e-07 $l=1.03078e-07 $layer=LI1_cond $X=8.16 $Y=1.2
+ $X2=8.075 $Y2=1.16
r208 61 63 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=8.16 $Y=1.2
+ $X2=8.485 $Y2=1.2
r209 59 73 4.32966 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=1.325
+ $X2=8.075 $Y2=1.16
r210 59 60 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.075 $Y=1.325
+ $X2=8.075 $Y2=1.915
r211 58 72 4.32966 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.9 $Y=0.995
+ $X2=7.9 $Y2=1.16
r212 57 71 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.465 $X2=7.9
+ $Y2=0.38
r213 57 58 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.9 $Y=0.465
+ $X2=7.9 $Y2=0.995
r214 55 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.99 $Y=2
+ $X2=8.075 $Y2=1.915
r215 55 56 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.99 $Y=2 $X2=7.53
+ $Y2=2
r216 51 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.53 $Y2=2
r217 51 53 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.445 $Y2=2.21
r218 49 71 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.9 $Y2=0.38
r219 49 50 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.235 $Y2=0.38
r220 48 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=0.695
+ $X2=7.15 $Y2=0.78
r221 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.235 $Y2=0.38
r222 47 48 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.15 $Y2=0.695
r223 45 75 17.8171 $w=2.57e-07 $l=9.5e-08 $layer=POLY_cond $X=6.79 $Y=0.98
+ $X2=6.695 $Y2=0.98
r224 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=0.98 $X2=6.79 $Y2=0.98
r225 42 68 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=0.78
+ $X2=7.15 $Y2=0.78
r226 42 44 6.02413 $w=2.18e-07 $l=1.15e-07 $layer=LI1_cond $X=6.815 $Y=0.865
+ $X2=6.815 $Y2=0.98
r227 39 40 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=9.115 $Y=1.16
+ $X2=9.575 $Y2=1.16
r228 35 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.575 $Y=1.325
+ $X2=9.575 $Y2=1.16
r229 35 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.575 $Y=1.325
+ $X2=9.575 $Y2=1.985
r230 32 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.575 $Y=0.995
+ $X2=9.575 $Y2=1.16
r231 32 34 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.575 $Y=0.995
+ $X2=9.575 $Y2=0.56
r232 28 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=1.325
+ $X2=9.115 $Y2=1.16
r233 28 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.115 $Y=1.325
+ $X2=9.115 $Y2=1.985
r234 25 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=0.995
+ $X2=9.115 $Y2=1.16
r235 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.115 $Y=0.995
+ $X2=9.115 $Y2=0.56
r236 24 79 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.705 $Y=1.16
+ $X2=8.63 $Y2=1.16
r237 23 39 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.04 $Y=1.16
+ $X2=9.115 $Y2=1.16
r238 23 24 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=9.04 $Y=1.16
+ $X2=8.705 $Y2=1.16
r239 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.325
+ $X2=8.63 $Y2=1.16
r240 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=8.63 $Y=1.325
+ $X2=8.63 $Y2=2.125
r241 15 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=0.995
+ $X2=8.63 $Y2=1.16
r242 15 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.63 $Y=0.995
+ $X2=8.63 $Y2=0.445
r243 11 75 15.359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=0.98
r244 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=2.275
r245 7 75 38.4475 $w=2.57e-07 $l=2.75409e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.695 $Y2=0.98
r246 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.49 $Y2=0.445
r247 2 53 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=2.065 $X2=7.445 $Y2=2.21
r248 1 71 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=7.765
+ $Y=0.235 $X2=7.9 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_1108_47# 1 2 9 13 15 19 24 25 26 29 30
c103 25 0 2.04429e-20 $X=6.685 $Y=1.745
c104 24 0 1.60161e-19 $X=6.45 $Y=1.315
c105 19 0 1.03533e-19 $X=6.6 $Y=2.295
c106 15 0 4.70414e-20 $X=6.365 $Y=0.395
c107 13 0 1.79199e-19 $X=7.69 $Y=0.445
r108 30 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.66
+ $X2=7.655 $Y2=1.495
r109 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.655
+ $Y=1.66 $X2=7.655 $Y2=1.66
r110 27 32 3.26844 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.77 $Y=1.66 $X2=6.6
+ $Y2=1.66
r111 27 29 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.77 $Y=1.66
+ $X2=7.655 $Y2=1.66
r112 25 32 5.45986 $w=2.62e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.6 $Y2=1.66
r113 25 26 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.685 $Y2=2.125
r114 24 32 17.5667 $w=2.62e-07 $l=4.13249e-07 $layer=LI1_cond $X=6.45 $Y=1.315
+ $X2=6.6 $Y2=1.66
r115 23 24 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.45 $Y=0.535
+ $X2=6.45 $Y2=1.315
r116 19 26 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.685 $Y2=2.125
r117 19 21 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.065 $Y2=2.295
r118 15 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=6.45 $Y2=0.535
r119 15 17 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=5.75 $Y2=0.395
r120 13 34 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=7.69 $Y=0.445
+ $X2=7.69 $Y2=1.495
r121 7 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=1.66
r122 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=2.275
r123 2 21 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=2.065 $X2=6.065 $Y2=2.335
r124 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.54
+ $Y=0.235 $X2=5.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_1659_47# 1 2 7 9 12 14 16 19 23 27 29 30
+ 32 33 36 38 39 43 48
c117 48 0 1.91378e-19 $X=10.415 $Y=1.16
r118 44 48 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=9.995 $Y=1.16
+ $X2=10.415 $Y2=1.16
r119 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.995
+ $Y=1.16 $X2=9.995 $Y2=1.16
r120 40 43 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=9.75 $Y=1.16
+ $X2=9.995 $Y2=1.16
r121 35 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.75 $Y=1.325
+ $X2=9.75 $Y2=1.16
r122 35 36 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=9.75 $Y=1.325
+ $X2=9.75 $Y2=1.865
r123 34 39 4.40882 $w=2.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=8.99 $Y=1.95
+ $X2=8.905 $Y2=1.915
r124 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.665 $Y=1.95
+ $X2=9.75 $Y2=1.865
r125 33 34 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=9.665 $Y=1.95
+ $X2=8.99 $Y2=1.95
r126 32 39 2.0246 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=8.905 $Y=1.795
+ $X2=8.905 $Y2=1.915
r127 31 32 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=8.905 $Y=0.885
+ $X2=8.905 $Y2=1.795
r128 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.82 $Y=0.8
+ $X2=8.905 $Y2=0.885
r129 29 30 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.82 $Y=0.8
+ $X2=8.585 $Y2=0.8
r130 28 38 3.31033 $w=2.4e-07 $l=1.13e-07 $layer=LI1_cond $X=8.56 $Y=1.915
+ $X2=8.447 $Y2=1.915
r131 27 39 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=1.915
+ $X2=8.905 $Y2=1.915
r132 27 28 12.4848 $w=2.38e-07 $l=2.6e-07 $layer=LI1_cond $X=8.82 $Y=1.915
+ $X2=8.56 $Y2=1.915
r133 21 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.46 $Y=0.715
+ $X2=8.585 $Y2=0.8
r134 21 23 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=8.46 $Y=0.715
+ $X2=8.46 $Y2=0.51
r135 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.415 $Y=1.325
+ $X2=10.415 $Y2=1.16
r136 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.415 $Y=1.325
+ $X2=10.415 $Y2=1.985
r137 14 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.415 $Y=0.995
+ $X2=10.415 $Y2=1.16
r138 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.415 $Y=0.995
+ $X2=10.415 $Y2=0.56
r139 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.995 $Y=1.325
+ $X2=9.995 $Y2=1.16
r140 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.995 $Y=1.325
+ $X2=9.995 $Y2=1.985
r141 7 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.995 $Y=0.995
+ $X2=9.995 $Y2=1.16
r142 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.995 $Y=0.995
+ $X2=9.995 $Y2=0.56
r143 2 38 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=1.805 $X2=8.42 $Y2=1.96
r144 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.235 $X2=8.42 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 58 62 67 68 70 71 73 74 76 77 78 79 80 81 83 88 97 108 121 123 126 129 132
r187 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r188 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r189 126 127 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r190 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r191 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r192 118 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r193 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r194 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r195 115 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r196 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r197 112 132 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.07 $Y=2.72
+ $X2=8.9 $Y2=2.72
r198 112 114 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.07 $Y=2.72
+ $X2=9.43 $Y2=2.72
r199 111 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r200 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r201 108 132 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.73 $Y=2.72
+ $X2=8.9 $Y2=2.72
r202 108 110 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.73 $Y=2.72
+ $X2=8.51 $Y2=2.72
r203 107 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r204 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r205 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r206 104 130 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.29 $Y2=2.72
r207 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r208 101 129 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.14 $Y2=2.72
r209 101 103 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=6.67 $Y2=2.72
r210 100 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r211 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r212 97 129 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=5.14 $Y2=2.72
r213 97 99 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=4.83 $Y2=2.72
r214 96 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r215 96 127 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.07 $Y2=2.72
r216 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r217 93 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=1.975 $Y2=2.72
r218 93 95 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=3.91 $Y2=2.72
r219 92 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r220 92 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r221 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r222 89 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r223 89 91 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r224 88 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.975 $Y2=2.72
r225 88 91 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r226 83 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r227 83 85 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r228 81 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r229 81 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r230 79 117 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.59 $Y=2.72
+ $X2=10.35 $Y2=2.72
r231 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.59 $Y=2.72
+ $X2=10.675 $Y2=2.72
r232 78 120 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=10.76 $Y=2.72
+ $X2=10.81 $Y2=2.72
r233 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.76 $Y=2.72
+ $X2=10.675 $Y2=2.72
r234 76 114 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.43 $Y2=2.72
r235 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.785 $Y2=2.72
r236 75 117 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.95 $Y=2.72
+ $X2=10.35 $Y2=2.72
r237 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.95 $Y=2.72
+ $X2=9.785 $Y2=2.72
r238 73 106 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.59 $Y2=2.72
r239 73 74 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.882 $Y2=2.72
r240 72 110 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=8.055 $Y=2.72
+ $X2=8.51 $Y2=2.72
r241 72 74 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=8.055 $Y=2.72
+ $X2=7.882 $Y2=2.72
r242 70 103 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=6.67 $Y2=2.72
r243 70 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=7.065 $Y2=2.72
r244 69 106 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.19 $Y=2.72
+ $X2=7.59 $Y2=2.72
r245 69 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.19 $Y=2.72
+ $X2=7.065 $Y2=2.72
r246 67 95 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.99 $Y=2.72 $X2=3.91
+ $Y2=2.72
r247 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=2.72
+ $X2=4.155 $Y2=2.72
r248 66 99 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.83 $Y2=2.72
r249 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.155 $Y2=2.72
r250 62 65 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=10.675 $Y=1.66
+ $X2=10.675 $Y2=2.34
r251 60 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.675 $Y=2.635
+ $X2=10.675 $Y2=2.72
r252 60 65 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.675 $Y=2.635
+ $X2=10.675 $Y2=2.34
r253 56 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.785 $Y=2.635
+ $X2=9.785 $Y2=2.72
r254 56 58 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.785 $Y=2.635
+ $X2=9.785 $Y2=2.34
r255 52 132 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=2.635
+ $X2=8.9 $Y2=2.72
r256 52 54 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=8.9 $Y=2.635
+ $X2=8.9 $Y2=2.29
r257 48 74 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=7.882 $Y=2.635
+ $X2=7.882 $Y2=2.72
r258 48 50 9.85422 $w=3.43e-07 $l=2.95e-07 $layer=LI1_cond $X=7.882 $Y=2.635
+ $X2=7.882 $Y2=2.34
r259 44 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.72
r260 44 46 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.34
r261 40 129 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.72
r262 40 42 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.34
r263 36 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.72
r264 36 38 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.29
r265 32 126 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.72
r266 32 34 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.34
r267 28 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r268 28 30 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r269 9 65 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=10.49
+ $Y=1.485 $X2=10.675 $Y2=2.34
r270 9 62 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=10.49
+ $Y=1.485 $X2=10.675 $Y2=1.66
r271 8 58 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.485 $X2=9.785 $Y2=2.34
r272 7 54 600 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.805 $X2=8.905 $Y2=2.29
r273 6 50 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=2.065 $X2=7.875 $Y2=2.34
r274 5 46 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=2.065 $X2=7.025 $Y2=2.34
r275 4 42 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=1.645 $X2=5.14 $Y2=2.34
r276 3 38 600 $w=1.7e-07 $l=3.09233e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=2.065 $X2=4.155 $Y2=2.29
r277 2 34 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=2.065 $X2=2.015 $Y2=2.34
r278 1 30 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_448_47# 1 2 8 9 11
c34 8 0 6.94938e-20 $X=2.13 $Y=1.835
r35 9 11 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.215 $Y=0.39
+ $X2=2.375 $Y2=0.39
r36 8 14 22.5629 $w=2.72e-07 $l=5.35635e-07 $layer=LI1_cond $X=2.13 $Y=1.835
+ $X2=2.282 $Y2=2.3
r37 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.215 $Y2=0.39
r38 7 8 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.13 $Y2=1.835
r39 2 14 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.065 $X2=2.435 $Y2=2.3
r40 1 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.375 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%A_651_413# 1 2 9 11 12 15
c36 12 0 1.58851e-19 $X=3.755 $Y=1.95
r37 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.035
+ $X2=4.575 $Y2=2.21
r38 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=4.575 $Y2=2.035
r39 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=3.755 $Y2=1.95
r40 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.755 $Y2=1.95
r41 7 9 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.67 $Y2=2.21
r42 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=2.065 $X2=4.575 $Y2=2.21
r43 1 9 600 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=2.065 $X2=3.67 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%Q 1 2 7 10
r19 7 15 15.6526 $w=3.33e-07 $l=4.55e-07 $layer=LI1_cond $X=9.327 $Y=1.155
+ $X2=9.327 $Y2=1.61
r20 7 10 18.0607 $w=3.33e-07 $l=5.25e-07 $layer=LI1_cond $X=9.327 $Y=1.155
+ $X2=9.327 $Y2=0.63
r21 2 15 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.485 $X2=9.325 $Y2=1.61
r22 1 10 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=9.19
+ $Y=0.235 $X2=9.325 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%Q_N 1 2 9 13 18 21 25
c31 21 0 6.54241e-20 $X=10.275 $Y=1.11
r32 21 25 0.195722 $w=1.68e-07 $l=3e-09 $layer=LI1_cond $X=10.335 $Y=1.197
+ $X2=10.335 $Y2=1.2
r33 20 21 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=10.335 $Y=0.825
+ $X2=10.335 $Y2=1.197
r34 18 20 16.4563 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=10.23 $Y=0.4
+ $X2=10.23 $Y2=0.825
r35 14 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.335 $Y=1.535
+ $X2=10.335 $Y2=1.2
r36 13 15 14.2361 $w=3.88e-07 $l=4.6e-07 $layer=LI1_cond $X=10.225 $Y=1.62
+ $X2=10.225 $Y2=2.08
r37 13 14 6.24364 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=10.225 $Y=1.62
+ $X2=10.225 $Y2=1.535
r38 9 15 8.45125 $w=2.98e-07 $l=2.2e-07 $layer=LI1_cond $X=10.27 $Y=2.3
+ $X2=10.27 $Y2=2.08
r39 2 13 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=10.07
+ $Y=1.485 $X2=10.205 $Y2=1.62
r40 2 9 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=10.07
+ $Y=1.485 $X2=10.205 $Y2=2.3
r41 1 18 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=10.07
+ $Y=0.235 $X2=10.205 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DFRBP_2%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 46 50
+ 53 54 56 57 59 60 62 63 64 65 66 67 69 101 103 106
c162 101 0 2.71124e-20 $X=10.81 $Y=0
c163 46 0 1.91378e-19 $X=9.785 $Y=0.565
r164 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r165 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r166 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r167 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r168 98 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r169 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r170 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r171 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r172 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r173 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r174 89 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.51 $Y2=0
r175 88 91 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.13 $Y=0 $X2=8.51
+ $Y2=0
r176 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r177 86 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r178 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r179 83 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.67 $Y2=0
r180 82 85 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.67
+ $Y2=0
r181 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r182 80 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r183 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r184 77 80 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r185 77 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r186 76 79 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r187 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r188 74 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.71 $Y2=0
r189 74 76 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.07 $Y2=0
r190 69 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r191 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r192 67 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r193 67 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r194 65 97 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.59 $Y=0
+ $X2=10.35 $Y2=0
r195 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.59 $Y=0
+ $X2=10.675 $Y2=0
r196 64 100 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=10.76 $Y=0 $X2=10.81
+ $Y2=0
r197 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.76 $Y=0
+ $X2=10.675 $Y2=0
r198 62 94 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.7 $Y=0 $X2=9.43
+ $Y2=0
r199 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.7 $Y=0 $X2=9.785
+ $Y2=0
r200 61 97 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.87 $Y=0 $X2=10.35
+ $Y2=0
r201 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.87 $Y=0 $X2=9.785
+ $Y2=0
r202 59 91 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=8.755 $Y=0 $X2=8.51
+ $Y2=0
r203 59 60 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=8.872 $Y2=0
r204 58 94 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=8.99 $Y=0 $X2=9.43
+ $Y2=0
r205 58 60 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=8.99 $Y=0 $X2=8.872
+ $Y2=0
r206 56 85 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.67
+ $Y2=0
r207 56 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.8
+ $Y2=0
r208 55 88 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.895 $Y=0
+ $X2=7.13 $Y2=0
r209 55 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.895 $Y=0 $X2=6.8
+ $Y2=0
r210 53 79 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r211 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.64
+ $Y2=0
r212 52 82 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.83
+ $Y2=0
r213 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.64
+ $Y2=0
r214 48 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.675 $Y=0.085
+ $X2=10.675 $Y2=0
r215 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.675 $Y=0.085
+ $X2=10.675 $Y2=0.4
r216 44 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.785 $Y=0.085
+ $X2=9.785 $Y2=0
r217 44 46 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.785 $Y=0.085
+ $X2=9.785 $Y2=0.565
r218 40 60 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.872 $Y=0.085
+ $X2=8.872 $Y2=0
r219 40 42 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=8.872 $Y=0.085
+ $X2=8.872 $Y2=0.38
r220 36 57 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0
r221 36 38 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0.36
r222 32 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r223 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.38
r224 28 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r225 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.36
r226 27 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r227 26 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0
+ $X2=1.71 $Y2=0
r228 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=0.845
+ $Y2=0
r229 22 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r230 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r231 7 50 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=10.49
+ $Y=0.235 $X2=10.675 $Y2=0.4
r232 6 46 182 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_NDIFF $count=1 $X=9.65
+ $Y=0.235 $X2=9.785 $Y2=0.565
r233 5 42 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=8.705
+ $Y=0.235 $X2=8.905 $Y2=0.38
r234 4 38 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.81 $Y2=0.36
r235 3 34 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.64 $Y2=0.38
r236 2 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.71 $Y2=0.36
r237 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


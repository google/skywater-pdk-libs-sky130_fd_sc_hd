* File: sky130_fd_sc_hd__o41a_2.pxi.spice
* Created: Thu Aug 27 14:41:51 2020
* 
x_PM_SKY130_FD_SC_HD__O41A_2%A_79_21# N_A_79_21#_M1002_s N_A_79_21#_M1005_d
+ N_A_79_21#_c_74_n N_A_79_21#_M1004_g N_A_79_21#_M1001_g N_A_79_21#_c_75_n
+ N_A_79_21#_M1012_g N_A_79_21#_M1008_g N_A_79_21#_c_76_n N_A_79_21#_c_77_n
+ N_A_79_21#_c_78_n N_A_79_21#_c_87_n N_A_79_21#_c_79_n N_A_79_21#_c_80_n
+ N_A_79_21#_c_90_p N_A_79_21#_c_81_n N_A_79_21#_c_92_p N_A_79_21#_c_82_n
+ PM_SKY130_FD_SC_HD__O41A_2%A_79_21#
x_PM_SKY130_FD_SC_HD__O41A_2%B1 N_B1_M1005_g N_B1_M1002_g B1 N_B1_c_151_n
+ PM_SKY130_FD_SC_HD__O41A_2%B1
x_PM_SKY130_FD_SC_HD__O41A_2%A4 N_A4_M1003_g N_A4_M1006_g A4 A4 N_A4_c_185_n
+ N_A4_c_186_n PM_SKY130_FD_SC_HD__O41A_2%A4
x_PM_SKY130_FD_SC_HD__O41A_2%A3 N_A3_M1013_g N_A3_M1007_g A3 A3 A3 A3
+ N_A3_c_219_n N_A3_c_220_n PM_SKY130_FD_SC_HD__O41A_2%A3
x_PM_SKY130_FD_SC_HD__O41A_2%A2 N_A2_M1010_g N_A2_M1011_g A2 A2 A2 A2
+ N_A2_c_253_n N_A2_c_254_n PM_SKY130_FD_SC_HD__O41A_2%A2
x_PM_SKY130_FD_SC_HD__O41A_2%A1 N_A1_M1009_g N_A1_M1000_g A1 N_A1_c_284_n
+ N_A1_c_285_n PM_SKY130_FD_SC_HD__O41A_2%A1
x_PM_SKY130_FD_SC_HD__O41A_2%VPWR N_VPWR_M1001_d N_VPWR_M1008_d N_VPWR_M1000_d
+ N_VPWR_c_308_n N_VPWR_c_309_n N_VPWR_c_320_n N_VPWR_c_310_n N_VPWR_c_311_n
+ N_VPWR_c_312_n N_VPWR_c_325_n VPWR N_VPWR_c_313_n N_VPWR_c_314_n
+ N_VPWR_c_315_n N_VPWR_c_307_n PM_SKY130_FD_SC_HD__O41A_2%VPWR
x_PM_SKY130_FD_SC_HD__O41A_2%X N_X_M1004_s N_X_M1001_s X X X X X X N_X_c_376_n X
+ X PM_SKY130_FD_SC_HD__O41A_2%X
x_PM_SKY130_FD_SC_HD__O41A_2%VGND N_VGND_M1004_d N_VGND_M1012_d N_VGND_M1003_d
+ N_VGND_M1010_d N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n
+ N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n VGND N_VGND_c_399_n
+ N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n
+ PM_SKY130_FD_SC_HD__O41A_2%VGND
x_PM_SKY130_FD_SC_HD__O41A_2%A_393_47# N_A_393_47#_M1002_d N_A_393_47#_M1013_d
+ N_A_393_47#_M1009_d N_A_393_47#_c_485_n N_A_393_47#_c_457_n
+ N_A_393_47#_c_458_n N_A_393_47#_c_468_n N_A_393_47#_c_459_n
+ N_A_393_47#_c_481_n N_A_393_47#_c_460_n PM_SKY130_FD_SC_HD__O41A_2%A_393_47#
cc_1 VNB N_A_79_21#_c_74_n 0.0199911f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.975
cc_2 VNB N_A_79_21#_c_75_n 0.0186136f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.975
cc_3 VNB N_A_79_21#_c_76_n 0.0424984f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.16
cc_4 VNB N_A_79_21#_c_77_n 0.00212527f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.2
cc_5 VNB N_A_79_21#_c_78_n 0.0326683f $X=-0.19 $Y=-0.24 $X2=1.13 $Y2=1.16
cc_6 VNB N_A_79_21#_c_79_n 0.00442673f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=0.38
cc_7 VNB N_A_79_21#_c_80_n 0.00368914f $X=-0.19 $Y=-0.24 $X2=1.515 $Y2=1.075
cc_8 VNB N_A_79_21#_c_81_n 0.00284214f $X=-0.19 $Y=-0.24 $X2=1.477 $Y2=1.2
cc_9 VNB N_A_79_21#_c_82_n 0.00166933f $X=-0.19 $Y=-0.24 $X2=1.607 $Y2=0.85
cc_10 VNB N_B1_M1005_g 5.93976e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B1_M1002_g 0.0222485f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.975
cc_12 VNB B1 0.00191567f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_B1_c_151_n 0.0433676f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_14 VNB A4 0.00311333f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB N_A4_c_185_n 0.0209152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A4_c_186_n 0.017817f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_17 VNB A3 0.00316579f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_18 VNB N_A3_c_219_n 0.0201295f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.345
cc_19 VNB N_A3_c_220_n 0.0176886f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_20 VNB A2 0.00317005f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_A2_c_253_n 0.0201408f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.345
cc_22 VNB N_A2_c_254_n 0.0176531f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_23 VNB A1 0.0194553f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_24 VNB N_A1_c_284_n 0.0271106f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_25 VNB N_A1_c_285_n 0.0224181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_307_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB X 8.37336e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_28 VNB N_VGND_c_392_n 0.00991007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_393_n 0.0334157f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_30 VNB N_VGND_c_394_n 0.0118265f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_31 VNB N_VGND_c_395_n 0.00526389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_396_n 0.00529257f $X=-0.19 $Y=-0.24 $X2=1.13 $Y2=1.16
cc_33 VNB N_VGND_c_397_n 0.0191191f $X=-0.19 $Y=-0.24 $X2=1.477 $Y2=1.325
cc_34 VNB N_VGND_c_398_n 0.00516539f $X=-0.19 $Y=-0.24 $X2=1.477 $Y2=1.495
cc_35 VNB N_VGND_c_399_n 0.017949f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=0.38
cc_36 VNB N_VGND_c_400_n 0.0318226f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=2.34
cc_37 VNB N_VGND_c_401_n 0.0242032f $X=-0.19 $Y=-0.24 $X2=1.13 $Y2=1.16
cc_38 VNB N_VGND_c_402_n 0.249316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_403_n 0.00470919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_404_n 0.00506925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_393_47#_c_457_n 0.00753369f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.975
cc_42 VNB N_A_393_47#_c_458_n 0.00783996f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_43 VNB N_A_393_47#_c_459_n 0.0198057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_393_47#_c_460_n 0.00636986f $X=-0.19 $Y=-0.24 $X2=1.13 $Y2=1.2
cc_45 VPB N_A_79_21#_M1001_g 0.0237845f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_46 VPB N_A_79_21#_M1008_g 0.0204668f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_47 VPB N_A_79_21#_c_76_n 0.00817633f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.16
cc_48 VPB N_A_79_21#_c_77_n 0.00587975f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.2
cc_49 VPB N_A_79_21#_c_87_n 0.0017079f $X=-0.19 $Y=1.305 $X2=1.477 $Y2=1.495
cc_50 VPB N_B1_M1005_g 0.0253404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB B1 0.00400048f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_52 VPB N_A4_M1006_g 0.0209754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB A4 0.00367227f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_54 VPB N_A4_c_185_n 0.00539889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A3_M1007_g 0.0190642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB A3 0.00227681f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_57 VPB N_A3_c_219_n 0.00500477f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.345
cc_58 VPB N_A2_M1011_g 0.0190148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB A2 0.00298484f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_60 VPB N_A2_c_253_n 0.00501495f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.345
cc_61 VPB N_A1_M1000_g 0.0271105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB A1 0.00824277f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_63 VPB N_A1_c_284_n 0.0069113f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_64 VPB N_VPWR_c_308_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.345
cc_65 VPB N_VPWR_c_309_n 0.0429874f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_66 VPB N_VPWR_c_310_n 0.00599881f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.16
cc_67 VPB N_VPWR_c_311_n 0.0150617f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_68 VPB N_VPWR_c_312_n 0.00564356f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_69 VPB N_VPWR_c_313_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.607 $Y2=0.38
cc_70 VPB N_VPWR_c_314_n 0.0691779f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.665
cc_71 VPB N_VPWR_c_315_n 0.00977718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_307_n 0.0476553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB X 0.00124663f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_74 N_A_79_21#_c_76_n N_B1_M1005_g 0.00700016f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_87_n N_B1_M1005_g 0.00963407f $X=1.477 $Y=1.495 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_90_p N_B1_M1005_g 0.0106364f $X=1.86 $Y=2.34 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_81_n N_B1_M1005_g 8.71877e-19 $X=1.477 $Y=1.2 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_92_p N_B1_M1005_g 0.0133932f $X=1.86 $Y=1.66 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_80_n N_B1_M1002_g 0.0044451f $X=1.515 $Y=1.075 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_81_n B1 0.0196221f $X=1.477 $Y=1.2 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_92_p B1 0.0279534f $X=1.86 $Y=1.66 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_78_n N_B1_c_151_n 0.0123372f $X=1.13 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_80_n N_B1_c_151_n 0.00311908f $X=1.515 $Y=1.075 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_81_n N_B1_c_151_n 0.00634063f $X=1.477 $Y=1.2 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_92_p N_B1_c_151_n 0.00211696f $X=1.86 $Y=1.66 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_82_n N_B1_c_151_n 0.0055885f $X=1.607 $Y=0.85 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_90_p N_A4_M1006_g 0.00653397f $X=1.86 $Y=2.34 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_92_p N_A4_M1006_g 8.22166e-19 $X=1.86 $Y=1.66 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_87_n N_VPWR_M1008_d 6.5584e-19 $X=1.477 $Y=1.495 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_92_p N_VPWR_M1008_d 0.00416673f $X=1.86 $Y=1.66 $X2=0 $Y2=0
cc_91 N_A_79_21#_M1001_g N_VPWR_c_309_n 0.00321781f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_77_n N_VPWR_c_320_n 0.0140054f $X=1.355 $Y=1.2 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_78_n N_VPWR_c_320_n 0.00121344f $X=1.13 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_90_p N_VPWR_c_320_n 0.00544399f $X=1.86 $Y=2.34 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_92_p N_VPWR_c_320_n 0.0136682f $X=1.86 $Y=1.66 $X2=0 $Y2=0
cc_96 N_A_79_21#_M1008_g N_VPWR_c_310_n 0.00205456f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_77_n N_VPWR_c_325_n 0.00652797f $X=1.355 $Y=1.2 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_78_n N_VPWR_c_325_n 6.98043e-19 $X=1.13 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_92_p N_VPWR_c_325_n 0.013225f $X=1.86 $Y=1.66 $X2=0 $Y2=0
cc_100 N_A_79_21#_M1001_g N_VPWR_c_313_n 0.00541359f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_101 N_A_79_21#_M1008_g N_VPWR_c_313_n 0.00541359f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_c_90_p N_VPWR_c_314_n 0.029423f $X=1.86 $Y=2.34 $X2=0 $Y2=0
cc_103 N_A_79_21#_M1005_d N_VPWR_c_307_n 0.0111774f $X=1.725 $Y=1.485 $X2=0
+ $Y2=0
cc_104 N_A_79_21#_M1001_g N_VPWR_c_307_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_79_21#_M1008_g N_VPWR_c_307_n 0.0101559f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_90_p N_VPWR_c_307_n 0.0170482f $X=1.86 $Y=2.34 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_74_n X 0.00645876f $X=0.47 $Y=0.975 $X2=0 $Y2=0
cc_108 N_A_79_21#_M1001_g X 0.00762851f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_75_n X 0.00385583f $X=0.89 $Y=0.975 $X2=0 $Y2=0
cc_110 N_A_79_21#_M1008_g X 0.00188164f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_76_n X 0.0349909f $X=0.965 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_77_n X 0.0194431f $X=1.355 $Y=1.2 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_87_n X 0.00558057f $X=1.477 $Y=1.495 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_80_n X 0.00541929f $X=1.515 $Y=1.075 $X2=0 $Y2=0
cc_115 N_A_79_21#_M1001_g X 0.00907982f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_79_21#_M1008_g X 0.00905475f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_74_n N_X_c_376_n 0.00528656f $X=0.47 $Y=0.975 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_75_n N_X_c_376_n 0.00528656f $X=0.89 $Y=0.975 $X2=0 $Y2=0
cc_119 N_A_79_21#_M1001_g X 0.00181417f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_79_21#_M1008_g X 0.00256288f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_74_n N_VGND_c_393_n 0.00321781f $X=0.47 $Y=0.975 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_75_n N_VGND_c_394_n 0.00321006f $X=0.89 $Y=0.975 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_77_n N_VGND_c_394_n 0.0178766f $X=1.355 $Y=1.2 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_78_n N_VGND_c_394_n 0.00570552f $X=1.13 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_79_n N_VGND_c_394_n 0.0513585f $X=1.62 $Y=0.38 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_74_n N_VGND_c_399_n 0.00541359f $X=0.47 $Y=0.975 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_75_n N_VGND_c_399_n 0.00541359f $X=0.89 $Y=0.975 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_79_n N_VGND_c_400_n 0.0238974f $X=1.62 $Y=0.38 $X2=0 $Y2=0
cc_129 N_A_79_21#_M1002_s N_VGND_c_402_n 0.00362654f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_130 N_A_79_21#_c_74_n N_VGND_c_402_n 0.0104557f $X=0.47 $Y=0.975 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_75_n N_VGND_c_402_n 0.0108276f $X=0.89 $Y=0.975 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_79_n N_VGND_c_402_n 0.01357f $X=1.62 $Y=0.38 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_80_n N_A_393_47#_c_458_n 0.00160504f $X=1.515 $Y=1.075 $X2=0
+ $Y2=0
cc_134 N_B1_M1005_g A4 0.0025977f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_135 B1 A4 0.0209621f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_136 N_B1_c_151_n A4 6.44399e-19 $X=1.94 $Y=1.16 $X2=0 $Y2=0
cc_137 N_B1_M1005_g N_A4_c_185_n 0.0117069f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_138 B1 N_A4_c_185_n 8.69828e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_139 N_B1_c_151_n N_A4_c_185_n 0.0167261f $X=1.94 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B1_M1002_g N_A4_c_186_n 0.0102304f $X=1.89 $Y=0.56 $X2=0 $Y2=0
cc_141 N_B1_M1005_g N_VPWR_c_320_n 0.00168221f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B1_M1005_g N_VPWR_c_310_n 0.00345545f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B1_M1005_g N_VPWR_c_314_n 0.00541359f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B1_M1005_g N_VPWR_c_307_n 0.0108036f $X=1.65 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B1_M1002_g N_VGND_c_394_n 0.0027998f $X=1.89 $Y=0.56 $X2=0 $Y2=0
cc_146 N_B1_M1002_g N_VGND_c_400_n 0.00585385f $X=1.89 $Y=0.56 $X2=0 $Y2=0
cc_147 N_B1_M1002_g N_VGND_c_402_n 0.012229f $X=1.89 $Y=0.56 $X2=0 $Y2=0
cc_148 N_B1_M1002_g N_A_393_47#_c_458_n 2.76254e-19 $X=1.89 $Y=0.56 $X2=0 $Y2=0
cc_149 B1 N_A_393_47#_c_458_n 0.0142146f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_150 N_B1_c_151_n N_A_393_47#_c_458_n 0.00284579f $X=1.94 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A4_M1006_g N_A3_M1007_g 0.0438296f $X=2.405 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A4_M1006_g A3 9.64167e-19 $X=2.405 $Y=1.985 $X2=0 $Y2=0
cc_153 A4 A3 0.0683765f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A4_c_185_n A3 7.6629e-19 $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_155 A4 N_A3_c_219_n 0.00452322f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A4_c_185_n N_A3_c_219_n 0.0220385f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A4_c_186_n N_A3_c_220_n 0.0235877f $X=2.477 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A4_M1006_g N_VPWR_c_314_n 0.00382445f $X=2.405 $Y=1.985 $X2=0 $Y2=0
cc_159 A4 N_VPWR_c_314_n 0.0113375f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_160 N_A4_M1006_g N_VPWR_c_307_n 0.00626406f $X=2.405 $Y=1.985 $X2=0 $Y2=0
cc_161 A4 N_VPWR_c_307_n 0.0110525f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_162 A4 A_496_297# 0.00879686f $X=2.445 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_163 N_A4_c_186_n N_VGND_c_395_n 0.00320758f $X=2.477 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A4_c_186_n N_VGND_c_400_n 0.00436487f $X=2.477 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A4_c_186_n N_VGND_c_402_n 0.00621427f $X=2.477 $Y=0.995 $X2=0 $Y2=0
cc_166 A4 N_A_393_47#_c_457_n 0.0260031f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A4_c_185_n N_A_393_47#_c_457_n 0.0035815f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A4_c_186_n N_A_393_47#_c_457_n 0.0113124f $X=2.477 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A4_c_186_n N_A_393_47#_c_468_n 5.4344e-19 $X=2.477 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A3_M1007_g N_A2_M1011_g 0.0450937f $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A3_M1007_g A2 9.6479e-19 $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_172 A3 A2 0.0681759f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_173 N_A3_c_219_n A2 7.6636e-19 $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_174 A3 N_A2_c_253_n 0.00449056f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_175 N_A3_c_219_n N_A2_c_253_n 0.0220295f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A3_c_220_n N_A2_c_254_n 0.0184483f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A3_M1007_g N_VPWR_c_314_n 0.00382445f $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_178 A3 N_VPWR_c_314_n 0.0112468f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A3_M1007_g N_VPWR_c_307_n 0.00581096f $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_180 A3 N_VPWR_c_307_n 0.0110525f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_181 A3 A_597_297# 0.0087545f $X=2.905 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_182 N_A3_c_220_n N_VGND_c_395_n 0.00560851f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A3_c_220_n N_VGND_c_397_n 0.00422241f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A3_c_220_n N_VGND_c_402_n 0.00627034f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_185 A3 N_A_393_47#_c_457_n 0.00994288f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_186 N_A3_c_220_n N_A_393_47#_c_457_n 0.00936929f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A3_c_220_n N_A_393_47#_c_468_n 0.00690761f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_188 A3 N_A_393_47#_c_460_n 0.0176752f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_189 N_A3_c_219_n N_A_393_47#_c_460_n 0.00358038f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A3_c_220_n N_A_393_47#_c_460_n 0.00120357f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_M1011_g N_A1_M1000_g 0.0408383f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_192 A2 A1 0.0219557f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_193 N_A2_c_253_n A1 8.68831e-19 $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_194 A2 N_A1_c_284_n 0.0128462f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_195 N_A2_c_253_n N_A1_c_284_n 0.0220307f $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A2_c_254_n N_A1_c_285_n 0.0197301f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_197 A2 N_VPWR_c_312_n 0.0351711f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_198 N_A2_M1011_g N_VPWR_c_314_n 0.00383378f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_199 A2 N_VPWR_c_314_n 0.0110432f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_200 N_A2_M1011_g N_VPWR_c_307_n 0.0058067f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_201 A2 N_VPWR_c_307_n 0.0110141f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_202 A2 A_697_297# 0.0119511f $X=3.365 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_203 N_A2_c_254_n N_VGND_c_396_n 0.00311271f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_c_254_n N_VGND_c_397_n 0.00436487f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_c_254_n N_VGND_c_402_n 0.00626202f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_206 A2 N_A_393_47#_c_459_n 0.0260258f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_207 N_A2_c_253_n N_A_393_47#_c_459_n 0.003458f $X=3.49 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A2_c_254_n N_A_393_47#_c_459_n 0.0137112f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_M1000_g N_VPWR_c_312_n 0.0316548f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_210 A1 N_VPWR_c_312_n 0.0276365f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_211 N_A1_c_284_n N_VPWR_c_312_n 0.00137444f $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A1_M1000_g N_VPWR_c_314_n 0.00585385f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A1_M1000_g N_VPWR_c_307_n 0.0121347f $X=3.91 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A1_c_285_n N_VGND_c_396_n 0.0046886f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A1_c_285_n N_VGND_c_401_n 0.00436487f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A1_c_285_n N_VGND_c_402_n 0.00729423f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_217 A1 N_A_393_47#_c_459_n 0.045529f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_218 N_A1_c_284_n N_A_393_47#_c_459_n 0.00351017f $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A1_c_285_n N_A_393_47#_c_459_n 0.0151622f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A1_c_285_n N_A_393_47#_c_481_n 0.0137756f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_221 N_VPWR_c_307_n N_X_M1001_s 0.00215201f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_313_n X 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_c_307_n X 0.0122113f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_c_307_n A_496_297# 0.00892712f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_225 N_VPWR_c_307_n A_597_297# 0.00888445f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_226 N_VPWR_c_307_n A_697_297# 0.00919816f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_227 N_VPWR_c_309_n N_VGND_c_393_n 0.00886897f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_228 N_X_c_376_n N_VGND_c_399_n 0.0188922f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_229 N_X_M1004_s N_VGND_c_402_n 0.00215201f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_230 N_X_c_376_n N_VGND_c_402_n 0.0122173f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_231 N_VGND_c_402_n N_A_393_47#_M1002_d 0.00366865f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_232 N_VGND_c_402_n N_A_393_47#_M1013_d 0.00303553f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_402_n N_A_393_47#_M1009_d 0.00370066f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_400_n N_A_393_47#_c_485_n 0.0203242f $X=2.485 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_402_n N_A_393_47#_c_485_n 0.0126169f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_M1003_d N_A_393_47#_c_457_n 0.00273793f $X=2.48 $Y=0.235 $X2=0
+ $Y2=0
cc_237 N_VGND_c_395_n N_A_393_47#_c_457_n 0.0166712f $X=2.615 $Y=0.38 $X2=0
+ $Y2=0
cc_238 N_VGND_c_397_n N_A_393_47#_c_457_n 0.00251009f $X=3.505 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_400_n N_A_393_47#_c_457_n 0.00221217f $X=2.485 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_402_n N_A_393_47#_c_457_n 0.00964759f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_395_n N_A_393_47#_c_468_n 0.0191649f $X=2.615 $Y=0.38 $X2=0
+ $Y2=0
cc_242 N_VGND_c_397_n N_A_393_47#_c_468_n 0.0207144f $X=3.505 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_402_n N_A_393_47#_c_468_n 0.0124119f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_M1010_d N_A_393_47#_c_459_n 0.00241143f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_VGND_c_396_n N_A_393_47#_c_459_n 0.0182439f $X=3.64 $Y=0.38 $X2=0 $Y2=0
cc_246 N_VGND_c_397_n N_A_393_47#_c_459_n 0.00261576f $X=3.505 $Y=0 $X2=0 $Y2=0
cc_247 N_VGND_c_401_n N_A_393_47#_c_459_n 0.00334601f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_402_n N_A_393_47#_c_459_n 0.0131375f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_396_n N_A_393_47#_c_481_n 0.0154643f $X=3.64 $Y=0.38 $X2=0 $Y2=0
cc_250 N_VGND_c_401_n N_A_393_47#_c_481_n 0.022989f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_251 N_VGND_c_402_n N_A_393_47#_c_481_n 0.0126169f $X=4.37 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dlymetal6s2s_1.pxi.spice
* Created: Tue Sep  1 19:06:49 2020
* 
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A N_A_M1005_g N_A_M1000_g A A N_A_c_88_n
+ N_A_c_89_n PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_62_47# N_A_62_47#_M1005_s
+ N_A_62_47#_M1000_s N_A_62_47#_M1003_g N_A_62_47#_M1001_g N_A_62_47#_c_118_n
+ N_A_62_47#_c_125_n N_A_62_47#_c_126_n N_A_62_47#_c_119_n N_A_62_47#_c_127_n
+ N_A_62_47#_c_120_n N_A_62_47#_c_121_n N_A_62_47#_c_122_n N_A_62_47#_c_123_n
+ PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_62_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%X N_X_M1003_d N_X_M1001_d N_X_M1011_g
+ N_X_M1007_g X X X X X X X X N_X_c_178_n N_X_c_179_n
+ PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%X
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_381_47# N_A_381_47#_M1011_s
+ N_A_381_47#_M1007_s N_A_381_47#_M1006_g N_A_381_47#_M1008_g
+ N_A_381_47#_c_233_n N_A_381_47#_c_226_n N_A_381_47#_c_227_n
+ N_A_381_47#_c_228_n N_A_381_47#_c_234_n N_A_381_47#_c_235_n
+ N_A_381_47#_c_229_n N_A_381_47#_c_236_n N_A_381_47#_c_230_n
+ N_A_381_47#_c_231_n PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_381_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_558_47# N_A_558_47#_M1006_d
+ N_A_558_47#_M1008_d N_A_558_47#_M1004_g N_A_558_47#_M1002_g
+ N_A_558_47#_c_294_n N_A_558_47#_c_295_n N_A_558_47#_c_301_n
+ N_A_558_47#_c_296_n N_A_558_47#_c_297_n N_A_558_47#_c_298_n
+ PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_558_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_664_47# N_A_664_47#_M1004_s
+ N_A_664_47#_M1002_s N_A_664_47#_M1009_g N_A_664_47#_M1010_g
+ N_A_664_47#_c_348_n N_A_664_47#_c_355_n N_A_664_47#_c_349_n
+ N_A_664_47#_c_350_n N_A_664_47#_c_356_n N_A_664_47#_c_357_n
+ N_A_664_47#_c_351_n N_A_664_47#_c_358_n N_A_664_47#_c_352_n
+ N_A_664_47#_c_353_n PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_664_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%VPWR N_VPWR_M1000_d N_VPWR_M1007_d
+ N_VPWR_M1002_d N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n VPWR
+ N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_414_n N_VPWR_c_422_n
+ N_VPWR_c_423_n N_VPWR_c_424_n VPWR PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%VPWR
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_841_47# N_A_841_47#_M1009_d
+ N_A_841_47#_M1010_d N_A_841_47#_c_476_n N_A_841_47#_c_479_n
+ N_A_841_47#_c_480_n N_A_841_47#_c_477_n N_A_841_47#_c_478_n
+ PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_841_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%VGND N_VGND_M1005_d N_VGND_M1011_d
+ N_VGND_M1004_d N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n VGND
+ N_VGND_c_496_n N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n
+ N_VGND_c_501_n N_VGND_c_502_n VGND PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%VGND
cc_1 VNB N_A_M1005_g 0.0375092f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.445
cc_2 VNB N_A_c_88_n 0.0168494f $X=-0.19 $Y=-0.24 $X2=0.42 $Y2=1.16
cc_3 VNB N_A_c_89_n 0.0364194f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_4 VNB N_A_62_47#_c_118_n 0.00223093f $X=-0.19 $Y=-0.24 $X2=0.42 $Y2=1.16
cc_5 VNB N_A_62_47#_c_119_n 0.0323229f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.53
cc_6 VNB N_A_62_47#_c_120_n 0.00181412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_62_47#_c_121_n 0.0247986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_62_47#_c_122_n 0.00164805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_62_47#_c_123_n 0.0190541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_X_M1011_g 0.0342839f $X=-0.19 $Y=-0.24 $X2=0.12 $Y2=1.105
cc_11 VNB N_X_c_178_n 0.0348303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_X_c_179_n 0.0315919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_381_47#_c_226_n 0.00416701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_381_47#_c_227_n 9.94839e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_381_47#_c_228_n 0.00373045f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.53
cc_16 VNB N_A_381_47#_c_229_n 0.00358937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_381_47#_c_230_n 0.0236222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_381_47#_c_231_n 0.0190552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_558_47#_M1004_g 0.0342872f $X=-0.19 $Y=-0.24 $X2=0.12 $Y2=1.105
cc_20 VNB N_A_558_47#_c_294_n 0.00413128f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_21 VNB N_A_558_47#_c_295_n 0.0144963f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_22 VNB N_A_558_47#_c_296_n 0.003435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_558_47#_c_297_n 0.0010532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_558_47#_c_298_n 0.0338076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_664_47#_c_348_n 0.00392805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_664_47#_c_349_n 9.94839e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_664_47#_c_350_n 0.00362699f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.53
cc_28 VNB N_A_664_47#_c_351_n 0.00359032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_664_47#_c_352_n 0.0227379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_664_47#_c_353_n 0.0190552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_414_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_841_47#_c_476_n 0.0170421f $X=-0.19 $Y=-0.24 $X2=0.12 $Y2=1.105
cc_33 VNB N_A_841_47#_c_477_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_34 VNB N_A_841_47#_c_478_n 0.0219921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_493_n 4.8975e-19 $X=-0.19 $Y=-0.24 $X2=0.42 $Y2=1.16
cc_36 VNB N_VGND_c_494_n 4.8975e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_495_n 4.8975e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_496_n 0.0292346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_497_n 0.0252189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_498_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_499_n 0.258137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_500_n 0.0233399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_501_n 0.00509417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_502_n 0.00509417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VPB N_A_M1000_g 0.0605617f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=2.275
cc_46 VPB N_A_c_88_n 0.025716f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.16
cc_47 VPB N_A_c_89_n 0.00991829f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_48 VPB N_A_62_47#_M1001_g 0.0216941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_62_47#_c_125_n 0.00279153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_62_47#_c_126_n 0.00421703f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.19
cc_51 VPB N_A_62_47#_c_127_n 0.0342336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_62_47#_c_121_n 0.00491423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_X_M1007_g 0.0573581f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.16
cc_54 VPB X 0.0143438f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.16
cc_55 VPB N_X_c_178_n 0.0099102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_X_c_179_n 0.0200645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_381_47#_M1008_g 0.0216941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_381_47#_c_233_n 0.00502651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_381_47#_c_234_n 0.00171281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_381_47#_c_235_n 0.00465697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_381_47#_c_236_n 0.00414885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_381_47#_c_230_n 0.00483834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_558_47#_M1002_g 0.0573581f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.16
cc_64 VPB N_A_558_47#_c_295_n 0.0182197f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.16
cc_65 VPB N_A_558_47#_c_301_n 0.00786923f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.19
cc_66 VPB N_A_558_47#_c_298_n 0.00984422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_664_47#_M1010_g 0.0216957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_664_47#_c_355_n 0.00444492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_664_47#_c_356_n 0.00171281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_664_47#_c_357_n 0.00427171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_664_47#_c_358_n 0.00414885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_664_47#_c_352_n 0.00478128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_415_n 4.8975e-19 $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.16
cc_74 VPB N_VPWR_c_416_n 4.8975e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_417_n 4.8975e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_418_n 0.0291003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_419_n 0.0252539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_420_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_414_n 0.0636833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_422_n 0.0233767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_423_n 0.00509586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_424_n 0.00509586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_841_47#_c_479_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_841_47#_c_480_n 0.0322452f $X=-0.19 $Y=1.305 $X2=0.42 $Y2=1.16
cc_85 VPB N_A_841_47#_c_478_n 0.00891602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 N_A_M1000_g N_A_62_47#_M1001_g 0.0332384f $X=0.645 $Y=2.275 $X2=0 $Y2=0
cc_87 N_A_M1005_g N_A_62_47#_c_118_n 0.0169506f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_c_88_n N_A_62_47#_c_118_n 0.00392725f $X=0.42 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_c_89_n N_A_62_47#_c_118_n 3.45424e-19 $X=0.645 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_M1000_g N_A_62_47#_c_125_n 0.017035f $X=0.645 $Y=2.275 $X2=0 $Y2=0
cc_91 N_A_c_88_n N_A_62_47#_c_125_n 0.00415099f $X=0.42 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_M1000_g N_A_62_47#_c_126_n 0.00523842f $X=0.645 $Y=2.275 $X2=0 $Y2=0
cc_93 N_A_M1005_g N_A_62_47#_c_119_n 0.00157466f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_c_88_n N_A_62_47#_c_119_n 0.0390823f $X=0.42 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_c_89_n N_A_62_47#_c_119_n 0.00181525f $X=0.645 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_M1000_g N_A_62_47#_c_127_n 0.0029776f $X=0.645 $Y=2.275 $X2=0 $Y2=0
cc_97 N_A_c_88_n N_A_62_47#_c_127_n 0.0402782f $X=0.42 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_c_89_n N_A_62_47#_c_127_n 8.36308e-19 $X=0.645 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_c_88_n N_A_62_47#_c_120_n 0.0594526f $X=0.42 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_c_89_n N_A_62_47#_c_120_n 0.00523842f $X=0.645 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_c_88_n N_A_62_47#_c_121_n 2.33019e-19 $X=0.42 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_c_89_n N_A_62_47#_c_121_n 0.0207322f $X=0.645 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_M1005_g N_A_62_47#_c_122_n 0.00523842f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_M1005_g N_A_62_47#_c_123_n 0.0194517f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_M1000_g N_VPWR_c_415_n 0.00906078f $X=0.645 $Y=2.275 $X2=0 $Y2=0
cc_106 N_A_M1000_g N_VPWR_c_414_n 0.0052023f $X=0.645 $Y=2.275 $X2=0 $Y2=0
cc_107 N_A_M1000_g N_VPWR_c_422_n 0.00344532f $X=0.645 $Y=2.275 $X2=0 $Y2=0
cc_108 N_A_M1005_g N_VGND_c_493_n 0.00878516f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_M1005_g N_VGND_c_499_n 0.00515284f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_M1005_g N_VGND_c_500_n 0.00341689f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_62_47#_c_121_n N_X_c_178_n 0.00328875f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_62_47#_M1001_g N_X_c_179_n 0.00379362f $X=1.12 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_62_47#_c_126_n N_X_c_179_n 0.0108745f $X=0.907 $Y=1.87 $X2=0 $Y2=0
cc_114 N_A_62_47#_c_120_n N_X_c_179_n 0.0282481f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_62_47#_c_121_n N_X_c_179_n 0.00401301f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_62_47#_c_122_n N_X_c_179_n 0.0101847f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_62_47#_c_123_n N_X_c_179_n 0.00367346f $X=1.065 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_62_47#_c_125_n N_VPWR_M1000_d 0.00207054f $X=0.74 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_62_47#_c_126_n N_VPWR_M1000_d 7.20661e-19 $X=0.907 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_62_47#_M1001_g N_VPWR_c_415_n 0.00905956f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_62_47#_c_125_n N_VPWR_c_415_n 0.0245954f $X=0.74 $Y=1.955 $X2=0 $Y2=0
cc_122 N_A_62_47#_M1001_g N_VPWR_c_418_n 0.0046653f $X=1.12 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_62_47#_M1000_s N_VPWR_c_414_n 0.00230841f $X=0.31 $Y=2.065 $X2=0
+ $Y2=0
cc_124 N_A_62_47#_M1001_g N_VPWR_c_414_n 0.00921786f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_62_47#_c_125_n N_VPWR_c_414_n 0.00581522f $X=0.74 $Y=1.955 $X2=0
+ $Y2=0
cc_126 N_A_62_47#_c_127_n N_VPWR_c_414_n 0.0166176f $X=0.302 $Y=1.955 $X2=0
+ $Y2=0
cc_127 N_A_62_47#_c_125_n N_VPWR_c_422_n 0.00259647f $X=0.74 $Y=1.955 $X2=0
+ $Y2=0
cc_128 N_A_62_47#_c_127_n N_VPWR_c_422_n 0.0302478f $X=0.302 $Y=1.955 $X2=0
+ $Y2=0
cc_129 N_A_62_47#_c_118_n N_VGND_M1005_d 0.00264964f $X=0.74 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_62_47#_c_118_n N_VGND_c_493_n 0.024366f $X=0.74 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_62_47#_c_121_n N_VGND_c_493_n 3.47021e-19 $X=1.065 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_62_47#_c_123_n N_VGND_c_493_n 0.00877802f $X=1.065 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_62_47#_c_123_n N_VGND_c_496_n 0.0046653f $X=1.065 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_62_47#_M1005_s N_VGND_c_499_n 0.00229009f $X=0.31 $Y=0.235 $X2=0
+ $Y2=0
cc_135 N_A_62_47#_c_118_n N_VGND_c_499_n 0.00598099f $X=0.74 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_62_47#_c_119_n N_VGND_c_499_n 0.0165992f $X=0.435 $Y=0.445 $X2=0
+ $Y2=0
cc_137 N_A_62_47#_c_123_n N_VGND_c_499_n 0.00934473f $X=1.065 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_A_62_47#_c_118_n N_VGND_c_500_n 0.00273399f $X=0.74 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_62_47#_c_119_n N_VGND_c_500_n 0.0301526f $X=0.435 $Y=0.445 $X2=0
+ $Y2=0
cc_140 N_X_M1007_g N_A_381_47#_M1008_g 0.0333474f $X=2.24 $Y=2.275 $X2=0 $Y2=0
cc_141 N_X_M1007_g N_A_381_47#_c_233_n 0.00127827f $X=2.24 $Y=2.275 $X2=0 $Y2=0
cc_142 X N_A_381_47#_c_233_n 0.0355571f $X=1.5 $Y=1.785 $X2=0 $Y2=0
cc_143 N_X_c_179_n N_A_381_47#_c_226_n 0.0309004f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_144 N_X_M1011_g N_A_381_47#_c_227_n 0.0178202f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_145 N_X_c_178_n N_A_381_47#_c_227_n 8.08044e-19 $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_146 N_X_c_179_n N_A_381_47#_c_227_n 0.00275926f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_147 N_X_c_178_n N_A_381_47#_c_228_n 0.00182316f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_148 N_X_c_179_n N_A_381_47#_c_228_n 0.0367289f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_149 N_X_M1007_g N_A_381_47#_c_234_n 0.0192581f $X=2.24 $Y=2.275 $X2=0 $Y2=0
cc_150 N_X_c_178_n N_A_381_47#_c_234_n 5.13753e-19 $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_151 N_X_c_179_n N_A_381_47#_c_234_n 0.00294539f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_152 X N_A_381_47#_c_235_n 0.0175677f $X=1.5 $Y=1.785 $X2=0 $Y2=0
cc_153 N_X_c_178_n N_A_381_47#_c_235_n 8.79705e-19 $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_154 N_X_c_179_n N_A_381_47#_c_235_n 0.0255903f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_155 N_X_M1011_g N_A_381_47#_c_229_n 0.00558618f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_156 N_X_c_179_n N_A_381_47#_c_229_n 0.0339191f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_157 N_X_M1007_g N_A_381_47#_c_236_n 0.00592384f $X=2.24 $Y=2.275 $X2=0 $Y2=0
cc_158 X N_A_381_47#_c_236_n 0.00558909f $X=1.5 $Y=1.785 $X2=0 $Y2=0
cc_159 N_X_c_179_n N_A_381_47#_c_236_n 0.0310274f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_160 N_X_c_178_n N_A_381_47#_c_230_n 0.0207275f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_161 N_X_c_179_n N_A_381_47#_c_230_n 2.21861e-19 $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_162 N_X_M1011_g N_A_381_47#_c_231_n 0.0194472f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_163 N_X_M1007_g N_VPWR_c_416_n 0.00906078f $X=2.24 $Y=2.275 $X2=0 $Y2=0
cc_164 N_X_M1007_g N_VPWR_c_418_n 0.00344532f $X=2.24 $Y=2.275 $X2=0 $Y2=0
cc_165 X N_VPWR_c_418_n 0.0298308f $X=1.5 $Y=1.785 $X2=0 $Y2=0
cc_166 N_X_M1001_d N_VPWR_c_414_n 0.00382897f $X=1.195 $Y=1.485 $X2=0 $Y2=0
cc_167 N_X_M1007_g N_VPWR_c_414_n 0.00545273f $X=2.24 $Y=2.275 $X2=0 $Y2=0
cc_168 X N_VPWR_c_414_n 0.0162905f $X=1.5 $Y=1.785 $X2=0 $Y2=0
cc_169 N_X_M1011_g N_VGND_c_494_n 0.00878516f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_170 N_X_M1011_g N_VGND_c_496_n 0.00341689f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_171 N_X_c_179_n N_VGND_c_496_n 0.0298767f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_172 N_X_M1003_d N_VGND_c_499_n 0.003837f $X=1.195 $Y=0.235 $X2=0 $Y2=0
cc_173 N_X_M1011_g N_VGND_c_499_n 0.00540327f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_174 N_X_c_179_n N_VGND_c_499_n 0.0163543f $X=1.457 $Y=1.675 $X2=0 $Y2=0
cc_175 N_A_381_47#_M1008_g N_A_558_47#_c_295_n 0.00377535f $X=2.715 $Y=1.985
+ $X2=0 $Y2=0
cc_176 N_A_381_47#_c_229_n N_A_558_47#_c_295_n 0.0283504f $X=2.495 $Y=1.325
+ $X2=0 $Y2=0
cc_177 N_A_381_47#_c_236_n N_A_558_47#_c_295_n 0.0108652f $X=2.495 $Y=1.845
+ $X2=0 $Y2=0
cc_178 N_A_381_47#_c_230_n N_A_558_47#_c_295_n 0.00336476f $X=2.66 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_381_47#_c_229_n N_A_558_47#_c_296_n 0.00962502f $X=2.495 $Y=1.325
+ $X2=0 $Y2=0
cc_180 N_A_381_47#_c_231_n N_A_558_47#_c_296_n 0.00355882f $X=2.66 $Y=0.995
+ $X2=0 $Y2=0
cc_181 N_A_381_47#_c_229_n N_A_558_47#_c_298_n 2.35222e-19 $X=2.495 $Y=1.325
+ $X2=0 $Y2=0
cc_182 N_A_381_47#_c_230_n N_A_558_47#_c_298_n 0.0058474f $X=2.66 $Y=1.16 $X2=0
+ $Y2=0
cc_183 N_A_381_47#_c_234_n N_VPWR_M1007_d 0.00207054f $X=2.32 $Y=1.942 $X2=0
+ $Y2=0
cc_184 N_A_381_47#_c_236_n N_VPWR_M1007_d 6.23798e-19 $X=2.495 $Y=1.845 $X2=0
+ $Y2=0
cc_185 N_A_381_47#_M1008_g N_VPWR_c_416_n 0.00905956f $X=2.715 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_381_47#_c_234_n N_VPWR_c_416_n 0.024785f $X=2.32 $Y=1.942 $X2=0 $Y2=0
cc_187 N_A_381_47#_c_233_n N_VPWR_c_418_n 0.0189483f $X=2.03 $Y=2.275 $X2=0
+ $Y2=0
cc_188 N_A_381_47#_c_234_n N_VPWR_c_418_n 0.00261227f $X=2.32 $Y=1.942 $X2=0
+ $Y2=0
cc_189 N_A_381_47#_M1008_g N_VPWR_c_419_n 0.0046653f $X=2.715 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_381_47#_M1007_s N_VPWR_c_414_n 0.00230841f $X=1.905 $Y=2.065 $X2=0
+ $Y2=0
cc_191 N_A_381_47#_M1008_g N_VPWR_c_414_n 0.00921786f $X=2.715 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_381_47#_c_233_n N_VPWR_c_414_n 0.0104883f $X=2.03 $Y=2.275 $X2=0
+ $Y2=0
cc_193 N_A_381_47#_c_234_n N_VPWR_c_414_n 0.005846f $X=2.32 $Y=1.942 $X2=0 $Y2=0
cc_194 N_A_381_47#_c_229_n N_VGND_M1011_d 0.0028099f $X=2.495 $Y=1.325 $X2=0
+ $Y2=0
cc_195 N_A_381_47#_c_227_n N_VGND_c_494_n 0.00217981f $X=2.32 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_381_47#_c_229_n N_VGND_c_494_n 0.0222857f $X=2.495 $Y=1.325 $X2=0
+ $Y2=0
cc_197 N_A_381_47#_c_230_n N_VGND_c_494_n 3.47021e-19 $X=2.66 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_381_47#_c_231_n N_VGND_c_494_n 0.00878394f $X=2.66 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_381_47#_c_226_n N_VGND_c_496_n 0.0174182f $X=2.03 $Y=0.44 $X2=0 $Y2=0
cc_200 N_A_381_47#_c_227_n N_VGND_c_496_n 0.00273399f $X=2.32 $Y=0.74 $X2=0
+ $Y2=0
cc_201 N_A_381_47#_c_231_n N_VGND_c_497_n 0.0046653f $X=2.66 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_381_47#_M1011_s N_VGND_c_499_n 0.00229009f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_203 N_A_381_47#_c_226_n N_VGND_c_499_n 0.00969887f $X=2.03 $Y=0.44 $X2=0
+ $Y2=0
cc_204 N_A_381_47#_c_227_n N_VGND_c_499_n 0.00430392f $X=2.32 $Y=0.74 $X2=0
+ $Y2=0
cc_205 N_A_381_47#_c_229_n N_VGND_c_499_n 0.00168578f $X=2.495 $Y=1.325 $X2=0
+ $Y2=0
cc_206 N_A_381_47#_c_231_n N_VGND_c_499_n 0.00934473f $X=2.66 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_558_47#_M1002_g N_A_664_47#_M1010_g 0.0333474f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_208 N_A_558_47#_c_294_n N_A_664_47#_c_348_n 0.0294952f $X=2.925 $Y=0.44 $X2=0
+ $Y2=0
cc_209 N_A_558_47#_M1002_g N_A_664_47#_c_355_n 0.00126954f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_210 N_A_558_47#_c_301_n N_A_664_47#_c_355_n 0.0313409f $X=2.925 $Y=1.96 $X2=0
+ $Y2=0
cc_211 N_A_558_47#_M1004_g N_A_664_47#_c_349_n 0.0178202f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_212 N_A_558_47#_c_295_n N_A_664_47#_c_349_n 0.00275926f $X=2.962 $Y=1.675
+ $X2=0 $Y2=0
cc_213 N_A_558_47#_c_298_n N_A_664_47#_c_349_n 8.08044e-19 $X=3.655 $Y=1.16
+ $X2=0 $Y2=0
cc_214 N_A_558_47#_c_294_n N_A_664_47#_c_350_n 0.0135733f $X=2.925 $Y=0.44 $X2=0
+ $Y2=0
cc_215 N_A_558_47#_c_295_n N_A_664_47#_c_350_n 0.0225151f $X=2.962 $Y=1.675
+ $X2=0 $Y2=0
cc_216 N_A_558_47#_c_298_n N_A_664_47#_c_350_n 0.00182316f $X=3.655 $Y=1.16
+ $X2=0 $Y2=0
cc_217 N_A_558_47#_M1002_g N_A_664_47#_c_356_n 0.0192005f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_218 N_A_558_47#_c_295_n N_A_664_47#_c_356_n 0.00294539f $X=2.962 $Y=1.675
+ $X2=0 $Y2=0
cc_219 N_A_558_47#_c_298_n N_A_664_47#_c_356_n 5.13753e-19 $X=3.655 $Y=1.16
+ $X2=0 $Y2=0
cc_220 N_A_558_47#_c_295_n N_A_664_47#_c_357_n 0.0237293f $X=2.962 $Y=1.675
+ $X2=0 $Y2=0
cc_221 N_A_558_47#_c_301_n N_A_664_47#_c_357_n 0.0156118f $X=2.925 $Y=1.96 $X2=0
+ $Y2=0
cc_222 N_A_558_47#_c_298_n N_A_664_47#_c_357_n 8.79705e-19 $X=3.655 $Y=1.16
+ $X2=0 $Y2=0
cc_223 N_A_558_47#_M1004_g N_A_664_47#_c_351_n 0.00558831f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_224 N_A_558_47#_c_295_n N_A_664_47#_c_351_n 0.0282667f $X=2.962 $Y=1.675
+ $X2=0 $Y2=0
cc_225 N_A_558_47#_c_296_n N_A_664_47#_c_351_n 0.00522819f $X=3 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_558_47#_M1002_g N_A_664_47#_c_358_n 0.00592384f $X=3.655 $Y=2.275
+ $X2=0 $Y2=0
cc_227 N_A_558_47#_c_295_n N_A_664_47#_c_358_n 0.0309738f $X=2.962 $Y=1.675
+ $X2=0 $Y2=0
cc_228 N_A_558_47#_c_301_n N_A_664_47#_c_358_n 0.00536031f $X=2.925 $Y=1.96
+ $X2=0 $Y2=0
cc_229 N_A_558_47#_c_295_n N_A_664_47#_c_352_n 2.22114e-19 $X=2.962 $Y=1.675
+ $X2=0 $Y2=0
cc_230 N_A_558_47#_c_298_n N_A_664_47#_c_352_n 0.0207275f $X=3.655 $Y=1.16 $X2=0
+ $Y2=0
cc_231 N_A_558_47#_M1004_g N_A_664_47#_c_353_n 0.0194472f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_232 N_A_558_47#_M1002_g N_VPWR_c_417_n 0.00906078f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_233 N_A_558_47#_M1002_g N_VPWR_c_419_n 0.00344532f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_234 N_A_558_47#_c_301_n N_VPWR_c_419_n 0.0169256f $X=2.925 $Y=1.96 $X2=0
+ $Y2=0
cc_235 N_A_558_47#_M1008_d N_VPWR_c_414_n 0.00382897f $X=2.79 $Y=1.485 $X2=0
+ $Y2=0
cc_236 N_A_558_47#_M1002_g N_VPWR_c_414_n 0.00545273f $X=3.655 $Y=2.275 $X2=0
+ $Y2=0
cc_237 N_A_558_47#_c_301_n N_VPWR_c_414_n 0.00935836f $X=2.925 $Y=1.96 $X2=0
+ $Y2=0
cc_238 N_A_558_47#_M1004_g N_VGND_c_495_n 0.00878516f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_239 N_A_558_47#_M1004_g N_VGND_c_497_n 0.00341689f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_240 N_A_558_47#_c_294_n N_VGND_c_497_n 0.0168644f $X=2.925 $Y=0.44 $X2=0
+ $Y2=0
cc_241 N_A_558_47#_M1006_d N_VGND_c_499_n 0.00387172f $X=2.79 $Y=0.235 $X2=0
+ $Y2=0
cc_242 N_A_558_47#_M1004_g N_VGND_c_499_n 0.00540327f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_243 N_A_558_47#_c_294_n N_VGND_c_499_n 0.00934531f $X=2.925 $Y=0.44 $X2=0
+ $Y2=0
cc_244 N_A_664_47#_c_356_n N_VPWR_M1002_d 0.00207054f $X=3.735 $Y=1.942 $X2=0
+ $Y2=0
cc_245 N_A_664_47#_c_358_n N_VPWR_M1002_d 6.23798e-19 $X=3.91 $Y=1.845 $X2=0
+ $Y2=0
cc_246 N_A_664_47#_M1010_g N_VPWR_c_417_n 0.00905956f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_664_47#_c_356_n N_VPWR_c_417_n 0.024785f $X=3.735 $Y=1.942 $X2=0
+ $Y2=0
cc_248 N_A_664_47#_c_355_n N_VPWR_c_419_n 0.0175244f $X=3.445 $Y=2.275 $X2=0
+ $Y2=0
cc_249 N_A_664_47#_c_356_n N_VPWR_c_419_n 0.00261227f $X=3.735 $Y=1.942 $X2=0
+ $Y2=0
cc_250 N_A_664_47#_M1010_g N_VPWR_c_420_n 0.0046653f $X=4.13 $Y=1.985 $X2=0
+ $Y2=0
cc_251 N_A_664_47#_M1002_s N_VPWR_c_414_n 0.00230841f $X=3.32 $Y=2.065 $X2=0
+ $Y2=0
cc_252 N_A_664_47#_M1010_g N_VPWR_c_414_n 0.008846f $X=4.13 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_664_47#_c_355_n N_VPWR_c_414_n 0.00971993f $X=3.445 $Y=2.275 $X2=0
+ $Y2=0
cc_254 N_A_664_47#_c_356_n N_VPWR_c_414_n 0.005846f $X=3.735 $Y=1.942 $X2=0
+ $Y2=0
cc_255 N_A_664_47#_M1010_g N_A_841_47#_c_478_n 0.00357537f $X=4.13 $Y=1.985
+ $X2=0 $Y2=0
cc_256 N_A_664_47#_c_351_n N_A_841_47#_c_478_n 0.0352893f $X=3.91 $Y=1.325 $X2=0
+ $Y2=0
cc_257 N_A_664_47#_c_358_n N_A_841_47#_c_478_n 0.0097546f $X=3.91 $Y=1.845 $X2=0
+ $Y2=0
cc_258 N_A_664_47#_c_352_n N_A_841_47#_c_478_n 0.00754383f $X=4.075 $Y=1.16
+ $X2=0 $Y2=0
cc_259 N_A_664_47#_c_353_n N_A_841_47#_c_478_n 0.00357326f $X=4.075 $Y=0.995
+ $X2=0 $Y2=0
cc_260 N_A_664_47#_c_351_n N_VGND_M1004_d 0.0028099f $X=3.91 $Y=1.325 $X2=0
+ $Y2=0
cc_261 N_A_664_47#_c_349_n N_VGND_c_495_n 0.00217981f $X=3.735 $Y=0.74 $X2=0
+ $Y2=0
cc_262 N_A_664_47#_c_351_n N_VGND_c_495_n 0.0222857f $X=3.91 $Y=1.325 $X2=0
+ $Y2=0
cc_263 N_A_664_47#_c_352_n N_VGND_c_495_n 3.47021e-19 $X=4.075 $Y=1.16 $X2=0
+ $Y2=0
cc_264 N_A_664_47#_c_353_n N_VGND_c_495_n 0.00878394f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_664_47#_c_348_n N_VGND_c_497_n 0.0174182f $X=3.445 $Y=0.44 $X2=0
+ $Y2=0
cc_266 N_A_664_47#_c_349_n N_VGND_c_497_n 0.00273399f $X=3.735 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_664_47#_c_353_n N_VGND_c_498_n 0.0046653f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_268 N_A_664_47#_M1004_s N_VGND_c_499_n 0.00229009f $X=3.32 $Y=0.235 $X2=0
+ $Y2=0
cc_269 N_A_664_47#_c_348_n N_VGND_c_499_n 0.00969887f $X=3.445 $Y=0.44 $X2=0
+ $Y2=0
cc_270 N_A_664_47#_c_349_n N_VGND_c_499_n 0.00430392f $X=3.735 $Y=0.74 $X2=0
+ $Y2=0
cc_271 N_A_664_47#_c_351_n N_VGND_c_499_n 0.00168578f $X=3.91 $Y=1.325 $X2=0
+ $Y2=0
cc_272 N_A_664_47#_c_353_n N_VGND_c_499_n 0.00895857f $X=4.075 $Y=0.995 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_414_n N_A_841_47#_M1010_d 0.00382897f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_420_n N_A_841_47#_c_480_n 0.018001f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_275 N_VPWR_c_414_n N_A_841_47#_c_480_n 0.00993603f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_A_841_47#_c_476_n N_VGND_c_498_n 0.0179398f $X=4.34 $Y=0.44 $X2=0 $Y2=0
cc_277 N_A_841_47#_M1009_d N_VGND_c_499_n 0.00387172f $X=4.205 $Y=0.235 $X2=0
+ $Y2=0
cc_278 N_A_841_47#_c_476_n N_VGND_c_499_n 0.00992299f $X=4.34 $Y=0.44 $X2=0
+ $Y2=0

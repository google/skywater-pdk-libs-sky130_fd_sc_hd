* File: sky130_fd_sc_hd__o32ai_4.pex.spice
* Created: Tue Sep  1 19:26:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O32AI_4%B2 3 7 11 15 19 23 27 31 33 34 35 48 49
r69 47 49 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.73 $Y2=1.16
r70 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r71 45 47 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r72 44 45 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r73 43 44 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r74 40 43 40.336 $w=2.9e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r75 35 48 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.52 $Y2=1.175
r76 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.155 $Y2=1.175
r77 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r78 33 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r79 29 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.73 $Y=1.305
+ $X2=1.73 $Y2=1.16
r80 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.73 $Y=1.305
+ $X2=1.73 $Y2=1.985
r81 25 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.73 $Y=1.015
+ $X2=1.73 $Y2=1.16
r82 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.73 $Y=1.015
+ $X2=1.73 $Y2=0.56
r83 21 45 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.31 $Y=1.305
+ $X2=1.31 $Y2=1.16
r84 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.31 $Y=1.305
+ $X2=1.31 $Y2=1.985
r85 17 45 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.31 $Y=1.015
+ $X2=1.31 $Y2=1.16
r86 17 19 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.31 $Y=1.015
+ $X2=1.31 $Y2=0.56
r87 13 44 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.89 $Y=1.305
+ $X2=0.89 $Y2=1.16
r88 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.89 $Y=1.305
+ $X2=0.89 $Y2=1.985
r89 9 44 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.89 $Y=1.015
+ $X2=0.89 $Y2=1.16
r90 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.89 $Y=1.015
+ $X2=0.89 $Y2=0.56
r91 5 43 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r92 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=1.985
r93 1 43 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r94 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%B1 3 7 11 15 19 23 27 31 33 34 35 49
c65 27 0 1.79953e-19 $X=3.425 $Y=0.56
r66 47 49 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=3.215 $Y=1.16
+ $X2=3.425 $Y2=1.16
r67 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=1.16 $X2=3.215 $Y2=1.16
r68 45 47 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=3.005 $Y=1.16
+ $X2=3.215 $Y2=1.16
r69 44 45 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=2.585 $Y=1.16
+ $X2=3.005 $Y2=1.16
r70 42 44 44.473 $w=2.9e-07 $l=2.15e-07 $layer=POLY_cond $X=2.37 $Y=1.16
+ $X2=2.585 $Y2=1.16
r71 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.16 $X2=2.37 $Y2=1.16
r72 39 42 42.4045 $w=2.9e-07 $l=2.05e-07 $layer=POLY_cond $X=2.165 $Y=1.16
+ $X2=2.37 $Y2=1.16
r73 35 48 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=3.455 $Y=1.175
+ $X2=3.215 $Y2=1.175
r74 34 48 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=3.215 $Y2=1.175
r75 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.995 $Y2=1.175
r76 33 43 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.37 $Y2=1.175
r77 29 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.425 $Y=1.305
+ $X2=3.425 $Y2=1.16
r78 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.425 $Y=1.305
+ $X2=3.425 $Y2=1.985
r79 25 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.425 $Y=1.015
+ $X2=3.425 $Y2=1.16
r80 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.425 $Y=1.015
+ $X2=3.425 $Y2=0.56
r81 21 45 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.005 $Y=1.305
+ $X2=3.005 $Y2=1.16
r82 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.005 $Y=1.305
+ $X2=3.005 $Y2=1.985
r83 17 45 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.005 $Y=1.015
+ $X2=3.005 $Y2=1.16
r84 17 19 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.005 $Y=1.015
+ $X2=3.005 $Y2=0.56
r85 13 44 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.585 $Y=1.305
+ $X2=2.585 $Y2=1.16
r86 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.585 $Y=1.305
+ $X2=2.585 $Y2=1.985
r87 9 44 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.585 $Y=1.015
+ $X2=2.585 $Y2=1.16
r88 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.585 $Y=1.015
+ $X2=2.585 $Y2=0.56
r89 5 39 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.165 $Y=1.305
+ $X2=2.165 $Y2=1.16
r90 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.165 $Y=1.305
+ $X2=2.165 $Y2=1.985
r91 1 39 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.165 $Y=1.015
+ $X2=2.165 $Y2=1.16
r92 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.165 $Y=1.015
+ $X2=2.165 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 55
c86 3 0 7.99167e-20 $X=3.845 $Y=0.56
r87 54 55 74.4665 $w=2.9e-07 $l=3.6e-07 $layer=POLY_cond $X=5.265 $Y=1.16
+ $X2=5.625 $Y2=1.16
r88 53 54 12.4111 $w=2.9e-07 $l=6e-08 $layer=POLY_cond $X=5.205 $Y=1.16
+ $X2=5.265 $Y2=1.16
r89 51 53 2.06851 $w=2.9e-07 $l=1e-08 $layer=POLY_cond $X=5.195 $Y=1.16
+ $X2=5.205 $Y2=1.16
r90 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.195
+ $Y=1.16 $X2=5.195 $Y2=1.16
r91 49 51 84.8091 $w=2.9e-07 $l=4.1e-07 $layer=POLY_cond $X=4.785 $Y=1.16
+ $X2=5.195 $Y2=1.16
r92 48 49 20.6851 $w=2.9e-07 $l=1e-07 $layer=POLY_cond $X=4.685 $Y=1.16
+ $X2=4.785 $Y2=1.16
r93 47 48 66.1924 $w=2.9e-07 $l=3.2e-07 $layer=POLY_cond $X=4.365 $Y=1.16
+ $X2=4.685 $Y2=1.16
r94 46 47 20.6851 $w=2.9e-07 $l=1e-07 $layer=POLY_cond $X=4.265 $Y=1.16
+ $X2=4.365 $Y2=1.16
r95 44 46 68.261 $w=2.9e-07 $l=3.3e-07 $layer=POLY_cond $X=3.935 $Y=1.16
+ $X2=4.265 $Y2=1.16
r96 41 44 18.6166 $w=2.9e-07 $l=9e-08 $layer=POLY_cond $X=3.845 $Y=1.16
+ $X2=3.935 $Y2=1.16
r97 36 52 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=5.295 $Y=1.175
+ $X2=5.195 $Y2=1.175
r98 35 52 19.9636 $w=1.98e-07 $l=3.6e-07 $layer=LI1_cond $X=4.835 $Y=1.175
+ $X2=5.195 $Y2=1.175
r99 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.375 $Y=1.175
+ $X2=4.835 $Y2=1.175
r100 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.915 $Y=1.175
+ $X2=4.375 $Y2=1.175
r101 33 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.935
+ $Y=1.16 $X2=3.935 $Y2=1.16
r102 29 55 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.625 $Y=1.305
+ $X2=5.625 $Y2=1.16
r103 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.625 $Y=1.305
+ $X2=5.625 $Y2=1.985
r104 25 54 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.265 $Y=1.015
+ $X2=5.265 $Y2=1.16
r105 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.265 $Y=1.015
+ $X2=5.265 $Y2=0.56
r106 21 53 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.205 $Y=1.305
+ $X2=5.205 $Y2=1.16
r107 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.205 $Y=1.305
+ $X2=5.205 $Y2=1.985
r108 17 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.785 $Y=1.305
+ $X2=4.785 $Y2=1.16
r109 17 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.785 $Y=1.305
+ $X2=4.785 $Y2=1.985
r110 13 48 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.685 $Y=1.015
+ $X2=4.685 $Y2=1.16
r111 13 15 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.685 $Y=1.015
+ $X2=4.685 $Y2=0.56
r112 9 47 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.365 $Y=1.305
+ $X2=4.365 $Y2=1.16
r113 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.365 $Y=1.305
+ $X2=4.365 $Y2=1.985
r114 5 46 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.265 $Y=1.015
+ $X2=4.265 $Y2=1.16
r115 5 7 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.265 $Y=1.015
+ $X2=4.265 $Y2=0.56
r116 1 41 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.845 $Y=1.015
+ $X2=3.845 $Y2=1.16
r117 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.845 $Y=1.015
+ $X2=3.845 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%A2 3 7 11 15 19 23 27 31 33 34 35 49
r76 47 49 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=7.095 $Y=1.16
+ $X2=7.305 $Y2=1.16
r77 45 47 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=6.885 $Y=1.16
+ $X2=7.095 $Y2=1.16
r78 44 45 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=6.465 $Y=1.16
+ $X2=6.885 $Y2=1.16
r79 42 44 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=6.255 $Y=1.16
+ $X2=6.465 $Y2=1.16
r80 39 42 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=6.045 $Y=1.16
+ $X2=6.255 $Y2=1.16
r81 35 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.095
+ $Y=1.16 $X2=7.095 $Y2=1.16
r82 34 35 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=6.675 $Y=1.175
+ $X2=7.095 $Y2=1.175
r83 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.215 $Y=1.175
+ $X2=6.675 $Y2=1.175
r84 33 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.255
+ $Y=1.16 $X2=6.255 $Y2=1.16
r85 29 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.305 $Y=1.305
+ $X2=7.305 $Y2=1.16
r86 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.305 $Y=1.305
+ $X2=7.305 $Y2=1.985
r87 25 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.305 $Y=1.015
+ $X2=7.305 $Y2=1.16
r88 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.305 $Y=1.015
+ $X2=7.305 $Y2=0.56
r89 21 45 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=6.885 $Y=1.305
+ $X2=6.885 $Y2=1.16
r90 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.885 $Y=1.305
+ $X2=6.885 $Y2=1.985
r91 17 45 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=6.885 $Y=1.015
+ $X2=6.885 $Y2=1.16
r92 17 19 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.885 $Y=1.015
+ $X2=6.885 $Y2=0.56
r93 13 44 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=6.465 $Y=1.305
+ $X2=6.465 $Y2=1.16
r94 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.465 $Y=1.305
+ $X2=6.465 $Y2=1.985
r95 9 44 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=6.465 $Y=1.015
+ $X2=6.465 $Y2=1.16
r96 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.465 $Y=1.015
+ $X2=6.465 $Y2=0.56
r97 5 39 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=6.045 $Y=1.305
+ $X2=6.045 $Y2=1.16
r98 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.045 $Y=1.305
+ $X2=6.045 $Y2=1.985
r99 1 39 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=6.045 $Y=1.015
+ $X2=6.045 $Y2=1.16
r100 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.045 $Y=1.015
+ $X2=6.045 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%A1 3 7 11 15 19 23 25 26 29 33 35 36 37 38
+ 52 64
r81 53 64 10.8136 $w=1.98e-07 $l=1.95e-07 $layer=LI1_cond $X=9.715 $Y=1.175
+ $X2=9.91 $Y2=1.175
r82 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.715
+ $Y=1.16 $X2=9.715 $Y2=1.16
r83 50 52 23.7879 $w=2.9e-07 $l=1.15e-07 $layer=POLY_cond $X=9.6 $Y=1.16
+ $X2=9.715 $Y2=1.16
r84 48 49 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=8.665 $Y=1.16
+ $X2=9.085 $Y2=1.16
r85 46 48 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=8.455 $Y=1.16
+ $X2=8.665 $Y2=1.16
r86 43 46 43.4388 $w=2.9e-07 $l=2.1e-07 $layer=POLY_cond $X=8.245 $Y=1.16
+ $X2=8.455 $Y2=1.16
r87 38 64 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=9.915 $Y=1.175
+ $X2=9.91 $Y2=1.175
r88 37 53 14.4182 $w=1.98e-07 $l=2.6e-07 $layer=LI1_cond $X=9.455 $Y=1.175
+ $X2=9.715 $Y2=1.175
r89 36 37 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=8.995 $Y=1.175
+ $X2=9.455 $Y2=1.175
r90 35 36 29.9455 $w=1.98e-07 $l=5.4e-07 $layer=LI1_cond $X=8.455 $Y=1.175
+ $X2=8.995 $Y2=1.175
r91 35 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.455
+ $Y=1.16 $X2=8.455 $Y2=1.16
r92 31 50 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=9.6 $Y=1.305
+ $X2=9.6 $Y2=1.16
r93 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.6 $Y=1.305 $X2=9.6
+ $Y2=1.985
r94 27 50 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=9.6 $Y=1.015
+ $X2=9.6 $Y2=1.16
r95 27 29 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.6 $Y=1.015
+ $X2=9.6 $Y2=0.56
r96 26 49 15.5139 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=9.16 $Y=1.16
+ $X2=9.085 $Y2=1.16
r97 25 50 15.5139 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=9.525 $Y=1.16
+ $X2=9.6 $Y2=1.16
r98 25 26 75.5008 $w=2.9e-07 $l=3.65e-07 $layer=POLY_cond $X=9.525 $Y=1.16
+ $X2=9.16 $Y2=1.16
r99 21 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=9.085 $Y=1.305
+ $X2=9.085 $Y2=1.16
r100 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.085 $Y=1.305
+ $X2=9.085 $Y2=1.985
r101 17 49 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=9.085 $Y=1.015
+ $X2=9.085 $Y2=1.16
r102 17 19 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.085 $Y=1.015
+ $X2=9.085 $Y2=0.56
r103 13 48 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.665 $Y=1.305
+ $X2=8.665 $Y2=1.16
r104 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.665 $Y=1.305
+ $X2=8.665 $Y2=1.985
r105 9 48 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.665 $Y=1.015
+ $X2=8.665 $Y2=1.16
r106 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=8.665 $Y=1.015
+ $X2=8.665 $Y2=0.56
r107 5 43 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.245 $Y=1.305
+ $X2=8.245 $Y2=1.16
r108 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.245 $Y=1.305
+ $X2=8.245 $Y2=1.985
r109 1 43 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.245 $Y=1.015
+ $X2=8.245 $Y2=1.16
r110 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=8.245 $Y=1.015
+ $X2=8.245 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 31 32 33
+ 36 38 40 42 47 49
r65 40 51 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=2.005
+ $X2=3.675 $Y2=1.92
r66 40 42 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.675 $Y=2.005
+ $X2=3.675 $Y2=2.26
r67 39 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=1.92
+ $X2=2.795 $Y2=1.92
r68 38 51 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.55 $Y=1.92
+ $X2=3.675 $Y2=1.92
r69 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.55 $Y=1.92
+ $X2=2.88 $Y2=1.92
r70 34 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=2.005
+ $X2=2.795 $Y2=1.92
r71 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.795 $Y=2.005
+ $X2=2.795 $Y2=2.26
r72 32 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=1.92
+ $X2=2.795 $Y2=1.92
r73 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.71 $Y=1.92
+ $X2=2.04 $Y2=1.92
r74 29 31 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=2.255
+ $X2=1.955 $Y2=2.17
r75 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=2.005
+ $X2=2.04 $Y2=1.92
r76 28 31 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=2.005
+ $X2=1.955 $Y2=2.17
r77 27 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.36 $X2=1.1
+ $Y2=2.36
r78 26 29 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.87 $Y=2.36
+ $X2=1.955 $Y2=2.255
r79 26 27 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=1.87 $Y=2.36
+ $X2=1.185 $Y2=2.36
r80 22 47 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.1 $Y=2.255 $X2=1.1
+ $Y2=2.36
r81 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.1 $Y=2.255
+ $X2=1.1 $Y2=2
r82 21 45 3.79048 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=2.36
+ $X2=0.217 $Y2=2.36
r83 20 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.36 $X2=1.1
+ $Y2=2.36
r84 20 21 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=2.36
+ $X2=0.345 $Y2=2.36
r85 16 45 3.10938 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=0.217 $Y=2.255
+ $X2=0.217 $Y2=2.36
r86 16 18 26.8903 $w=2.53e-07 $l=5.95e-07 $layer=LI1_cond $X=0.217 $Y=2.255
+ $X2=0.217 $Y2=1.66
r87 5 51 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.485 $X2=3.635 $Y2=1.92
r88 5 42 600 $w=1.7e-07 $l=8.39792e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.485 $X2=3.635 $Y2=2.26
r89 4 49 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.485 $X2=2.795 $Y2=1.92
r90 4 36 600 $w=1.7e-07 $l=8.39792e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.485 $X2=2.795 $Y2=2.26
r91 3 31 600 $w=1.7e-07 $l=7.5629e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.955 $Y2=2.17
r92 2 47 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r93 2 24 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r94 1 45 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r95 1 18 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%Y 1 2 3 4 5 6 7 8 25 33 36 41 43 44 47 52 57
+ 59 61 62
c116 41 0 7.99167e-20 $X=3.215 $Y=0.74
r117 54 62 6.84785 $w=3.43e-07 $l=2.05e-07 $layer=LI1_cond $X=1.527 $Y=1.665
+ $X2=1.527 $Y2=1.87
r118 54 56 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.52 $Y=1.58
+ $X2=1.945 $Y2=1.58
r119 48 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=1.58
+ $X2=4.575 $Y2=1.58
r120 47 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.25 $Y=1.58
+ $X2=5.415 $Y2=1.58
r121 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.25 $Y=1.58
+ $X2=4.74 $Y2=1.58
r122 44 56 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.035 $Y=1.58
+ $X2=1.945 $Y2=1.58
r123 43 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=1.58
+ $X2=4.575 $Y2=1.58
r124 43 44 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=4.41 $Y=1.58
+ $X2=2.035 $Y2=1.58
r125 39 41 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=2.375 $Y=0.78
+ $X2=3.215 $Y2=0.78
r126 37 57 3.89906 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.035 $Y=0.78
+ $X2=1.945 $Y2=0.78
r127 37 39 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.035 $Y=0.78
+ $X2=2.375 $Y2=0.78
r128 36 56 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=1.495
+ $X2=1.945 $Y2=1.58
r129 35 57 2.54814 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.945 $Y=0.905
+ $X2=1.945 $Y2=0.78
r130 35 36 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=1.945 $Y=0.905
+ $X2=1.945 $Y2=1.495
r131 34 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.58
+ $X2=0.68 $Y2=1.58
r132 33 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.58
+ $X2=1.52 $Y2=1.58
r133 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.58
+ $X2=0.845 $Y2=1.58
r134 27 30 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=0.68 $Y=0.78
+ $X2=1.52 $Y2=0.78
r135 25 57 3.89906 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.855 $Y=0.78
+ $X2=1.945 $Y2=0.78
r136 25 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.855 $Y=0.78
+ $X2=1.52 $Y2=0.78
r137 8 61 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=5.28
+ $Y=1.485 $X2=5.415 $Y2=1.66
r138 7 59 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=1.485 $X2=4.575 $Y2=1.66
r139 6 54 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r140 5 52 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r141 4 41 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.235 $X2=3.215 $Y2=0.74
r142 3 39 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.375 $Y2=0.74
r143 2 30 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.74
r144 1 27 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%VPWR 1 2 3 4 5 18 22 26 30 32 34 39 40 42 43
+ 45 46 48 49 50 71 77
r144 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r145 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r146 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r147 71 76 5.52694 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=9.63 $Y=2.72
+ $X2=9.875 $Y2=2.72
r148 71 73 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.63 $Y=2.72 $X2=9.43
+ $Y2=2.72
r149 70 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r150 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r151 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r152 66 67 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r153 64 67 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=7.59 $Y2=2.72
r154 63 66 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=7.59 $Y2=2.72
r155 63 64 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r156 61 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r157 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r158 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r159 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r160 53 57 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r161 50 58 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r162 50 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r163 48 69 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.79 $Y=2.72
+ $X2=8.51 $Y2=2.72
r164 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.79 $Y=2.72
+ $X2=8.875 $Y2=2.72
r165 47 73 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=8.96 $Y=2.72
+ $X2=9.43 $Y2=2.72
r166 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=2.72
+ $X2=8.875 $Y2=2.72
r167 45 66 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.87 $Y=2.72
+ $X2=7.59 $Y2=2.72
r168 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.87 $Y=2.72
+ $X2=7.995 $Y2=2.72
r169 44 69 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.12 $Y=2.72
+ $X2=8.51 $Y2=2.72
r170 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.12 $Y=2.72
+ $X2=7.995 $Y2=2.72
r171 42 60 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.05 $Y=2.72 $X2=2.99
+ $Y2=2.72
r172 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=2.72
+ $X2=3.215 $Y2=2.72
r173 41 63 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.38 $Y=2.72 $X2=3.45
+ $Y2=2.72
r174 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=2.72
+ $X2=3.215 $Y2=2.72
r175 39 57 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.07 $Y2=2.72
r176 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.72
+ $X2=2.375 $Y2=2.72
r177 38 60 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.54 $Y=2.72
+ $X2=2.99 $Y2=2.72
r178 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=2.72
+ $X2=2.375 $Y2=2.72
r179 34 37 19.3497 $w=4.03e-07 $l=6.8e-07 $layer=LI1_cond $X=9.832 $Y=1.66
+ $X2=9.832 $Y2=2.34
r180 32 76 2.88754 $w=4.05e-07 $l=1.04307e-07 $layer=LI1_cond $X=9.832 $Y=2.635
+ $X2=9.875 $Y2=2.72
r181 32 37 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=9.832 $Y=2.635
+ $X2=9.832 $Y2=2.34
r182 28 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.875 $Y=2.635
+ $X2=8.875 $Y2=2.72
r183 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.875 $Y=2.635
+ $X2=8.875 $Y2=2
r184 24 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.995 $Y=2.635
+ $X2=7.995 $Y2=2.72
r185 24 26 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.995 $Y=2.635
+ $X2=7.995 $Y2=2
r186 20 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.635
+ $X2=3.215 $Y2=2.72
r187 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.215 $Y=2.635
+ $X2=3.215 $Y2=2.34
r188 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.635
+ $X2=2.375 $Y2=2.72
r189 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.375 $Y=2.635
+ $X2=2.375 $Y2=2.34
r190 5 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=1.485 $X2=9.81 $Y2=2.34
r191 5 34 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=1.485 $X2=9.81 $Y2=1.66
r192 4 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.74
+ $Y=1.485 $X2=8.875 $Y2=2
r193 3 26 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=7.91
+ $Y=1.485 $X2=8.035 $Y2=2
r194 2 22 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.485 $X2=3.215 $Y2=2.34
r195 1 18 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.485 $X2=2.375 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%A_806_297# 1 2 3 4 5 16 18 20 24 26 32 36 38
+ 40 42 47 49 51
r62 40 53 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.555 $Y=2.255
+ $X2=7.555 $Y2=2.36
r63 40 42 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.555 $Y=2.255
+ $X2=7.555 $Y2=2
r64 39 51 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=2.36 $X2=6.675
+ $Y2=2.36
r65 38 53 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=7.43 $Y=2.36
+ $X2=7.555 $Y2=2.36
r66 38 39 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=7.43 $Y=2.36
+ $X2=6.76 $Y2=2.36
r67 34 51 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.675 $Y=2.255
+ $X2=6.675 $Y2=2.36
r68 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.675 $Y=2.255
+ $X2=6.675 $Y2=2
r69 33 49 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.36 $X2=5.835
+ $Y2=2.36
r70 32 51 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=2.36 $X2=6.675
+ $Y2=2.36
r71 32 33 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=6.59 $Y=2.36
+ $X2=5.92 $Y2=2.36
r72 28 49 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.835 $Y=2.255
+ $X2=5.835 $Y2=2.36
r73 28 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.835 $Y=2.255
+ $X2=5.835 $Y2=2
r74 27 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=2.36 $X2=4.995
+ $Y2=2.36
r75 26 49 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.75 $Y=2.36 $X2=5.835
+ $Y2=2.36
r76 26 27 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=5.75 $Y=2.36
+ $X2=5.08 $Y2=2.36
r77 22 47 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.995 $Y=2.255
+ $X2=4.995 $Y2=2.36
r78 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.995 $Y=2.255
+ $X2=4.995 $Y2=2
r79 21 45 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.24 $Y=2.36
+ $X2=4.115 $Y2=2.36
r80 20 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=2.36 $X2=4.995
+ $Y2=2.36
r81 20 21 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=4.91 $Y=2.36
+ $X2=4.24 $Y2=2.36
r82 16 45 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.115 $Y=2.255
+ $X2=4.115 $Y2=2.36
r83 16 18 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.115 $Y=2.255
+ $X2=4.115 $Y2=2
r84 5 53 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.38
+ $Y=1.485 $X2=7.515 $Y2=2.34
r85 5 42 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=7.38
+ $Y=1.485 $X2=7.515 $Y2=2
r86 4 51 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.54
+ $Y=1.485 $X2=6.675 $Y2=2.34
r87 4 36 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=6.54
+ $Y=1.485 $X2=6.675 $Y2=2
r88 3 49 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.485 $X2=5.835 $Y2=2.34
r89 3 30 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.485 $X2=5.835 $Y2=2
r90 2 47 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.86
+ $Y=1.485 $X2=4.995 $Y2=2.34
r91 2 24 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=4.86
+ $Y=1.485 $X2=4.995 $Y2=2
r92 1 45 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.485 $X2=4.155 $Y2=2.34
r93 1 18 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.485 $X2=4.155 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%A_1224_297# 1 2 3 4 15 19 23 25 27 29 32 34
+ 36
r63 27 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=1.665
+ $X2=9.295 $Y2=1.58
r64 27 29 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.295 $Y=1.665
+ $X2=9.295 $Y2=2.34
r65 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=1.58
+ $X2=8.455 $Y2=1.58
r66 25 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.13 $Y=1.58
+ $X2=9.295 $Y2=1.58
r67 25 26 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.13 $Y=1.58
+ $X2=8.62 $Y2=1.58
r68 21 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.455 $Y=1.665
+ $X2=8.455 $Y2=1.58
r69 21 23 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.455 $Y=1.665
+ $X2=8.455 $Y2=2.34
r70 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=1.58
+ $X2=7.095 $Y2=1.58
r71 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.29 $Y=1.58
+ $X2=8.455 $Y2=1.58
r72 19 20 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=8.29 $Y=1.58
+ $X2=7.26 $Y2=1.58
r73 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.42 $Y=1.58
+ $X2=6.255 $Y2=1.58
r74 15 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=1.58
+ $X2=7.095 $Y2=1.58
r75 15 16 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.93 $Y=1.58
+ $X2=6.42 $Y2=1.58
r76 4 38 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.485 $X2=9.295 $Y2=1.66
r77 4 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.485 $X2=9.295 $Y2=2.34
r78 3 36 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.32
+ $Y=1.485 $X2=8.455 $Y2=1.66
r79 3 23 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.32
+ $Y=1.485 $X2=8.455 $Y2=2.34
r80 2 34 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=6.96
+ $Y=1.485 $X2=7.095 $Y2=1.66
r81 1 32 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=6.12
+ $Y=1.485 $X2=6.255 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%A_27_47# 1 2 3 4 5 6 7 8 9 10 11 34 36 38 46
+ 47 48 52 56 60 64 68 70 74 82 85 86 87 90 91 92
c166 47 0 1.79953e-19 $X=3.675 $Y=0.735
r167 89 91 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=0.58
+ $X2=8.04 $Y2=0.58
r168 89 90 17.1064 $w=6.48e-07 $l=5.25e-07 $layer=LI1_cond $X=7.875 $Y=0.58
+ $X2=7.35 $Y2=0.58
r169 84 86 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0.58
+ $X2=5.98 $Y2=0.58
r170 84 85 16.7383 $w=6.48e-07 $l=5.05e-07 $layer=LI1_cond $X=5.815 $Y=0.58
+ $X2=5.31 $Y2=0.58
r171 72 74 10.4902 $w=3.88e-07 $l=3.55e-07 $layer=LI1_cond $X=9.84 $Y=0.735
+ $X2=9.84 $Y2=0.38
r172 71 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.04 $Y=0.82
+ $X2=8.875 $Y2=0.82
r173 70 72 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=9.645 $Y=0.82
+ $X2=9.84 $Y2=0.735
r174 70 71 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.645 $Y=0.82
+ $X2=9.04 $Y2=0.82
r175 66 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.875 $Y=0.735
+ $X2=8.875 $Y2=0.82
r176 66 68 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=8.875 $Y=0.735
+ $X2=8.875 $Y2=0.38
r177 64 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.71 $Y=0.82
+ $X2=8.875 $Y2=0.82
r178 64 91 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.71 $Y=0.82
+ $X2=8.04 $Y2=0.82
r179 63 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.84 $Y=0.82
+ $X2=6.675 $Y2=0.82
r180 63 90 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.84 $Y=0.82
+ $X2=7.35 $Y2=0.82
r181 58 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=0.735
+ $X2=6.675 $Y2=0.82
r182 58 60 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.675 $Y=0.735
+ $X2=6.675 $Y2=0.38
r183 56 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.51 $Y=0.82
+ $X2=6.675 $Y2=0.82
r184 56 86 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.51 $Y=0.82
+ $X2=5.98 $Y2=0.82
r185 55 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=0.82
+ $X2=4.475 $Y2=0.82
r186 55 85 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.64 $Y=0.82
+ $X2=5.31 $Y2=0.82
r187 50 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.735
+ $X2=4.475 $Y2=0.82
r188 50 52 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.475 $Y=0.735
+ $X2=4.475 $Y2=0.38
r189 49 81 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.8 $Y=0.82
+ $X2=3.675 $Y2=0.82
r190 48 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=0.82
+ $X2=4.475 $Y2=0.82
r191 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.31 $Y=0.82
+ $X2=3.8 $Y2=0.82
r192 47 81 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=0.735
+ $X2=3.675 $Y2=0.82
r193 46 79 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.675 $Y=0.465
+ $X2=3.675 $Y2=0.36
r194 46 47 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=3.675 $Y=0.465
+ $X2=3.675 $Y2=0.735
r195 43 45 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=1.94 $Y=0.36
+ $X2=2.795 $Y2=0.36
r196 41 43 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=0.36
+ $X2=1.94 $Y2=0.36
r197 39 77 3.79048 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.36
+ $X2=0.217 $Y2=0.36
r198 39 41 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=0.345 $Y=0.36
+ $X2=1.1 $Y2=0.36
r199 38 79 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.55 $Y=0.36
+ $X2=3.675 $Y2=0.36
r200 38 45 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=3.55 $Y=0.36
+ $X2=2.795 $Y2=0.36
r201 34 77 3.10938 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.217 $Y2=0.36
r202 34 36 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.217 $Y2=0.72
r203 11 74 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=9.675
+ $Y=0.235 $X2=9.81 $Y2=0.38
r204 10 68 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=8.74
+ $Y=0.235 $X2=8.875 $Y2=0.38
r205 9 89 45.5 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=4 $X=7.38
+ $Y=0.235 $X2=7.875 $Y2=0.38
r206 8 60 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.54
+ $Y=0.235 $X2=6.675 $Y2=0.38
r207 7 84 45.5 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_NDIFF $count=4 $X=5.34
+ $Y=0.235 $X2=5.815 $Y2=0.38
r208 6 52 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.34
+ $Y=0.235 $X2=4.475 $Y2=0.38
r209 5 81 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.235 $X2=3.635 $Y2=0.74
r210 5 79 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.235 $X2=3.635 $Y2=0.38
r211 4 45 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.66
+ $Y=0.235 $X2=2.795 $Y2=0.38
r212 3 43 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r213 2 41 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r214 1 77 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r215 1 36 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_4%VGND 1 2 3 4 5 6 21 23 27 31 35 39 43 45 46
+ 48 49 51 52 53 62 67 80 81 84 87 90
r135 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r136 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r137 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r138 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r139 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r140 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r141 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r142 75 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=7.13
+ $Y2=0
r143 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r144 72 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=0 $X2=7.095
+ $Y2=0
r145 72 74 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=7.18 $Y=0 $X2=8.05
+ $Y2=0
r146 71 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r147 71 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r148 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r149 68 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.34 $Y=0 $X2=6.255
+ $Y2=0
r150 68 70 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=6.67
+ $Y2=0
r151 67 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=0 $X2=7.095
+ $Y2=0
r152 67 70 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=0 $X2=6.67
+ $Y2=0
r153 66 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r154 66 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r155 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r156 63 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=4.975
+ $Y2=0
r157 63 65 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.29
+ $Y2=0
r158 62 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=0 $X2=6.255
+ $Y2=0
r159 62 65 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=6.17 $Y=0 $X2=5.29
+ $Y2=0
r160 61 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r161 60 61 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r162 56 60 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=3.91
+ $Y2=0
r163 53 61 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=3.91
+ $Y2=0
r164 53 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r165 51 77 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.21 $Y=0 $X2=8.97
+ $Y2=0
r166 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.21 $Y=0 $X2=9.34
+ $Y2=0
r167 50 80 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.89
+ $Y2=0
r168 50 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.34
+ $Y2=0
r169 48 74 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.37 $Y=0 $X2=8.05
+ $Y2=0
r170 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.37 $Y=0 $X2=8.455
+ $Y2=0
r171 47 77 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.54 $Y=0 $X2=8.97
+ $Y2=0
r172 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.54 $Y=0 $X2=8.455
+ $Y2=0
r173 45 60 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.91
+ $Y2=0
r174 45 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.055
+ $Y2=0
r175 41 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=0.085
+ $X2=9.34 $Y2=0
r176 41 43 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=9.34 $Y=0.085
+ $X2=9.34 $Y2=0.38
r177 37 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.455 $Y=0.085
+ $X2=8.455 $Y2=0
r178 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.455 $Y=0.085
+ $X2=8.455 $Y2=0.38
r179 33 90 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.095 $Y2=0
r180 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.095 $Y2=0.38
r181 29 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0
r182 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0.38
r183 25 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=0.085
+ $X2=4.975 $Y2=0
r184 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.975 $Y=0.085
+ $X2=4.975 $Y2=0.38
r185 24 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.055
+ $Y2=0
r186 23 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.81 $Y=0 $X2=4.975
+ $Y2=0
r187 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.81 $Y=0 $X2=4.14
+ $Y2=0
r188 19 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0
r189 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0.38
r190 6 43 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.235 $X2=9.34 $Y2=0.38
r191 5 39 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.32
+ $Y=0.235 $X2=8.455 $Y2=0.38
r192 4 35 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.96
+ $Y=0.235 $X2=7.095 $Y2=0.38
r193 3 31 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.235 $X2=6.255 $Y2=0.38
r194 2 27 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=4.76
+ $Y=0.235 $X2=4.975 $Y2=0.38
r195 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.235 $X2=4.055 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__a32o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 VPWR A3 a_299_297# VPB phighvt w=1e+06u l=150000u
+  ad=9.6e+11p pd=7.92e+06u as=8e+11p ps=7.6e+06u
M1001 a_299_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_21_199# B1 a_352_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.3075e+11p ps=2.01e+06u
M1003 a_665_47# A2 a_549_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=2.795e+11p ps=2.16e+06u
M1004 X a_21_199# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.2e+11p pd=5.04e+06u as=0p ps=0u
M1005 VGND A3 a_665_47# VNB nshort w=650000u l=150000u
+  ad=7.5725e+11p pd=6.23e+06u as=0p ps=0u
M1006 VGND a_21_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1007 a_549_47# A1 a_21_199# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_352_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_299_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_21_199# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_299_297# B1 a_21_199# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1012 a_21_199# B2 a_299_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_21_199# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


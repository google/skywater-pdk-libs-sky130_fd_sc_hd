* File: sky130_fd_sc_hd__and4b_4.spice
* Created: Thu Aug 27 14:08:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and4b_4.spice.pex"
.subckt sky130_fd_sc_hd__and4b_4  VNB VPB A_N D C B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_A_N_M1016_g N_A_27_47#_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_174_21#_M1002_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11785 PD=0.92 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1002_d N_A_174_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_174_21#_M1007_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.3
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1017 N_X_M1007_d N_A_174_21#_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.212875 PD=0.92 PS=1.305 NRD=0 NRS=5.532 M=1 R=4.33333
+ SA=75001.7 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1011 A_617_47# N_D_M1011_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.212875 PD=0.92 PS=1.305 NRD=14.76 NRS=63.684 M=1 R=4.33333 SA=75002.6
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1008 A_701_47# N_C_M1008_g A_617_47# VNB NSHORT L=0.15 W=0.65 AD=0.1365
+ AS=0.08775 PD=1.07 PS=0.92 NRD=28.608 NRS=14.76 M=1 R=4.33333 SA=75003
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1015 A_815_47# N_B_M1015_g A_701_47# VNB NSHORT L=0.15 W=0.65 AD=0.143
+ AS=0.1365 PD=1.09 PS=1.07 NRD=30.456 NRS=28.608 M=1 R=4.33333 SA=75003.5
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_174_21#_M1005_d N_A_27_47#_M1005_g A_815_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.143 PD=1.82 PS=1.09 NRD=0 NRS=30.456 M=1 R=4.33333 SA=75004.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VPWR_M1009_d N_A_N_M1009_g N_A_27_47#_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0832606 AS=0.1092 PD=0.783803 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004.3 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1009_d N_A_174_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.198239 AS=0.135 PD=1.8662 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75000.4 SB=75003.8 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_174_21#_M1003_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1003_d N_A_174_21#_M1013_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75003 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A_174_21#_M1014_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3275 AS=0.135 PD=1.655 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75002.6 A=0.15 P=2.3 MULT=1
MM1012 N_A_174_21#_M1012_d N_D_M1012_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.3275 PD=1.27 PS=1.655 NRD=0 NRS=74.8403 M=1 R=6.66667 SA=75002.4
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_C_M1010_g N_A_174_21#_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.135 PD=1.42 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1006 N_A_174_21#_M1006_d N_B_M1006_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.22 AS=0.21 PD=1.44 PS=1.42 NRD=32.4853 NRS=28.565 M=1 R=6.66667
+ SA=75003.4 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_27_47#_M1000_g N_A_174_21#_M1006_d VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.22 PD=2.52 PS=1.44 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=8.7312 P=14.09
c_81 VPB 0 1.34065e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__and4b_4.spice.SKY130_FD_SC_HD__AND4B_4.pxi"
*
.ends
*
*

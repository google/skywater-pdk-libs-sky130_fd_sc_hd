* File: sky130_fd_sc_hd__einvn_8.pxi.spice
* Created: Tue Sep  1 19:08:07 2020
* 
x_PM_SKY130_FD_SC_HD__EINVN_8%TE_B N_TE_B_c_143_n N_TE_B_M1030_g N_TE_B_M1023_g
+ N_TE_B_c_144_n N_TE_B_c_150_n N_TE_B_M1000_g N_TE_B_c_151_n N_TE_B_c_152_n
+ N_TE_B_M1005_g N_TE_B_c_153_n N_TE_B_c_154_n N_TE_B_M1006_g N_TE_B_c_155_n
+ N_TE_B_c_156_n N_TE_B_M1010_g N_TE_B_c_157_n N_TE_B_c_158_n N_TE_B_M1013_g
+ N_TE_B_c_159_n N_TE_B_c_160_n N_TE_B_M1016_g N_TE_B_c_161_n N_TE_B_c_162_n
+ N_TE_B_M1024_g N_TE_B_c_163_n N_TE_B_c_164_n N_TE_B_M1028_g N_TE_B_c_145_n
+ N_TE_B_c_166_n N_TE_B_c_167_n N_TE_B_c_168_n N_TE_B_c_169_n N_TE_B_c_170_n
+ N_TE_B_c_171_n TE_B N_TE_B_c_147_n PM_SKY130_FD_SC_HD__EINVN_8%TE_B
x_PM_SKY130_FD_SC_HD__EINVN_8%A_27_47# N_A_27_47#_M1030_s N_A_27_47#_M1023_s
+ N_A_27_47#_c_274_n N_A_27_47#_M1008_g N_A_27_47#_c_275_n N_A_27_47#_c_276_n
+ N_A_27_47#_c_277_n N_A_27_47#_M1009_g N_A_27_47#_c_278_n N_A_27_47#_c_279_n
+ N_A_27_47#_M1012_g N_A_27_47#_c_280_n N_A_27_47#_c_281_n N_A_27_47#_M1014_g
+ N_A_27_47#_c_282_n N_A_27_47#_c_283_n N_A_27_47#_M1015_g N_A_27_47#_c_284_n
+ N_A_27_47#_c_285_n N_A_27_47#_M1017_g N_A_27_47#_c_286_n N_A_27_47#_c_287_n
+ N_A_27_47#_M1018_g N_A_27_47#_c_288_n N_A_27_47#_c_289_n N_A_27_47#_M1021_g
+ N_A_27_47#_c_290_n N_A_27_47#_c_291_n N_A_27_47#_c_292_n N_A_27_47#_c_293_n
+ N_A_27_47#_c_294_n N_A_27_47#_c_295_n N_A_27_47#_c_296_n N_A_27_47#_c_301_n
+ N_A_27_47#_c_297_n N_A_27_47#_c_298_n N_A_27_47#_c_302_n N_A_27_47#_c_299_n
+ N_A_27_47#_c_343_n N_A_27_47#_c_300_n PM_SKY130_FD_SC_HD__EINVN_8%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVN_8%A N_A_c_438_n N_A_M1002_g N_A_M1001_g N_A_c_439_n
+ N_A_M1003_g N_A_M1007_g N_A_c_440_n N_A_M1004_g N_A_M1019_g N_A_c_441_n
+ N_A_M1011_g N_A_M1020_g N_A_c_442_n N_A_M1027_g N_A_M1022_g N_A_c_443_n
+ N_A_M1031_g N_A_M1025_g N_A_c_444_n N_A_M1032_g N_A_M1026_g N_A_c_445_n
+ N_A_M1033_g N_A_M1029_g A A A A A A A N_A_c_447_n
+ PM_SKY130_FD_SC_HD__EINVN_8%A
x_PM_SKY130_FD_SC_HD__EINVN_8%VPWR N_VPWR_M1023_d N_VPWR_M1005_d N_VPWR_M1010_d
+ N_VPWR_M1016_d N_VPWR_M1028_d N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n
+ N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n
+ N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n VPWR N_VPWR_c_583_n
+ N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_571_n N_VPWR_c_587_n N_VPWR_c_588_n
+ PM_SKY130_FD_SC_HD__EINVN_8%VPWR
x_PM_SKY130_FD_SC_HD__EINVN_8%A_204_309# N_A_204_309#_M1000_s
+ N_A_204_309#_M1006_s N_A_204_309#_M1013_s N_A_204_309#_M1024_s
+ N_A_204_309#_M1001_s N_A_204_309#_M1007_s N_A_204_309#_M1020_s
+ N_A_204_309#_M1025_s N_A_204_309#_M1029_s N_A_204_309#_c_704_n
+ N_A_204_309#_c_692_n N_A_204_309#_c_693_n N_A_204_309#_c_761_n
+ N_A_204_309#_c_694_n N_A_204_309#_c_765_n N_A_204_309#_c_695_n
+ N_A_204_309#_c_769_n N_A_204_309#_c_696_n N_A_204_309#_c_697_n
+ N_A_204_309#_c_740_n N_A_204_309#_c_698_n N_A_204_309#_c_798_p
+ N_A_204_309#_c_742_n N_A_204_309#_c_803_p N_A_204_309#_c_744_n
+ N_A_204_309#_c_807_p N_A_204_309#_c_699_n N_A_204_309#_c_700_n
+ N_A_204_309#_c_701_n N_A_204_309#_c_702_n N_A_204_309#_c_703_n
+ N_A_204_309#_c_785_n N_A_204_309#_c_787_n N_A_204_309#_c_789_n
+ PM_SKY130_FD_SC_HD__EINVN_8%A_204_309#
x_PM_SKY130_FD_SC_HD__EINVN_8%Z N_Z_M1002_s N_Z_M1004_s N_Z_M1027_s N_Z_M1032_s
+ N_Z_M1001_d N_Z_M1019_d N_Z_M1022_d N_Z_M1026_d N_Z_c_826_n N_Z_c_817_n
+ N_Z_c_818_n N_Z_c_837_n N_Z_c_819_n N_Z_c_820_n N_Z_c_821_n N_Z_c_822_n
+ N_Z_c_823_n N_Z_c_824_n Z Z Z Z N_Z_c_873_n N_Z_c_877_n N_Z_c_815_n Z
+ PM_SKY130_FD_SC_HD__EINVN_8%Z
x_PM_SKY130_FD_SC_HD__EINVN_8%VGND N_VGND_M1030_d N_VGND_M1008_s N_VGND_M1012_s
+ N_VGND_M1015_s N_VGND_M1018_s N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n
+ N_VGND_c_928_n N_VGND_c_929_n N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n
+ N_VGND_c_933_n VGND N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n
+ N_VGND_c_937_n N_VGND_c_938_n N_VGND_c_939_n N_VGND_c_940_n N_VGND_c_941_n
+ PM_SKY130_FD_SC_HD__EINVN_8%VGND
x_PM_SKY130_FD_SC_HD__EINVN_8%A_215_47# N_A_215_47#_M1008_d N_A_215_47#_M1009_d
+ N_A_215_47#_M1014_d N_A_215_47#_M1017_d N_A_215_47#_M1021_d
+ N_A_215_47#_M1003_d N_A_215_47#_M1011_d N_A_215_47#_M1031_d
+ N_A_215_47#_M1033_d N_A_215_47#_c_1049_n N_A_215_47#_c_1055_n
+ N_A_215_47#_c_1050_n N_A_215_47#_c_1120_n N_A_215_47#_c_1061_n
+ N_A_215_47#_c_1127_n N_A_215_47#_c_1065_n N_A_215_47#_c_1134_n
+ N_A_215_47#_c_1069_n N_A_215_47#_c_1141_n N_A_215_47#_c_1073_n
+ N_A_215_47#_c_1051_n N_A_215_47#_c_1074_n N_A_215_47#_c_1076_n
+ N_A_215_47#_c_1078_n PM_SKY130_FD_SC_HD__EINVN_8%A_215_47#
cc_1 VNB N_TE_B_c_143_n 0.0250205f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_TE_B_c_144_n 0.0136319f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.25
cc_3 VNB N_TE_B_c_145_n 0.0100604f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.25
cc_4 VNB TE_B 0.0135404f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_TE_B_c_147_n 0.0362295f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_6 VNB N_A_27_47#_c_274_n 0.0175424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_275_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.47
cc_8 VNB N_A_27_47#_c_276_n 0.00831588f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=2.015
cc_9 VNB N_A_27_47#_c_277_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=2.015
cc_10 VNB N_A_27_47#_c_278_n 0.00891962f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.47
cc_11 VNB N_A_27_47#_c_279_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_12 VNB N_A_27_47#_c_280_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.47
cc_13 VNB N_A_27_47#_c_281_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=2.015
cc_14 VNB N_A_27_47#_c_282_n 0.00891962f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=1.47
cc_15 VNB N_A_27_47#_c_283_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=2.015
cc_16 VNB N_A_27_47#_c_284_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=1.47
cc_17 VNB N_A_27_47#_c_285_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=2.015
cc_18 VNB N_A_27_47#_c_286_n 0.00891962f $X=-0.19 $Y=-0.24 $X2=3.045 $Y2=1.47
cc_19 VNB N_A_27_47#_c_287_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=3.045 $Y2=2.015
cc_20 VNB N_A_27_47#_c_288_n 0.00887388f $X=-0.19 $Y=-0.24 $X2=3.465 $Y2=1.47
cc_21 VNB N_A_27_47#_c_289_n 0.014583f $X=-0.19 $Y=-0.24 $X2=3.465 $Y2=2.015
cc_22 VNB N_A_27_47#_c_290_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=3.885 $Y2=1.47
cc_23 VNB N_A_27_47#_c_291_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=3.885 $Y2=2.015
cc_24 VNB N_A_27_47#_c_292_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=3.885 $Y2=2.015
cc_25 VNB N_A_27_47#_c_293_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.25
cc_26 VNB N_A_27_47#_c_294_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_295_n 0.00473803f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.395
cc_28 VNB N_A_27_47#_c_296_n 0.0155191f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.395
cc_29 VNB N_A_27_47#_c_297_n 0.00942441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_298_n 0.0030044f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_31 VNB N_A_27_47#_c_299_n 0.0117143f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_32 VNB N_A_27_47#_c_300_n 0.0213763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_c_438_n 0.0167495f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_34 VNB N_A_c_439_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.25
cc_35 VNB N_A_c_440_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.47
cc_36 VNB N_A_c_441_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=2.015
cc_37 VNB N_A_c_442_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=2.28 $Y2=1.395
cc_38 VNB N_A_c_443_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=3.045 $Y2=2.015
cc_39 VNB N_A_c_444_n 0.0160026f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=1.395
cc_40 VNB N_A_c_445_n 0.0192291f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.395
cc_41 VNB A 0.00545171f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_42 VNB N_A_c_447_n 0.129445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VPWR_c_571_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Z_c_815_n 0.00954692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB Z 0.0232765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_925_n 0.00474451f $X=-0.19 $Y=-0.24 $X2=1.71 $Y2=1.395
cc_47 VNB N_VGND_c_926_n 3.18775e-19 $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=2.015
cc_48 VNB N_VGND_c_927_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=2.015
cc_49 VNB N_VGND_c_928_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=1.47
cc_50 VNB N_VGND_c_929_n 3.95505e-19 $X=-0.19 $Y=-0.24 $X2=2.7 $Y2=1.395
cc_51 VNB N_VGND_c_930_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=3.045 $Y2=2.015
cc_52 VNB N_VGND_c_931_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=3.39 $Y2=1.395
cc_53 VNB N_VGND_c_932_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=3.465 $Y2=1.47
cc_54 VNB N_VGND_c_933_n 0.00449573f $X=-0.19 $Y=-0.24 $X2=3.465 $Y2=2.015
cc_55 VNB N_VGND_c_934_n 0.014366f $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=1.395
cc_56 VNB N_VGND_c_935_n 0.0150454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_936_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=1.395
cc_58 VNB N_VGND_c_937_n 0.0906903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_938_n 0.397812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_939_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_940_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_941_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_215_47#_c_1049_n 0.00496433f $X=-0.19 $Y=-0.24 $X2=2.55 $Y2=1.395
cc_64 VNB N_A_215_47#_c_1050_n 0.00198743f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=2.015
cc_65 VNB N_A_215_47#_c_1051_n 0.00962047f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_66 VPB N_TE_B_M1023_g 0.0257066f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_TE_B_c_144_n 0.00483829f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.25
cc_68 VPB N_TE_B_c_150_n 0.0144321f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.47
cc_69 VPB N_TE_B_c_151_n 0.013715f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.395
cc_70 VPB N_TE_B_c_152_n 0.0135568f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.47
cc_71 VPB N_TE_B_c_153_n 0.0088967f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=1.395
cc_72 VPB N_TE_B_c_154_n 0.013575f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.47
cc_73 VPB N_TE_B_c_155_n 0.00885591f $X=-0.19 $Y=1.305 $X2=2.13 $Y2=1.395
cc_74 VPB N_TE_B_c_156_n 0.013575f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=1.47
cc_75 VPB N_TE_B_c_157_n 0.0088967f $X=-0.19 $Y=1.305 $X2=2.55 $Y2=1.395
cc_76 VPB N_TE_B_c_158_n 0.013575f $X=-0.19 $Y=1.305 $X2=2.625 $Y2=1.47
cc_77 VPB N_TE_B_c_159_n 0.00885591f $X=-0.19 $Y=1.305 $X2=2.97 $Y2=1.395
cc_78 VPB N_TE_B_c_160_n 0.013575f $X=-0.19 $Y=1.305 $X2=3.045 $Y2=1.47
cc_79 VPB N_TE_B_c_161_n 0.0088967f $X=-0.19 $Y=1.305 $X2=3.39 $Y2=1.395
cc_80 VPB N_TE_B_c_162_n 0.013575f $X=-0.19 $Y=1.305 $X2=3.465 $Y2=1.47
cc_81 VPB N_TE_B_c_163_n 0.0207809f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=1.395
cc_82 VPB N_TE_B_c_164_n 0.0171184f $X=-0.19 $Y=1.305 $X2=3.885 $Y2=1.47
cc_83 VPB N_TE_B_c_145_n 0.00578605f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.25
cc_84 VPB N_TE_B_c_166_n 0.00473803f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.395
cc_85 VPB N_TE_B_c_167_n 0.00391059f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.395
cc_86 VPB N_TE_B_c_168_n 0.00391059f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=1.395
cc_87 VPB N_TE_B_c_169_n 0.00391059f $X=-0.19 $Y=1.305 $X2=2.625 $Y2=1.395
cc_88 VPB N_TE_B_c_170_n 0.00391059f $X=-0.19 $Y=1.305 $X2=3.045 $Y2=1.395
cc_89 VPB N_TE_B_c_171_n 0.00391059f $X=-0.19 $Y=1.305 $X2=3.465 $Y2=1.395
cc_90 VPB TE_B 0.00306878f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_91 VPB N_TE_B_c_147_n 0.00941639f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_92 VPB N_A_27_47#_c_301_n 0.0306167f $X=-0.19 $Y=1.305 $X2=3.465 $Y2=1.395
cc_93 VPB N_A_27_47#_c_302_n 0.00983295f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_94 VPB N_A_27_47#_c_299_n 0.00251088f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_95 VPB N_A_27_47#_c_300_n 0.00828812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_M1001_g 0.0258424f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_97 VPB N_A_M1007_g 0.0182176f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.395
cc_98 VPB N_A_M1019_g 0.0182176f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.47
cc_99 VPB N_A_M1020_g 0.0182176f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=2.015
cc_100 VPB N_A_M1022_g 0.0182176f $X=-0.19 $Y=1.305 $X2=2.7 $Y2=1.395
cc_101 VPB N_A_M1025_g 0.0182176f $X=-0.19 $Y=1.305 $X2=3.465 $Y2=2.015
cc_102 VPB N_A_M1026_g 0.0182145f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.25
cc_103 VPB N_A_M1029_g 0.0219619f $X=-0.19 $Y=1.305 $X2=3.045 $Y2=1.395
cc_104 VPB N_A_c_447_n 0.0223781f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_572_n 0.00210688f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=1.395
cc_106 VPB N_VPWR_c_573_n 3.11529e-19 $X=-0.19 $Y=1.305 $X2=1.785 $Y2=2.015
cc_107 VPB N_VPWR_c_574_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=2.205 $Y2=2.015
cc_108 VPB N_VPWR_c_575_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=2.625 $Y2=1.47
cc_109 VPB N_VPWR_c_576_n 0.00944386f $X=-0.19 $Y=1.305 $X2=2.7 $Y2=1.395
cc_110 VPB N_VPWR_c_577_n 0.0124915f $X=-0.19 $Y=1.305 $X2=3.045 $Y2=2.015
cc_111 VPB N_VPWR_c_578_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.39 $Y2=1.395
cc_112 VPB N_VPWR_c_579_n 0.0124915f $X=-0.19 $Y=1.305 $X2=3.465 $Y2=1.47
cc_113 VPB N_VPWR_c_580_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.465 $Y2=2.015
cc_114 VPB N_VPWR_c_581_n 0.0124915f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=1.395
cc_115 VPB N_VPWR_c_582_n 0.00546352f $X=-0.19 $Y=1.305 $X2=3.54 $Y2=1.395
cc_116 VPB N_VPWR_c_583_n 0.0151047f $X=-0.19 $Y=1.305 $X2=3.885 $Y2=2.015
cc_117 VPB N_VPWR_c_584_n 0.0146397f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.395
cc_118 VPB N_VPWR_c_585_n 0.0932248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_571_n 0.0521487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_587_n 0.0050755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_588_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_204_309#_c_692_n 0.00251378f $X=-0.19 $Y=1.305 $X2=2.625
+ $Y2=2.015
cc_123 VPB N_A_204_309#_c_693_n 0.0017513f $X=-0.19 $Y=1.305 $X2=2.97 $Y2=1.395
cc_124 VPB N_A_204_309#_c_694_n 0.00239417f $X=-0.19 $Y=1.305 $X2=3.39 $Y2=1.395
cc_125 VPB N_A_204_309#_c_695_n 0.00239417f $X=-0.19 $Y=1.305 $X2=3.54 $Y2=1.395
cc_126 VPB N_A_204_309#_c_696_n 0.0120425f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.395
cc_127 VPB N_A_204_309#_c_697_n 0.00645359f $X=-0.19 $Y=1.305 $X2=3.045
+ $Y2=1.395
cc_128 VPB N_A_204_309#_c_698_n 0.00178145f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_129 VPB N_A_204_309#_c_699_n 0.00820528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_204_309#_c_700_n 0.021034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_204_309#_c_701_n 0.00108194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_204_309#_c_702_n 0.00108194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_204_309#_c_703_n 0.00108194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_Z_c_817_n 0.00218546f $X=-0.19 $Y=1.305 $X2=2.28 $Y2=1.395
cc_135 VPB N_Z_c_818_n 0.00223333f $X=-0.19 $Y=1.305 $X2=2.625 $Y2=1.47
cc_136 VPB N_Z_c_819_n 0.00218546f $X=-0.19 $Y=1.305 $X2=3.045 $Y2=1.47
cc_137 VPB N_Z_c_820_n 0.00218546f $X=-0.19 $Y=1.305 $X2=3.045 $Y2=2.015
cc_138 VPB N_Z_c_821_n 0.0103765f $X=-0.19 $Y=1.305 $X2=3.12 $Y2=1.395
cc_139 VPB N_Z_c_822_n 0.00223333f $X=-0.19 $Y=1.305 $X2=3.465 $Y2=2.015
cc_140 VPB N_Z_c_823_n 0.00223333f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=1.395
cc_141 VPB N_Z_c_824_n 0.00223333f $X=-0.19 $Y=1.305 $X2=3.885 $Y2=1.47
cc_142 VPB Z 0.00770139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 N_TE_B_c_153_n N_A_27_47#_c_275_n 0.0141957f $X=1.71 $Y=1.395 $X2=0 $Y2=0
cc_144 N_TE_B_c_166_n N_A_27_47#_c_276_n 0.0141957f $X=1.365 $Y=1.395 $X2=0
+ $Y2=0
cc_145 N_TE_B_c_155_n N_A_27_47#_c_278_n 0.0141957f $X=2.13 $Y=1.395 $X2=0 $Y2=0
cc_146 N_TE_B_c_157_n N_A_27_47#_c_280_n 0.0141957f $X=2.55 $Y=1.395 $X2=0 $Y2=0
cc_147 N_TE_B_c_159_n N_A_27_47#_c_282_n 0.0141957f $X=2.97 $Y=1.395 $X2=0 $Y2=0
cc_148 N_TE_B_c_161_n N_A_27_47#_c_284_n 0.0141957f $X=3.39 $Y=1.395 $X2=0 $Y2=0
cc_149 N_TE_B_c_163_n N_A_27_47#_c_286_n 0.0141957f $X=3.81 $Y=1.395 $X2=0 $Y2=0
cc_150 N_TE_B_c_167_n N_A_27_47#_c_290_n 0.0141957f $X=1.785 $Y=1.395 $X2=0
+ $Y2=0
cc_151 N_TE_B_c_168_n N_A_27_47#_c_291_n 0.0141957f $X=2.205 $Y=1.395 $X2=0
+ $Y2=0
cc_152 N_TE_B_c_169_n N_A_27_47#_c_292_n 0.0141957f $X=2.625 $Y=1.395 $X2=0
+ $Y2=0
cc_153 N_TE_B_c_170_n N_A_27_47#_c_293_n 0.0141957f $X=3.045 $Y=1.395 $X2=0
+ $Y2=0
cc_154 N_TE_B_c_171_n N_A_27_47#_c_294_n 0.0141957f $X=3.465 $Y=1.395 $X2=0
+ $Y2=0
cc_155 N_TE_B_c_143_n N_A_27_47#_c_297_n 0.0138539f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_156 N_TE_B_c_144_n N_A_27_47#_c_297_n 9.15163e-19 $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_157 TE_B N_A_27_47#_c_297_n 0.0186928f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_158 N_TE_B_c_147_n N_A_27_47#_c_297_n 0.00163649f $X=0.545 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_TE_B_c_143_n N_A_27_47#_c_298_n 0.0108991f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_160 N_TE_B_M1023_g N_A_27_47#_c_302_n 0.0254542f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_161 N_TE_B_c_144_n N_A_27_47#_c_302_n 7.21838e-19 $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_162 N_TE_B_c_150_n N_A_27_47#_c_302_n 0.00105498f $X=0.945 $Y=1.47 $X2=0
+ $Y2=0
cc_163 N_TE_B_c_145_n N_A_27_47#_c_302_n 0.00517984f $X=0.945 $Y=1.25 $X2=0
+ $Y2=0
cc_164 TE_B N_A_27_47#_c_302_n 0.0186928f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_165 N_TE_B_c_147_n N_A_27_47#_c_302_n 0.00163649f $X=0.545 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_TE_B_c_144_n N_A_27_47#_c_299_n 0.00183428f $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_167 N_TE_B_c_151_n N_A_27_47#_c_299_n 0.00881838f $X=1.29 $Y=1.395 $X2=0
+ $Y2=0
cc_168 N_TE_B_c_153_n N_A_27_47#_c_299_n 0.0058575f $X=1.71 $Y=1.395 $X2=0 $Y2=0
cc_169 N_TE_B_c_155_n N_A_27_47#_c_299_n 0.00581507f $X=2.13 $Y=1.395 $X2=0
+ $Y2=0
cc_170 N_TE_B_c_157_n N_A_27_47#_c_299_n 0.0058575f $X=2.55 $Y=1.395 $X2=0 $Y2=0
cc_171 N_TE_B_c_159_n N_A_27_47#_c_299_n 0.00581507f $X=2.97 $Y=1.395 $X2=0
+ $Y2=0
cc_172 N_TE_B_c_161_n N_A_27_47#_c_299_n 0.0058575f $X=3.39 $Y=1.395 $X2=0 $Y2=0
cc_173 N_TE_B_c_163_n N_A_27_47#_c_299_n 0.00936175f $X=3.81 $Y=1.395 $X2=0
+ $Y2=0
cc_174 N_TE_B_c_145_n N_A_27_47#_c_299_n 0.0154391f $X=0.945 $Y=1.25 $X2=0 $Y2=0
cc_175 N_TE_B_c_166_n N_A_27_47#_c_299_n 0.00405558f $X=1.365 $Y=1.395 $X2=0
+ $Y2=0
cc_176 N_TE_B_c_167_n N_A_27_47#_c_299_n 0.00354669f $X=1.785 $Y=1.395 $X2=0
+ $Y2=0
cc_177 N_TE_B_c_168_n N_A_27_47#_c_299_n 0.00354669f $X=2.205 $Y=1.395 $X2=0
+ $Y2=0
cc_178 N_TE_B_c_169_n N_A_27_47#_c_299_n 0.00354669f $X=2.625 $Y=1.395 $X2=0
+ $Y2=0
cc_179 N_TE_B_c_170_n N_A_27_47#_c_299_n 0.00354669f $X=3.045 $Y=1.395 $X2=0
+ $Y2=0
cc_180 N_TE_B_c_171_n N_A_27_47#_c_299_n 0.00354669f $X=3.465 $Y=1.395 $X2=0
+ $Y2=0
cc_181 N_TE_B_c_144_n N_A_27_47#_c_343_n 0.0130163f $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_182 TE_B N_A_27_47#_c_343_n 0.0258602f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_183 N_TE_B_c_147_n N_A_27_47#_c_343_n 0.0101792f $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_184 N_TE_B_c_163_n N_A_27_47#_c_300_n 3.38171e-19 $X=3.81 $Y=1.395 $X2=0
+ $Y2=0
cc_185 N_TE_B_M1023_g N_VPWR_c_572_n 0.0129471f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_186 N_TE_B_c_150_n N_VPWR_c_572_n 0.0016047f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_187 N_TE_B_c_150_n N_VPWR_c_573_n 7.4754e-19 $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_188 N_TE_B_c_152_n N_VPWR_c_573_n 0.0111574f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_189 N_TE_B_c_154_n N_VPWR_c_573_n 0.0110282f $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_190 N_TE_B_c_156_n N_VPWR_c_573_n 6.72101e-19 $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_191 N_TE_B_c_154_n N_VPWR_c_574_n 6.72101e-19 $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_192 N_TE_B_c_156_n N_VPWR_c_574_n 0.0110282f $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_193 N_TE_B_c_158_n N_VPWR_c_574_n 0.0110282f $X=2.625 $Y=1.47 $X2=0 $Y2=0
cc_194 N_TE_B_c_160_n N_VPWR_c_574_n 6.72101e-19 $X=3.045 $Y=1.47 $X2=0 $Y2=0
cc_195 N_TE_B_c_158_n N_VPWR_c_575_n 6.72101e-19 $X=2.625 $Y=1.47 $X2=0 $Y2=0
cc_196 N_TE_B_c_160_n N_VPWR_c_575_n 0.0110282f $X=3.045 $Y=1.47 $X2=0 $Y2=0
cc_197 N_TE_B_c_162_n N_VPWR_c_575_n 0.0110282f $X=3.465 $Y=1.47 $X2=0 $Y2=0
cc_198 N_TE_B_c_164_n N_VPWR_c_575_n 6.72101e-19 $X=3.885 $Y=1.47 $X2=0 $Y2=0
cc_199 N_TE_B_c_162_n N_VPWR_c_576_n 6.73128e-19 $X=3.465 $Y=1.47 $X2=0 $Y2=0
cc_200 N_TE_B_c_164_n N_VPWR_c_576_n 0.0121688f $X=3.885 $Y=1.47 $X2=0 $Y2=0
cc_201 N_TE_B_c_154_n N_VPWR_c_577_n 0.0046653f $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_202 N_TE_B_c_156_n N_VPWR_c_577_n 0.0046653f $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_203 N_TE_B_c_158_n N_VPWR_c_579_n 0.0046653f $X=2.625 $Y=1.47 $X2=0 $Y2=0
cc_204 N_TE_B_c_160_n N_VPWR_c_579_n 0.0046653f $X=3.045 $Y=1.47 $X2=0 $Y2=0
cc_205 N_TE_B_c_162_n N_VPWR_c_581_n 0.0046653f $X=3.465 $Y=1.47 $X2=0 $Y2=0
cc_206 N_TE_B_c_164_n N_VPWR_c_581_n 0.0046653f $X=3.885 $Y=1.47 $X2=0 $Y2=0
cc_207 N_TE_B_M1023_g N_VPWR_c_583_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_208 N_TE_B_c_150_n N_VPWR_c_584_n 0.00579312f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_209 N_TE_B_c_152_n N_VPWR_c_584_n 0.0046653f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_210 N_TE_B_M1023_g N_VPWR_c_571_n 0.00895857f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_211 N_TE_B_c_150_n N_VPWR_c_571_n 0.010505f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_212 N_TE_B_c_152_n N_VPWR_c_571_n 0.00796766f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_213 N_TE_B_c_154_n N_VPWR_c_571_n 0.00796766f $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_214 N_TE_B_c_156_n N_VPWR_c_571_n 0.00796766f $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_215 N_TE_B_c_158_n N_VPWR_c_571_n 0.00796766f $X=2.625 $Y=1.47 $X2=0 $Y2=0
cc_216 N_TE_B_c_160_n N_VPWR_c_571_n 0.00796766f $X=3.045 $Y=1.47 $X2=0 $Y2=0
cc_217 N_TE_B_c_162_n N_VPWR_c_571_n 0.00796766f $X=3.465 $Y=1.47 $X2=0 $Y2=0
cc_218 N_TE_B_c_164_n N_VPWR_c_571_n 0.00796766f $X=3.885 $Y=1.47 $X2=0 $Y2=0
cc_219 N_TE_B_M1023_g N_A_204_309#_c_704_n 4.91309e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_TE_B_c_150_n N_A_204_309#_c_704_n 0.00967786f $X=0.945 $Y=1.47 $X2=0
+ $Y2=0
cc_221 N_TE_B_c_152_n N_A_204_309#_c_692_n 0.0134056f $X=1.365 $Y=1.47 $X2=0
+ $Y2=0
cc_222 N_TE_B_c_153_n N_A_204_309#_c_692_n 0.0020486f $X=1.71 $Y=1.395 $X2=0
+ $Y2=0
cc_223 N_TE_B_c_154_n N_A_204_309#_c_692_n 0.0133633f $X=1.785 $Y=1.47 $X2=0
+ $Y2=0
cc_224 N_TE_B_c_150_n N_A_204_309#_c_693_n 0.00301378f $X=0.945 $Y=1.47 $X2=0
+ $Y2=0
cc_225 N_TE_B_c_151_n N_A_204_309#_c_693_n 0.00215435f $X=1.29 $Y=1.395 $X2=0
+ $Y2=0
cc_226 N_TE_B_c_156_n N_A_204_309#_c_694_n 0.0133633f $X=2.205 $Y=1.47 $X2=0
+ $Y2=0
cc_227 N_TE_B_c_157_n N_A_204_309#_c_694_n 0.0020486f $X=2.55 $Y=1.395 $X2=0
+ $Y2=0
cc_228 N_TE_B_c_158_n N_A_204_309#_c_694_n 0.0133633f $X=2.625 $Y=1.47 $X2=0
+ $Y2=0
cc_229 N_TE_B_c_160_n N_A_204_309#_c_695_n 0.0133633f $X=3.045 $Y=1.47 $X2=0
+ $Y2=0
cc_230 N_TE_B_c_161_n N_A_204_309#_c_695_n 0.0020486f $X=3.39 $Y=1.395 $X2=0
+ $Y2=0
cc_231 N_TE_B_c_162_n N_A_204_309#_c_695_n 0.0133633f $X=3.465 $Y=1.47 $X2=0
+ $Y2=0
cc_232 N_TE_B_c_164_n N_A_204_309#_c_696_n 0.0154663f $X=3.885 $Y=1.47 $X2=0
+ $Y2=0
cc_233 N_TE_B_c_164_n N_A_204_309#_c_697_n 0.00397974f $X=3.885 $Y=1.47 $X2=0
+ $Y2=0
cc_234 N_TE_B_c_155_n N_A_204_309#_c_701_n 0.00215435f $X=2.13 $Y=1.395 $X2=0
+ $Y2=0
cc_235 N_TE_B_c_159_n N_A_204_309#_c_702_n 0.00215435f $X=2.97 $Y=1.395 $X2=0
+ $Y2=0
cc_236 N_TE_B_c_163_n N_A_204_309#_c_703_n 0.00215435f $X=3.81 $Y=1.395 $X2=0
+ $Y2=0
cc_237 N_TE_B_c_143_n N_VGND_c_925_n 0.00966951f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_238 N_TE_B_c_143_n N_VGND_c_934_n 0.00341689f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_239 N_TE_B_c_143_n N_VGND_c_938_n 0.0050171f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_240 N_TE_B_c_143_n N_A_215_47#_c_1049_n 0.00178374f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_TE_B_c_143_n N_A_215_47#_c_1050_n 7.04009e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_TE_B_c_151_n N_A_215_47#_c_1050_n 0.00101297f $X=1.29 $Y=1.395 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_289_n N_A_c_438_n 0.0199259f $X=4.35 $Y=0.96 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_27_47#_c_299_n A 0.0269779f $X=4.305 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_300_n A 0.00107743f $X=4.305 $Y=1.035 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_299_n N_A_c_447_n 0.00195057f $X=4.305 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_300_n N_A_c_447_n 0.0132663f $X=4.305 $Y=1.035 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_302_n N_VPWR_M1023_d 0.00404069f $X=0.68 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_249 N_A_27_47#_c_302_n N_VPWR_c_572_n 0.0193336f $X=0.68 $Y=1.495 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_301_n N_VPWR_c_583_n 0.0176426f $X=0.26 $Y=1.815 $X2=0 $Y2=0
cc_251 N_A_27_47#_M1023_s N_VPWR_c_571_n 0.00387172f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_301_n N_VPWR_c_571_n 0.00974347f $X=0.26 $Y=1.815 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_276_n N_A_204_309#_c_692_n 4.28192e-19 $X=1.485 $Y=1.035
+ $X2=0 $Y2=0
cc_254 N_A_27_47#_c_299_n N_A_204_309#_c_692_n 0.0490093f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_302_n N_A_204_309#_c_693_n 0.0093578f $X=0.68 $Y=1.495 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_299_n N_A_204_309#_c_693_n 0.0189161f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_291_n N_A_204_309#_c_694_n 3.59173e-19 $X=2.25 $Y=1.035
+ $X2=0 $Y2=0
cc_258 N_A_27_47#_c_299_n N_A_204_309#_c_694_n 0.0490092f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_293_n N_A_204_309#_c_695_n 3.59173e-19 $X=3.09 $Y=1.035
+ $X2=0 $Y2=0
cc_260 N_A_27_47#_c_299_n N_A_204_309#_c_695_n 0.0490092f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_295_n N_A_204_309#_c_696_n 8.9107e-19 $X=3.93 $Y=1.035 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_299_n N_A_204_309#_c_696_n 0.0543037f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_300_n N_A_204_309#_c_696_n 0.00700619f $X=4.305 $Y=1.035
+ $X2=0 $Y2=0
cc_264 N_A_27_47#_c_278_n N_A_204_309#_c_701_n 2.23657e-19 $X=2.175 $Y=1.035
+ $X2=0 $Y2=0
cc_265 N_A_27_47#_c_299_n N_A_204_309#_c_701_n 0.0143368f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_282_n N_A_204_309#_c_702_n 2.23657e-19 $X=3.015 $Y=1.035
+ $X2=0 $Y2=0
cc_267 N_A_27_47#_c_299_n N_A_204_309#_c_702_n 0.0143368f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_286_n N_A_204_309#_c_703_n 2.23657e-19 $X=3.855 $Y=1.035
+ $X2=0 $Y2=0
cc_269 N_A_27_47#_c_299_n N_A_204_309#_c_703_n 0.0143368f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_297_n N_VGND_M1030_d 0.00334969f $X=0.68 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_271 N_A_27_47#_c_298_n N_VGND_M1030_d 8.61564e-19 $X=0.68 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_272 N_A_27_47#_c_274_n N_VGND_c_925_n 0.00195572f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_297_n N_VGND_c_925_n 0.0207342f $X=0.68 $Y=0.825 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_274_n N_VGND_c_926_n 0.00725083f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_277_n N_VGND_c_926_n 0.00685342f $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_279_n N_VGND_c_926_n 5.54209e-19 $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_277_n N_VGND_c_927_n 5.54209e-19 $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_279_n N_VGND_c_927_n 0.00685342f $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_281_n N_VGND_c_927_n 0.00685342f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_283_n N_VGND_c_927_n 5.54209e-19 $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_281_n N_VGND_c_928_n 5.54209e-19 $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_283_n N_VGND_c_928_n 0.00685342f $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_285_n N_VGND_c_928_n 0.00685342f $X=3.51 $Y=0.96 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_287_n N_VGND_c_928_n 5.54209e-19 $X=3.93 $Y=0.96 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_285_n N_VGND_c_929_n 5.54817e-19 $X=3.51 $Y=0.96 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_287_n N_VGND_c_929_n 0.00685342f $X=3.93 $Y=0.96 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_289_n N_VGND_c_929_n 0.00866947f $X=4.35 $Y=0.96 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_281_n N_VGND_c_930_n 0.00341689f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_283_n N_VGND_c_930_n 0.00341689f $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_285_n N_VGND_c_932_n 0.00341689f $X=3.51 $Y=0.96 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_287_n N_VGND_c_932_n 0.00341689f $X=3.93 $Y=0.96 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_296_n N_VGND_c_934_n 0.0169851f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_297_n N_VGND_c_934_n 0.00235077f $X=0.68 $Y=0.825 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_274_n N_VGND_c_935_n 0.00341689f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_277_n N_VGND_c_936_n 0.00341689f $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_279_n N_VGND_c_936_n 0.00341689f $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_289_n N_VGND_c_937_n 0.00313154f $X=4.35 $Y=0.96 $X2=0 $Y2=0
cc_298 N_A_27_47#_M1030_s N_VGND_c_938_n 0.00230206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_274_n N_VGND_c_938_n 0.00540327f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_277_n N_VGND_c_938_n 0.0040262f $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_279_n N_VGND_c_938_n 0.0040262f $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_281_n N_VGND_c_938_n 0.0040262f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_283_n N_VGND_c_938_n 0.0040262f $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_285_n N_VGND_c_938_n 0.0040262f $X=3.51 $Y=0.96 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_287_n N_VGND_c_938_n 0.0040262f $X=3.93 $Y=0.96 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_289_n N_VGND_c_938_n 0.00390035f $X=4.35 $Y=0.96 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_296_n N_VGND_c_938_n 0.00961382f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_297_n N_VGND_c_938_n 0.00561958f $X=0.68 $Y=0.825 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_274_n N_A_215_47#_c_1055_n 0.0108561f $X=1.41 $Y=0.96 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_275_n N_A_215_47#_c_1055_n 0.00179137f $X=1.755 $Y=1.035
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_277_n N_A_215_47#_c_1055_n 0.010245f $X=1.83 $Y=0.96 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_299_n N_A_215_47#_c_1055_n 0.0410653f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_297_n N_A_215_47#_c_1050_n 0.0157409f $X=0.68 $Y=0.825 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_299_n N_A_215_47#_c_1050_n 0.0228911f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_279_n N_A_215_47#_c_1061_n 0.010245f $X=2.25 $Y=0.96 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_280_n N_A_215_47#_c_1061_n 0.00179137f $X=2.595 $Y=1.035
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_c_281_n N_A_215_47#_c_1061_n 0.010245f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_299_n N_A_215_47#_c_1061_n 0.0408222f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_283_n N_A_215_47#_c_1065_n 0.010245f $X=3.09 $Y=0.96 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_284_n N_A_215_47#_c_1065_n 0.00179137f $X=3.435 $Y=1.035
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_285_n N_A_215_47#_c_1065_n 0.010245f $X=3.51 $Y=0.96 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_299_n N_A_215_47#_c_1065_n 0.0408222f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_287_n N_A_215_47#_c_1069_n 0.0102303f $X=3.93 $Y=0.96 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_288_n N_A_215_47#_c_1069_n 0.00183302f $X=4.17 $Y=1.035
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_c_289_n N_A_215_47#_c_1069_n 0.0102044f $X=4.35 $Y=0.96 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_299_n N_A_215_47#_c_1069_n 0.0410036f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_289_n N_A_215_47#_c_1073_n 0.00126767f $X=4.35 $Y=0.96 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_278_n N_A_215_47#_c_1074_n 0.00186022f $X=2.175 $Y=1.035
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_299_n N_A_215_47#_c_1074_n 0.0132296f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_282_n N_A_215_47#_c_1076_n 0.00186022f $X=3.015 $Y=1.035
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_299_n N_A_215_47#_c_1076_n 0.0132296f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_286_n N_A_215_47#_c_1078_n 0.00186022f $X=3.855 $Y=1.035
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_299_n N_A_215_47#_c_1078_n 0.0132296f $X=4.305 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A_M1001_g N_VPWR_c_576_n 0.00320814f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A_M1001_g N_VPWR_c_585_n 0.00357877f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_M1007_g N_VPWR_c_585_n 0.00357877f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_M1019_g N_VPWR_c_585_n 0.00357877f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A_M1020_g N_VPWR_c_585_n 0.00357877f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A_M1022_g N_VPWR_c_585_n 0.00357877f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_340 N_A_M1025_g N_VPWR_c_585_n 0.00357877f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A_M1026_g N_VPWR_c_585_n 0.00357877f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A_M1029_g N_VPWR_c_585_n 0.00357877f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_343 N_A_M1001_g N_VPWR_c_571_n 0.00664112f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A_M1007_g N_VPWR_c_571_n 0.00522516f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A_M1019_g N_VPWR_c_571_n 0.00522516f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A_M1020_g N_VPWR_c_571_n 0.00522516f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A_M1022_g N_VPWR_c_571_n 0.00522516f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A_M1025_g N_VPWR_c_571_n 0.00522516f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A_M1026_g N_VPWR_c_571_n 0.00522516f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A_M1029_g N_VPWR_c_571_n 0.00621986f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_351 A N_A_204_309#_c_696_n 0.00378383f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_352 N_A_M1001_g N_A_204_309#_c_740_n 0.0136016f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A_M1007_g N_A_204_309#_c_740_n 0.00941684f $X=5.245 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_M1019_g N_A_204_309#_c_742_n 0.00941684f $X=5.665 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A_M1020_g N_A_204_309#_c_742_n 0.00941684f $X=6.085 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A_M1022_g N_A_204_309#_c_744_n 0.00941684f $X=6.505 $Y=1.985 $X2=0
+ $Y2=0
cc_357 N_A_M1025_g N_A_204_309#_c_744_n 0.00941684f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_358 N_A_M1026_g N_A_204_309#_c_699_n 0.00941684f $X=7.345 $Y=1.985 $X2=0
+ $Y2=0
cc_359 N_A_M1029_g N_A_204_309#_c_699_n 0.00941684f $X=7.765 $Y=1.985 $X2=0
+ $Y2=0
cc_360 N_A_M1001_g N_Z_c_826_n 0.00588511f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A_M1007_g N_Z_c_826_n 0.00678236f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A_M1019_g N_Z_c_826_n 5.3107e-19 $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A_M1007_g N_Z_c_817_n 0.00889211f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_364 N_A_M1019_g N_Z_c_817_n 0.00889211f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_365 A N_Z_c_817_n 0.0369911f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_366 N_A_c_447_n N_Z_c_817_n 0.00211509f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_367 N_A_M1001_g N_Z_c_818_n 0.00433405f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A_M1007_g N_Z_c_818_n 0.00146767f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_369 A N_Z_c_818_n 0.0272853f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_370 N_A_c_447_n N_Z_c_818_n 0.00219557f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_371 N_A_M1007_g N_Z_c_837_n 5.3107e-19 $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_372 N_A_M1019_g N_Z_c_837_n 0.00678236f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_373 N_A_M1020_g N_Z_c_837_n 0.00678236f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A_M1022_g N_Z_c_837_n 5.3107e-19 $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_375 N_A_M1020_g N_Z_c_819_n 0.00889211f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_376 N_A_M1022_g N_Z_c_819_n 0.00889211f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_377 A N_Z_c_819_n 0.0369911f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_378 N_A_c_447_n N_Z_c_819_n 0.00211509f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A_M1025_g N_Z_c_820_n 0.00889211f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A_M1026_g N_Z_c_820_n 0.00889211f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_381 A N_Z_c_820_n 0.0369911f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_382 N_A_c_447_n N_Z_c_820_n 0.00211509f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_M1029_g N_Z_c_821_n 0.0110139f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_384 A N_Z_c_821_n 0.00562029f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_385 N_A_M1019_g N_Z_c_822_n 0.00146767f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_386 N_A_M1020_g N_Z_c_822_n 0.00146767f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_387 A N_Z_c_822_n 0.0272853f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_388 N_A_c_447_n N_Z_c_822_n 0.00219557f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_M1022_g N_Z_c_823_n 0.00146767f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_390 N_A_M1025_g N_Z_c_823_n 0.00146767f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_391 A N_Z_c_823_n 0.0272853f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_392 N_A_c_447_n N_Z_c_823_n 0.00219557f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_393 N_A_M1026_g N_Z_c_824_n 0.00146767f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A_M1029_g N_Z_c_824_n 0.00146767f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_395 A N_Z_c_824_n 0.0272853f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_396 N_A_c_447_n N_Z_c_824_n 0.00219557f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_397 N_A_c_438_n Z 0.0029286f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A_c_439_n Z 0.00928392f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A_c_440_n Z 0.00928392f $X=5.665 $Y=0.995 $X2=0 $Y2=0
cc_400 N_A_c_441_n Z 0.00928392f $X=6.085 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_c_442_n Z 0.00928392f $X=6.505 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A_c_443_n Z 0.00928392f $X=6.925 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A_c_444_n Z 0.00928392f $X=7.345 $Y=0.995 $X2=0 $Y2=0
cc_404 N_A_c_445_n Z 0.0117284f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_405 A Z 0.184568f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_406 N_A_c_447_n Z 0.0141859f $X=7.765 $Y=1.16 $X2=0 $Y2=0
cc_407 N_A_M1020_g N_Z_c_873_n 5.3107e-19 $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A_M1022_g N_Z_c_873_n 0.00678236f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_409 N_A_M1025_g N_Z_c_873_n 0.00678236f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_410 N_A_M1026_g N_Z_c_873_n 5.3107e-19 $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_411 N_A_M1025_g N_Z_c_877_n 5.3107e-19 $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_412 N_A_M1026_g N_Z_c_877_n 0.00678236f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_413 N_A_M1029_g N_Z_c_877_n 0.011421f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_414 N_A_c_445_n Z 0.0208811f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_415 A Z 0.023488f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_416 N_A_c_438_n N_VGND_c_929_n 0.00119014f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_417 N_A_c_438_n N_VGND_c_937_n 0.00357877f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_418 N_A_c_439_n N_VGND_c_937_n 0.00357877f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_419 N_A_c_440_n N_VGND_c_937_n 0.00357877f $X=5.665 $Y=0.995 $X2=0 $Y2=0
cc_420 N_A_c_441_n N_VGND_c_937_n 0.00357877f $X=6.085 $Y=0.995 $X2=0 $Y2=0
cc_421 N_A_c_442_n N_VGND_c_937_n 0.00357877f $X=6.505 $Y=0.995 $X2=0 $Y2=0
cc_422 N_A_c_443_n N_VGND_c_937_n 0.00357877f $X=6.925 $Y=0.995 $X2=0 $Y2=0
cc_423 N_A_c_444_n N_VGND_c_937_n 0.00357877f $X=7.345 $Y=0.995 $X2=0 $Y2=0
cc_424 N_A_c_445_n N_VGND_c_937_n 0.00357877f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_425 N_A_c_438_n N_VGND_c_938_n 0.00542674f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A_c_439_n N_VGND_c_938_n 0.00522516f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_427 N_A_c_440_n N_VGND_c_938_n 0.00522516f $X=5.665 $Y=0.995 $X2=0 $Y2=0
cc_428 N_A_c_441_n N_VGND_c_938_n 0.00522516f $X=6.085 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A_c_442_n N_VGND_c_938_n 0.00522516f $X=6.505 $Y=0.995 $X2=0 $Y2=0
cc_430 N_A_c_443_n N_VGND_c_938_n 0.00522516f $X=6.925 $Y=0.995 $X2=0 $Y2=0
cc_431 N_A_c_444_n N_VGND_c_938_n 0.00522516f $X=7.345 $Y=0.995 $X2=0 $Y2=0
cc_432 N_A_c_445_n N_VGND_c_938_n 0.00621986f $X=7.765 $Y=0.995 $X2=0 $Y2=0
cc_433 A N_A_215_47#_c_1069_n 0.00435364f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_434 N_A_c_438_n N_A_215_47#_c_1051_n 0.0109439f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_435 N_A_c_439_n N_A_215_47#_c_1051_n 0.00822564f $X=5.245 $Y=0.995 $X2=0
+ $Y2=0
cc_436 N_A_c_440_n N_A_215_47#_c_1051_n 0.00827637f $X=5.665 $Y=0.995 $X2=0
+ $Y2=0
cc_437 N_A_c_441_n N_A_215_47#_c_1051_n 0.00827637f $X=6.085 $Y=0.995 $X2=0
+ $Y2=0
cc_438 N_A_c_442_n N_A_215_47#_c_1051_n 0.00827637f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_439 N_A_c_443_n N_A_215_47#_c_1051_n 0.00827637f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_440 N_A_c_444_n N_A_215_47#_c_1051_n 0.00827637f $X=7.345 $Y=0.995 $X2=0
+ $Y2=0
cc_441 N_A_c_445_n N_A_215_47#_c_1051_n 0.00827637f $X=7.765 $Y=0.995 $X2=0
+ $Y2=0
cc_442 A N_A_215_47#_c_1051_n 0.00419156f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_443 N_VPWR_c_571_n N_A_204_309#_M1000_s 0.00393857f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_444 N_VPWR_c_571_n N_A_204_309#_M1006_s 0.00570907f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_571_n N_A_204_309#_M1013_s 0.00570907f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_571_n N_A_204_309#_M1024_s 0.00570907f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_571_n N_A_204_309#_M1001_s 0.00210127f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_571_n N_A_204_309#_M1007_s 0.0021521f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_571_n N_A_204_309#_M1020_s 0.0021521f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_571_n N_A_204_309#_M1025_s 0.0021521f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_571_n N_A_204_309#_M1029_s 0.00209324f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_584_n N_A_204_309#_c_704_n 0.0134781f $X=1.41 $Y=2.72 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_571_n N_A_204_309#_c_704_n 0.00856983f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_454 N_VPWR_M1005_d N_A_204_309#_c_692_n 0.00165831f $X=1.44 $Y=1.545 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_573_n N_A_204_309#_c_692_n 0.0170258f $X=1.575 $Y=2.02 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_577_n N_A_204_309#_c_761_n 0.0113958f $X=2.25 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_571_n N_A_204_309#_c_761_n 0.00646998f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_458 N_VPWR_M1010_d N_A_204_309#_c_694_n 0.00165831f $X=2.28 $Y=1.545 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_574_n N_A_204_309#_c_694_n 0.0170258f $X=2.415 $Y=2.02 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_579_n N_A_204_309#_c_765_n 0.0113958f $X=3.09 $Y=2.72 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_571_n N_A_204_309#_c_765_n 0.00646998f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_462 N_VPWR_M1016_d N_A_204_309#_c_695_n 0.00165831f $X=3.12 $Y=1.545 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_575_n N_A_204_309#_c_695_n 0.0170258f $X=3.255 $Y=2.02 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_581_n N_A_204_309#_c_769_n 0.0113958f $X=3.93 $Y=2.72 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_571_n N_A_204_309#_c_769_n 0.00646998f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_M1028_d N_A_204_309#_c_696_n 0.00268486f $X=3.96 $Y=1.545 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_576_n N_A_204_309#_c_696_n 0.0236659f $X=4.095 $Y=2 $X2=0 $Y2=0
cc_468 N_VPWR_c_576_n N_A_204_309#_c_697_n 0.0376463f $X=4.095 $Y=2 $X2=0 $Y2=0
cc_469 N_VPWR_c_585_n N_A_204_309#_c_740_n 0.0358653f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_571_n N_A_204_309#_c_740_n 0.0235123f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_576_n N_A_204_309#_c_698_n 0.0151017f $X=4.095 $Y=2 $X2=0 $Y2=0
cc_472 N_VPWR_c_585_n N_A_204_309#_c_698_n 0.0173913f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_571_n N_A_204_309#_c_698_n 0.00962794f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_585_n N_A_204_309#_c_742_n 0.0358391f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_571_n N_A_204_309#_c_742_n 0.0234424f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_585_n N_A_204_309#_c_744_n 0.0358391f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_571_n N_A_204_309#_c_744_n 0.0234424f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_585_n N_A_204_309#_c_699_n 0.0571143f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_571_n N_A_204_309#_c_699_n 0.0351787f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_585_n N_A_204_309#_c_785_n 0.0114548f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_571_n N_A_204_309#_c_785_n 0.00654447f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_585_n N_A_204_309#_c_787_n 0.0114548f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_571_n N_A_204_309#_c_787_n 0.00654447f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_585_n N_A_204_309#_c_789_n 0.0114548f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_571_n N_A_204_309#_c_789_n 0.00654447f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_571_n N_Z_M1001_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_487 N_VPWR_c_571_n N_Z_M1019_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_488 N_VPWR_c_571_n N_Z_M1022_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_489 N_VPWR_c_571_n N_Z_M1026_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_490 N_A_204_309#_c_740_n N_Z_M1001_d 0.00312348f $X=5.37 $Y=2.38 $X2=0 $Y2=0
cc_491 N_A_204_309#_c_742_n N_Z_M1019_d 0.00312348f $X=6.21 $Y=2.38 $X2=0 $Y2=0
cc_492 N_A_204_309#_c_744_n N_Z_M1022_d 0.00312348f $X=7.05 $Y=2.38 $X2=0 $Y2=0
cc_493 N_A_204_309#_c_699_n N_Z_M1026_d 0.00312348f $X=7.89 $Y=2.38 $X2=0 $Y2=0
cc_494 N_A_204_309#_c_740_n N_Z_c_826_n 0.0159307f $X=5.37 $Y=2.38 $X2=0 $Y2=0
cc_495 N_A_204_309#_M1007_s N_Z_c_817_n 0.00165831f $X=5.32 $Y=1.485 $X2=0 $Y2=0
cc_496 N_A_204_309#_c_740_n N_Z_c_817_n 0.00256303f $X=5.37 $Y=2.38 $X2=0 $Y2=0
cc_497 N_A_204_309#_c_798_p N_Z_c_817_n 0.0126766f $X=5.455 $Y=1.96 $X2=0 $Y2=0
cc_498 N_A_204_309#_c_742_n N_Z_c_817_n 0.00256303f $X=6.21 $Y=2.38 $X2=0 $Y2=0
cc_499 N_A_204_309#_c_742_n N_Z_c_837_n 0.0159307f $X=6.21 $Y=2.38 $X2=0 $Y2=0
cc_500 N_A_204_309#_M1020_s N_Z_c_819_n 0.00165831f $X=6.16 $Y=1.485 $X2=0 $Y2=0
cc_501 N_A_204_309#_c_742_n N_Z_c_819_n 0.00256303f $X=6.21 $Y=2.38 $X2=0 $Y2=0
cc_502 N_A_204_309#_c_803_p N_Z_c_819_n 0.0126766f $X=6.295 $Y=1.96 $X2=0 $Y2=0
cc_503 N_A_204_309#_c_744_n N_Z_c_819_n 0.00256303f $X=7.05 $Y=2.38 $X2=0 $Y2=0
cc_504 N_A_204_309#_M1025_s N_Z_c_820_n 0.00165831f $X=7 $Y=1.485 $X2=0 $Y2=0
cc_505 N_A_204_309#_c_744_n N_Z_c_820_n 0.00256303f $X=7.05 $Y=2.38 $X2=0 $Y2=0
cc_506 N_A_204_309#_c_807_p N_Z_c_820_n 0.0126766f $X=7.135 $Y=1.96 $X2=0 $Y2=0
cc_507 N_A_204_309#_c_699_n N_Z_c_820_n 0.00256303f $X=7.89 $Y=2.38 $X2=0 $Y2=0
cc_508 N_A_204_309#_M1029_s N_Z_c_821_n 0.00282391f $X=7.84 $Y=1.485 $X2=0 $Y2=0
cc_509 N_A_204_309#_c_699_n N_Z_c_821_n 0.00256303f $X=7.89 $Y=2.38 $X2=0 $Y2=0
cc_510 N_A_204_309#_c_700_n N_Z_c_821_n 0.0264014f $X=7.975 $Y=1.96 $X2=0 $Y2=0
cc_511 N_A_204_309#_c_744_n N_Z_c_873_n 0.0159307f $X=7.05 $Y=2.38 $X2=0 $Y2=0
cc_512 N_A_204_309#_c_699_n N_Z_c_877_n 0.0159307f $X=7.89 $Y=2.38 $X2=0 $Y2=0
cc_513 N_A_204_309#_c_696_n N_A_215_47#_c_1069_n 0.00504579f $X=4.45 $Y=1.58
+ $X2=0 $Y2=0
cc_514 N_Z_M1002_s N_VGND_c_938_n 0.00216833f $X=4.9 $Y=0.235 $X2=0 $Y2=0
cc_515 N_Z_M1004_s N_VGND_c_938_n 0.00216833f $X=5.74 $Y=0.235 $X2=0 $Y2=0
cc_516 N_Z_M1027_s N_VGND_c_938_n 0.00216833f $X=6.58 $Y=0.235 $X2=0 $Y2=0
cc_517 N_Z_M1032_s N_VGND_c_938_n 0.00216833f $X=7.42 $Y=0.235 $X2=0 $Y2=0
cc_518 Z N_A_215_47#_M1003_d 0.00306867f $X=7.97 $Y=0.765 $X2=0 $Y2=0
cc_519 Z N_A_215_47#_M1011_d 0.00306867f $X=7.97 $Y=0.765 $X2=0 $Y2=0
cc_520 Z N_A_215_47#_M1031_d 0.00306867f $X=7.97 $Y=0.765 $X2=0 $Y2=0
cc_521 Z N_A_215_47#_M1033_d 0.00212897f $X=7.97 $Y=0.765 $X2=0 $Y2=0
cc_522 N_Z_c_815_n N_A_215_47#_M1033_d 0.00273062f $X=8.082 $Y=0.825 $X2=0 $Y2=0
cc_523 Z N_A_215_47#_M1033_d 0.00101757f $X=8.055 $Y=0.85 $X2=0 $Y2=0
cc_524 N_Z_M1002_s N_A_215_47#_c_1051_n 0.00304533f $X=4.9 $Y=0.235 $X2=0 $Y2=0
cc_525 N_Z_M1004_s N_A_215_47#_c_1051_n 0.00304533f $X=5.74 $Y=0.235 $X2=0 $Y2=0
cc_526 N_Z_M1027_s N_A_215_47#_c_1051_n 0.00304533f $X=6.58 $Y=0.235 $X2=0 $Y2=0
cc_527 N_Z_M1032_s N_A_215_47#_c_1051_n 0.00304533f $X=7.42 $Y=0.235 $X2=0 $Y2=0
cc_528 Z N_A_215_47#_c_1051_n 0.15253f $X=7.97 $Y=0.765 $X2=0 $Y2=0
cc_529 N_Z_c_815_n N_A_215_47#_c_1051_n 0.0176261f $X=8.082 $Y=0.825 $X2=0 $Y2=0
cc_530 N_VGND_c_938_n N_A_215_47#_M1008_d 0.00229009f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_531 N_VGND_c_938_n N_A_215_47#_M1009_d 0.00254582f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_938_n N_A_215_47#_M1014_d 0.00254582f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_c_938_n N_A_215_47#_M1017_d 0.00254582f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_938_n N_A_215_47#_M1021_d 0.00284605f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_938_n N_A_215_47#_M1003_d 0.00215227f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_938_n N_A_215_47#_M1011_d 0.00215227f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_938_n N_A_215_47#_M1031_d 0.00215227f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_938_n N_A_215_47#_M1033_d 0.00225742f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_c_925_n N_A_215_47#_c_1049_n 0.0188652f $X=0.68 $Y=0.38 $X2=0
+ $Y2=0
cc_540 N_VGND_c_935_n N_A_215_47#_c_1049_n 0.0184794f $X=1.455 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_938_n N_A_215_47#_c_1049_n 0.0102739f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_542 N_VGND_M1008_s N_A_215_47#_c_1055_n 0.00297022f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_543 N_VGND_c_926_n N_A_215_47#_c_1055_n 0.0160613f $X=1.62 $Y=0.36 $X2=0
+ $Y2=0
cc_544 N_VGND_c_935_n N_A_215_47#_c_1055_n 0.00232396f $X=1.455 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_936_n N_A_215_47#_c_1055_n 0.00232396f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_546 N_VGND_c_938_n N_A_215_47#_c_1055_n 0.00970544f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_547 N_VGND_c_936_n N_A_215_47#_c_1120_n 0.0112554f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_548 N_VGND_c_938_n N_A_215_47#_c_1120_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_549 N_VGND_M1012_s N_A_215_47#_c_1061_n 0.00297022f $X=2.325 $Y=0.235 $X2=0
+ $Y2=0
cc_550 N_VGND_c_927_n N_A_215_47#_c_1061_n 0.0160613f $X=2.46 $Y=0.36 $X2=0
+ $Y2=0
cc_551 N_VGND_c_930_n N_A_215_47#_c_1061_n 0.00232396f $X=3.135 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_936_n N_A_215_47#_c_1061_n 0.00232396f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_938_n N_A_215_47#_c_1061_n 0.00970544f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_554 N_VGND_c_930_n N_A_215_47#_c_1127_n 0.0112554f $X=3.135 $Y=0 $X2=0 $Y2=0
cc_555 N_VGND_c_938_n N_A_215_47#_c_1127_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_M1015_s N_A_215_47#_c_1065_n 0.00297022f $X=3.165 $Y=0.235 $X2=0
+ $Y2=0
cc_557 N_VGND_c_928_n N_A_215_47#_c_1065_n 0.0160613f $X=3.3 $Y=0.36 $X2=0 $Y2=0
cc_558 N_VGND_c_930_n N_A_215_47#_c_1065_n 0.00232396f $X=3.135 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_932_n N_A_215_47#_c_1065_n 0.00232396f $X=3.975 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_c_938_n N_A_215_47#_c_1065_n 0.00970544f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_932_n N_A_215_47#_c_1134_n 0.0112554f $X=3.975 $Y=0 $X2=0 $Y2=0
cc_562 N_VGND_c_938_n N_A_215_47#_c_1134_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_563 N_VGND_M1018_s N_A_215_47#_c_1069_n 0.00304947f $X=4.005 $Y=0.235 $X2=0
+ $Y2=0
cc_564 N_VGND_c_929_n N_A_215_47#_c_1069_n 0.0167799f $X=4.14 $Y=0.36 $X2=0
+ $Y2=0
cc_565 N_VGND_c_932_n N_A_215_47#_c_1069_n 0.00232396f $X=3.975 $Y=0 $X2=0 $Y2=0
cc_566 N_VGND_c_937_n N_A_215_47#_c_1069_n 0.00226054f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_938_n N_A_215_47#_c_1069_n 0.00978344f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_c_929_n N_A_215_47#_c_1141_n 0.0025982f $X=4.14 $Y=0.36 $X2=0
+ $Y2=0
cc_569 N_VGND_c_929_n N_A_215_47#_c_1073_n 0.0161366f $X=4.14 $Y=0.36 $X2=0
+ $Y2=0
cc_570 N_VGND_c_937_n N_A_215_47#_c_1073_n 0.0146879f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_938_n N_A_215_47#_c_1073_n 0.00824212f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_937_n N_A_215_47#_c_1051_n 0.19523f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_938_n N_A_215_47#_c_1051_n 0.124598f $X=8.05 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__xnor2_2.spice
* Created: Tue Sep  1 19:32:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__xnor2_2.pex.spice"
.subckt sky130_fd_sc_hd__xnor2_2  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1008 N_A_27_47#_M1008_d N_B_M1008_g N_A_27_297#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.17875 AS=0.08775 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1015 N_A_27_47#_M1015_d N_B_M1015_g N_A_27_297#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_27_47#_M1015_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1007_d N_A_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_A_560_47#_M1014_d N_A_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1019 N_A_560_47#_M1014_d N_A_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1019_s N_B_M1010_g N_A_560_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.099125 PD=0.92 PS=0.955 NRD=0 NRS=5.532 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_B_M1016_g N_A_560_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.099125 PD=1.82 PS=0.955 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A_27_297#_M1000_g N_A_560_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A_27_297#_M1004_g N_A_560_47#_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1003_d N_B_M1018_g N_A_27_297#_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1009 N_A_27_297#_M1018_s N_A_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_A_27_297#_M1011_d N_A_M1011_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_474_297#_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 N_A_474_297#_M1005_d N_A_M1005_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1012_d N_B_M1012_g N_A_474_297#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.135 PD=1.305 PS=1.27 NRD=5.8903 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_Y_M1012_d N_B_M1017_g N_A_474_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.26 PD=1.305 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_27_297#_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_297#_M1006_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__xnor2_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o221ai_4.spice
* Created: Tue Sep  1 19:22:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o221ai_4.pex.spice"
.subckt sky130_fd_sc_hd__o221ai_4  VNB VPB C1 B1 B2 A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1013 N_Y_M1013_d N_C1_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1013_d N_C1_M1018_g N_A_27_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1026 N_Y_M1026_d N_C1_M1026_g N_A_27_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1027 N_Y_M1026_d N_C1_M1027_g N_A_27_47#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_27_47#_M1003_d N_B1_M1003_g N_A_471_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75006.6 A=0.0975 P=1.6 MULT=1
MM1011 N_A_27_47#_M1003_d N_B1_M1011_g N_A_471_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75006.1 A=0.0975 P=1.6 MULT=1
MM1019 N_A_27_47#_M1019_d N_B1_M1019_g N_A_471_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75005.7 A=0.0975 P=1.6 MULT=1
MM1004 N_A_471_47#_M1004_d N_B2_M1004_g N_A_27_47#_M1019_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1014 N_A_471_47#_M1004_d N_B2_M1014_g N_A_27_47#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1016 N_A_471_47#_M1016_d N_B2_M1016_g N_A_27_47#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1020 N_A_471_47#_M1016_d N_B2_M1020_g N_A_27_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75004 A=0.0975 P=1.6 MULT=1
MM1038 N_A_27_47#_M1020_s N_B1_M1038_g N_A_471_47#_M1038_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75003.1 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_471_47#_M1038_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1000 N_A_471_47#_M1000_d N_A2_M1000_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1006 N_A_471_47#_M1000_d N_A2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1009 N_A_471_47#_M1009_d N_A2_M1009_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1021 N_A_471_47#_M1009_d N_A2_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1021_s N_A1_M1017_g N_A_471_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_A1_M1022_g N_A_471_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1028 N_VGND_M1022_d N_A1_M1028_g N_A_471_47#_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1010_d N_C1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75008.8 A=0.15
+ P=2.3 MULT=1
MM1029 N_Y_M1010_d N_C1_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75008.4
+ A=0.15 P=2.3 MULT=1
MM1032 N_Y_M1032_d N_C1_M1032_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75008 A=0.15
+ P=2.3 MULT=1
MM1036 N_Y_M1032_d N_C1_M1036_g N_VPWR_M1036_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.395 PD=1.27 PS=1.79 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75007.5
+ A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1036_s N_B1_M1001_g N_A_553_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.395 AS=0.135 PD=1.79 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75006.6 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_A_553_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75006.2 A=0.15 P=2.3 MULT=1
MM1023 N_VPWR_M1007_d N_B1_M1023_g N_A_553_297#_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75005.8 A=0.15 P=2.3 MULT=1
MM1008 N_A_553_297#_M1023_s N_B2_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.7
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1012 N_A_553_297#_M1012_d N_B2_M1012_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1033 N_A_553_297#_M1012_d N_B2_M1033_g N_Y_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1037 N_A_553_297#_M1037_d N_B2_M1037_g N_Y_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.9
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1025 N_VPWR_M1025_d N_B1_M1025_g N_A_553_297#_M1037_d VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.135 PD=1.35 PS=1.27 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75005.3
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1015 N_A_1241_297#_M1015_d N_A1_M1015_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.175 PD=1.27 PS=1.35 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75005.8
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1002_d N_A2_M1002_g N_A_1241_297#_M1015_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.3
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1031 N_Y_M1002_d N_A2_M1031_g N_A_1241_297#_M1031_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.7
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1034 N_Y_M1034_d N_A2_M1034_g N_A_1241_297#_M1031_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.1
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1039 N_Y_M1034_d N_A2_M1039_g N_A_1241_297#_M1039_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.5
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1024 N_A_1241_297#_M1039_s N_A1_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.9
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1030 N_A_1241_297#_M1030_d N_A1_M1030_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1035 N_A_1241_297#_M1030_d N_A1_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_124 VPB 0 1.20766e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__o221ai_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdfbbn_2.pex.spice
* Created: Thu Aug 27 14:45:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%CLK_N 4 5 7 8 10 13 17 19 20 24 26
c45 13 0 2.71124e-20 $X=0.47 $Y=0.805
r46 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r47 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r48 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r49 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r50 15 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=1.665
+ $X2=0.47 $Y2=1.665
r51 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.47 $Y2=0.805
r52 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r53 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r54 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r55 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r56 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r57 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r58 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r59 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_27_47# 1 2 9 13 17 19 20 23 26 27 29 32
+ 36 40 41 42 46 47 49 51 52 55 58 59 61 62 63 66 70 74 81 84 85
c278 61 0 9.71454e-20 $X=5.327 $Y=1.12
c279 49 0 1.20913e-19 $X=8.937 $Y=1.305
c280 47 0 1.7288e-19 $X=8.62 $Y=0.87
c281 17 0 4.43992e-20 $X=4.59 $Y=2.275
r282 84 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.93
+ $X2=5.19 $Y2=1.095
r283 84 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.93
+ $X2=5.19 $Y2=0.765
r284 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.19
+ $Y=0.93 $X2=5.19 $Y2=0.93
r285 78 81 31.1043 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=0.75 $Y=1.235
+ $X2=0.89 $Y2=1.235
r286 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.235 $X2=0.75 $Y2=1.235
r287 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=1.19
+ $X2=8.51 $Y2=1.19
r288 70 72 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=5.29 $Y=0.85
+ $X2=5.29 $Y2=0.965
r289 70 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0.85
+ $X2=5.29 $Y2=0.85
r290 66 79 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.72 $Y=0.85
+ $X2=0.72 $Y2=1.235
r291 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0.85
+ $X2=0.69 $Y2=0.85
r292 62 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=8.51 $Y2=1.19
r293 62 63 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=5.435 $Y2=1.19
r294 61 63 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=5.327 $Y=1.12
+ $X2=5.435 $Y2=1.19
r295 61 72 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=5.327 $Y=1.12
+ $X2=5.327 $Y2=0.965
r296 59 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=0.85
+ $X2=0.69 $Y2=0.85
r297 58 70 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=0.85
+ $X2=5.29 $Y2=0.85
r298 58 59 5.33415 $w=1.4e-07 $l=4.31e-06 $layer=MET1_cond $X=5.145 $Y=0.85
+ $X2=0.835 $Y2=0.85
r299 57 79 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.72 $Y=1.795
+ $X2=0.72 $Y2=1.235
r300 56 66 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.72 $Y=0.805
+ $X2=0.72 $Y2=0.85
r301 52 94 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.955 $Y=1.74
+ $X2=8.955 $Y2=1.875
r302 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.955
+ $Y=1.74 $X2=8.955 $Y2=1.74
r303 49 75 26.3101 $w=1.78e-07 $l=4.27e-07 $layer=LI1_cond $X=8.937 $Y=1.215
+ $X2=8.51 $Y2=1.215
r304 49 51 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=8.937 $Y=1.305
+ $X2=8.937 $Y2=1.74
r305 47 88 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=8.62 $Y=0.87
+ $X2=8.495 $Y2=0.87
r306 46 75 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=8.562 $Y=0.87
+ $X2=8.562 $Y2=1.125
r307 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.62
+ $Y=0.87 $X2=8.62 $Y2=0.87
r308 43 55 3.4683 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.257 $Y2=1.88
r309 42 57 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.72 $Y2=1.795
r310 42 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.345 $Y2=1.88
r311 40 56 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.72 $Y2=0.805
r312 40 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.345 $Y2=0.72
r313 34 41 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.345 $Y2=0.72
r314 34 36 7.92208 $w=1.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.257 $Y2=0.51
r315 32 94 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=8.925 $Y=2.275
+ $X2=8.925 $Y2=1.875
r316 27 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.495 $Y=0.705
+ $X2=8.495 $Y2=0.87
r317 27 29 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.495 $Y=0.705
+ $X2=8.495 $Y2=0.415
r318 26 87 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.13 $Y=1.245
+ $X2=5.13 $Y2=1.095
r319 23 86 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.13 $Y=0.415
+ $X2=5.13 $Y2=0.765
r320 19 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.055 $Y=1.32
+ $X2=5.13 $Y2=1.245
r321 19 20 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=5.055 $Y=1.32
+ $X2=4.665 $Y2=1.32
r322 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.59 $Y=1.395
+ $X2=4.665 $Y2=1.32
r323 15 17 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=4.59 $Y=1.395
+ $X2=4.59 $Y2=2.275
r324 11 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r325 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r326 7 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r327 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r328 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r329 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%SCD 3 7 9 10 17
c38 9 0 5.57791e-20 $X=1.61 $Y=1.19
c39 7 0 1.50346e-19 $X=1.83 $Y=2.135
c40 3 0 6.18549e-20 $X=1.83 $Y=0.445
r41 14 17 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.61 $Y=1.49
+ $X2=1.83 $Y2=1.49
r42 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.49 $X2=1.61 $Y2=1.49
r43 9 10 12.3476 $w=2.78e-07 $l=3e-07 $layer=LI1_cond $X=1.555 $Y=1.19 $X2=1.555
+ $Y2=1.49
r44 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.655
+ $X2=1.83 $Y2=1.49
r45 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.83 $Y=1.655 $X2=1.83
+ $Y2=2.135
r46 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.49
r47 1 3 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.83 $Y=1.325 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_423_315# 1 2 7 9 10 11 14 17 21 23 25 26
+ 30 31 33 34 40 46
c103 25 0 2.25267e-19 $X=3.475 $Y=0.71
c104 11 0 5.57791e-20 $X=2.265 $Y=1.65
r105 37 39 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=1.74
+ $X2=2.905 $Y2=1.905
r106 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.74 $X2=2.845 $Y2=1.74
r107 34 37 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=2.905 $Y=1.66
+ $X2=2.905 $Y2=1.74
r108 33 40 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.56 $Y=1.575
+ $X2=3.56 $Y2=1.095
r109 31 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=0.93
+ $X2=3.685 $Y2=0.765
r110 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=0.93 $X2=3.685 $Y2=0.93
r111 28 40 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=3.622 $Y=0.948
+ $X2=3.622 $Y2=1.095
r112 28 30 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=3.622 $Y=0.948
+ $X2=3.622 $Y2=0.93
r113 27 30 5.27389 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=3.622 $Y=0.795
+ $X2=3.622 $Y2=0.93
r114 25 27 19.9305 $w=8.7e-08 $l=1.84673e-07 $layer=LI1_cond $X=3.475 $Y=0.71
+ $X2=3.622 $Y2=0.795
r115 25 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.475 $Y=0.71
+ $X2=3.125 $Y2=0.71
r116 24 34 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.065 $Y=1.66
+ $X2=2.905 $Y2=1.66
r117 23 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.475 $Y=1.66
+ $X2=3.56 $Y2=1.575
r118 23 24 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.475 $Y=1.66
+ $X2=3.065 $Y2=1.66
r119 19 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.04 $Y=0.625
+ $X2=3.125 $Y2=0.71
r120 19 21 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.04 $Y=0.625
+ $X2=3.04 $Y2=0.47
r121 17 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.98 $Y=2.3
+ $X2=2.98 $Y2=1.905
r122 14 46 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.745 $Y=0.445
+ $X2=3.745 $Y2=0.765
r123 10 38 18.9432 $w=2.85e-07 $l=9e-08 $layer=POLY_cond $X=2.837 $Y=1.65
+ $X2=2.837 $Y2=1.74
r124 10 11 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.695 $Y=1.65
+ $X2=2.265 $Y2=1.65
r125 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.19 $Y=1.725
+ $X2=2.265 $Y2=1.65
r126 7 9 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.19 $Y=1.725
+ $X2=2.19 $Y2=2.135
r127 2 17 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=2.065 $X2=2.98 $Y2=2.3
r128 1 21 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%SCE 1 3 4 6 8 10 11 13 14 16 18 19 20 27 30
+ 31 32 39
c98 27 0 7.41594e-20 $X=2.25 $Y=0.93
c99 19 0 4.83365e-20 $X=3.257 $Y=0.81
r100 31 32 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.045 $Y=1.19
+ $X2=2.045 $Y2=1.53
r101 28 39 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=0.915
+ $X2=2.415 $Y2=0.915
r102 28 36 9.61737 $w=3.6e-07 $l=6e-08 $layer=POLY_cond $X=2.25 $Y=0.915
+ $X2=2.19 $Y2=0.915
r103 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=0.93 $X2=2.25 $Y2=0.93
r104 25 31 4.97646 $w=2.18e-07 $l=9.5e-08 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=2.045 $Y2=1.19
r105 24 27 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.045 $Y=0.93
+ $X2=2.25 $Y2=0.93
r106 24 25 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0.93
+ $X2=2.045 $Y2=1.095
r107 22 30 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=2.04 $Y=0.765
+ $X2=2.04 $Y2=0.51
r108 21 24 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.04 $Y=0.93
+ $X2=2.045 $Y2=0.93
r109 21 22 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.93
+ $X2=2.04 $Y2=0.765
r110 16 18 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.685 $Y=1.985
+ $X2=3.685 $Y2=2.275
r111 15 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=1.91
+ $X2=3.265 $Y2=1.91
r112 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.61 $Y=1.91
+ $X2=3.685 $Y2=1.985
r113 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.61 $Y=1.91
+ $X2=3.34 $Y2=1.91
r114 11 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.985
+ $X2=3.265 $Y2=1.91
r115 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.265 $Y=1.985
+ $X2=3.265 $Y2=2.275
r116 10 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.835
+ $X2=3.265 $Y2=1.91
r117 9 19 20.4101 $w=1.5e-07 $l=7.88987e-08 $layer=POLY_cond $X=3.265 $Y=0.885
+ $X2=3.257 $Y2=0.81
r118 9 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.265 $Y=0.885
+ $X2=3.265 $Y2=1.835
r119 6 19 20.4101 $w=1.5e-07 $l=7.84219e-08 $layer=POLY_cond $X=3.25 $Y=0.735
+ $X2=3.257 $Y2=0.81
r120 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.25 $Y=0.735
+ $X2=3.25 $Y2=0.445
r121 4 19 5.30422 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=3.175 $Y=0.81
+ $X2=3.257 $Y2=0.81
r122 4 39 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.175 $Y=0.81
+ $X2=2.415 $Y2=0.81
r123 1 36 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.19 $Y=0.735
+ $X2=2.19 $Y2=0.915
r124 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.19 $Y=0.735
+ $X2=2.19 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%D 3 7 9 10 17
c42 3 0 1.09936e-19 $X=4.105 $Y=0.445
r43 14 17 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.94 $Y=1.49
+ $X2=4.105 $Y2=1.49
r44 9 10 39.9273 $w=1.98e-07 $l=7.2e-07 $layer=LI1_cond $X=3.925 $Y=1.49
+ $X2=3.925 $Y2=2.21
r45 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.49 $X2=3.94 $Y2=1.49
r46 5 17 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=1.49
r47 5 7 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=2.275
r48 1 17 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.105 $Y=1.355
+ $X2=4.105 $Y2=1.49
r49 1 3 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.105 $Y=1.355
+ $X2=4.105 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_193_47# 1 2 7 9 12 18 20 21 24 28 29 31
+ 32 33 34 43 51 52 56 57 58 61
c214 56 0 2.05666e-19 $X=8.445 $Y=1.74
c215 29 0 9.71454e-20 $X=4.71 $Y=0.87
c216 18 0 3.84972e-20 $X=8.505 $Y=2.275
r217 56 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.74
+ $X2=8.445 $Y2=1.905
r218 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.74
+ $X2=8.445 $Y2=1.575
r219 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.445
+ $Y=1.74 $X2=8.445 $Y2=1.74
r220 51 54 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.04 $Y=1.74
+ $X2=5.04 $Y2=1.875
r221 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=1.74 $X2=5.04 $Y2=1.74
r222 43 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=1.87
+ $X2=8.51 $Y2=1.87
r223 41 52 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=1.765
+ $X2=5.04 $Y2=1.765
r224 41 69 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=4.83 $Y=1.765
+ $X2=4.735 $Y2=1.765
r225 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.87
+ $X2=4.83 $Y2=1.87
r226 37 61 71.2419 $w=2.18e-07 $l=1.36e-06 $layer=LI1_cond $X=1.125 $Y=1.87
+ $X2=1.125 $Y2=0.51
r227 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.87
+ $X2=1.15 $Y2=1.87
r228 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=1.87
+ $X2=4.83 $Y2=1.87
r229 33 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.365 $Y=1.87
+ $X2=8.51 $Y2=1.87
r230 33 34 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=8.365 $Y=1.87
+ $X2=4.975 $Y2=1.87
r231 32 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.87
+ $X2=1.15 $Y2=1.87
r232 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=4.83 $Y2=1.87
r233 31 32 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=1.295 $Y2=1.87
r234 29 46 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=4.71 $Y=0.87
+ $X2=4.58 $Y2=0.87
r235 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.71
+ $Y=0.87 $X2=4.71 $Y2=0.87
r236 26 69 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.735 $Y=1.575
+ $X2=4.735 $Y2=1.765
r237 26 28 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=4.735 $Y=1.575
+ $X2=4.735 $Y2=0.87
r238 22 24 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.04 $Y=1.245
+ $X2=9.04 $Y2=0.415
r239 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.965 $Y=1.32
+ $X2=9.04 $Y2=1.245
r240 20 21 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=8.965 $Y=1.32
+ $X2=8.58 $Y2=1.32
r241 18 59 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.505 $Y=2.275
+ $X2=8.505 $Y2=1.905
r242 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.505 $Y=1.395
+ $X2=8.58 $Y2=1.32
r243 14 58 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.505 $Y=1.395
+ $X2=8.505 $Y2=1.575
r244 12 54 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.01 $Y=2.275
+ $X2=5.01 $Y2=1.875
r245 7 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.58 $Y=0.705
+ $X2=4.58 $Y2=0.87
r246 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.58 $Y=0.705
+ $X2=4.58 $Y2=0.415
r247 2 37 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r248 1 61 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_1107_21# 1 2 9 13 17 19 21 22 26 28 30 31
+ 32 35 36 41 45 49
c146 45 0 9.81116e-20 $X=7.96 $Y=0.98
r147 49 56 10.4783 $w=2.76e-07 $l=6e-08 $layer=POLY_cond $X=7.96 $Y=1.15
+ $X2=8.02 $Y2=1.15
r148 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.96
+ $Y=1.15 $X2=7.96 $Y2=1.15
r149 45 48 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.96 $Y=0.98
+ $X2=7.96 $Y2=1.15
r150 43 44 14.1313 $w=2.59e-07 $l=3e-07 $layer=LI1_cond $X=6.87 $Y=0.68 $X2=6.87
+ $Y2=0.98
r151 36 53 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.74
+ $X2=5.695 $Y2=1.905
r152 36 52 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.74
+ $X2=5.695 $Y2=1.575
r153 35 38 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.76 $Y=1.74
+ $X2=5.76 $Y2=1.91
r154 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.72
+ $Y=1.74 $X2=5.72 $Y2=1.74
r155 33 44 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.035 $Y=0.98
+ $X2=6.87 $Y2=0.98
r156 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=0.98
+ $X2=7.96 $Y2=0.98
r157 32 33 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.795 $Y=0.98
+ $X2=7.035 $Y2=0.98
r158 30 44 5.44435 $w=2.59e-07 $l=9.88686e-08 $layer=LI1_cond $X=6.9 $Y=1.065
+ $X2=6.87 $Y2=0.98
r159 30 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.9 $Y=1.065
+ $X2=6.9 $Y2=1.785
r160 29 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.91
+ $X2=6.47 $Y2=1.91
r161 28 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.815 $Y=1.91
+ $X2=6.9 $Y2=1.785
r162 28 29 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=6.815 $Y=1.91
+ $X2=6.555 $Y2=1.91
r163 24 41 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.47 $Y=2.035
+ $X2=6.47 $Y2=1.91
r164 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.47 $Y=2.035
+ $X2=6.47 $Y2=2.21
r165 23 38 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=1.91
+ $X2=5.76 $Y2=1.91
r166 22 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=1.91
+ $X2=6.47 $Y2=1.91
r167 22 23 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=6.385 $Y=1.91
+ $X2=5.885 $Y2=1.91
r168 19 56 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.02 $Y=0.985
+ $X2=8.02 $Y2=1.15
r169 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.02 $Y=0.985
+ $X2=8.02 $Y2=0.555
r170 15 49 30.5616 $w=2.76e-07 $l=2.43926e-07 $layer=POLY_cond $X=7.785 $Y=1.315
+ $X2=7.96 $Y2=1.15
r171 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=7.785 $Y=1.315
+ $X2=7.785 $Y2=2.065
r172 13 53 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.61 $Y=2.275
+ $X2=5.61 $Y2=1.905
r173 9 52 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=5.61 $Y=0.445
+ $X2=5.61 $Y2=1.575
r174 2 41 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.065 $X2=6.47 $Y2=1.87
r175 2 26 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.065 $X2=6.47 $Y2=2.21
r176 1 43 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=6.735
+ $Y=0.235 $X2=6.87 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%SET_B 1 3 7 11 15 17 19 20 26 27 33
c131 33 0 1.0279e-19 $X=9.935 $Y=0.98
c132 19 0 1.0411e-19 $X=9.745 $Y=0.85
c133 15 0 1.0852e-19 $X=10.055 $Y=2.275
r134 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.965 $Y=0.98
+ $X2=9.965 $Y2=1.145
r135 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.965 $Y=0.98
+ $X2=9.965 $Y2=0.815
r136 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.935
+ $Y=0.98 $X2=9.935 $Y2=0.98
r137 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0.85
+ $X2=9.89 $Y2=0.85
r138 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.355 $Y=0.85
+ $X2=6.21 $Y2=0.85
r139 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.745 $Y=0.85
+ $X2=9.89 $Y2=0.85
r140 19 20 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=9.745 $Y=0.85
+ $X2=6.355 $Y2=0.85
r141 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.05
+ $Y=0.98 $X2=6.05 $Y2=0.98
r142 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0.85
+ $X2=6.21 $Y2=0.85
r143 15 36 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=10.055 $Y=2.275
+ $X2=10.055 $Y2=1.145
r144 11 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.945 $Y=0.445
+ $X2=9.945 $Y2=0.815
r145 5 30 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=6.18 $Y=0.815
+ $X2=6.085 $Y2=0.98
r146 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.18 $Y=0.815
+ $X2=6.18 $Y2=0.445
r147 1 30 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=6.14 $Y=1.145
+ $X2=6.085 $Y2=0.98
r148 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.14 $Y=1.145
+ $X2=6.14 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_931_47# 1 2 9 13 15 19 24 26 27 32 35
c106 35 0 1.0411e-19 $X=6.56 $Y=1.32
c107 32 0 4.43992e-20 $X=5.715 $Y=1.3
r108 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=1.32
+ $X2=6.59 $Y2=1.485
r109 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=1.32
+ $X2=6.59 $Y2=1.155
r110 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.56
+ $Y=1.32 $X2=6.56 $Y2=1.32
r111 31 32 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=5.63 $Y=1.3
+ $X2=5.715 $Y2=1.3
r112 29 31 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=5.38 $Y=1.3
+ $X2=5.63 $Y2=1.3
r113 27 34 8.9562 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=1.32
+ $X2=6.56 $Y2=1.32
r114 27 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.395 $Y=1.32
+ $X2=5.715 $Y2=1.32
r115 26 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.63 $Y=1.195
+ $X2=5.63 $Y2=1.3
r116 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.63 $Y=0.465
+ $X2=5.63 $Y2=1.195
r117 23 29 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.38 $Y=1.405
+ $X2=5.38 $Y2=1.3
r118 23 24 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.38 $Y=1.405
+ $X2=5.38 $Y2=2.25
r119 19 25 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.545 $Y=0.365
+ $X2=5.63 $Y2=0.465
r120 19 21 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=5.545 $Y=0.365
+ $X2=4.865 $Y2=0.365
r121 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.295 $Y=2.335
+ $X2=5.38 $Y2=2.25
r122 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.295 $Y=2.335
+ $X2=4.8 $Y2=2.335
r123 13 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.68 $Y=2.065
+ $X2=6.68 $Y2=1.485
r124 9 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.66 $Y=0.555 $X2=6.66
+ $Y2=1.155
r125 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=2.065 $X2=4.8 $Y2=2.335
r126 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.235 $X2=4.865 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_1401_21# 1 2 7 9 10 12 16 20 22 23 24 26
+ 30 33 41 42 45 48 53 56
c156 53 0 1.89563e-19 $X=10.955 $Y=1.32
c157 41 0 2.58372e-20 $X=11.125 $Y=1.53
c158 26 0 1.511e-19 $X=11.76 $Y=1.66
c159 7 0 9.81116e-20 $X=7.08 $Y=0.95
r160 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.165
+ $Y=1.32 $X2=11.165 $Y2=1.32
r161 53 55 32.9707 $w=3.07e-07 $l=2.1e-07 $layer=POLY_cond $X=10.955 $Y=1.32
+ $X2=11.165 $Y2=1.32
r162 52 53 9.4202 $w=3.07e-07 $l=6e-08 $layer=POLY_cond $X=10.895 $Y=1.32
+ $X2=10.955 $Y2=1.32
r163 49 56 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=11.217 $Y=1.53
+ $X2=11.217 $Y2=1.32
r164 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=1.53
+ $X2=11.27 $Y2=1.53
r165 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=1.53
+ $X2=8.05 $Y2=1.53
r166 42 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.195 $Y=1.53
+ $X2=8.05 $Y2=1.53
r167 41 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.125 $Y=1.53
+ $X2=11.27 $Y2=1.53
r168 41 42 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.125 $Y=1.53
+ $X2=8.195 $Y2=1.53
r169 40 49 1.88582 $w=2.73e-07 $l=4.5e-08 $layer=LI1_cond $X=11.217 $Y=1.575
+ $X2=11.217 $Y2=1.53
r170 39 56 16.5533 $w=2.73e-07 $l=3.95e-07 $layer=LI1_cond $X=11.217 $Y=0.925
+ $X2=11.217 $Y2=1.32
r171 37 45 27.1304 $w=2.38e-07 $l=5.65e-07 $layer=LI1_cond $X=7.485 $Y=1.535
+ $X2=8.05 $Y2=1.535
r172 36 37 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=7.32 $Y=1.535
+ $X2=7.485 $Y2=1.535
r173 33 36 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.32 $Y=1.32
+ $X2=7.32 $Y2=1.535
r174 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.32
+ $Y=1.32 $X2=7.32 $Y2=1.32
r175 28 30 16.6464 $w=2.23e-07 $l=3.25e-07 $layer=LI1_cond $X=11.732 $Y=0.755
+ $X2=11.732 $Y2=0.43
r176 24 40 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=11.355 $Y=1.66
+ $X2=11.217 $Y2=1.575
r177 24 26 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=11.355 $Y=1.66
+ $X2=11.76 $Y2=1.66
r178 23 39 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=11.355 $Y=0.84
+ $X2=11.217 $Y2=0.925
r179 22 28 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=11.62 $Y=0.84
+ $X2=11.732 $Y2=0.755
r180 22 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.62 $Y=0.84
+ $X2=11.355 $Y2=0.84
r181 18 53 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.955 $Y=1.155
+ $X2=10.955 $Y2=1.32
r182 18 20 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=10.955 $Y=1.155
+ $X2=10.955 $Y2=0.555
r183 14 52 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.895 $Y=1.485
+ $X2=10.895 $Y2=1.32
r184 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.895 $Y=1.485
+ $X2=10.895 $Y2=2.065
r185 10 34 38.5876 $w=3.28e-07 $l=2.20624e-07 $layer=POLY_cond $X=7.1 $Y=1.485
+ $X2=7.23 $Y2=1.32
r186 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.1 $Y=1.485
+ $X2=7.1 $Y2=2.065
r187 7 34 68.7126 $w=3.28e-07 $l=4.38634e-07 $layer=POLY_cond $X=7.08 $Y=0.95
+ $X2=7.23 $Y2=1.32
r188 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.08 $Y=0.95
+ $X2=7.08 $Y2=0.555
r189 2 26 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=11.635
+ $Y=1.505 $X2=11.76 $Y2=1.66
r190 1 30 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=11.635
+ $Y=0.235 $X2=11.76 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_1888_21# 1 2 9 13 15 17 20 24 28 30 31 33
+ 35 36 38 39 41 44 46 49 53 54 56 57 60 62 65 66 69 70 74 76 78
c195 78 0 1.15981e-19 $X=12.395 $Y=1.16
c196 74 0 1.22108e-19 $X=10.82 $Y=0.687
c197 20 0 1.511e-19 $X=12.455 $Y=1.985
c198 9 0 8.81272e-20 $X=9.515 $Y=0.445
r199 79 86 9.87031 $w=2.93e-07 $l=6e-08 $layer=POLY_cond $X=12.395 $Y=1.16
+ $X2=12.455 $Y2=1.16
r200 78 81 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=12.36 $Y=1.16
+ $X2=12.36 $Y2=1.325
r201 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.395
+ $Y=1.16 $X2=12.395 $Y2=1.16
r202 72 74 4.49631 $w=1.83e-07 $l=7.5e-08 $layer=LI1_cond $X=10.745 $Y=0.687
+ $X2=10.82 $Y2=0.687
r203 69 81 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.325 $Y=1.915
+ $X2=12.325 $Y2=1.325
r204 67 76 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=10.91 $Y=2 $X2=10.82
+ $Y2=2
r205 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.24 $Y=2
+ $X2=12.325 $Y2=1.915
r206 66 67 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=12.24 $Y=2
+ $X2=10.91 $Y2=2
r207 65 76 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.82 $Y=1.915
+ $X2=10.82 $Y2=2
r208 64 74 0.88302 $w=1.8e-07 $l=9.3e-08 $layer=LI1_cond $X=10.82 $Y=0.78
+ $X2=10.82 $Y2=0.687
r209 64 65 69.9343 $w=1.78e-07 $l=1.135e-06 $layer=LI1_cond $X=10.82 $Y=0.78
+ $X2=10.82 $Y2=1.915
r210 63 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.41 $Y=2
+ $X2=10.325 $Y2=2
r211 62 76 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=10.73 $Y=2 $X2=10.82
+ $Y2=2
r212 62 63 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.73 $Y=2 $X2=10.41
+ $Y2=2
r213 58 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.325 $Y=2.085
+ $X2=10.325 $Y2=2
r214 58 60 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.325 $Y=2.085
+ $X2=10.325 $Y2=2.21
r215 56 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.24 $Y=2
+ $X2=10.325 $Y2=2
r216 56 57 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=10.24 $Y=2 $X2=9.8
+ $Y2=2
r217 54 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.74
+ $X2=9.605 $Y2=1.905
r218 54 83 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.74
+ $X2=9.605 $Y2=1.575
r219 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.635
+ $Y=1.74 $X2=9.635 $Y2=1.74
r220 51 57 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.675 $Y=1.915
+ $X2=9.8 $Y2=2
r221 51 53 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=9.675 $Y=1.915
+ $X2=9.675 $Y2=1.74
r222 47 49 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=13.685 $Y=1.61
+ $X2=13.815 $Y2=1.61
r223 42 44 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=13.685 $Y=0.805
+ $X2=13.815 $Y2=0.805
r224 39 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.815 $Y=1.685
+ $X2=13.815 $Y2=1.61
r225 39 41 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=13.815 $Y=1.685
+ $X2=13.815 $Y2=2.085
r226 36 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.815 $Y=0.73
+ $X2=13.815 $Y2=0.805
r227 36 38 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.815 $Y=0.73
+ $X2=13.815 $Y2=0.445
r228 35 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.685 $Y=1.535
+ $X2=13.685 $Y2=1.61
r229 34 46 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.685 $Y=1.295
+ $X2=13.685 $Y2=1.16
r230 34 35 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=13.685 $Y=1.295
+ $X2=13.685 $Y2=1.535
r231 33 46 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.685 $Y=1.025
+ $X2=13.685 $Y2=1.16
r232 32 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.685 $Y=0.88
+ $X2=13.685 $Y2=0.805
r233 32 33 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=13.685 $Y=0.88
+ $X2=13.685 $Y2=1.025
r234 30 46 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=13.61 $Y=1.16
+ $X2=13.685 $Y2=1.16
r235 30 31 146.635 $w=2.7e-07 $l=6.6e-07 $layer=POLY_cond $X=13.61 $Y=1.16
+ $X2=12.95 $Y2=1.16
r236 22 31 12.7172 $w=2.93e-07 $l=7.5e-08 $layer=POLY_cond $X=12.875 $Y=1.16
+ $X2=12.95 $Y2=1.16
r237 22 86 69.0921 $w=2.93e-07 $l=4.2e-07 $layer=POLY_cond $X=12.875 $Y=1.16
+ $X2=12.455 $Y2=1.16
r238 22 28 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=12.875 $Y=1.295
+ $X2=12.875 $Y2=1.985
r239 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.875 $Y=1.025
+ $X2=12.875 $Y2=0.56
r240 18 86 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.455 $Y=1.325
+ $X2=12.455 $Y2=1.16
r241 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.455 $Y=1.325
+ $X2=12.455 $Y2=1.985
r242 15 86 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.455 $Y=0.995
+ $X2=12.455 $Y2=1.16
r243 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.455 $Y=0.995
+ $X2=12.455 $Y2=0.56
r244 13 84 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.515 $Y=2.275
+ $X2=9.515 $Y2=1.905
r245 9 83 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=9.515 $Y=0.445
+ $X2=9.515 $Y2=1.575
r246 2 60 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=2.065 $X2=10.325 $Y2=2.21
r247 1 72 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=10.61
+ $Y=0.235 $X2=10.745 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_1714_47# 1 2 9 13 15 19 24 26 27 29 31 32
c99 32 0 2.58372e-20 $X=10.475 $Y=1.24
c100 31 0 1.75976e-19 $X=10.475 $Y=1.24
c101 26 0 3.84972e-20 $X=9.295 $Y=2.25
r102 32 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.475 $Y=1.24
+ $X2=10.475 $Y2=1.405
r103 32 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.475 $Y=1.24
+ $X2=10.475 $Y2=1.075
r104 31 34 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=10.45 $Y=1.24
+ $X2=10.45 $Y2=1.32
r105 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.475
+ $Y=1.24 $X2=10.475 $Y2=1.24
r106 28 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.38 $Y=1.32
+ $X2=9.295 $Y2=1.32
r107 27 34 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=10.34 $Y=1.32
+ $X2=10.45 $Y2=1.32
r108 27 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.34 $Y=1.32
+ $X2=9.38 $Y2=1.32
r109 25 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=1.405
+ $X2=9.295 $Y2=1.32
r110 25 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=9.295 $Y=1.405
+ $X2=9.295 $Y2=2.25
r111 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=1.235
+ $X2=9.295 $Y2=1.32
r112 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=9.295 $Y=0.465
+ $X2=9.295 $Y2=1.235
r113 19 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.21 $Y=0.365
+ $X2=9.295 $Y2=0.465
r114 19 21 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=9.21 $Y=0.365
+ $X2=8.78 $Y2=0.365
r115 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.21 $Y=2.335
+ $X2=9.295 $Y2=2.25
r116 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.21 $Y=2.335
+ $X2=8.715 $Y2=2.335
r117 13 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.535 $Y=2.065
+ $X2=10.535 $Y2=1.405
r118 9 37 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=10.535 $Y=0.555
+ $X2=10.535 $Y2=1.075
r119 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=8.58
+ $Y=2.065 $X2=8.715 $Y2=2.335
r120 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.57
+ $Y=0.235 $X2=8.78 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%RESET_B 3 7 9 15
r36 12 15 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.755 $Y=1.18
+ $X2=11.97 $Y2=1.18
r37 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.755
+ $Y=1.18 $X2=11.755 $Y2=1.18
r38 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.97 $Y=1.345
+ $X2=11.97 $Y2=1.18
r39 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.97 $Y=1.345
+ $X2=11.97 $Y2=1.825
r40 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.97 $Y=1.015
+ $X2=11.97 $Y2=1.18
r41 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=11.97 $Y=1.015
+ $X2=11.97 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_2696_47# 1 2 7 9 12 14 16 19 23 27 31 34
+ 38
c75 38 0 3.03687e-19 $X=14.71 $Y=1.16
r76 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=14.29 $Y=1.16
+ $X2=14.71 $Y2=1.16
r77 32 37 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=14.205 $Y=1.16
+ $X2=14.29 $Y2=1.16
r78 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.205
+ $Y=1.16 $X2=14.205 $Y2=1.16
r79 29 34 1.17559 $w=3.3e-07 $l=1.58e-07 $layer=LI1_cond $X=13.77 $Y=1.16
+ $X2=13.612 $Y2=1.16
r80 29 31 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=13.77 $Y=1.16
+ $X2=14.205 $Y2=1.16
r81 25 34 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=13.612 $Y=1.325
+ $X2=13.612 $Y2=1.16
r82 25 27 21.4025 $w=3.13e-07 $l=5.85e-07 $layer=LI1_cond $X=13.612 $Y=1.325
+ $X2=13.612 $Y2=1.91
r83 21 34 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=13.612 $Y=0.995
+ $X2=13.612 $Y2=1.16
r84 21 23 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=13.612 $Y=0.995
+ $X2=13.612 $Y2=0.51
r85 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.71 $Y=1.325
+ $X2=14.71 $Y2=1.16
r86 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.71 $Y=1.325
+ $X2=14.71 $Y2=1.985
r87 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.71 $Y=0.995
+ $X2=14.71 $Y2=1.16
r88 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.71 $Y=0.995
+ $X2=14.71 $Y2=0.56
r89 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.29 $Y=1.325
+ $X2=14.29 $Y2=1.16
r90 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.29 $Y=1.325
+ $X2=14.29 $Y2=1.985
r91 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.29 $Y=0.995
+ $X2=14.29 $Y2=1.16
r92 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.29 $Y=0.995
+ $X2=14.29 $Y2=0.56
r93 2 27 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=13.48
+ $Y=1.765 $X2=13.605 $Y2=1.91
r94 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=13.48
+ $Y=0.235 $X2=13.605 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48 52
+ 56 60 64 66 68 73 74 75 79 80 82 84 90 95 103 115 126 130 135 141 144 147 150
+ 153 164 166 169 173
r226 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r227 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r228 167 170 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=14.03 $Y2=2.72
r229 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r230 163 164 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=2.53
+ $X2=12.41 $Y2=2.53
r231 160 163 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=12.19 $Y=2.53
+ $X2=12.245 $Y2=2.53
r232 160 161 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r233 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r234 153 156 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=9.81 $Y=2.34
+ $X2=9.81 $Y2=2.72
r235 150 151 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r236 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r237 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r238 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r239 139 173 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.95 $Y2=2.72
r240 139 170 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.03 $Y2=2.72
r241 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r242 136 169 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=14.245 $Y=2.72
+ $X2=14.097 $Y2=2.72
r243 136 138 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=14.245 $Y=2.72
+ $X2=14.49 $Y2=2.72
r244 135 172 3.93994 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=14.835 $Y=2.72
+ $X2=15.007 $Y2=2.72
r245 135 138 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.835 $Y=2.72
+ $X2=14.49 $Y2=2.72
r246 134 167 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r247 134 161 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r248 133 164 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=12.65 $Y=2.72
+ $X2=12.41 $Y2=2.72
r249 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r250 130 166 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=13 $Y=2.72
+ $X2=13.117 $Y2=2.72
r251 130 133 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=13 $Y=2.72
+ $X2=12.65 $Y2=2.72
r252 129 161 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r253 128 129 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r254 126 160 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=12.135 $Y=2.53
+ $X2=12.19 $Y2=2.53
r255 126 128 18.8111 $w=5.48e-07 $l=8.65e-07 $layer=LI1_cond $X=12.135 $Y=2.53
+ $X2=11.27 $Y2=2.53
r256 125 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r257 125 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=9.89 $Y2=2.72
r258 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r259 122 156 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10 $Y=2.72
+ $X2=9.81 $Y2=2.72
r260 122 124 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=10 $Y=2.72
+ $X2=10.81 $Y2=2.72
r261 121 157 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r262 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r263 118 121 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r264 117 120 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r265 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r266 115 156 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.81 $Y2=2.72
r267 115 120 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.43 $Y2=2.72
r268 114 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r269 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r270 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r271 111 151 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r272 110 113 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r273 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r274 108 150 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=5.895 $Y2=2.72
r275 108 110 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=6.21 $Y2=2.72
r276 107 151 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.75 $Y2=2.72
r277 107 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r278 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r279 104 147 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.64 $Y=2.72
+ $X2=3.467 $Y2=2.72
r280 104 106 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.64 $Y=2.72
+ $X2=3.91 $Y2=2.72
r281 103 150 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=5.895 $Y2=2.72
r282 103 106 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=3.91 $Y2=2.72
r283 102 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r284 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r285 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r286 99 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r287 98 101 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r288 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r289 96 144 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.607 $Y2=2.72
r290 96 98 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r291 95 147 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.467 $Y2=2.72
r292 95 101 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=2.99 $Y2=2.72
r293 94 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r294 94 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r295 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r296 91 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r297 91 93 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r298 90 144 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.607 $Y2=2.72
r299 90 93 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.15 $Y2=2.72
r300 84 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r301 82 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r302 80 84 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r303 80 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r304 79 124 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=10.94 $Y=2.72
+ $X2=10.81 $Y2=2.72
r305 78 79 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=11.105 $Y=2.53
+ $X2=10.94 $Y2=2.53
r306 75 128 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=11.215 $Y=2.53
+ $X2=11.27 $Y2=2.53
r307 75 78 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=11.215 $Y=2.53
+ $X2=11.105 $Y2=2.53
r308 73 113 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.13 $Y2=2.72
r309 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.34 $Y2=2.72
r310 72 117 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=7.59 $Y2=2.72
r311 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=7.34 $Y2=2.72
r312 68 71 32.6526 $w=2.38e-07 $l=6.8e-07 $layer=LI1_cond $X=14.955 $Y=1.66
+ $X2=14.955 $Y2=2.34
r313 66 172 3.13821 $w=2.4e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.955 $Y=2.635
+ $X2=15.007 $Y2=2.72
r314 66 71 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=14.955 $Y=2.635
+ $X2=14.955 $Y2=2.34
r315 62 169 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=14.097 $Y=2.635
+ $X2=14.097 $Y2=2.72
r316 62 64 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=14.097 $Y=2.635
+ $X2=14.097 $Y2=1.94
r317 61 166 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=13.235 $Y=2.72
+ $X2=13.117 $Y2=2.72
r318 60 169 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=13.95 $Y=2.72
+ $X2=14.097 $Y2=2.72
r319 60 61 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=13.95 $Y=2.72
+ $X2=13.235 $Y2=2.72
r320 56 59 33.3473 $w=2.33e-07 $l=6.8e-07 $layer=LI1_cond $X=13.117 $Y=1.66
+ $X2=13.117 $Y2=2.34
r321 54 166 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=13.117 $Y=2.635
+ $X2=13.117 $Y2=2.72
r322 54 59 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=13.117 $Y=2.635
+ $X2=13.117 $Y2=2.34
r323 50 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.34 $Y=2.635
+ $X2=7.34 $Y2=2.72
r324 50 52 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.34 $Y=2.635
+ $X2=7.34 $Y2=2
r325 46 150 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.895 $Y=2.635
+ $X2=5.895 $Y2=2.72
r326 46 48 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=5.895 $Y=2.635
+ $X2=5.895 $Y2=2.29
r327 42 147 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.467 $Y=2.635
+ $X2=3.467 $Y2=2.72
r328 42 44 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=3.467 $Y=2.635
+ $X2=3.467 $Y2=2.3
r329 38 144 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.72
r330 38 40 21.588 $w=3.53e-07 $l=6.65e-07 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=1.97
r331 34 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r332 34 36 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r333 11 71 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=14.785
+ $Y=1.485 $X2=14.92 $Y2=2.34
r334 11 68 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=14.785
+ $Y=1.485 $X2=14.92 $Y2=1.66
r335 10 64 300 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=2 $X=13.89
+ $Y=1.765 $X2=14.08 $Y2=1.94
r336 9 59 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.95
+ $Y=1.485 $X2=13.085 $Y2=2.34
r337 9 56 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=12.95
+ $Y=1.485 $X2=13.085 $Y2=1.66
r338 8 163 600 $w=1.7e-07 $l=9.29637e-07 $layer=licon1_PDIFF $count=1 $X=12.045
+ $Y=1.505 $X2=12.245 $Y2=2.34
r339 7 78 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=10.97
+ $Y=1.645 $X2=11.105 $Y2=2.34
r340 6 153 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=9.59
+ $Y=2.065 $X2=9.785 $Y2=2.34
r341 5 52 300 $w=1.7e-07 $l=4.29651e-07 $layer=licon1_PDIFF $count=2 $X=7.175
+ $Y=1.645 $X2=7.34 $Y2=2
r342 4 48 600 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=2.065 $X2=5.87 $Y2=2.29
r343 3 44 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.065 $X2=3.475 $Y2=2.3
r344 2 40 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.815 $X2=1.62 $Y2=1.97
r345 1 36 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_453_47# 1 2 3 4 13 16 18 19 24 28 29 32
+ 35 41
c114 29 0 1.89491e-19 $X=3.135 $Y=1.19
c115 19 0 1.50346e-19 $X=2.395 $Y=1.875
c116 16 0 6.18549e-20 $X=2.645 $Y=1.075
r117 36 45 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=4.342 $Y=1.19
+ $X2=4.342 $Y2=2.3
r118 36 41 36.8782 $w=2.23e-07 $l=7.2e-07 $layer=LI1_cond $X=4.342 $Y=1.19
+ $X2=4.342 $Y2=0.47
r119 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=1.19
+ $X2=4.37 $Y2=1.19
r120 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.19
+ $X2=2.99 $Y2=1.19
r121 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.19
+ $X2=2.99 $Y2=1.19
r122 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.19
+ $X2=4.37 $Y2=1.19
r123 28 29 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=4.225 $Y=1.19
+ $X2=3.135 $Y2=1.19
r124 27 32 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.73 $Y=1.24
+ $X2=2.99 $Y2=1.24
r125 22 24 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.4 $Y=0.43
+ $X2=2.645 $Y2=0.43
r126 18 19 5.95004 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=1.96
+ $X2=2.395 $Y2=1.875
r127 16 27 9.33298 $w=2.48e-07 $l=2.00237e-07 $layer=LI1_cond $X=2.645 $Y=1.075
+ $X2=2.567 $Y2=1.24
r128 15 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0.595
+ $X2=2.645 $Y2=0.43
r129 15 16 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.645 $Y=0.595
+ $X2=2.645 $Y2=1.075
r130 13 27 9.33298 $w=2.48e-07 $l=1.99825e-07 $layer=LI1_cond $X=2.49 $Y=1.405
+ $X2=2.567 $Y2=1.24
r131 13 19 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.49 $Y=1.405
+ $X2=2.49 $Y2=1.875
r132 4 45 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=2.065 $X2=4.315 $Y2=2.3
r133 3 18 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.815 $X2=2.4 $Y2=1.96
r134 2 41 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.235 $X2=4.315 $Y2=0.47
r135 1 22 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%Q_N 1 2 9 10 11 12 13 18 21
r24 18 21 3.904 $w=2.5e-07 $l=8e-08 $layer=LI1_cond $X=12.705 $Y=0.59 $X2=12.705
+ $Y2=0.51
r25 12 13 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=12.705 $Y=1.815
+ $X2=12.705 $Y2=2.21
r26 11 30 6.85717 $w=2.48e-07 $l=1.23e-07 $layer=LI1_cond $X=12.705 $Y=0.592
+ $X2=12.705 $Y2=0.715
r27 11 18 0.0921954 $w=2.48e-07 $l=2e-09 $layer=LI1_cond $X=12.705 $Y=0.592
+ $X2=12.705 $Y2=0.59
r28 11 21 0.1464 $w=2.5e-07 $l=3e-09 $layer=LI1_cond $X=12.705 $Y=0.507
+ $X2=12.705 $Y2=0.51
r29 10 30 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=12.745 $Y=1.63
+ $X2=12.745 $Y2=0.715
r30 9 12 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=12.705 $Y=1.755
+ $X2=12.705 $Y2=1.815
r31 9 10 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=12.705 $Y=1.755
+ $X2=12.705 $Y2=1.63
r32 2 12 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=12.53
+ $Y=1.485 $X2=12.665 $Y2=1.815
r33 1 21 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=12.53
+ $Y=0.235 $X2=12.665 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%Q 1 2 10 11 12 13 14 15
c21 11 0 1.58152e-19 $X=14.54 $Y=1.57
c22 10 0 1.45535e-19 $X=14.54 $Y=0.825
r23 14 15 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=14.54 $Y=1.82
+ $X2=14.54 $Y2=2.21
r24 11 14 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=14.54 $Y=1.57
+ $X2=14.54 $Y2=1.82
r25 11 12 6.16968 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=14.54 $Y=1.57
+ $X2=14.54 $Y2=1.445
r26 10 12 33.5432 $w=2.03e-07 $l=6.2e-07 $layer=LI1_cond $X=14.562 $Y=0.825
+ $X2=14.562 $Y2=1.445
r27 9 13 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=14.54 $Y=0.7
+ $X2=14.54 $Y2=0.51
r28 9 10 6.16968 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=14.54 $Y=0.7
+ $X2=14.54 $Y2=0.825
r29 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=14.365
+ $Y=1.485 $X2=14.5 $Y2=1.82
r30 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=14.365
+ $Y=0.235 $X2=14.5 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 61 63 67 69 71 74 75 77 78 80 81 82 84 86 92 97 121 128 133 139 142 145 148
+ 151 154 158
c232 158 0 2.71124e-20 $X=14.95 $Y=0
c233 97 0 4.83365e-20 $X=3.37 $Y=0
c234 53 0 1.0279e-19 $X=9.735 $Y=0.36
r235 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r236 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r237 152 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=14.03 $Y2=0
r238 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r239 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r240 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r241 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r242 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r243 137 158 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.95 $Y2=0
r244 137 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.03 $Y2=0
r245 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r246 134 154 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=14.245 $Y=0
+ $X2=14.097 $Y2=0
r247 134 136 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=14.245 $Y=0
+ $X2=14.49 $Y2=0
r248 133 157 3.93994 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=14.835 $Y=0
+ $X2=15.007 $Y2=0
r249 133 136 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.835 $Y=0
+ $X2=14.49 $Y2=0
r250 132 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r251 132 149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r252 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r253 129 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.41 $Y=0
+ $X2=12.245 $Y2=0
r254 129 131 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=12.41 $Y=0
+ $X2=12.65 $Y2=0
r255 128 151 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=13 $Y=0
+ $X2=13.117 $Y2=0
r256 128 131 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=13 $Y=0 $X2=12.65
+ $Y2=0
r257 127 149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r258 126 127 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r259 124 127 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r260 123 126 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r261 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r262 121 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.08 $Y=0
+ $X2=12.245 $Y2=0
r263 121 126 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.08 $Y=0
+ $X2=11.73 $Y2=0
r264 120 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r265 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r266 117 120 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.43 $Y2=0
r267 116 119 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=9.43 $Y2=0
r268 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r269 114 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r270 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r271 111 114 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r272 110 113 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r273 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r274 108 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r275 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r276 105 108 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r277 105 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=3.45 $Y2=0
r278 104 107 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r279 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r280 102 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.7 $Y=0
+ $X2=3.535 $Y2=0
r281 102 104 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.91
+ $Y2=0
r282 101 146 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r283 101 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r284 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r285 98 142 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=1.567 $Y2=0
r286 98 100 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r287 97 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.37 $Y=0
+ $X2=3.535 $Y2=0
r288 97 100 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=3.37 $Y=0 $X2=2.07
+ $Y2=0
r289 96 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r290 96 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r291 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r292 93 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r293 93 95 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r294 92 142 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.43 $Y=0
+ $X2=1.567 $Y2=0
r295 92 95 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.43 $Y=0 $X2=1.15
+ $Y2=0
r296 86 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r297 84 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r298 82 86 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r299 82 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r300 80 119 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=9.56 $Y=0 $X2=9.43
+ $Y2=0
r301 80 81 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.56 $Y=0 $X2=9.69
+ $Y2=0
r302 79 123 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=9.82 $Y=0 $X2=9.89
+ $Y2=0
r303 79 81 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.82 $Y=0 $X2=9.69
+ $Y2=0
r304 77 113 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.645 $Y=0
+ $X2=7.59 $Y2=0
r305 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.645 $Y=0 $X2=7.81
+ $Y2=0
r306 76 116 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.975 $Y=0
+ $X2=8.05 $Y2=0
r307 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=7.81
+ $Y2=0
r308 74 107 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.885 $Y=0
+ $X2=5.75 $Y2=0
r309 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=0 $X2=5.97
+ $Y2=0
r310 73 110 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.055 $Y=0
+ $X2=6.21 $Y2=0
r311 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=0 $X2=5.97
+ $Y2=0
r312 69 157 3.13821 $w=2.4e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.955 $Y=0.085
+ $X2=15.007 $Y2=0
r313 69 71 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=14.955 $Y=0.085
+ $X2=14.955 $Y2=0.38
r314 65 154 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=14.097 $Y=0.085
+ $X2=14.097 $Y2=0
r315 65 67 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=14.097 $Y=0.085
+ $X2=14.097 $Y2=0.38
r316 64 151 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=13.235 $Y=0
+ $X2=13.117 $Y2=0
r317 63 154 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=13.95 $Y=0
+ $X2=14.097 $Y2=0
r318 63 64 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=13.95 $Y=0
+ $X2=13.235 $Y2=0
r319 59 151 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=13.117 $Y=0.085
+ $X2=13.117 $Y2=0
r320 59 61 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=13.117 $Y=0.085
+ $X2=13.117 $Y2=0.38
r321 55 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.245 $Y=0.085
+ $X2=12.245 $Y2=0
r322 55 57 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=12.245 $Y=0.085
+ $X2=12.245 $Y2=0.38
r323 51 81 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=0.085
+ $X2=9.69 $Y2=0
r324 51 53 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=9.69 $Y=0.085
+ $X2=9.69 $Y2=0.36
r325 47 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0
r326 47 49 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0.38
r327 43 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0
r328 43 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0.36
r329 39 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0
r330 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0.36
r331 35 142 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.567 $Y=0.085
+ $X2=1.567 $Y2=0
r332 35 37 16.1342 $w=2.73e-07 $l=3.85e-07 $layer=LI1_cond $X=1.567 $Y=0.085
+ $X2=1.567 $Y2=0.47
r333 31 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r334 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r335 10 71 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=14.785
+ $Y=0.235 $X2=14.92 $Y2=0.38
r336 9 67 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=13.89
+ $Y=0.235 $X2=14.08 $Y2=0.38
r337 8 61 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.95
+ $Y=0.235 $X2=13.085 $Y2=0.38
r338 7 57 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=12.045
+ $Y=0.235 $X2=12.245 $Y2=0.38
r339 6 53 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=9.59
+ $Y=0.235 $X2=9.735 $Y2=0.36
r340 5 49 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.235 $X2=7.81 $Y2=0.38
r341 4 45 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.97 $Y2=0.36
r342 3 41 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.535 $Y2=0.36
r343 2 37 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.47
r344 1 33 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_1251_47# 1 2 7 11 16
r26 14 16 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.39 $Y=0.38
+ $X2=6.555 $Y2=0.38
r27 9 11 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.29 $Y=0.425
+ $X2=7.29 $Y2=0.55
r28 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.205 $Y=0.34
+ $X2=7.29 $Y2=0.425
r29 7 16 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.205 $Y=0.34
+ $X2=6.555 $Y2=0.34
r30 2 11 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=7.155
+ $Y=0.235 $X2=7.29 $Y2=0.55
r31 1 14 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.235 $X2=6.39 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBN_2%A_2004_47# 1 2 7 9 16
r22 9 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=10.245 $Y=0.34
+ $X2=10.245 $Y2=0.46
r23 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.41 $Y=0.34
+ $X2=10.245 $Y2=0.34
r24 7 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.08 $Y=0.34
+ $X2=11.165 $Y2=0.34
r25 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.08 $Y=0.34
+ $X2=10.41 $Y2=0.34
r26 2 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=11.03
+ $Y=0.235 $X2=11.165 $Y2=0.42
r27 1 12 182 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=1 $X=10.02
+ $Y=0.235 $X2=10.245 $Y2=0.46
.ends


* File: sky130_fd_sc_hd__nand4_2.pxi.spice
* Created: Tue Sep  1 19:16:45 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4_2%D N_D_M1004_g N_D_M1002_g N_D_c_73_n N_D_M1013_g
+ N_D_M1008_g D D PM_SKY130_FD_SC_HD__NAND4_2%D
x_PM_SKY130_FD_SC_HD__NAND4_2%C N_C_M1006_g N_C_M1001_g N_C_M1007_g N_C_M1011_g
+ C C N_C_c_124_n PM_SKY130_FD_SC_HD__NAND4_2%C
x_PM_SKY130_FD_SC_HD__NAND4_2%B N_B_M1003_g N_B_M1010_g N_B_M1005_g N_B_M1014_g
+ B B N_B_c_172_n PM_SKY130_FD_SC_HD__NAND4_2%B
x_PM_SKY130_FD_SC_HD__NAND4_2%A N_A_M1009_g N_A_M1000_g N_A_M1015_g N_A_M1012_g
+ N_A_c_218_n A N_A_c_220_n PM_SKY130_FD_SC_HD__NAND4_2%A
x_PM_SKY130_FD_SC_HD__NAND4_2%VPWR N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_M1011_s
+ N_VPWR_M1005_d N_VPWR_M1012_s N_VPWR_c_256_n N_VPWR_c_257_n N_VPWR_c_258_n
+ N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_263_n
+ N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n VPWR N_VPWR_c_267_n
+ N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_255_n PM_SKY130_FD_SC_HD__NAND4_2%VPWR
x_PM_SKY130_FD_SC_HD__NAND4_2%Y N_Y_M1009_d N_Y_M1002_s N_Y_M1001_d N_Y_M1003_s
+ N_Y_M1000_d N_Y_c_324_n N_Y_c_335_n N_Y_c_325_n N_Y_c_338_n N_Y_c_326_n
+ N_Y_c_346_n N_Y_c_356_n N_Y_c_370_n N_Y_c_327_n Y Y Y Y
+ PM_SKY130_FD_SC_HD__NAND4_2%Y
x_PM_SKY130_FD_SC_HD__NAND4_2%A_27_47# N_A_27_47#_M1004_d N_A_27_47#_M1013_d
+ N_A_27_47#_M1007_d N_A_27_47#_c_409_n N_A_27_47#_c_410_n N_A_27_47#_c_411_n
+ N_A_27_47#_c_422_n N_A_27_47#_c_423_n N_A_27_47#_c_412_n
+ PM_SKY130_FD_SC_HD__NAND4_2%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND4_2%VGND N_VGND_M1004_s N_VGND_c_450_n VGND
+ N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n
+ PM_SKY130_FD_SC_HD__NAND4_2%VGND
x_PM_SKY130_FD_SC_HD__NAND4_2%A_277_47# N_A_277_47#_M1006_s N_A_277_47#_M1010_s
+ N_A_277_47#_c_503_n PM_SKY130_FD_SC_HD__NAND4_2%A_277_47#
x_PM_SKY130_FD_SC_HD__NAND4_2%A_471_47# N_A_471_47#_M1010_d N_A_471_47#_M1014_d
+ N_A_471_47#_M1015_s N_A_471_47#_c_525_n N_A_471_47#_c_526_n
+ N_A_471_47#_c_531_n N_A_471_47#_c_527_n N_A_471_47#_c_528_n
+ N_A_471_47#_c_554_n PM_SKY130_FD_SC_HD__NAND4_2%A_471_47#
cc_1 VNB N_D_M1004_g 0.0230765f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_D_c_73_n 0.052468f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_3 VNB N_D_M1013_g 0.017551f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_4 VNB N_D_M1008_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_5 VNB D 0.00806404f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_6 VNB N_C_M1006_g 0.0176998f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_7 VNB N_C_M1001_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_8 VNB N_C_M1007_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_9 VNB N_C_M1011_g 5.16172e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_10 VNB C 0.00467413f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_11 VNB N_C_c_124_n 0.031284f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_12 VNB N_B_M1003_g 5.16172e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_B_M1010_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_14 VNB N_B_M1005_g 5.71338e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_15 VNB N_B_M1014_g 0.017695f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_16 VNB B 0.00215636f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_17 VNB N_B_c_172_n 0.0628192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_M1009_g 0.017202f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_19 VNB N_A_M1000_g 4.69403e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_20 VNB N_A_M1015_g 0.0225092f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_21 VNB N_A_c_218_n 0.0257393f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB A 0.00738464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_c_220_n 0.0372336f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_24 VNB N_VPWR_c_255_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB Y 0.00337456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_409_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_410_n 0.00500854f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_28 VNB N_A_27_47#_c_411_n 0.00924038f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_29 VNB N_A_27_47#_c_412_n 0.00254525f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_30 VNB N_VGND_c_450_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_31 VNB N_VGND_c_451_n 0.0171909f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_32 VNB N_VGND_c_452_n 0.0908251f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_33 VNB N_VGND_c_453_n 0.244463f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_34 VNB N_VGND_c_454_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_35 VNB N_A_277_47#_c_503_n 0.0191566f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_36 VNB N_A_471_47#_c_525_n 0.00247236f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_37 VNB N_A_471_47#_c_526_n 0.00214417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_471_47#_c_527_n 0.00884635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_471_47#_c_528_n 0.0190796f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_40 VPB N_D_M1002_g 0.0274016f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_41 VPB N_D_c_73_n 0.00821255f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.025
cc_42 VPB N_D_M1008_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_43 VPB N_C_M1001_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_C_M1011_g 0.0212126f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_45 VPB N_B_M1003_g 0.0212126f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_46 VPB N_B_M1005_g 0.023005f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_47 VPB N_A_M1000_g 0.0214122f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_48 VPB N_A_M1012_g 0.0257859f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_49 VPB N_A_c_220_n 0.0137892f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_50 VPB N_VPWR_c_256_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_257_n 0.0423592f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_52 VPB N_VPWR_c_258_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_53 VPB N_VPWR_c_259_n 0.0050002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_260_n 0.00564356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_261_n 0.0141015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_262_n 0.00988115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_263_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_264_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_265_n 0.0224008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_266_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_267_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_268_n 0.0211279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_269_n 0.00631492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_255_n 0.0446751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_Y_c_324_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_Y_c_325_n 0.00311143f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_Y_c_326_n 0.00661385f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_68 VPB N_Y_c_327_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB Y 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB Y 0.0023066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB Y 0.00686935f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 N_D_M1013_g N_C_M1006_g 0.0196359f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_73 N_D_M1008_g N_C_M1001_g 0.0196359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_74 N_D_c_73_n C 0.00190331f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_75 D C 0.0141957f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_76 N_D_c_73_n N_C_c_124_n 0.0196359f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_77 N_D_M1002_g N_VPWR_c_257_n 0.00321527f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_78 N_D_c_73_n N_VPWR_c_257_n 0.00534919f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_79 D N_VPWR_c_257_n 0.0151342f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_80 N_D_M1008_g N_VPWR_c_258_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_81 N_D_M1002_g N_VPWR_c_263_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_82 N_D_M1008_g N_VPWR_c_263_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_83 N_D_M1002_g N_VPWR_c_255_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_84 N_D_M1008_g N_VPWR_c_255_n 0.00952874f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_85 N_D_M1002_g N_Y_c_324_n 0.00514019f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_86 N_D_c_73_n N_Y_c_324_n 0.00206439f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_87 N_D_M1008_g N_Y_c_324_n 0.00149073f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_88 D N_Y_c_324_n 0.026643f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_89 N_D_M1002_g N_Y_c_335_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_90 N_D_M1008_g N_Y_c_335_n 0.00975139f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_91 N_D_M1008_g N_Y_c_325_n 0.013439f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_92 N_D_M1008_g N_Y_c_338_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 N_D_M1004_g N_A_27_47#_c_409_n 0.00655349f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_94 N_D_M1013_g N_A_27_47#_c_409_n 5.77896e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_95 N_D_M1004_g N_A_27_47#_c_410_n 0.00845772f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_96 N_D_c_73_n N_A_27_47#_c_410_n 0.00205431f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_97 N_D_M1013_g N_A_27_47#_c_410_n 0.0110274f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_98 D N_A_27_47#_c_410_n 0.0298076f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_99 N_D_M1004_g N_A_27_47#_c_411_n 0.00126954f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_100 N_D_c_73_n N_A_27_47#_c_411_n 0.00693855f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_101 D N_A_27_47#_c_411_n 0.0254514f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_102 N_D_M1013_g N_A_27_47#_c_422_n 0.00244813f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_103 N_D_M1004_g N_A_27_47#_c_423_n 5.17008e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_104 N_D_M1013_g N_A_27_47#_c_423_n 0.00411304f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_105 N_D_M1004_g N_VGND_c_450_n 0.00268723f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_106 N_D_M1013_g N_VGND_c_450_n 0.00268723f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_107 N_D_M1004_g N_VGND_c_451_n 0.00424416f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_108 N_D_M1013_g N_VGND_c_452_n 0.00422898f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_109 N_D_M1004_g N_VGND_c_453_n 0.00669028f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_110 N_D_M1013_g N_VGND_c_453_n 0.00577235f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_111 N_C_M1011_g N_B_M1003_g 0.0194789f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_112 C B 0.00647256f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_113 N_C_c_124_n B 9.59916e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_114 C N_B_c_172_n 2.03866e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_115 N_C_c_124_n N_B_c_172_n 0.0194789f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C_M1001_g N_VPWR_c_258_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_117 N_C_M1011_g N_VPWR_c_259_n 0.00575644f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_118 N_C_M1001_g N_VPWR_c_267_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_119 N_C_M1011_g N_VPWR_c_267_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_120 N_C_M1001_g N_VPWR_c_255_n 0.00952874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_121 N_C_M1011_g N_VPWR_c_255_n 0.00996204f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_122 N_C_M1001_g N_Y_c_335_n 6.1949e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_123 N_C_M1001_g N_Y_c_325_n 0.0119784f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_124 C N_Y_c_325_n 0.021194f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_125 N_C_M1001_g N_Y_c_338_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C_M1011_g N_Y_c_338_n 0.0104675f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_127 N_C_M1011_g N_Y_c_326_n 0.0143001f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_128 C N_Y_c_326_n 0.00101487f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_129 N_C_M1011_g N_Y_c_346_n 6.59253e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_130 N_C_M1001_g N_Y_c_327_n 0.00149073f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_131 N_C_M1011_g N_Y_c_327_n 0.00149073f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_132 C N_Y_c_327_n 0.026643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_133 N_C_c_124_n N_Y_c_327_n 0.00206439f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_134 C N_A_27_47#_c_410_n 0.00978542f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_135 N_C_M1006_g N_A_27_47#_c_412_n 0.0103313f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_136 N_C_M1007_g N_A_27_47#_c_412_n 0.00866705f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_137 C N_A_27_47#_c_412_n 0.00368637f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_138 N_C_M1006_g N_VGND_c_452_n 0.00357877f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_139 N_C_M1007_g N_VGND_c_452_n 0.00357877f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_140 N_C_M1006_g N_VGND_c_453_n 0.00525237f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_141 N_C_M1007_g N_VGND_c_453_n 0.00655123f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_142 N_C_M1006_g N_A_277_47#_c_503_n 0.00383287f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_143 N_C_M1007_g N_A_277_47#_c_503_n 0.015881f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_144 C N_A_277_47#_c_503_n 0.0256202f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_145 N_C_c_124_n N_A_277_47#_c_503_n 0.00207887f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B_M1014_g N_A_M1009_g 0.0133029f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_147 N_B_M1005_g N_A_M1000_g 0.0160214f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B_c_172_n N_A_c_218_n 0.0133029f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_149 N_B_M1003_g N_VPWR_c_259_n 0.00708399f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B_M1005_g N_VPWR_c_260_n 0.00990358f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B_M1003_g N_VPWR_c_265_n 0.00541359f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B_M1005_g N_VPWR_c_265_n 0.00541359f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B_M1003_g N_VPWR_c_255_n 0.00996204f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B_M1005_g N_VPWR_c_255_n 0.0104583f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B_M1003_g N_Y_c_338_n 6.59253e-19 $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B_M1003_g N_Y_c_326_n 0.0130107f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_157 B N_Y_c_326_n 0.00836582f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_158 N_B_M1003_g N_Y_c_346_n 0.0104675f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B_M1005_g N_Y_c_346_n 0.016848f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B_M1014_g N_Y_c_356_n 8.95831e-19 $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_161 N_B_M1003_g Y 0.00149073f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_162 N_B_M1005_g Y 0.00149073f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_163 B Y 0.026643f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_164 N_B_c_172_n Y 0.00206439f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B_M1005_g Y 0.00295344f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_166 B Y 0.0115915f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_167 N_B_c_172_n Y 0.00301214f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B_M1005_g Y 0.0137699f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_169 B Y 0.0286839f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_170 N_B_c_172_n Y 0.0123886f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B_M1010_g N_VGND_c_452_n 0.00357877f $X=2.71 $Y=0.56 $X2=0 $Y2=0
cc_172 N_B_M1014_g N_VGND_c_452_n 0.00357877f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_173 N_B_M1010_g N_VGND_c_453_n 0.00655123f $X=2.71 $Y=0.56 $X2=0 $Y2=0
cc_174 N_B_M1014_g N_VGND_c_453_n 0.00525237f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_175 N_B_M1010_g N_A_277_47#_c_503_n 0.0145787f $X=2.71 $Y=0.56 $X2=0 $Y2=0
cc_176 N_B_M1014_g N_A_277_47#_c_503_n 0.00401078f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_177 B N_A_277_47#_c_503_n 0.0627795f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_178 N_B_c_172_n N_A_277_47#_c_503_n 0.0129039f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B_M1010_g N_A_471_47#_c_525_n 0.00866705f $X=2.71 $Y=0.56 $X2=0 $Y2=0
cc_180 N_B_M1014_g N_A_471_47#_c_525_n 0.0124168f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_M1000_g N_VPWR_c_260_n 0.010343f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_M1012_g N_VPWR_c_262_n 0.0247226f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_183 A N_VPWR_c_262_n 0.0211194f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A_c_220_n N_VPWR_c_262_n 0.00811148f $X=4.33 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_M1000_g N_VPWR_c_268_n 0.00541359f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_M1012_g N_VPWR_c_268_n 0.00541359f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_M1000_g N_VPWR_c_255_n 0.0104583f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_M1012_g N_VPWR_c_255_n 0.0106948f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_M1009_g N_Y_c_356_n 0.00716109f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A_M1015_g N_Y_c_356_n 0.00963157f $X=3.97 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_c_218_n N_Y_c_356_n 0.00519633f $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_M1000_g N_Y_c_370_n 0.016201f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_M1012_g N_Y_c_370_n 0.00902485f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_M1000_g Y 0.0181424f $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_M1012_g Y 0.0108883f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_c_218_n Y 0.0232981f $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_197 A Y 0.0117914f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_198 N_A_M1000_g Y 6.15761e-19 $X=3.55 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_M1009_g N_VGND_c_452_n 0.00357877f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_M1015_g N_VGND_c_452_n 0.00357877f $X=3.97 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_M1009_g N_VGND_c_453_n 0.00525237f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A_M1015_g N_VGND_c_453_n 0.00638167f $X=3.97 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_M1009_g N_A_471_47#_c_531_n 0.0102564f $X=3.55 $Y=0.56 $X2=0 $Y2=0
cc_204 N_A_M1015_g N_A_471_47#_c_531_n 0.01694f $X=3.97 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A_c_218_n N_A_471_47#_c_531_n 2.87379e-19 $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_M1015_g N_A_471_47#_c_528_n 0.0085369f $X=3.97 $Y=0.56 $X2=0 $Y2=0
cc_207 A N_A_471_47#_c_528_n 0.0210369f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_208 N_A_c_220_n N_A_471_47#_c_528_n 0.00838601f $X=4.33 $Y=1.16 $X2=0 $Y2=0
cc_209 N_VPWR_c_255_n N_Y_M1002_s 0.00215201f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_210 N_VPWR_c_255_n N_Y_M1001_d 0.00215201f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_211 N_VPWR_c_255_n N_Y_M1003_s 0.00215201f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_212 N_VPWR_c_255_n N_Y_M1000_d 0.00215201f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_263_n N_Y_c_335_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_255_n N_Y_c_335_n 0.0122217f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_M1008_d N_Y_c_325_n 0.00167154f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_216 N_VPWR_c_258_n N_Y_c_325_n 0.0129161f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_217 N_VPWR_c_267_n N_Y_c_338_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_255_n N_Y_c_338_n 0.0122217f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_M1011_s N_Y_c_326_n 0.00407949f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_220 N_VPWR_c_259_n N_Y_c_326_n 0.0261634f $X=2.02 $Y=2 $X2=0 $Y2=0
cc_221 N_VPWR_c_260_n N_Y_c_346_n 0.0308572f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_222 N_VPWR_c_265_n N_Y_c_346_n 0.0189039f $X=2.995 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_c_255_n N_Y_c_346_n 0.0122217f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_c_260_n N_Y_c_370_n 0.034303f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_225 N_VPWR_c_268_n N_Y_c_370_n 0.0189039f $X=4.095 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_c_255_n N_Y_c_370_n 0.0122217f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_M1005_d Y 0.00258327f $X=2.805 $Y=1.485 $X2=0 $Y2=0
cc_228 N_VPWR_c_262_n Y 0.0405409f $X=4.26 $Y=1.66 $X2=0 $Y2=0
cc_229 N_VPWR_M1005_d Y 0.0140969f $X=2.805 $Y=1.485 $X2=0 $Y2=0
cc_230 N_VPWR_c_260_n Y 0.027157f $X=3.16 $Y=2 $X2=0 $Y2=0
cc_231 N_VPWR_c_257_n N_A_27_47#_c_411_n 7.42972e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_232 N_VPWR_c_262_n N_A_471_47#_c_528_n 0.00284499f $X=4.26 $Y=1.66 $X2=0
+ $Y2=0
cc_233 N_Y_c_325_n N_A_27_47#_c_410_n 0.00730782f $X=1.355 $Y=1.555 $X2=0 $Y2=0
cc_234 N_Y_M1009_d N_VGND_c_453_n 0.00216833f $X=3.625 $Y=0.235 $X2=0 $Y2=0
cc_235 N_Y_c_326_n N_A_277_47#_c_503_n 0.0182712f $X=2.355 $Y=1.555 $X2=0 $Y2=0
cc_236 N_Y_c_356_n N_A_277_47#_c_503_n 6.16413e-19 $X=3.76 $Y=0.72 $X2=0 $Y2=0
cc_237 Y N_A_471_47#_c_526_n 0.0045377f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_238 Y N_A_471_47#_c_526_n 0.00392188f $X=3.37 $Y=1.445 $X2=0 $Y2=0
cc_239 N_Y_M1009_d N_A_471_47#_c_531_n 0.00305226f $X=3.625 $Y=0.235 $X2=0 $Y2=0
cc_240 N_Y_c_356_n N_A_471_47#_c_531_n 0.016329f $X=3.76 $Y=0.72 $X2=0 $Y2=0
cc_241 Y N_A_471_47#_c_531_n 0.00423076f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_242 N_Y_c_356_n N_A_471_47#_c_528_n 0.0109215f $X=3.76 $Y=0.72 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_410_n N_VGND_M1004_s 0.00169589f $X=0.935 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_27_47#_c_410_n N_VGND_c_450_n 0.0111177f $X=0.935 $Y=0.82 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_409_n N_VGND_c_451_n 0.0213324f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_410_n N_VGND_c_451_n 0.00193763f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_410_n N_VGND_c_452_n 0.00193763f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_422_n N_VGND_c_452_n 0.0152108f $X=1.06 $Y=0.465 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_412_n N_VGND_c_452_n 0.053439f $X=1.96 $Y=0.38 $X2=0 $Y2=0
cc_250 N_A_27_47#_M1004_d N_VGND_c_453_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1013_d N_VGND_c_453_n 0.00215206f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1007_d N_VGND_c_453_n 0.00225742f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_409_n N_VGND_c_453_n 0.0126042f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_410_n N_VGND_c_453_n 0.00828806f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_422_n N_VGND_c_453_n 0.00940698f $X=1.06 $Y=0.465 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_412_n N_VGND_c_453_n 0.0336592f $X=1.96 $Y=0.38 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_412_n N_A_277_47#_M1006_s 0.00305599f $X=1.96 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_258 N_A_27_47#_M1007_d N_A_277_47#_c_503_n 0.00369694f $X=1.805 $Y=0.235
+ $X2=0 $Y2=0
cc_259 N_A_27_47#_c_410_n N_A_277_47#_c_503_n 0.00799569f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_412_n N_A_277_47#_c_503_n 0.0425424f $X=1.96 $Y=0.38 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_412_n N_A_471_47#_c_525_n 0.0180052f $X=1.96 $Y=0.38 $X2=0
+ $Y2=0
cc_262 N_VGND_c_453_n N_A_277_47#_M1006_s 0.00216833f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_263 N_VGND_c_453_n N_A_277_47#_M1010_s 0.00216833f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_264 N_VGND_c_452_n N_A_277_47#_c_503_n 0.00358979f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_453_n N_A_277_47#_c_503_n 0.00861284f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_453_n N_A_471_47#_M1010_d 0.00225742f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_267 N_VGND_c_453_n N_A_471_47#_M1014_d 0.0021521f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_453_n N_A_471_47#_M1015_s 0.00292107f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_452_n N_A_471_47#_c_525_n 0.053439f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_270 N_VGND_c_453_n N_A_471_47#_c_525_n 0.0336592f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_271 N_VGND_c_452_n N_A_471_47#_c_531_n 0.0362657f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_453_n N_A_471_47#_c_531_n 0.0236233f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_273 N_VGND_c_452_n N_A_471_47#_c_527_n 0.0229144f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_274 N_VGND_c_453_n N_A_471_47#_c_527_n 0.0126939f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_452_n N_A_471_47#_c_554_n 0.0114055f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_453_n N_A_471_47#_c_554_n 0.00653405f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_277 N_A_277_47#_c_503_n N_A_471_47#_M1010_d 0.00369694f $X=2.92 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_278 N_A_277_47#_M1010_s N_A_471_47#_c_525_n 0.00305599f $X=2.785 $Y=0.235
+ $X2=0 $Y2=0
cc_279 N_A_277_47#_c_503_n N_A_471_47#_c_525_n 0.0425424f $X=2.92 $Y=0.72 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__a2bb2oi_4.pxi.spice
* Created: Tue Sep  1 18:54:20 2020
* 
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%B1 N_B1_c_154_n N_B1_M1014_g N_B1_M1004_g
+ N_B1_c_155_n N_B1_M1023_g N_B1_M1007_g N_B1_c_156_n N_B1_M1034_g N_B1_M1024_g
+ N_B1_c_157_n N_B1_M1038_g N_B1_M1036_g N_B1_c_158_n N_B1_c_168_n N_B1_c_207_p
+ N_B1_c_159_n N_B1_c_160_n N_B1_c_161_n B1 N_B1_c_162_n B1
+ PM_SKY130_FD_SC_HD__A2BB2OI_4%B1
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%B2 N_B2_c_279_n N_B2_M1018_g N_B2_M1001_g
+ N_B2_c_280_n N_B2_M1019_g N_B2_M1008_g N_B2_c_281_n N_B2_M1025_g N_B2_M1027_g
+ N_B2_c_282_n N_B2_M1033_g N_B2_M1035_g B2 N_B2_c_283_n N_B2_c_284_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_4%B2
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%A_751_21# N_A_751_21#_M1010_d
+ N_A_751_21#_M1016_d N_A_751_21#_M1017_d N_A_751_21#_M1031_d
+ N_A_751_21#_M1012_s N_A_751_21#_M1029_s N_A_751_21#_c_344_n
+ N_A_751_21#_M1000_g N_A_751_21#_M1003_g N_A_751_21#_c_345_n
+ N_A_751_21#_M1006_g N_A_751_21#_M1011_g N_A_751_21#_c_346_n
+ N_A_751_21#_M1030_g N_A_751_21#_M1015_g N_A_751_21#_c_347_n
+ N_A_751_21#_M1039_g N_A_751_21#_M1021_g N_A_751_21#_c_348_n
+ N_A_751_21#_c_349_n N_A_751_21#_c_350_n N_A_751_21#_c_351_n
+ N_A_751_21#_c_379_p N_A_751_21#_c_352_n N_A_751_21#_c_383_p
+ N_A_751_21#_c_353_n N_A_751_21#_c_391_p N_A_751_21#_c_366_n
+ N_A_751_21#_c_354_n N_A_751_21#_c_410_p N_A_751_21#_c_367_n
+ N_A_751_21#_c_355_n N_A_751_21#_c_356_n N_A_751_21#_c_357_n
+ N_A_751_21#_c_358_n N_A_751_21#_c_359_n N_A_751_21#_c_369_n
+ N_A_751_21#_c_360_n N_A_751_21#_c_370_n N_A_751_21#_c_361_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_4%A_751_21#
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%A1_N N_A1_N_c_559_n N_A1_N_M1010_g
+ N_A1_N_M1002_g N_A1_N_c_560_n N_A1_N_M1013_g N_A1_N_M1005_g N_A1_N_c_561_n
+ N_A1_N_M1016_g N_A1_N_M1009_g N_A1_N_c_562_n N_A1_N_M1020_g N_A1_N_M1028_g
+ A1_N N_A1_N_c_563_n N_A1_N_c_564_n PM_SKY130_FD_SC_HD__A2BB2OI_4%A1_N
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%A2_N N_A2_N_c_641_n N_A2_N_M1017_g
+ N_A2_N_M1012_g N_A2_N_c_642_n N_A2_N_M1026_g N_A2_N_M1022_g N_A2_N_c_643_n
+ N_A2_N_M1031_g N_A2_N_M1029_g N_A2_N_c_644_n N_A2_N_M1032_g N_A2_N_M1037_g
+ A2_N N_A2_N_c_645_n N_A2_N_c_646_n PM_SKY130_FD_SC_HD__A2BB2OI_4%A2_N
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%A_27_297# N_A_27_297#_M1004_s
+ N_A_27_297#_M1007_s N_A_27_297#_M1001_s N_A_27_297#_M1027_s
+ N_A_27_297#_M1036_s N_A_27_297#_M1011_d N_A_27_297#_M1021_d
+ N_A_27_297#_c_721_n N_A_27_297#_c_722_n N_A_27_297#_c_723_n
+ N_A_27_297#_c_724_n N_A_27_297#_c_742_n N_A_27_297#_c_746_n
+ N_A_27_297#_c_747_n N_A_27_297#_c_749_n N_A_27_297#_c_756_n
+ N_A_27_297#_c_784_p N_A_27_297#_c_811_p N_A_27_297#_c_758_n
+ N_A_27_297#_c_725_n N_A_27_297#_c_726_n N_A_27_297#_c_774_p
+ N_A_27_297#_c_750_n N_A_27_297#_c_751_n N_A_27_297#_c_787_p
+ PM_SKY130_FD_SC_HD__A2BB2OI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%VPWR N_VPWR_M1004_d N_VPWR_M1024_d
+ N_VPWR_M1008_d N_VPWR_M1035_d N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_c_818_n
+ N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n
+ N_VPWR_c_824_n N_VPWR_c_825_n N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n
+ N_VPWR_c_829_n VPWR N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_832_n
+ N_VPWR_c_833_n N_VPWR_c_817_n N_VPWR_c_835_n N_VPWR_c_836_n N_VPWR_c_837_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%Y N_Y_M1018_d N_Y_M1025_d N_Y_M1000_s
+ N_Y_M1030_s N_Y_M1003_s N_Y_M1015_s N_Y_c_961_n N_Y_c_962_n N_Y_c_963_n
+ N_Y_c_979_n N_Y_c_1025_n N_Y_c_968_n N_Y_c_969_n N_Y_c_964_n N_Y_c_1012_n
+ N_Y_c_965_n N_Y_c_966_n Y Y N_Y_c_1029_n PM_SKY130_FD_SC_HD__A2BB2OI_4%Y
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%A_1139_297# N_A_1139_297#_M1002_s
+ N_A_1139_297#_M1005_s N_A_1139_297#_M1028_s N_A_1139_297#_M1022_d
+ N_A_1139_297#_M1037_d N_A_1139_297#_c_1058_n N_A_1139_297#_c_1059_n
+ N_A_1139_297#_c_1060_n N_A_1139_297#_c_1113_n N_A_1139_297#_c_1061_n
+ N_A_1139_297#_c_1062_n N_A_1139_297#_c_1117_n N_A_1139_297#_c_1072_n
+ N_A_1139_297#_c_1075_n N_A_1139_297#_c_1079_n N_A_1139_297#_c_1063_n
+ N_A_1139_297#_c_1080_n PM_SKY130_FD_SC_HD__A2BB2OI_4%A_1139_297#
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%VGND N_VGND_M1014_d N_VGND_M1023_d
+ N_VGND_M1038_d N_VGND_M1006_d N_VGND_M1039_d N_VGND_M1013_s N_VGND_M1020_s
+ N_VGND_M1026_s N_VGND_M1032_s N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n
+ N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n N_VGND_c_1131_n
+ N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n
+ N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n N_VGND_c_1139_n
+ N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n N_VGND_c_1143_n
+ N_VGND_c_1144_n N_VGND_c_1145_n VGND N_VGND_c_1146_n N_VGND_c_1147_n
+ N_VGND_c_1148_n N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_4%VGND
x_PM_SKY130_FD_SC_HD__A2BB2OI_4%A_109_47# N_A_109_47#_M1014_s
+ N_A_109_47#_M1034_s N_A_109_47#_M1019_s N_A_109_47#_M1033_s
+ N_A_109_47#_c_1287_n N_A_109_47#_c_1284_n N_A_109_47#_c_1285_n
+ N_A_109_47#_c_1298_n N_A_109_47#_c_1286_n N_A_109_47#_c_1303_n
+ PM_SKY130_FD_SC_HD__A2BB2OI_4%A_109_47#
cc_1 VNB N_B1_c_154_n 0.0216231f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B1_c_155_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_B1_c_156_n 0.0159983f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_B1_c_157_n 0.0161959f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.995
cc_5 VNB N_B1_c_158_n 3.4661e-19 $X=-0.19 $Y=-0.24 $X2=1.47 $Y2=1.445
cc_6 VNB N_B1_c_159_n 0.00347218f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.16
cc_7 VNB N_B1_c_160_n 0.0189915f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.16
cc_8 VNB N_B1_c_161_n 0.0210139f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=1.18
cc_9 VNB N_B1_c_162_n 0.0529737f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_10 VNB N_B2_c_279_n 0.0161471f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_11 VNB N_B2_c_280_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_12 VNB N_B2_c_281_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_13 VNB N_B2_c_282_n 0.0159974f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.995
cc_14 VNB N_B2_c_283_n 0.0014172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B2_c_284_n 0.0626151f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_16 VNB N_A_751_21#_c_344_n 0.0150886f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_17 VNB N_A_751_21#_c_345_n 0.0157866f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.985
cc_18 VNB N_A_751_21#_c_346_n 0.0157824f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.445
cc_19 VNB N_A_751_21#_c_347_n 0.0195882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_751_21#_c_348_n 0.0209354f $X=-0.19 $Y=-0.24 $X2=1.235 $Y2=1.16
cc_21 VNB N_A_751_21#_c_349_n 0.00467747f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_22 VNB N_A_751_21#_c_350_n 0.00345181f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.18
cc_23 VNB N_A_751_21#_c_351_n 3.34189e-19 $X=-0.19 $Y=-0.24 $X2=1.235 $Y2=1.18
cc_24 VNB N_A_751_21#_c_352_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_751_21#_c_353_n 0.00386497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_751_21#_c_354_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_751_21#_c_355_n 0.014973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_751_21#_c_356_n 0.0234981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_751_21#_c_357_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_751_21#_c_358_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_751_21#_c_359_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_751_21#_c_360_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_751_21#_c_361_n 0.0664243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A1_N_c_559_n 0.0193125f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_35 VNB N_A1_N_c_560_n 0.0157992f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_36 VNB N_A1_N_c_561_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_37 VNB N_A1_N_c_562_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.995
cc_38 VNB N_A1_N_c_563_n 0.00310534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A1_N_c_564_n 0.0682635f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_40 VNB N_A2_N_c_641_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_41 VNB N_A2_N_c_642_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_42 VNB N_A2_N_c_643_n 0.0157986f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_43 VNB N_A2_N_c_644_n 0.0192362f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.995
cc_44 VNB N_A2_N_c_645_n 0.00432859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A2_N_c_646_n 0.0660089f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_46 VNB N_VPWR_c_817_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_Y_c_961_n 0.00611208f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_48 VNB N_Y_c_962_n 0.00976856f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.325
cc_49 VNB N_Y_c_963_n 0.00401215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_964_n 0.00440484f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_51 VNB N_Y_c_965_n 4.62713e-19 $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.16
cc_52 VNB N_Y_c_966_n 0.00254034f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_53 VNB N_VGND_c_1125_n 0.0110498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1126_n 0.00622824f $X=-0.19 $Y=-0.24 $X2=1.47 $Y2=1.445
cc_55 VNB N_VGND_c_1127_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.16
cc_56 VNB N_VGND_c_1128_n 0.0041055f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=1.18
cc_57 VNB N_VGND_c_1129_n 0.00359327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1130_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=1.235 $Y2=1.16
cc_59 VNB N_VGND_c_1131_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.16
cc_60 VNB N_VGND_c_1132_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_61 VNB N_VGND_c_1133_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1134_n 0.0538772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1135_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1136_n 0.0170081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1137_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1138_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1139_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1140_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1141_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1142_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1143_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1144_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1145_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1146_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1147_n 0.0135861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1148_n 0.451309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1149_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1150_n 0.0176493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1151_n 0.019738f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_109_47#_c_1284_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_81 VNB N_A_109_47#_c_1285_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_82 VNB N_A_109_47#_c_1286_n 0.00248542f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_83 VPB N_B1_M1004_g 0.0252519f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_84 VPB N_B1_M1007_g 0.0182139f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_85 VPB N_B1_M1024_g 0.0185416f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_86 VPB N_B1_M1036_g 0.0172299f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_87 VPB N_B1_c_158_n 0.00253572f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=1.445
cc_88 VPB N_B1_c_168_n 0.0118888f $X=-0.19 $Y=1.305 $X2=3.245 $Y2=1.53
cc_89 VPB N_B1_c_159_n 0.00229947f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.16
cc_90 VPB N_B1_c_160_n 0.00441099f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.16
cc_91 VPB N_B1_c_162_n 0.0078521f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_92 VPB N_B2_M1001_g 0.0183498f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_93 VPB N_B2_M1008_g 0.0181173f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_94 VPB N_B2_M1027_g 0.018119f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_95 VPB N_B2_M1035_g 0.0183386f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_96 VPB N_B2_c_284_n 0.0100802f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_97 VPB N_A_751_21#_M1003_g 0.0171748f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=0.56
cc_98 VPB N_A_751_21#_M1011_g 0.0178559f $X=-0.19 $Y=1.305 $X2=3.245 $Y2=1.53
cc_99 VPB N_A_751_21#_M1015_g 0.0178517f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=1.18
cc_100 VPB N_A_751_21#_M1021_g 0.0253782f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.16
cc_101 VPB N_A_751_21#_c_366_n 0.0023954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_751_21#_c_367_n 0.0210962f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_751_21#_c_356_n 0.00910387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_751_21#_c_369_n 0.00231717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_751_21#_c_370_n 0.00206552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_751_21#_c_361_n 0.0105881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A1_N_M1002_g 0.0252519f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_108 VPB N_A1_N_M1005_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_109 VPB N_A1_N_M1009_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_110 VPB N_A1_N_M1028_g 0.0185045f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_111 VPB N_A1_N_c_564_n 0.0108808f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_112 VPB N_A2_N_M1012_g 0.018818f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_113 VPB N_A2_N_M1022_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_114 VPB N_A2_N_M1029_g 0.0182024f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_115 VPB N_A2_N_M1037_g 0.0220253f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_116 VPB N_A2_N_c_646_n 0.0102978f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_117 VPB N_A_27_297#_c_721_n 0.0332602f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=0.56
cc_118 VPB N_A_27_297#_c_722_n 0.00226814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_297#_c_723_n 0.0107079f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=1.285
cc_120 VPB N_A_27_297#_c_724_n 0.00217577f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=1.445
cc_121 VPB N_A_27_297#_c_725_n 0.00182586f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_122 VPB N_A_27_297#_c_726_n 0.0105904f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.18
cc_123 VPB N_VPWR_c_818_n 0.00428214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_819_n 0.00393015f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.325
cc_125 VPB N_VPWR_c_820_n 0.00393015f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=1.285
cc_126 VPB N_VPWR_c_821_n 0.00454762f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.445
cc_127 VPB N_VPWR_c_822_n 0.00428214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_823_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_129 VPB N_VPWR_c_824_n 0.0158243f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.16
cc_130 VPB N_VPWR_c_825_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.16
cc_131 VPB N_VPWR_c_826_n 0.0151708f $X=-0.19 $Y=1.305 $X2=1.235 $Y2=1.16
cc_132 VPB N_VPWR_c_827_n 0.00478242f $X=-0.19 $Y=1.305 $X2=1.235 $Y2=1.16
cc_133 VPB N_VPWR_c_828_n 0.0151708f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_134 VPB N_VPWR_c_829_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_830_n 0.0177718f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_136 VPB N_VPWR_c_831_n 0.0671338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_832_n 0.0164723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_833_n 0.0615611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_817_n 0.0631827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_835_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_836_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_837_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_Y_c_963_n 0.00166564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_Y_c_968_n 0.00226767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_Y_c_969_n 0.00291497f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=1.18
cc_146 VPB Y 0.00241364f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_147 VPB N_A_1139_297#_c_1058_n 0.00775861f $X=-0.19 $Y=1.305 $X2=1.31
+ $Y2=1.325
cc_148 VPB N_A_1139_297#_c_1059_n 0.00235794f $X=-0.19 $Y=1.305 $X2=3.41
+ $Y2=0.995
cc_149 VPB N_A_1139_297#_c_1060_n 0.00587207f $X=-0.19 $Y=1.305 $X2=3.41
+ $Y2=0.56
cc_150 VPB N_A_1139_297#_c_1061_n 0.00249473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_1139_297#_c_1062_n 0.00398447f $X=-0.19 $Y=1.305 $X2=1.47
+ $Y2=1.445
cc_152 VPB N_A_1139_297#_c_1063_n 0.00198944f $X=-0.19 $Y=1.305 $X2=0.555
+ $Y2=1.16
cc_153 N_B1_c_156_n N_B2_c_279_n 0.0237807f $X=1.31 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_154 N_B1_M1024_g N_B2_M1001_g 0.0237807f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B1_c_168_n N_B2_M1001_g 0.0125227f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B1_c_168_n N_B2_M1008_g 0.0103848f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_157 N_B1_c_168_n N_B2_M1027_g 0.010429f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_158 N_B1_c_157_n N_B2_c_282_n 0.0266272f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B1_M1036_g N_B2_M1035_g 0.0433771f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B1_c_168_n N_B2_M1035_g 0.0103848f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_161 N_B1_c_168_n N_B2_c_283_n 0.095778f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_162 N_B1_c_159_n N_B2_c_283_n 0.0175089f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_163 N_B1_c_160_n N_B2_c_283_n 6.99391e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B1_c_161_n N_B2_c_283_n 0.0176509f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_165 N_B1_c_158_n N_B2_c_284_n 0.00361105f $X=1.47 $Y=1.445 $X2=0 $Y2=0
cc_166 N_B1_c_168_n N_B2_c_284_n 0.00642092f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_167 N_B1_c_159_n N_B2_c_284_n 0.00458937f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B1_c_160_n N_B2_c_284_n 0.0223811f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B1_c_161_n N_B2_c_284_n 0.00212345f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_170 N_B1_c_162_n N_B2_c_284_n 0.0237807f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B1_c_157_n N_A_751_21#_c_344_n 0.0257803f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_M1036_g N_A_751_21#_M1003_g 0.0275835f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B1_c_168_n N_A_751_21#_M1003_g 6.56566e-19 $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_174 N_B1_c_159_n N_A_751_21#_c_361_n 0.00110695f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B1_c_160_n N_A_751_21#_c_361_n 0.0212433f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B1_c_168_n N_A_27_297#_M1001_s 0.00169858f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_177 N_B1_c_168_n N_A_27_297#_M1027_s 0.00169858f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_178 N_B1_c_168_n N_A_27_297#_M1036_s 0.00148539f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_179 N_B1_M1004_g N_A_27_297#_c_721_n 0.0102794f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B1_M1007_g N_A_27_297#_c_721_n 6.39698e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B1_M1004_g N_A_27_297#_c_722_n 0.0106747f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B1_M1007_g N_A_27_297#_c_722_n 0.0132081f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_c_161_n N_A_27_297#_c_722_n 0.0388745f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_184 N_B1_c_162_n N_A_27_297#_c_722_n 0.00211509f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_185 N_B1_M1004_g N_A_27_297#_c_723_n 0.00149004f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_c_161_n N_A_27_297#_c_723_n 0.0275988f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_187 N_B1_M1024_g N_A_27_297#_c_724_n 2.51853e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B1_c_207_p N_A_27_297#_c_724_n 0.00812971f $X=1.555 $Y=1.53 $X2=0 $Y2=0
cc_189 N_B1_c_161_n N_A_27_297#_c_724_n 0.0196366f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_190 N_B1_c_162_n N_A_27_297#_c_724_n 0.00220041f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B1_M1024_g N_A_27_297#_c_742_n 0.0118746f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B1_c_168_n N_A_27_297#_c_742_n 0.0126377f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_193 N_B1_c_207_p N_A_27_297#_c_742_n 0.00864541f $X=1.555 $Y=1.53 $X2=0 $Y2=0
cc_194 N_B1_c_161_n N_A_27_297#_c_742_n 0.00447207f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_195 N_B1_c_168_n N_A_27_297#_c_746_n 0.0302178f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_196 N_B1_M1036_g N_A_27_297#_c_747_n 0.0102393f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B1_c_168_n N_A_27_297#_c_747_n 0.0314037f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_198 N_B1_c_168_n N_A_27_297#_c_749_n 0.00280049f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_199 N_B1_c_168_n N_A_27_297#_c_750_n 0.012146f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_200 N_B1_c_168_n N_A_27_297#_c_751_n 0.012146f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_201 N_B1_c_168_n N_VPWR_M1024_d 4.58388e-19 $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_202 N_B1_c_207_p N_VPWR_M1024_d 0.00151261f $X=1.555 $Y=1.53 $X2=0 $Y2=0
cc_203 N_B1_c_168_n N_VPWR_M1008_d 0.00170258f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_204 N_B1_c_168_n N_VPWR_M1035_d 0.00169261f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_205 N_B1_M1004_g N_VPWR_c_818_n 0.00274642f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B1_M1007_g N_VPWR_c_818_n 0.00155565f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1024_g N_VPWR_c_819_n 0.00157837f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_M1036_g N_VPWR_c_821_n 0.00302074f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1007_g N_VPWR_c_824_n 0.00585385f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_M1024_g N_VPWR_c_824_n 0.00441875f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1004_g N_VPWR_c_830_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1036_g N_VPWR_c_831_n 0.00441875f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1004_g N_VPWR_c_817_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1007_g N_VPWR_c_817_n 0.0104367f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1024_g N_VPWR_c_817_n 0.00588739f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B1_M1036_g N_VPWR_c_817_n 0.00591459f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B1_c_157_n N_Y_c_962_n 0.0121351f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_168_n N_Y_c_962_n 0.00575485f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_219 N_B1_c_159_n N_Y_c_962_n 0.0255336f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B1_c_160_n N_Y_c_962_n 0.00296008f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_221 N_B1_c_157_n N_Y_c_963_n 0.00164339f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_M1036_g N_Y_c_963_n 2.25871e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B1_c_159_n N_Y_c_963_n 0.0269473f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_224 N_B1_c_160_n N_Y_c_963_n 0.00224632f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_225 N_B1_c_157_n N_Y_c_979_n 8.55715e-19 $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B1_M1036_g N_Y_c_969_n 3.09709e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B1_c_168_n N_Y_c_969_n 0.00951514f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_228 N_B1_c_159_n N_Y_c_969_n 0.00252282f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_229 N_B1_c_157_n N_Y_c_965_n 4.26631e-19 $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B1_c_154_n N_VGND_c_1126_n 0.00338128f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B1_c_161_n N_VGND_c_1126_n 0.0138247f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_232 N_B1_c_155_n N_VGND_c_1127_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B1_c_156_n N_VGND_c_1127_n 0.00268723f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B1_c_157_n N_VGND_c_1128_n 0.00268723f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B1_c_156_n N_VGND_c_1134_n 0.00421816f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B1_c_157_n N_VGND_c_1134_n 0.00421857f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B1_c_154_n N_VGND_c_1146_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B1_c_155_n N_VGND_c_1146_n 0.00423334f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B1_c_154_n N_VGND_c_1148_n 0.0104557f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B1_c_155_n N_VGND_c_1148_n 0.0057163f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B1_c_156_n N_VGND_c_1148_n 0.00575258f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B1_c_157_n N_VGND_c_1148_n 0.00577981f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_243 N_B1_c_154_n N_A_109_47#_c_1287_n 0.00539651f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_B1_c_155_n N_A_109_47#_c_1287_n 0.00630972f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_B1_c_156_n N_A_109_47#_c_1287_n 5.22228e-19 $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_B1_c_155_n N_A_109_47#_c_1284_n 0.00865686f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_B1_c_156_n N_A_109_47#_c_1284_n 0.00870364f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_B1_c_161_n N_A_109_47#_c_1284_n 0.0362443f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_249 N_B1_c_162_n N_A_109_47#_c_1284_n 0.00222133f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B1_c_154_n N_A_109_47#_c_1285_n 0.00299247f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_B1_c_155_n N_A_109_47#_c_1285_n 0.00113286f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_B1_c_161_n N_A_109_47#_c_1285_n 0.0266272f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_253 N_B1_c_162_n N_A_109_47#_c_1285_n 0.00230339f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_c_156_n N_A_109_47#_c_1298_n 0.00255288f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_255 N_B1_c_155_n N_A_109_47#_c_1286_n 4.58193e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_256 N_B1_c_156_n N_A_109_47#_c_1286_n 0.0048497f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B1_c_168_n N_A_109_47#_c_1286_n 0.00186641f $X=3.245 $Y=1.53 $X2=0
+ $Y2=0
cc_258 N_B1_c_161_n N_A_109_47#_c_1286_n 0.0178786f $X=1.385 $Y=1.18 $X2=0 $Y2=0
cc_259 N_B1_c_157_n N_A_109_47#_c_1303_n 0.00302655f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_B2_M1001_g N_A_27_297#_c_742_n 0.0102454f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_261 N_B2_M1008_g N_A_27_297#_c_746_n 0.0102895f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_262 N_B2_M1027_g N_A_27_297#_c_746_n 0.0102895f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_263 N_B2_M1035_g N_A_27_297#_c_747_n 0.0102454f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_264 N_B2_M1001_g N_VPWR_c_819_n 0.00157837f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B2_M1008_g N_VPWR_c_820_n 0.00157837f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_266 N_B2_M1027_g N_VPWR_c_820_n 0.00157837f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_267 N_B2_M1035_g N_VPWR_c_821_n 0.00157837f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_268 N_B2_M1001_g N_VPWR_c_826_n 0.00441875f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B2_M1008_g N_VPWR_c_826_n 0.00441875f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_270 N_B2_M1027_g N_VPWR_c_828_n 0.00441875f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B2_M1035_g N_VPWR_c_828_n 0.00441875f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B2_M1001_g N_VPWR_c_817_n 0.00588739f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B2_M1008_g N_VPWR_c_817_n 0.00586018f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B2_M1027_g N_VPWR_c_817_n 0.00586018f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B2_M1035_g N_VPWR_c_817_n 0.00588739f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B2_c_279_n N_Y_c_961_n 0.00372684f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B2_c_280_n N_Y_c_961_n 0.0109625f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B2_c_281_n N_Y_c_961_n 0.0109625f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B2_c_283_n N_Y_c_961_n 0.0952641f $X=2.91 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B2_c_284_n N_Y_c_961_n 0.00672641f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_281 N_B2_c_282_n N_Y_c_962_n 0.00526882f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B2_c_282_n N_Y_c_965_n 0.00561677f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B2_c_279_n N_VGND_c_1134_n 0.00357877f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B2_c_280_n N_VGND_c_1134_n 0.00357877f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B2_c_281_n N_VGND_c_1134_n 0.00357877f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B2_c_282_n N_VGND_c_1134_n 0.00357877f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B2_c_279_n N_VGND_c_1148_n 0.00525237f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B2_c_280_n N_VGND_c_1148_n 0.00522516f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B2_c_281_n N_VGND_c_1148_n 0.00522516f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B2_c_282_n N_VGND_c_1148_n 0.00525237f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B2_c_279_n N_A_109_47#_c_1303_n 0.0118054f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B2_c_280_n N_A_109_47#_c_1303_n 0.00892725f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_B2_c_281_n N_A_109_47#_c_1303_n 0.00892725f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_B2_c_282_n N_A_109_47#_c_1303_n 0.00914579f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_B2_c_283_n N_A_109_47#_c_1303_n 0.00123352f $X=2.91 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_751_21#_c_349_n N_A1_N_c_559_n 0.00595356f $X=5.64 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_297 N_A_751_21#_c_350_n N_A1_N_c_559_n 0.0101683f $X=6.075 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_298 N_A_751_21#_c_379_p N_A1_N_c_559_n 0.0109565f $X=6.24 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_751_21#_c_357_n N_A1_N_c_559_n 0.00158032f $X=6.24 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_751_21#_c_379_p N_A1_N_c_560_n 0.00630972f $X=6.24 $Y=0.39 $X2=0
+ $Y2=0
cc_301 N_A_751_21#_c_352_n N_A1_N_c_560_n 0.00870364f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_302 N_A_751_21#_c_383_p N_A1_N_c_560_n 5.22228e-19 $X=7.08 $Y=0.39 $X2=0
+ $Y2=0
cc_303 N_A_751_21#_c_357_n N_A1_N_c_560_n 0.00113286f $X=6.24 $Y=0.815 $X2=0
+ $Y2=0
cc_304 N_A_751_21#_c_379_p N_A1_N_c_561_n 5.22228e-19 $X=6.24 $Y=0.39 $X2=0
+ $Y2=0
cc_305 N_A_751_21#_c_352_n N_A1_N_c_561_n 0.00870364f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_306 N_A_751_21#_c_383_p N_A1_N_c_561_n 0.00630972f $X=7.08 $Y=0.39 $X2=0
+ $Y2=0
cc_307 N_A_751_21#_c_358_n N_A1_N_c_561_n 0.00113286f $X=7.08 $Y=0.815 $X2=0
+ $Y2=0
cc_308 N_A_751_21#_c_383_p N_A1_N_c_562_n 0.00630972f $X=7.08 $Y=0.39 $X2=0
+ $Y2=0
cc_309 N_A_751_21#_c_353_n N_A1_N_c_562_n 0.00921556f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_310 N_A_751_21#_c_391_p N_A1_N_c_562_n 5.22228e-19 $X=7.92 $Y=0.39 $X2=0
+ $Y2=0
cc_311 N_A_751_21#_c_358_n N_A1_N_c_562_n 0.00113286f $X=7.08 $Y=0.815 $X2=0
+ $Y2=0
cc_312 N_A_751_21#_c_348_n N_A1_N_c_563_n 0.0131912f $X=5.555 $Y=1.16 $X2=0
+ $Y2=0
cc_313 N_A_751_21#_c_350_n N_A1_N_c_563_n 0.00896514f $X=6.075 $Y=0.82 $X2=0
+ $Y2=0
cc_314 N_A_751_21#_c_352_n N_A1_N_c_563_n 0.036111f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_315 N_A_751_21#_c_353_n N_A1_N_c_563_n 0.00513615f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_316 N_A_751_21#_c_357_n N_A1_N_c_563_n 0.0265405f $X=6.24 $Y=0.815 $X2=0
+ $Y2=0
cc_317 N_A_751_21#_c_358_n N_A1_N_c_563_n 0.0265405f $X=7.08 $Y=0.815 $X2=0
+ $Y2=0
cc_318 N_A_751_21#_c_348_n N_A1_N_c_564_n 0.00125151f $X=5.555 $Y=1.16 $X2=0
+ $Y2=0
cc_319 N_A_751_21#_c_352_n N_A1_N_c_564_n 0.00222133f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_320 N_A_751_21#_c_357_n N_A1_N_c_564_n 0.00230339f $X=6.24 $Y=0.815 $X2=0
+ $Y2=0
cc_321 N_A_751_21#_c_358_n N_A1_N_c_564_n 0.00230339f $X=7.08 $Y=0.815 $X2=0
+ $Y2=0
cc_322 N_A_751_21#_c_383_p N_A2_N_c_641_n 5.22228e-19 $X=7.08 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_323 N_A_751_21#_c_353_n N_A2_N_c_641_n 0.00865686f $X=7.755 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_324 N_A_751_21#_c_391_p N_A2_N_c_641_n 0.00630972f $X=7.92 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_325 N_A_751_21#_c_359_n N_A2_N_c_641_n 0.00113286f $X=7.92 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_326 N_A_751_21#_c_369_n N_A2_N_M1012_g 2.57315e-19 $X=7.92 $Y=1.62 $X2=0
+ $Y2=0
cc_327 N_A_751_21#_c_391_p N_A2_N_c_642_n 0.00630972f $X=7.92 $Y=0.39 $X2=0
+ $Y2=0
cc_328 N_A_751_21#_c_354_n N_A2_N_c_642_n 0.00870364f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_329 N_A_751_21#_c_410_p N_A2_N_c_642_n 5.22228e-19 $X=8.76 $Y=0.39 $X2=0
+ $Y2=0
cc_330 N_A_751_21#_c_359_n N_A2_N_c_642_n 0.00113286f $X=7.92 $Y=0.815 $X2=0
+ $Y2=0
cc_331 N_A_751_21#_c_366_n N_A2_N_M1022_g 0.0109871f $X=8.635 $Y=1.54 $X2=0
+ $Y2=0
cc_332 N_A_751_21#_c_391_p N_A2_N_c_643_n 5.22228e-19 $X=7.92 $Y=0.39 $X2=0
+ $Y2=0
cc_333 N_A_751_21#_c_354_n N_A2_N_c_643_n 0.00870364f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_334 N_A_751_21#_c_410_p N_A2_N_c_643_n 0.00630972f $X=8.76 $Y=0.39 $X2=0
+ $Y2=0
cc_335 N_A_751_21#_c_360_n N_A2_N_c_643_n 0.00113286f $X=8.76 $Y=0.815 $X2=0
+ $Y2=0
cc_336 N_A_751_21#_c_366_n N_A2_N_M1029_g 0.0110013f $X=8.635 $Y=1.54 $X2=0
+ $Y2=0
cc_337 N_A_751_21#_c_410_p N_A2_N_c_644_n 0.0109314f $X=8.76 $Y=0.39 $X2=0 $Y2=0
cc_338 N_A_751_21#_c_355_n N_A2_N_c_644_n 0.0103835f $X=9.215 $Y=0.82 $X2=0
+ $Y2=0
cc_339 N_A_751_21#_c_356_n N_A2_N_c_644_n 0.00696435f $X=9.395 $Y=1.455 $X2=0
+ $Y2=0
cc_340 N_A_751_21#_c_360_n N_A2_N_c_644_n 0.00158032f $X=8.76 $Y=0.815 $X2=0
+ $Y2=0
cc_341 N_A_751_21#_c_367_n N_A2_N_M1037_g 0.0129271f $X=9.215 $Y=1.54 $X2=0
+ $Y2=0
cc_342 N_A_751_21#_c_353_n N_A2_N_c_645_n 0.0113012f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_343 N_A_751_21#_c_366_n N_A2_N_c_645_n 0.0397077f $X=8.635 $Y=1.54 $X2=0
+ $Y2=0
cc_344 N_A_751_21#_c_354_n N_A2_N_c_645_n 0.036111f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_345 N_A_751_21#_c_367_n N_A2_N_c_645_n 0.0104919f $X=9.215 $Y=1.54 $X2=0
+ $Y2=0
cc_346 N_A_751_21#_c_355_n N_A2_N_c_645_n 0.00820272f $X=9.215 $Y=0.82 $X2=0
+ $Y2=0
cc_347 N_A_751_21#_c_356_n N_A2_N_c_645_n 0.0167248f $X=9.395 $Y=1.455 $X2=0
+ $Y2=0
cc_348 N_A_751_21#_c_359_n N_A2_N_c_645_n 0.0265405f $X=7.92 $Y=0.815 $X2=0
+ $Y2=0
cc_349 N_A_751_21#_c_369_n N_A2_N_c_645_n 0.0195077f $X=7.92 $Y=1.62 $X2=0 $Y2=0
cc_350 N_A_751_21#_c_360_n N_A2_N_c_645_n 0.0265405f $X=8.76 $Y=0.815 $X2=0
+ $Y2=0
cc_351 N_A_751_21#_c_370_n N_A2_N_c_645_n 0.0195077f $X=8.76 $Y=1.62 $X2=0 $Y2=0
cc_352 N_A_751_21#_c_366_n N_A2_N_c_646_n 0.00212663f $X=8.635 $Y=1.54 $X2=0
+ $Y2=0
cc_353 N_A_751_21#_c_354_n N_A2_N_c_646_n 0.00222133f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_354 N_A_751_21#_c_356_n N_A2_N_c_646_n 0.00857983f $X=9.395 $Y=1.455 $X2=0
+ $Y2=0
cc_355 N_A_751_21#_c_359_n N_A2_N_c_646_n 0.00230339f $X=7.92 $Y=0.815 $X2=0
+ $Y2=0
cc_356 N_A_751_21#_c_369_n N_A2_N_c_646_n 0.00221143f $X=7.92 $Y=1.62 $X2=0
+ $Y2=0
cc_357 N_A_751_21#_c_360_n N_A2_N_c_646_n 0.00230339f $X=8.76 $Y=0.815 $X2=0
+ $Y2=0
cc_358 N_A_751_21#_c_370_n N_A2_N_c_646_n 0.00221143f $X=8.76 $Y=1.62 $X2=0
+ $Y2=0
cc_359 N_A_751_21#_M1003_g N_A_27_297#_c_756_n 0.0121747f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_360 N_A_751_21#_M1011_g N_A_27_297#_c_756_n 0.0121306f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_361 N_A_751_21#_M1015_g N_A_27_297#_c_758_n 0.0121747f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_362 N_A_751_21#_M1021_g N_A_27_297#_c_758_n 0.0101149f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_363 N_A_751_21#_M1021_g N_A_27_297#_c_725_n 7.12665e-19 $X=5.09 $Y=1.985
+ $X2=0 $Y2=0
cc_364 N_A_751_21#_M1015_g N_A_27_297#_c_726_n 6.55258e-19 $X=4.67 $Y=1.985
+ $X2=0 $Y2=0
cc_365 N_A_751_21#_M1021_g N_A_27_297#_c_726_n 0.011111f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_366 N_A_751_21#_c_348_n N_A_27_297#_c_726_n 0.0236235f $X=5.555 $Y=1.16 $X2=0
+ $Y2=0
cc_367 N_A_751_21#_M1003_g N_VPWR_c_831_n 0.00357877f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_368 N_A_751_21#_M1011_g N_VPWR_c_831_n 0.00357877f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_A_751_21#_M1015_g N_VPWR_c_831_n 0.00357877f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A_751_21#_M1021_g N_VPWR_c_831_n 0.00357835f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_371 N_A_751_21#_M1012_s N_VPWR_c_817_n 0.00216833f $X=7.785 $Y=1.485 $X2=0
+ $Y2=0
cc_372 N_A_751_21#_M1029_s N_VPWR_c_817_n 0.00216833f $X=8.625 $Y=1.485 $X2=0
+ $Y2=0
cc_373 N_A_751_21#_M1003_g N_VPWR_c_817_n 0.00525237f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_374 N_A_751_21#_M1011_g N_VPWR_c_817_n 0.00522516f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_375 N_A_751_21#_M1015_g N_VPWR_c_817_n 0.00522516f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_376 N_A_751_21#_M1021_g N_VPWR_c_817_n 0.0065512f $X=5.09 $Y=1.985 $X2=0
+ $Y2=0
cc_377 N_A_751_21#_c_344_n N_Y_c_963_n 0.00175435f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A_751_21#_M1003_g N_Y_c_963_n 0.00224717f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A_751_21#_c_345_n N_Y_c_963_n 0.00164339f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_751_21#_M1011_g N_Y_c_963_n 0.00165913f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A_751_21#_c_348_n N_Y_c_963_n 0.0127974f $X=5.555 $Y=1.16 $X2=0 $Y2=0
cc_382 N_A_751_21#_c_361_n N_Y_c_963_n 0.0148574f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_751_21#_c_344_n N_Y_c_979_n 0.00631188f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A_751_21#_c_345_n N_Y_c_979_n 0.00612654f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_385 N_A_751_21#_c_346_n N_Y_c_979_n 5.16334e-19 $X=4.67 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A_751_21#_M1011_g N_Y_c_968_n 0.0145761f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_387 N_A_751_21#_M1015_g N_Y_c_968_n 0.0138388f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_388 N_A_751_21#_c_361_n N_Y_c_968_n 0.00222712f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_751_21#_M1003_g N_Y_c_969_n 0.0113424f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_390 N_A_751_21#_c_348_n N_Y_c_969_n 0.0466096f $X=5.555 $Y=1.16 $X2=0 $Y2=0
cc_391 N_A_751_21#_c_361_n N_Y_c_969_n 0.00261044f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_392 N_A_751_21#_c_345_n N_Y_c_964_n 0.00870364f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_393 N_A_751_21#_c_346_n N_Y_c_964_n 0.00983594f $X=4.67 $Y=0.995 $X2=0 $Y2=0
cc_394 N_A_751_21#_c_347_n N_Y_c_964_n 0.00441657f $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_395 N_A_751_21#_c_348_n N_Y_c_964_n 0.0618592f $X=5.555 $Y=1.16 $X2=0 $Y2=0
cc_396 N_A_751_21#_c_351_n N_Y_c_964_n 0.0063267f $X=5.725 $Y=0.82 $X2=0 $Y2=0
cc_397 N_A_751_21#_c_361_n N_Y_c_964_n 0.00452248f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_398 N_A_751_21#_c_345_n N_Y_c_1012_n 5.16334e-19 $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A_751_21#_c_346_n N_Y_c_1012_n 0.00612654f $X=4.67 $Y=0.995 $X2=0 $Y2=0
cc_400 N_A_751_21#_c_347_n N_Y_c_1012_n 0.0107625f $X=5.09 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_751_21#_c_344_n N_Y_c_966_n 0.00782147f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A_751_21#_c_345_n N_Y_c_966_n 0.00113229f $X=4.25 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A_751_21#_c_348_n N_Y_c_966_n 0.00948654f $X=5.555 $Y=1.16 $X2=0 $Y2=0
cc_404 N_A_751_21#_c_361_n N_Y_c_966_n 0.00280293f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_405 N_A_751_21#_M1015_g Y 5.94088e-19 $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_406 N_A_751_21#_M1021_g Y 0.00150511f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_407 N_A_751_21#_c_348_n Y 0.0178184f $X=5.555 $Y=1.16 $X2=0 $Y2=0
cc_408 N_A_751_21#_c_361_n Y 0.0023098f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_409 N_A_751_21#_c_366_n N_A_1139_297#_M1022_d 0.00165831f $X=8.635 $Y=1.54
+ $X2=0 $Y2=0
cc_410 N_A_751_21#_c_367_n N_A_1139_297#_M1037_d 0.00372748f $X=9.215 $Y=1.54
+ $X2=0 $Y2=0
cc_411 N_A_751_21#_M1021_g N_A_1139_297#_c_1060_n 3.89135e-19 $X=5.09 $Y=1.985
+ $X2=0 $Y2=0
cc_412 N_A_751_21#_c_348_n N_A_1139_297#_c_1060_n 0.00552702f $X=5.555 $Y=1.16
+ $X2=0 $Y2=0
cc_413 N_A_751_21#_c_350_n N_A_1139_297#_c_1060_n 0.0081926f $X=6.075 $Y=0.82
+ $X2=0 $Y2=0
cc_414 N_A_751_21#_c_353_n N_A_1139_297#_c_1061_n 0.00148678f $X=7.755 $Y=0.815
+ $X2=0 $Y2=0
cc_415 N_A_751_21#_c_353_n N_A_1139_297#_c_1062_n 0.00824139f $X=7.755 $Y=0.815
+ $X2=0 $Y2=0
cc_416 N_A_751_21#_c_369_n N_A_1139_297#_c_1062_n 0.00271526f $X=7.92 $Y=1.62
+ $X2=0 $Y2=0
cc_417 N_A_751_21#_M1012_s N_A_1139_297#_c_1072_n 0.00312348f $X=7.785 $Y=1.485
+ $X2=0 $Y2=0
cc_418 N_A_751_21#_c_366_n N_A_1139_297#_c_1072_n 0.00320918f $X=8.635 $Y=1.54
+ $X2=0 $Y2=0
cc_419 N_A_751_21#_c_369_n N_A_1139_297#_c_1072_n 0.0118729f $X=7.92 $Y=1.62
+ $X2=0 $Y2=0
cc_420 N_A_751_21#_M1029_s N_A_1139_297#_c_1075_n 0.00312348f $X=8.625 $Y=1.485
+ $X2=0 $Y2=0
cc_421 N_A_751_21#_c_366_n N_A_1139_297#_c_1075_n 0.00320918f $X=8.635 $Y=1.54
+ $X2=0 $Y2=0
cc_422 N_A_751_21#_c_367_n N_A_1139_297#_c_1075_n 0.00320918f $X=9.215 $Y=1.54
+ $X2=0 $Y2=0
cc_423 N_A_751_21#_c_370_n N_A_1139_297#_c_1075_n 0.0118729f $X=8.76 $Y=1.62
+ $X2=0 $Y2=0
cc_424 N_A_751_21#_c_367_n N_A_1139_297#_c_1079_n 0.0176118f $X=9.215 $Y=1.54
+ $X2=0 $Y2=0
cc_425 N_A_751_21#_c_366_n N_A_1139_297#_c_1080_n 0.0126766f $X=8.635 $Y=1.54
+ $X2=0 $Y2=0
cc_426 N_A_751_21#_c_350_n N_VGND_M1039_d 0.00223655f $X=6.075 $Y=0.82 $X2=0
+ $Y2=0
cc_427 N_A_751_21#_c_351_n N_VGND_M1039_d 0.00558189f $X=5.725 $Y=0.82 $X2=0
+ $Y2=0
cc_428 N_A_751_21#_c_352_n N_VGND_M1013_s 0.00162089f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_429 N_A_751_21#_c_353_n N_VGND_M1020_s 0.00162089f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_430 N_A_751_21#_c_354_n N_VGND_M1026_s 0.00162089f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_431 N_A_751_21#_c_355_n N_VGND_M1032_s 0.00321114f $X=9.215 $Y=0.82 $X2=0
+ $Y2=0
cc_432 N_A_751_21#_c_344_n N_VGND_c_1128_n 0.00146448f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_433 N_A_751_21#_c_345_n N_VGND_c_1129_n 0.00146448f $X=4.25 $Y=0.995 $X2=0
+ $Y2=0
cc_434 N_A_751_21#_c_346_n N_VGND_c_1129_n 0.00146339f $X=4.67 $Y=0.995 $X2=0
+ $Y2=0
cc_435 N_A_751_21#_c_352_n N_VGND_c_1130_n 0.0122559f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_436 N_A_751_21#_c_353_n N_VGND_c_1131_n 0.0122559f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_437 N_A_751_21#_c_354_n N_VGND_c_1132_n 0.0122559f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_438 N_A_751_21#_c_355_n N_VGND_c_1133_n 0.0124497f $X=9.215 $Y=0.82 $X2=0
+ $Y2=0
cc_439 N_A_751_21#_c_344_n N_VGND_c_1136_n 0.00424029f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_440 N_A_751_21#_c_345_n N_VGND_c_1136_n 0.00424138f $X=4.25 $Y=0.995 $X2=0
+ $Y2=0
cc_441 N_A_751_21#_c_350_n N_VGND_c_1138_n 0.00193763f $X=6.075 $Y=0.82 $X2=0
+ $Y2=0
cc_442 N_A_751_21#_c_379_p N_VGND_c_1138_n 0.0188551f $X=6.24 $Y=0.39 $X2=0
+ $Y2=0
cc_443 N_A_751_21#_c_352_n N_VGND_c_1138_n 0.00198695f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_444 N_A_751_21#_c_352_n N_VGND_c_1140_n 0.00198695f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_445 N_A_751_21#_c_383_p N_VGND_c_1140_n 0.0188551f $X=7.08 $Y=0.39 $X2=0
+ $Y2=0
cc_446 N_A_751_21#_c_353_n N_VGND_c_1140_n 0.00198695f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_447 N_A_751_21#_c_353_n N_VGND_c_1142_n 0.00198695f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_448 N_A_751_21#_c_391_p N_VGND_c_1142_n 0.0188551f $X=7.92 $Y=0.39 $X2=0
+ $Y2=0
cc_449 N_A_751_21#_c_354_n N_VGND_c_1142_n 0.00198695f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_450 N_A_751_21#_c_354_n N_VGND_c_1144_n 0.00198695f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_451 N_A_751_21#_c_410_p N_VGND_c_1144_n 0.0188551f $X=8.76 $Y=0.39 $X2=0
+ $Y2=0
cc_452 N_A_751_21#_c_355_n N_VGND_c_1144_n 0.00193763f $X=9.215 $Y=0.82 $X2=0
+ $Y2=0
cc_453 N_A_751_21#_c_355_n N_VGND_c_1147_n 0.00513476f $X=9.215 $Y=0.82 $X2=0
+ $Y2=0
cc_454 N_A_751_21#_M1010_d N_VGND_c_1148_n 0.00215201f $X=6.105 $Y=0.235 $X2=0
+ $Y2=0
cc_455 N_A_751_21#_M1016_d N_VGND_c_1148_n 0.00215201f $X=6.945 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_A_751_21#_M1017_d N_VGND_c_1148_n 0.00215201f $X=7.785 $Y=0.235 $X2=0
+ $Y2=0
cc_457 N_A_751_21#_M1031_d N_VGND_c_1148_n 0.00215201f $X=8.625 $Y=0.235 $X2=0
+ $Y2=0
cc_458 N_A_751_21#_c_344_n N_VGND_c_1148_n 0.0057425f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_A_751_21#_c_345_n N_VGND_c_1148_n 0.00571728f $X=4.25 $Y=0.995 $X2=0
+ $Y2=0
cc_460 N_A_751_21#_c_346_n N_VGND_c_1148_n 0.00571728f $X=4.67 $Y=0.995 $X2=0
+ $Y2=0
cc_461 N_A_751_21#_c_347_n N_VGND_c_1148_n 0.0108261f $X=5.09 $Y=0.995 $X2=0
+ $Y2=0
cc_462 N_A_751_21#_c_350_n N_VGND_c_1148_n 0.0044874f $X=6.075 $Y=0.82 $X2=0
+ $Y2=0
cc_463 N_A_751_21#_c_351_n N_VGND_c_1148_n 7.23891e-19 $X=5.725 $Y=0.82 $X2=0
+ $Y2=0
cc_464 N_A_751_21#_c_379_p N_VGND_c_1148_n 0.0122069f $X=6.24 $Y=0.39 $X2=0
+ $Y2=0
cc_465 N_A_751_21#_c_352_n N_VGND_c_1148_n 0.00835832f $X=6.915 $Y=0.815 $X2=0
+ $Y2=0
cc_466 N_A_751_21#_c_383_p N_VGND_c_1148_n 0.0122069f $X=7.08 $Y=0.39 $X2=0
+ $Y2=0
cc_467 N_A_751_21#_c_353_n N_VGND_c_1148_n 0.00835832f $X=7.755 $Y=0.815 $X2=0
+ $Y2=0
cc_468 N_A_751_21#_c_391_p N_VGND_c_1148_n 0.0122069f $X=7.92 $Y=0.39 $X2=0
+ $Y2=0
cc_469 N_A_751_21#_c_354_n N_VGND_c_1148_n 0.00835832f $X=8.595 $Y=0.815 $X2=0
+ $Y2=0
cc_470 N_A_751_21#_c_410_p N_VGND_c_1148_n 0.0122069f $X=8.76 $Y=0.39 $X2=0
+ $Y2=0
cc_471 N_A_751_21#_c_355_n N_VGND_c_1148_n 0.0131896f $X=9.215 $Y=0.82 $X2=0
+ $Y2=0
cc_472 N_A_751_21#_c_346_n N_VGND_c_1150_n 0.00424138f $X=4.67 $Y=0.995 $X2=0
+ $Y2=0
cc_473 N_A_751_21#_c_347_n N_VGND_c_1150_n 0.00542163f $X=5.09 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_751_21#_c_347_n N_VGND_c_1151_n 0.00335921f $X=5.09 $Y=0.995 $X2=0
+ $Y2=0
cc_475 N_A_751_21#_c_348_n N_VGND_c_1151_n 0.0123169f $X=5.555 $Y=1.16 $X2=0
+ $Y2=0
cc_476 N_A_751_21#_c_350_n N_VGND_c_1151_n 0.0128272f $X=6.075 $Y=0.82 $X2=0
+ $Y2=0
cc_477 N_A_751_21#_c_351_n N_VGND_c_1151_n 0.0136696f $X=5.725 $Y=0.82 $X2=0
+ $Y2=0
cc_478 N_A1_N_c_562_n N_A2_N_c_641_n 0.0197107f $X=7.29 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_479 N_A1_N_M1028_g N_A2_N_M1012_g 0.0197107f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_480 N_A1_N_c_563_n N_A2_N_c_645_n 0.0122976f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_481 N_A1_N_c_564_n N_A2_N_c_645_n 0.00164744f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_482 N_A1_N_c_563_n N_A2_N_c_646_n 2.18547e-19 $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_483 N_A1_N_c_564_n N_A2_N_c_646_n 0.0197107f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_484 N_A1_N_M1002_g N_A_27_297#_c_726_n 0.00138578f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_A1_N_M1002_g N_VPWR_c_822_n 0.00274642f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_486 N_A1_N_M1005_g N_VPWR_c_822_n 0.00155565f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_487 N_A1_N_M1009_g N_VPWR_c_823_n 0.00157837f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_488 N_A1_N_M1028_g N_VPWR_c_823_n 0.00302074f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_489 N_A1_N_M1002_g N_VPWR_c_831_n 0.00541359f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_490 N_A1_N_M1005_g N_VPWR_c_832_n 0.00585385f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_491 N_A1_N_M1009_g N_VPWR_c_832_n 0.00585385f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_492 N_A1_N_M1028_g N_VPWR_c_833_n 0.00585385f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_493 N_A1_N_M1002_g N_VPWR_c_817_n 0.0108276f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_494 N_A1_N_M1005_g N_VPWR_c_817_n 0.0104367f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_495 N_A1_N_M1009_g N_VPWR_c_817_n 0.0104367f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_496 N_A1_N_M1028_g N_VPWR_c_817_n 0.010464f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_497 N_A1_N_M1002_g N_A_1139_297#_c_1058_n 0.0102929f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_498 N_A1_N_M1005_g N_A_1139_297#_c_1058_n 6.41022e-19 $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A1_N_M1002_g N_A_1139_297#_c_1059_n 0.0107675f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_500 N_A1_N_M1005_g N_A_1139_297#_c_1059_n 0.0133328f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_501 N_A1_N_c_563_n N_A_1139_297#_c_1059_n 0.0373978f $X=7.155 $Y=1.16 $X2=0
+ $Y2=0
cc_502 N_A1_N_c_564_n N_A_1139_297#_c_1059_n 0.00212663f $X=7.29 $Y=1.16 $X2=0
+ $Y2=0
cc_503 N_A1_N_M1002_g N_A_1139_297#_c_1060_n 0.00149869f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_504 N_A1_N_c_563_n N_A_1139_297#_c_1060_n 0.00302711f $X=7.155 $Y=1.16 $X2=0
+ $Y2=0
cc_505 N_A1_N_M1009_g N_A_1139_297#_c_1061_n 0.0132886f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_506 N_A1_N_M1028_g N_A_1139_297#_c_1061_n 0.0138132f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_507 N_A1_N_c_563_n N_A_1139_297#_c_1061_n 0.0364467f $X=7.155 $Y=1.16 $X2=0
+ $Y2=0
cc_508 N_A1_N_c_564_n N_A_1139_297#_c_1061_n 0.00212663f $X=7.29 $Y=1.16 $X2=0
+ $Y2=0
cc_509 N_A1_N_c_563_n N_A_1139_297#_c_1063_n 0.018751f $X=7.155 $Y=1.16 $X2=0
+ $Y2=0
cc_510 N_A1_N_c_564_n N_A_1139_297#_c_1063_n 0.00221654f $X=7.29 $Y=1.16 $X2=0
+ $Y2=0
cc_511 N_A1_N_c_560_n N_VGND_c_1130_n 0.00146339f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_512 N_A1_N_c_561_n N_VGND_c_1130_n 0.00146448f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_513 N_A1_N_c_562_n N_VGND_c_1131_n 0.00146448f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_514 N_A1_N_c_559_n N_VGND_c_1138_n 0.00424416f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_515 N_A1_N_c_560_n N_VGND_c_1138_n 0.00423334f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_516 N_A1_N_c_561_n N_VGND_c_1140_n 0.00423334f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_517 N_A1_N_c_562_n N_VGND_c_1140_n 0.00423334f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_518 N_A1_N_c_559_n N_VGND_c_1148_n 0.00705967f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_519 N_A1_N_c_560_n N_VGND_c_1148_n 0.0057163f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_520 N_A1_N_c_561_n N_VGND_c_1148_n 0.0057163f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_521 N_A1_N_c_562_n N_VGND_c_1148_n 0.0057435f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_522 N_A1_N_c_559_n N_VGND_c_1151_n 0.00335921f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_523 N_A2_N_M1012_g N_VPWR_c_833_n 0.00357877f $X=7.71 $Y=1.985 $X2=0 $Y2=0
cc_524 N_A2_N_M1022_g N_VPWR_c_833_n 0.00357877f $X=8.13 $Y=1.985 $X2=0 $Y2=0
cc_525 N_A2_N_M1029_g N_VPWR_c_833_n 0.00357877f $X=8.55 $Y=1.985 $X2=0 $Y2=0
cc_526 N_A2_N_M1037_g N_VPWR_c_833_n 0.00357877f $X=8.97 $Y=1.985 $X2=0 $Y2=0
cc_527 N_A2_N_M1012_g N_VPWR_c_817_n 0.00525237f $X=7.71 $Y=1.985 $X2=0 $Y2=0
cc_528 N_A2_N_M1022_g N_VPWR_c_817_n 0.00522516f $X=8.13 $Y=1.985 $X2=0 $Y2=0
cc_529 N_A2_N_M1029_g N_VPWR_c_817_n 0.00522516f $X=8.55 $Y=1.985 $X2=0 $Y2=0
cc_530 N_A2_N_M1037_g N_VPWR_c_817_n 0.00633386f $X=8.97 $Y=1.985 $X2=0 $Y2=0
cc_531 N_A2_N_M1012_g N_A_1139_297#_c_1062_n 2.57315e-19 $X=7.71 $Y=1.985 $X2=0
+ $Y2=0
cc_532 N_A2_N_c_645_n N_A_1139_297#_c_1062_n 0.0024604f $X=8.855 $Y=1.16 $X2=0
+ $Y2=0
cc_533 N_A2_N_M1012_g N_A_1139_297#_c_1072_n 0.0121747f $X=7.71 $Y=1.985 $X2=0
+ $Y2=0
cc_534 N_A2_N_M1022_g N_A_1139_297#_c_1072_n 0.00984328f $X=8.13 $Y=1.985 $X2=0
+ $Y2=0
cc_535 N_A2_N_M1029_g N_A_1139_297#_c_1075_n 0.00984328f $X=8.55 $Y=1.985 $X2=0
+ $Y2=0
cc_536 N_A2_N_M1037_g N_A_1139_297#_c_1075_n 0.00988743f $X=8.97 $Y=1.985 $X2=0
+ $Y2=0
cc_537 N_A2_N_c_641_n N_VGND_c_1131_n 0.00146448f $X=7.71 $Y=0.995 $X2=0 $Y2=0
cc_538 N_A2_N_c_642_n N_VGND_c_1132_n 0.00146448f $X=8.13 $Y=0.995 $X2=0 $Y2=0
cc_539 N_A2_N_c_643_n N_VGND_c_1132_n 0.00146448f $X=8.55 $Y=0.995 $X2=0 $Y2=0
cc_540 N_A2_N_c_644_n N_VGND_c_1133_n 0.00316354f $X=8.97 $Y=0.995 $X2=0 $Y2=0
cc_541 N_A2_N_c_641_n N_VGND_c_1142_n 0.00423334f $X=7.71 $Y=0.995 $X2=0 $Y2=0
cc_542 N_A2_N_c_642_n N_VGND_c_1142_n 0.00423334f $X=8.13 $Y=0.995 $X2=0 $Y2=0
cc_543 N_A2_N_c_643_n N_VGND_c_1144_n 0.00423334f $X=8.55 $Y=0.995 $X2=0 $Y2=0
cc_544 N_A2_N_c_644_n N_VGND_c_1144_n 0.00424416f $X=8.97 $Y=0.995 $X2=0 $Y2=0
cc_545 N_A2_N_c_641_n N_VGND_c_1148_n 0.0057435f $X=7.71 $Y=0.995 $X2=0 $Y2=0
cc_546 N_A2_N_c_642_n N_VGND_c_1148_n 0.0057163f $X=8.13 $Y=0.995 $X2=0 $Y2=0
cc_547 N_A2_N_c_643_n N_VGND_c_1148_n 0.0057163f $X=8.55 $Y=0.995 $X2=0 $Y2=0
cc_548 N_A2_N_c_644_n N_VGND_c_1148_n 0.00684476f $X=8.97 $Y=0.995 $X2=0 $Y2=0
cc_549 N_A_27_297#_c_722_n N_VPWR_M1004_d 0.00165831f $X=0.975 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_550 N_A_27_297#_c_742_n N_VPWR_M1024_d 0.00332352f $X=1.815 $Y=1.88 $X2=0
+ $Y2=0
cc_551 N_A_27_297#_c_746_n N_VPWR_M1008_d 0.00320726f $X=2.655 $Y=1.88 $X2=0
+ $Y2=0
cc_552 N_A_27_297#_c_747_n N_VPWR_M1035_d 0.00329291f $X=3.495 $Y=1.88 $X2=0
+ $Y2=0
cc_553 N_A_27_297#_c_722_n N_VPWR_c_818_n 0.0126919f $X=0.975 $Y=1.54 $X2=0
+ $Y2=0
cc_554 N_A_27_297#_c_742_n N_VPWR_c_819_n 0.0123012f $X=1.815 $Y=1.88 $X2=0
+ $Y2=0
cc_555 N_A_27_297#_c_746_n N_VPWR_c_820_n 0.0123012f $X=2.655 $Y=1.88 $X2=0
+ $Y2=0
cc_556 N_A_27_297#_c_747_n N_VPWR_c_821_n 0.0123012f $X=3.495 $Y=1.88 $X2=0
+ $Y2=0
cc_557 N_A_27_297#_c_742_n N_VPWR_c_824_n 0.00208769f $X=1.815 $Y=1.88 $X2=0
+ $Y2=0
cc_558 N_A_27_297#_c_774_p N_VPWR_c_824_n 0.0138795f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_559 N_A_27_297#_c_742_n N_VPWR_c_826_n 0.00201582f $X=1.815 $Y=1.88 $X2=0
+ $Y2=0
cc_560 N_A_27_297#_c_746_n N_VPWR_c_826_n 0.00201582f $X=2.655 $Y=1.88 $X2=0
+ $Y2=0
cc_561 N_A_27_297#_c_750_n N_VPWR_c_826_n 0.0142224f $X=1.94 $Y=1.96 $X2=0 $Y2=0
cc_562 N_A_27_297#_c_746_n N_VPWR_c_828_n 0.00201582f $X=2.655 $Y=1.88 $X2=0
+ $Y2=0
cc_563 N_A_27_297#_c_747_n N_VPWR_c_828_n 0.00201582f $X=3.495 $Y=1.88 $X2=0
+ $Y2=0
cc_564 N_A_27_297#_c_751_n N_VPWR_c_828_n 0.0142224f $X=2.78 $Y=1.96 $X2=0 $Y2=0
cc_565 N_A_27_297#_c_721_n N_VPWR_c_830_n 0.0217551f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_566 N_A_27_297#_c_747_n N_VPWR_c_831_n 0.00201582f $X=3.495 $Y=1.88 $X2=0
+ $Y2=0
cc_567 N_A_27_297#_c_756_n N_VPWR_c_831_n 0.0330174f $X=4.335 $Y=2.38 $X2=0
+ $Y2=0
cc_568 N_A_27_297#_c_784_p N_VPWR_c_831_n 0.0142933f $X=3.745 $Y=2.38 $X2=0
+ $Y2=0
cc_569 N_A_27_297#_c_758_n N_VPWR_c_831_n 0.031172f $X=5.135 $Y=2.38 $X2=0 $Y2=0
cc_570 N_A_27_297#_c_725_n N_VPWR_c_831_n 0.021178f $X=5.3 $Y=2.295 $X2=0 $Y2=0
cc_571 N_A_27_297#_c_787_p N_VPWR_c_831_n 0.0139385f $X=4.455 $Y=2.38 $X2=0
+ $Y2=0
cc_572 N_A_27_297#_M1004_s N_VPWR_c_817_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_573 N_A_27_297#_M1007_s N_VPWR_c_817_n 0.00259411f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_574 N_A_27_297#_M1001_s N_VPWR_c_817_n 0.0022335f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_575 N_A_27_297#_M1027_s N_VPWR_c_817_n 0.0022335f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_576 N_A_27_297#_M1036_s N_VPWR_c_817_n 0.00220079f $X=3.485 $Y=1.485 $X2=0
+ $Y2=0
cc_577 N_A_27_297#_M1011_d N_VPWR_c_817_n 0.00215204f $X=4.325 $Y=1.485 $X2=0
+ $Y2=0
cc_578 N_A_27_297#_M1021_d N_VPWR_c_817_n 0.00209319f $X=5.165 $Y=1.485 $X2=0
+ $Y2=0
cc_579 N_A_27_297#_c_721_n N_VPWR_c_817_n 0.0128119f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_580 N_A_27_297#_c_742_n N_VPWR_c_817_n 0.00825891f $X=1.815 $Y=1.88 $X2=0
+ $Y2=0
cc_581 N_A_27_297#_c_746_n N_VPWR_c_817_n 0.00800071f $X=2.655 $Y=1.88 $X2=0
+ $Y2=0
cc_582 N_A_27_297#_c_747_n N_VPWR_c_817_n 0.00800071f $X=3.495 $Y=1.88 $X2=0
+ $Y2=0
cc_583 N_A_27_297#_c_756_n N_VPWR_c_817_n 0.0204627f $X=4.335 $Y=2.38 $X2=0
+ $Y2=0
cc_584 N_A_27_297#_c_784_p N_VPWR_c_817_n 0.00962418f $X=3.745 $Y=2.38 $X2=0
+ $Y2=0
cc_585 N_A_27_297#_c_758_n N_VPWR_c_817_n 0.0195523f $X=5.135 $Y=2.38 $X2=0
+ $Y2=0
cc_586 N_A_27_297#_c_725_n N_VPWR_c_817_n 0.0124992f $X=5.3 $Y=2.295 $X2=0 $Y2=0
cc_587 N_A_27_297#_c_774_p N_VPWR_c_817_n 0.0091658f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_588 N_A_27_297#_c_750_n N_VPWR_c_817_n 0.00954719f $X=1.94 $Y=1.96 $X2=0
+ $Y2=0
cc_589 N_A_27_297#_c_751_n N_VPWR_c_817_n 0.00954719f $X=2.78 $Y=1.96 $X2=0
+ $Y2=0
cc_590 N_A_27_297#_c_787_p N_VPWR_c_817_n 0.00923924f $X=4.455 $Y=2.38 $X2=0
+ $Y2=0
cc_591 N_A_27_297#_c_756_n N_Y_M1003_s 0.00312348f $X=4.335 $Y=2.38 $X2=0 $Y2=0
cc_592 N_A_27_297#_c_758_n N_Y_M1015_s 0.00312348f $X=5.135 $Y=2.38 $X2=0 $Y2=0
cc_593 N_A_27_297#_c_756_n N_Y_c_1025_n 0.0116277f $X=4.335 $Y=2.38 $X2=0 $Y2=0
cc_594 N_A_27_297#_M1011_d N_Y_c_968_n 0.00170714f $X=4.325 $Y=1.485 $X2=0 $Y2=0
cc_595 N_A_27_297#_c_811_p N_Y_c_968_n 0.0122805f $X=4.46 $Y=1.96 $X2=0 $Y2=0
cc_596 N_A_27_297#_c_726_n Y 0.00738407f $X=5.3 $Y=1.65 $X2=0 $Y2=0
cc_597 N_A_27_297#_c_758_n N_Y_c_1029_n 0.0119263f $X=5.135 $Y=2.38 $X2=0 $Y2=0
cc_598 N_A_27_297#_c_725_n N_A_1139_297#_c_1058_n 0.0139f $X=5.3 $Y=2.295 $X2=0
+ $Y2=0
cc_599 N_A_27_297#_c_726_n N_A_1139_297#_c_1058_n 0.0515145f $X=5.3 $Y=1.65
+ $X2=0 $Y2=0
cc_600 N_A_27_297#_c_726_n N_A_1139_297#_c_1060_n 0.0139f $X=5.3 $Y=1.65 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_817_n N_Y_M1003_s 0.00216833f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_602 N_VPWR_c_817_n N_Y_M1015_s 0.0021603f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_603 N_VPWR_c_817_n N_A_1139_297#_M1002_s 0.00209319f $X=9.43 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_604 N_VPWR_c_817_n N_A_1139_297#_M1005_s 0.00319348f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_605 N_VPWR_c_817_n N_A_1139_297#_M1028_s 0.00246446f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_606 N_VPWR_c_817_n N_A_1139_297#_M1022_d 0.00215203f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_607 N_VPWR_c_817_n N_A_1139_297#_M1037_d 0.0027779f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_608 N_VPWR_c_831_n N_A_1139_297#_c_1058_n 0.0210382f $X=6.155 $Y=2.72 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_817_n N_A_1139_297#_c_1058_n 0.0124268f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_610 N_VPWR_M1002_d N_A_1139_297#_c_1059_n 0.00165831f $X=6.105 $Y=1.485 $X2=0
+ $Y2=0
cc_611 N_VPWR_c_822_n N_A_1139_297#_c_1059_n 0.0126919f $X=6.24 $Y=1.96 $X2=0
+ $Y2=0
cc_612 N_VPWR_c_832_n N_A_1139_297#_c_1113_n 0.0138795f $X=6.955 $Y=2.72 $X2=0
+ $Y2=0
cc_613 N_VPWR_c_817_n N_A_1139_297#_c_1113_n 0.0091658f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_614 N_VPWR_M1009_d N_A_1139_297#_c_1061_n 0.00165831f $X=6.945 $Y=1.485 $X2=0
+ $Y2=0
cc_615 N_VPWR_c_823_n N_A_1139_297#_c_1061_n 0.0126919f $X=7.08 $Y=1.96 $X2=0
+ $Y2=0
cc_616 N_VPWR_c_833_n N_A_1139_297#_c_1117_n 0.0143053f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_617 N_VPWR_c_817_n N_A_1139_297#_c_1117_n 0.00962794f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_618 N_VPWR_c_833_n N_A_1139_297#_c_1072_n 0.0330174f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_619 N_VPWR_c_817_n N_A_1139_297#_c_1072_n 0.0204627f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_620 N_VPWR_c_833_n N_A_1139_297#_c_1075_n 0.0492948f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_621 N_VPWR_c_817_n N_A_1139_297#_c_1075_n 0.0302732f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_622 N_VPWR_c_833_n N_A_1139_297#_c_1080_n 0.0142933f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_623 N_VPWR_c_817_n N_A_1139_297#_c_1080_n 0.00962421f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_624 N_Y_c_962_n N_VGND_M1038_d 0.00162089f $X=3.745 $Y=0.815 $X2=0 $Y2=0
cc_625 N_Y_c_964_n N_VGND_M1006_d 0.00162089f $X=4.715 $Y=0.815 $X2=0 $Y2=0
cc_626 N_Y_c_962_n N_VGND_c_1128_n 0.0122559f $X=3.745 $Y=0.815 $X2=0 $Y2=0
cc_627 N_Y_c_964_n N_VGND_c_1129_n 0.0122559f $X=4.715 $Y=0.815 $X2=0 $Y2=0
cc_628 N_Y_c_962_n N_VGND_c_1134_n 0.00199263f $X=3.745 $Y=0.815 $X2=0 $Y2=0
cc_629 N_Y_c_979_n N_VGND_c_1136_n 0.0167138f $X=4.04 $Y=0.39 $X2=0 $Y2=0
cc_630 N_Y_c_964_n N_VGND_c_1136_n 0.00198695f $X=4.715 $Y=0.815 $X2=0 $Y2=0
cc_631 N_Y_c_966_n N_VGND_c_1136_n 0.00185026f $X=3.975 $Y=0.815 $X2=0 $Y2=0
cc_632 N_Y_M1018_d N_VGND_c_1148_n 0.00216833f $X=1.805 $Y=0.235 $X2=0 $Y2=0
cc_633 N_Y_M1025_d N_VGND_c_1148_n 0.00216833f $X=2.645 $Y=0.235 $X2=0 $Y2=0
cc_634 N_Y_M1000_s N_VGND_c_1148_n 0.00216035f $X=3.905 $Y=0.235 $X2=0 $Y2=0
cc_635 N_Y_M1030_s N_VGND_c_1148_n 0.00216035f $X=4.745 $Y=0.235 $X2=0 $Y2=0
cc_636 N_Y_c_962_n N_VGND_c_1148_n 0.00640255f $X=3.745 $Y=0.815 $X2=0 $Y2=0
cc_637 N_Y_c_979_n N_VGND_c_1148_n 0.0120751f $X=4.04 $Y=0.39 $X2=0 $Y2=0
cc_638 N_Y_c_964_n N_VGND_c_1148_n 0.00835832f $X=4.715 $Y=0.815 $X2=0 $Y2=0
cc_639 N_Y_c_1012_n N_VGND_c_1148_n 0.0120721f $X=4.88 $Y=0.39 $X2=0 $Y2=0
cc_640 N_Y_c_966_n N_VGND_c_1148_n 0.00300741f $X=3.975 $Y=0.815 $X2=0 $Y2=0
cc_641 N_Y_c_964_n N_VGND_c_1150_n 0.00198695f $X=4.715 $Y=0.815 $X2=0 $Y2=0
cc_642 N_Y_c_1012_n N_VGND_c_1150_n 0.0167046f $X=4.88 $Y=0.39 $X2=0 $Y2=0
cc_643 N_Y_c_961_n N_A_109_47#_M1019_s 0.00162317f $X=2.865 $Y=0.775 $X2=0 $Y2=0
cc_644 N_Y_c_962_n N_A_109_47#_M1033_s 0.00191752f $X=3.745 $Y=0.815 $X2=0 $Y2=0
cc_645 N_Y_c_961_n N_A_109_47#_c_1286_n 0.00841895f $X=2.865 $Y=0.775 $X2=0
+ $Y2=0
cc_646 N_Y_M1018_d N_A_109_47#_c_1303_n 0.00305026f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_647 N_Y_M1025_d N_A_109_47#_c_1303_n 0.00305026f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_648 N_Y_c_961_n N_A_109_47#_c_1303_n 0.0616167f $X=2.865 $Y=0.775 $X2=0 $Y2=0
cc_649 N_Y_c_962_n N_A_109_47#_c_1303_n 0.0126031f $X=3.745 $Y=0.815 $X2=0 $Y2=0
cc_650 N_VGND_c_1148_n N_A_109_47#_M1014_s 0.00215201f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_651 N_VGND_c_1148_n N_A_109_47#_M1034_s 0.00215206f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_c_1148_n N_A_109_47#_M1019_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_653 N_VGND_c_1148_n N_A_109_47#_M1033_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_654 N_VGND_c_1146_n N_A_109_47#_c_1287_n 0.0188551f $X=1.015 $Y=0 $X2=0 $Y2=0
cc_655 N_VGND_c_1148_n N_A_109_47#_c_1287_n 0.0122069f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_656 N_VGND_M1023_d N_A_109_47#_c_1284_n 0.00162089f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_657 N_VGND_c_1127_n N_A_109_47#_c_1284_n 0.0122559f $X=1.1 $Y=0.39 $X2=0
+ $Y2=0
cc_658 N_VGND_c_1134_n N_A_109_47#_c_1284_n 0.00198695f $X=3.535 $Y=0 $X2=0
+ $Y2=0
cc_659 N_VGND_c_1146_n N_A_109_47#_c_1284_n 0.00198695f $X=1.015 $Y=0 $X2=0
+ $Y2=0
cc_660 N_VGND_c_1148_n N_A_109_47#_c_1284_n 0.00835832f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_661 N_VGND_c_1126_n N_A_109_47#_c_1285_n 0.00750114f $X=0.26 $Y=0.39 $X2=0
+ $Y2=0
cc_662 N_VGND_c_1134_n N_A_109_47#_c_1298_n 0.0152108f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_663 N_VGND_c_1148_n N_A_109_47#_c_1298_n 0.00940698f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_664 N_VGND_c_1134_n N_A_109_47#_c_1303_n 0.0973818f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1148_n N_A_109_47#_c_1303_n 0.0626919f $X=9.43 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a2bb2oi_1.pex.spice
* Created: Tue Sep  1 18:54:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%A1_N 3 6 8 9 13 14 15
r27 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=1.325
r28 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=0.995
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r30 8 9 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.335 $Y=1.19 $X2=0.335
+ $Y2=1.53
r31 8 14 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=0.335 $Y=1.19
+ $X2=0.335 $Y2=1.16
r32 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r33 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%A2_N 3 5 7 8 11 17
r34 12 17 11.307 $w=2.63e-07 $l=2.6e-07 $layer=LI1_cond $X=0.89 $Y=1.142
+ $X2=1.15 $Y2=1.142
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=1.325
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r37 8 17 0.217442 $w=2.63e-07 $l=5e-09 $layer=LI1_cond $X=1.155 $Y=1.142
+ $X2=1.15 $Y2=1.142
r38 5 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r39 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
r40 3 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.83 $Y=1.985
+ $X2=0.83 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%A_109_47# 1 2 7 9 12 14 15 16 19 20 23 27
+ 28 32
r70 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r71 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.495 $Y=1.445
+ $X2=1.495 $Y2=1.16
r72 29 32 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.495 $Y=0.83
+ $X2=1.495 $Y2=1.16
r73 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.41 $Y=1.53
+ $X2=1.495 $Y2=1.445
r74 27 28 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.41 $Y=1.53
+ $X2=1.205 $Y2=1.53
r75 23 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.04 $Y=1.64
+ $X2=1.04 $Y2=2.32
r76 21 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.04 $Y=1.615
+ $X2=1.205 $Y2=1.53
r77 21 23 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.04 $Y=1.615
+ $X2=1.04 $Y2=1.64
r78 19 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.41 $Y=0.745
+ $X2=1.495 $Y2=0.83
r79 19 20 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.41 $Y=0.745
+ $X2=0.765 $Y2=0.745
r80 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=0.66
+ $X2=0.765 $Y2=0.745
r81 16 18 7.17647 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.68 $Y=0.66 $X2=0.68
+ $Y2=0.56
r82 14 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.835 $Y=1.16
+ $X2=1.495 $Y2=1.16
r83 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.835 $Y=1.16
+ $X2=1.91 $Y2=1.16
r84 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.325
+ $X2=1.91 $Y2=1.16
r85 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.91 $Y=1.325
+ $X2=1.91 $Y2=1.985
r86 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=0.995
+ $X2=1.91 $Y2=1.16
r87 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.91 $Y=0.995 $X2=1.91
+ $Y2=0.56
r88 2 25 400 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.485 $X2=1.04 $Y2=2.32
r89 2 23 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.485 $X2=1.04 $Y2=1.64
r90 1 18 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%B2 1 3 6 8 9 10 11 18 28
c46 18 0 1.50675e-19 $X=2.33 $Y=1.16
c47 6 0 1.60266e-19 $X=2.33 $Y=1.985
r48 26 28 0.410459 $w=3.63e-07 $l=1.3e-08 $layer=LI1_cond $X=2.427 $Y=1.177
+ $X2=2.427 $Y2=1.19
r49 19 26 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=2.427 $Y=1.16
+ $X2=2.427 $Y2=1.177
r50 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.16 $X2=2.33 $Y2=1.16
r51 10 19 0.599902 $w=3.63e-07 $l=1.9e-08 $layer=LI1_cond $X=2.427 $Y=1.141
+ $X2=2.427 $Y2=1.16
r52 10 34 7.9244 $w=3.63e-07 $l=1.46e-07 $layer=LI1_cond $X=2.427 $Y=1.141
+ $X2=2.427 $Y2=0.995
r53 10 11 9.59843 $w=3.63e-07 $l=3.04e-07 $layer=LI1_cond $X=2.427 $Y=1.226
+ $X2=2.427 $Y2=1.53
r54 10 28 1.13666 $w=3.63e-07 $l=3.6e-08 $layer=LI1_cond $X=2.427 $Y=1.226
+ $X2=2.427 $Y2=1.19
r55 9 34 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.525 $Y=0.85
+ $X2=2.525 $Y2=0.995
r56 8 9 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.525 $Y=0.51
+ $X2=2.525 $Y2=0.85
r57 4 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.325
+ $X2=2.33 $Y2=1.16
r58 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.33 $Y=1.325 $X2=2.33
+ $Y2=1.985
r59 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=0.995
+ $X2=2.33 $Y2=1.16
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.33 $Y=0.995 $X2=2.33
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%B1 3 6 8 11 13
r29 11 14 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.837 $Y=1.16
+ $X2=2.837 $Y2=1.325
r30 11 13 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.837 $Y=1.16
+ $X2=2.837 $Y2=0.995
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.16 $X2=2.865 $Y2=1.16
r32 8 12 2.31499 $w=6.18e-07 $l=1.2e-07 $layer=LI1_cond $X=2.985 $Y=1.305
+ $X2=2.865 $Y2=1.305
r33 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.75 $Y=1.985
+ $X2=2.75 $Y2=1.325
r34 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.56 $X2=2.75
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%VPWR 1 2 9 11 14 16 23 24 32 35
r43 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 24 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 21 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.58 $Y2=2.72
r47 21 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 20 33 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 19 20 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 16 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=2.58 $Y2=2.72
r52 16 19 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 14 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 11 35 16.8131 $w=4.98e-07 $l=6.45e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=1.99
r55 11 17 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.212 $Y=2.72
+ $X2=0.425 $Y2=2.72
r56 11 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 7 32 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.635
+ $X2=2.58 $Y2=2.72
r58 7 9 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.58 $Y=2.635
+ $X2=2.58 $Y2=2.36
r59 2 9 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.485 $X2=2.54 $Y2=2.36
r60 1 35 300 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%Y 1 2 8 9 10 11
c33 10 0 1.60266e-19 $X=1.605 $Y=2.21
r34 11 25 12.805 $w=4.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.99 $Y=0.51
+ $X2=1.99 $Y2=0.825
r35 10 18 6.9284 $w=4.05e-07 $l=2.3e-07 $layer=LI1_cond $X=1.682 $Y=2.21
+ $X2=1.682 $Y2=1.98
r36 9 18 3.31358 $w=4.05e-07 $l=1.1e-07 $layer=LI1_cond $X=1.682 $Y=1.87
+ $X2=1.682 $Y2=1.98
r37 8 9 6.7671 $w=4.05e-07 $l=2.16365e-07 $layer=LI1_cond $X=1.86 $Y=1.785
+ $X2=1.682 $Y2=1.87
r38 8 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.86 $Y=1.785 $X2=1.86
+ $Y2=0.825
r39 2 18 300 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.485 $X2=1.7 $Y2=1.98
r40 1 11 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.235 $X2=2.12 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%A_397_297# 1 2 8 9 10 11 13 16
c28 9 0 1.50675e-19 $X=2.875 $Y=1.87
r29 11 20 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.002 $Y=1.955
+ $X2=3.002 $Y2=1.87
r30 11 13 15.5919 $w=2.53e-07 $l=3.45e-07 $layer=LI1_cond $X=3.002 $Y=1.955
+ $X2=3.002 $Y2=2.3
r31 9 20 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.875 $Y=1.87
+ $X2=3.002 $Y2=1.87
r32 9 10 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.875 $Y=1.87
+ $X2=2.285 $Y2=1.87
r33 8 16 2.50919 $w=1.7e-07 $l=1.4975e-07 $layer=LI1_cond $X=2.2 $Y=2.235
+ $X2=2.12 $Y2=2.35
r34 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.2 $Y=1.955
+ $X2=2.285 $Y2=1.87
r35 7 8 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.2 $Y=1.955 $X2=2.2
+ $Y2=2.235
r36 2 20 600 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.87
r37 2 13 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=2.3
r38 1 16 600 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.485 $X2=2.12 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_1%VGND 1 2 3 10 12 14 17 24 40 43 46 48
r48 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r49 42 43 9.99343 $w=5.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.44 $Y=0.202
+ $X2=1.605 $Y2=0.202
r50 38 42 6.0324 $w=5.73e-07 $l=2.9e-07 $layer=LI1_cond $X=1.15 $Y=0.202
+ $X2=1.44 $Y2=0.202
r51 38 40 11.0335 $w=5.73e-07 $l=2.15e-07 $layer=LI1_cond $X=1.15 $Y=0.202
+ $X2=0.935 $Y2=0.202
r52 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r53 31 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r54 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r55 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r56 28 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r57 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r58 27 43 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.605
+ $Y2=0
r59 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r60 24 45 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.007
+ $Y2=0
r61 24 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.53
+ $Y2=0
r62 23 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r63 22 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=0.935
+ $Y2=0
r64 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r65 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r66 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r67 14 48 8.44056 $w=4.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r68 14 20 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.212 $Y=0 $X2=0.425
+ $Y2=0
r69 14 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 10 45 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=3.007 $Y2=0
r71 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=0.085
+ $X2=2.96 $Y2=0.38
r72 3 12 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.38
r73 2 42 91 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.44 $Y2=0.38
r74 1 48 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__or2b_2.pxi.spice
* Created: Thu Aug 27 14:43:03 2020
* 
x_PM_SKY130_FD_SC_HD__OR2B_2%B_N N_B_N_M1002_g N_B_N_M1007_g B_N N_B_N_c_59_n
+ B_N PM_SKY130_FD_SC_HD__OR2B_2%B_N
x_PM_SKY130_FD_SC_HD__OR2B_2%A_27_53# N_A_27_53#_M1002_s N_A_27_53#_M1007_d
+ N_A_27_53#_M1004_g N_A_27_53#_M1006_g N_A_27_53#_c_82_n N_A_27_53#_c_83_n
+ N_A_27_53#_c_84_n N_A_27_53#_c_89_n N_A_27_53#_c_85_n N_A_27_53#_c_86_n
+ PM_SKY130_FD_SC_HD__OR2B_2%A_27_53#
x_PM_SKY130_FD_SC_HD__OR2B_2%A N_A_c_126_n N_A_M1003_g N_A_M1008_g A N_A_c_129_n
+ PM_SKY130_FD_SC_HD__OR2B_2%A
x_PM_SKY130_FD_SC_HD__OR2B_2%A_218_297# N_A_218_297#_M1004_d
+ N_A_218_297#_M1006_s N_A_218_297#_c_161_n N_A_218_297#_M1005_g
+ N_A_218_297#_M1000_g N_A_218_297#_c_162_n N_A_218_297#_M1009_g
+ N_A_218_297#_M1001_g N_A_218_297#_c_175_n N_A_218_297#_c_228_p
+ N_A_218_297#_c_163_n N_A_218_297#_c_164_n N_A_218_297#_c_170_n
+ N_A_218_297#_c_171_n N_A_218_297#_c_165_n N_A_218_297#_c_166_n
+ N_A_218_297#_c_167_n PM_SKY130_FD_SC_HD__OR2B_2%A_218_297#
x_PM_SKY130_FD_SC_HD__OR2B_2%VPWR N_VPWR_M1007_s N_VPWR_M1008_d N_VPWR_M1001_d
+ N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n
+ VPWR N_VPWR_c_243_n N_VPWR_c_244_n N_VPWR_c_245_n N_VPWR_c_237_n
+ PM_SKY130_FD_SC_HD__OR2B_2%VPWR
x_PM_SKY130_FD_SC_HD__OR2B_2%X N_X_M1005_d N_X_M1000_s N_X_c_279_n N_X_c_281_n
+ N_X_c_277_n X PM_SKY130_FD_SC_HD__OR2B_2%X
x_PM_SKY130_FD_SC_HD__OR2B_2%VGND N_VGND_M1002_d N_VGND_M1003_d N_VGND_M1009_s
+ N_VGND_c_301_n N_VGND_c_302_n N_VGND_c_303_n VGND N_VGND_c_304_n
+ N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n
+ PM_SKY130_FD_SC_HD__OR2B_2%VGND
cc_1 VNB N_B_N_M1002_g 0.0404018f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB B_N 0.00929235f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_B_N_c_59_n 0.0403913f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_53#_M1004_g 0.0326337f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_53#_c_82_n 0.0197455f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_6 VNB N_A_27_53#_c_83_n 0.0154532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_53#_c_84_n 0.00895122f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_8 VNB N_A_27_53#_c_85_n 0.00459903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_53#_c_86_n 0.0346441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_M1003_g 0.041529f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_11 VNB N_A_218_297#_c_161_n 0.0164367f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.695
cc_12 VNB N_A_218_297#_c_162_n 0.0204745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_218_297#_c_163_n 0.00188528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_218_297#_c_164_n 0.00407348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_218_297#_c_165_n 0.00315488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_218_297#_c_166_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_218_297#_c_167_n 0.0494546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_237_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_277_n 7.1028e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_301_n 5.53369e-19 $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_21 VNB N_VGND_c_302_n 0.0123691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_303_n 0.0105265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_304_n 0.0122945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_305_n 0.0160155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_306_n 0.0174027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_307_n 0.019064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_308_n 0.0052385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_309_n 0.188783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_B_N_M1007_g 0.0294126f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_30 VPB B_N 8.86575e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_31 VPB N_B_N_c_59_n 0.0103665f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_32 VPB N_A_27_53#_M1006_g 0.0226372f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_33 VPB N_A_27_53#_c_83_n 0.00328375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_53#_c_89_n 0.00456577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_53#_c_85_n 0.00639431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_53#_c_86_n 0.00826773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_c_126_n 0.043427f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_38 VPB N_A_M1003_g 0.0314341f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_39 VPB A 0.0261628f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_40 VPB N_A_c_129_n 0.0371693f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_41 VPB N_A_218_297#_M1000_g 0.0209233f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_42 VPB N_A_218_297#_M1001_g 0.0246565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_218_297#_c_170_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_218_297#_c_171_n 0.00812057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_218_297#_c_165_n 2.03541e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_218_297#_c_167_n 0.00896334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_238_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_239_n 0.0557125f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_VPWR_c_240_n 0.0113766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_241_n 0.0123399f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_51 VPB N_VPWR_c_242_n 0.00974244f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_52 VPB N_VPWR_c_243_n 0.0395879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_244_n 0.0170833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_245_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_237_n 0.0634504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_X_c_277_n 0.00103314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 N_B_N_M1002_g N_A_27_53#_c_82_n 0.0125834f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_58 N_B_N_M1002_g N_A_27_53#_c_83_n 0.0228336f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_59 B_N N_A_27_53#_c_83_n 0.0196208f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_60 N_B_N_M1002_g N_A_27_53#_c_84_n 0.00414204f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_61 B_N N_A_27_53#_c_84_n 0.0258233f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_62 N_B_N_c_59_n N_A_27_53#_c_84_n 0.00741854f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_63 N_B_N_c_59_n N_A_27_53#_c_89_n 0.0083141f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B_N_c_59_n N_A_27_53#_c_86_n 0.00533699f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_65 N_B_N_M1007_g A 2.52857e-19 $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_66 N_B_N_M1007_g N_A_218_297#_c_171_n 0.00134798f $X=0.47 $Y=1.695 $X2=0
+ $Y2=0
cc_67 N_B_N_M1007_g N_VPWR_c_239_n 0.00616807f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_68 B_N N_VPWR_c_239_n 0.0207928f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_69 N_B_N_c_59_n N_VPWR_c_239_n 0.00554938f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_70 N_B_N_M1007_g N_VPWR_c_243_n 0.00317366f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_71 N_B_N_M1007_g N_VPWR_c_237_n 0.00403572f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_72 N_B_N_M1002_g N_VGND_c_306_n 0.00402941f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_73 N_B_N_M1002_g N_VGND_c_307_n 0.00505351f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_74 N_B_N_M1002_g N_VGND_c_309_n 0.0073571f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_75 N_A_27_53#_M1006_g N_A_c_126_n 0.00868417f $X=1.425 $Y=1.695 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_27_53#_M1004_g N_A_M1003_g 0.022046f $X=1.365 $Y=0.475 $X2=0 $Y2=0
cc_77 N_A_27_53#_c_85_n N_A_M1003_g 0.0014977f $X=1.215 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_27_53#_c_86_n N_A_M1003_g 0.0652533f $X=1.425 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_27_53#_M1006_g A 0.00164982f $X=1.425 $Y=1.695 $X2=0 $Y2=0
cc_80 N_A_27_53#_c_89_n A 0.0122083f $X=0.68 $Y=1.63 $X2=0 $Y2=0
cc_81 N_A_27_53#_M1006_g N_A_218_297#_c_175_n 0.00917186f $X=1.425 $Y=1.695
+ $X2=0 $Y2=0
cc_82 N_A_27_53#_M1004_g N_A_218_297#_c_164_n 0.00310482f $X=1.365 $Y=0.475
+ $X2=0 $Y2=0
cc_83 N_A_27_53#_c_83_n N_A_218_297#_c_164_n 0.00301169f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_84 N_A_27_53#_c_86_n N_A_218_297#_c_164_n 3.34812e-19 $X=1.425 $Y=1.16 $X2=0
+ $Y2=0
cc_85 N_A_27_53#_M1006_g N_A_218_297#_c_171_n 0.0100132f $X=1.425 $Y=1.695 $X2=0
+ $Y2=0
cc_86 N_A_27_53#_c_89_n N_A_218_297#_c_171_n 0.0257662f $X=0.68 $Y=1.63 $X2=0
+ $Y2=0
cc_87 N_A_27_53#_c_85_n N_A_218_297#_c_171_n 0.0263501f $X=1.215 $Y=1.16 $X2=0
+ $Y2=0
cc_88 N_A_27_53#_c_86_n N_A_218_297#_c_171_n 0.0062777f $X=1.425 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A_27_53#_M1004_g N_VGND_c_301_n 5.2524e-19 $X=1.365 $Y=0.475 $X2=0 $Y2=0
cc_90 N_A_27_53#_M1004_g N_VGND_c_304_n 0.00442511f $X=1.365 $Y=0.475 $X2=0
+ $Y2=0
cc_91 N_A_27_53#_c_82_n N_VGND_c_306_n 0.0187097f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_53#_c_83_n N_VGND_c_306_n 0.00229799f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_93 N_A_27_53#_M1004_g N_VGND_c_307_n 0.00956695f $X=1.365 $Y=0.475 $X2=0
+ $Y2=0
cc_94 N_A_27_53#_c_83_n N_VGND_c_307_n 0.0210226f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_95 N_A_27_53#_c_85_n N_VGND_c_307_n 0.0188842f $X=1.215 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_27_53#_c_86_n N_VGND_c_307_n 0.00387909f $X=1.425 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_27_53#_M1004_g N_VGND_c_309_n 0.00779323f $X=1.365 $Y=0.475 $X2=0
+ $Y2=0
cc_98 N_A_27_53#_c_82_n N_VGND_c_309_n 0.0118569f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_27_53#_c_83_n N_VGND_c_309_n 0.00488127f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_100 N_A_M1003_g N_A_218_297#_c_161_n 0.0172583f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_101 N_A_M1003_g N_A_218_297#_M1000_g 0.0251997f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_102 N_A_c_126_n N_A_218_297#_c_175_n 6.94119e-19 $X=1.71 $Y=2.34 $X2=0 $Y2=0
cc_103 N_A_M1003_g N_A_218_297#_c_175_n 0.0166311f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_104 A N_A_218_297#_c_175_n 0.0108145f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_105 N_A_M1003_g N_A_218_297#_c_163_n 0.0134701f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_106 N_A_c_126_n N_A_218_297#_c_171_n 9.41055e-19 $X=1.71 $Y=2.34 $X2=0 $Y2=0
cc_107 N_A_M1003_g N_A_218_297#_c_171_n 0.00122623f $X=1.785 $Y=0.475 $X2=0
+ $Y2=0
cc_108 A N_A_218_297#_c_171_n 0.034396f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_109 N_A_c_129_n N_A_218_297#_c_171_n 0.00119166f $X=1.17 $Y=2.28 $X2=0 $Y2=0
cc_110 N_A_M1003_g N_A_218_297#_c_166_n 0.0136533f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_111 N_A_M1003_g N_A_218_297#_c_167_n 0.0196839f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_112 A N_VPWR_c_239_n 0.0258923f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_113 N_A_c_129_n N_VPWR_c_239_n 0.00101565f $X=1.17 $Y=2.28 $X2=0 $Y2=0
cc_114 N_A_M1003_g N_VPWR_c_240_n 0.00820852f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_115 A N_VPWR_c_240_n 0.0259888f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_116 A N_VPWR_c_243_n 0.0584919f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_117 N_A_c_129_n N_VPWR_c_243_n 0.0214212f $X=1.17 $Y=2.28 $X2=0 $Y2=0
cc_118 A N_VPWR_c_237_n 0.043085f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_119 N_A_c_129_n N_VPWR_c_237_n 0.0300519f $X=1.17 $Y=2.28 $X2=0 $Y2=0
cc_120 N_A_M1003_g N_VGND_c_301_n 0.00709022f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_121 N_A_M1003_g N_VGND_c_304_n 0.00322006f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_122 N_A_M1003_g N_VGND_c_307_n 5.59171e-19 $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_123 N_A_M1003_g N_VGND_c_309_n 0.00390029f $X=1.785 $Y=0.475 $X2=0 $Y2=0
cc_124 N_A_218_297#_c_175_n N_VPWR_M1008_d 0.00526233f $X=2.06 $Y=1.58 $X2=0
+ $Y2=0
cc_125 N_A_218_297#_c_171_n N_VPWR_c_239_n 6.52973e-19 $X=1.195 $Y=1.58 $X2=0
+ $Y2=0
cc_126 N_A_218_297#_M1000_g N_VPWR_c_240_n 0.00342332f $X=2.275 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_218_297#_c_175_n N_VPWR_c_240_n 0.0190361f $X=2.06 $Y=1.58 $X2=0
+ $Y2=0
cc_128 N_A_218_297#_c_171_n N_VPWR_c_240_n 0.00145048f $X=1.195 $Y=1.58 $X2=0
+ $Y2=0
cc_129 N_A_218_297#_c_167_n N_VPWR_c_240_n 3.85151e-19 $X=2.695 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A_218_297#_M1001_g N_VPWR_c_242_n 0.00384418f $X=2.695 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_218_297#_M1000_g N_VPWR_c_244_n 0.00585385f $X=2.275 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_218_297#_M1001_g N_VPWR_c_244_n 0.00571722f $X=2.695 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_218_297#_M1000_g N_VPWR_c_237_n 0.0118387f $X=2.275 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_218_297#_M1001_g N_VPWR_c_237_n 0.0112329f $X=2.695 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_218_297#_c_175_n A_300_297# 0.0033195f $X=2.06 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_218_297#_c_162_n N_X_c_279_n 0.00344035f $X=2.695 $Y=0.995 $X2=0
+ $Y2=0
cc_137 N_A_218_297#_c_167_n N_X_c_279_n 7.59141e-19 $X=2.695 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_218_297#_M1001_g N_X_c_281_n 0.00211913f $X=2.695 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_218_297#_c_167_n N_X_c_281_n 8.88826e-19 $X=2.695 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_218_297#_c_161_n N_X_c_277_n 0.00152341f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_218_297#_M1000_g N_X_c_277_n 0.00116659f $X=2.275 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_218_297#_c_162_n N_X_c_277_n 0.00583782f $X=2.695 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_218_297#_M1001_g N_X_c_277_n 0.00681792f $X=2.695 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_218_297#_c_163_n N_X_c_277_n 0.00401263f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_218_297#_c_170_n N_X_c_277_n 0.0096046f $X=2.145 $Y=1.495 $X2=0 $Y2=0
cc_146 N_A_218_297#_c_165_n N_X_c_277_n 0.0228995f $X=2.205 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_218_297#_c_166_n N_X_c_277_n 0.0095636f $X=2.175 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_218_297#_c_167_n N_X_c_277_n 0.0255199f $X=2.695 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_218_297#_M1001_g X 0.00938209f $X=2.695 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_218_297#_c_163_n N_VGND_M1003_d 0.00482895f $X=2.06 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_218_297#_c_166_n N_VGND_M1003_d 6.98847e-19 $X=2.175 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_218_297#_c_161_n N_VGND_c_301_n 0.00770036f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_218_297#_c_162_n N_VGND_c_301_n 9.22792e-19 $X=2.695 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_A_218_297#_c_163_n N_VGND_c_301_n 0.020701f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_218_297#_c_167_n N_VGND_c_301_n 4.03696e-19 $X=2.695 $Y=1.16 $X2=0
+ $Y2=0
cc_156 N_A_218_297#_c_162_n N_VGND_c_303_n 0.00416229f $X=2.695 $Y=0.995 $X2=0
+ $Y2=0
cc_157 N_A_218_297#_c_228_p N_VGND_c_304_n 0.00846569f $X=1.575 $Y=0.47 $X2=0
+ $Y2=0
cc_158 N_A_218_297#_c_163_n N_VGND_c_304_n 0.00232396f $X=2.06 $Y=0.74 $X2=0
+ $Y2=0
cc_159 N_A_218_297#_c_161_n N_VGND_c_305_n 0.00524631f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_218_297#_c_162_n N_VGND_c_305_n 0.00573595f $X=2.695 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A_218_297#_c_163_n N_VGND_c_305_n 3.34073e-19 $X=2.06 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_218_297#_c_161_n N_VGND_c_309_n 0.00851181f $X=2.275 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_218_297#_c_162_n N_VGND_c_309_n 0.0112418f $X=2.695 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_218_297#_c_228_p N_VGND_c_309_n 0.00625722f $X=1.575 $Y=0.47 $X2=0
+ $Y2=0
cc_165 N_A_218_297#_c_163_n N_VGND_c_309_n 0.00637905f $X=2.06 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_VPWR_c_237_n N_X_M1000_s 0.00393857f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_167 N_VPWR_c_242_n N_X_c_277_n 0.0365142f $X=2.905 $Y=1.65 $X2=0 $Y2=0
cc_168 N_VPWR_c_244_n X 0.013819f $X=2.8 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_c_237_n X 0.00873952f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_170 N_VPWR_c_242_n N_VGND_c_303_n 0.0106517f $X=2.905 $Y=1.65 $X2=0 $Y2=0
cc_171 N_X_c_279_n N_VGND_c_303_n 0.0193667f $X=2.485 $Y=0.59 $X2=0 $Y2=0
cc_172 N_X_c_279_n N_VGND_c_305_n 0.00670356f $X=2.485 $Y=0.59 $X2=0 $Y2=0
cc_173 N_X_M1005_d N_VGND_c_309_n 0.0041316f $X=2.35 $Y=0.235 $X2=0 $Y2=0
cc_174 N_X_c_279_n N_VGND_c_309_n 0.00790197f $X=2.485 $Y=0.59 $X2=0 $Y2=0

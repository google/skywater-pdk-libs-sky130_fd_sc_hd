# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nand2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.315000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.085000 1.315000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 1.835000 2.170000 2.005000 ;
        RECT 1.000000 2.005000 1.330000 2.465000 ;
        RECT 1.420000 0.255000 2.170000 0.545000 ;
        RECT 1.800000 0.545000 2.170000 1.835000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.300000 0.085000 ;
        RECT 0.580000  0.085000 0.910000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.300000 2.805000 ;
        RECT 0.580000 1.835000 0.830000 2.635000 ;
        RECT 1.500000 2.175000 1.715000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.525000 0.360000 0.735000 ;
      RECT 0.090000 0.735000 1.425000 0.905000 ;
      RECT 0.090000 1.495000 1.425000 1.665000 ;
      RECT 0.090000 1.665000 0.370000 1.825000 ;
      RECT 1.255000 0.905000 1.425000 1.075000 ;
      RECT 1.255000 1.075000 1.630000 1.325000 ;
      RECT 1.255000 1.325000 1.425000 1.495000 ;
  END
END sky130_fd_sc_hd__nand2b_1

* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_1.spice.pex
* Created: Thu Aug 27 14:23:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%A_75_212# 1 2 9 13 18 19 20 21
+ 22 25 29 32 33 34
c73 22 0 4.19985e-20 $X=0.71 $Y=1.62
c74 19 0 1.55858e-19 $X=1.035 $Y=0.72
c75 9 0 6.6635e-20 $X=0.47 $Y=0.495
r76 33 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.225
+ $X2=0.51 $Y2=1.39
r77 33 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.225
+ $X2=0.51 $Y2=1.06
r78 32 35 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=1.225
+ $X2=0.567 $Y2=1.39
r79 32 34 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.567 $Y=1.225
+ $X2=0.567 $Y2=1.06
r80 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.225 $X2=0.51 $Y2=1.225
r81 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.12 $Y=1.705
+ $X2=1.12 $Y2=1.96
r82 23 25 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.12 $Y=0.635
+ $X2=1.12 $Y2=0.445
r83 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.62
+ $X2=1.12 $Y2=1.705
r84 21 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.035 $Y=1.62
+ $X2=0.71 $Y2=1.62
r85 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=0.72
+ $X2=1.12 $Y2=0.635
r86 19 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.035 $Y=0.72
+ $X2=0.71 $Y2=0.72
r87 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.535
+ $X2=0.71 $Y2=1.62
r88 18 35 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.625 $Y=1.535
+ $X2=0.625 $Y2=1.39
r89 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=0.805
+ $X2=0.71 $Y2=0.72
r90 15 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.625 $Y=0.805
+ $X2=0.625 $Y2=1.06
r91 13 38 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.47 $Y=2.09 $X2=0.47
+ $Y2=1.39
r92 9 37 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.47 $Y=0.495
+ $X2=0.47 $Y2=1.06
r93 2 29 300 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.695 $X2=1.12 $Y2=1.96
r94 1 25 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%A 1 3 6 7 9 10 11
c32 11 0 6.6635e-20 $X=1.15 $Y=1.19
c33 10 0 1.55858e-19 $X=0.925 $Y=1.62
r34 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.16 $X2=1.11 $Y2=1.16
r35 9 10 46.6452 $w=1.8e-07 $l=1.2e-07 $layer=POLY_cond $X=0.925 $Y=1.5
+ $X2=0.925 $Y2=1.62
r36 7 14 38.5318 $w=3.1e-07 $l=2.09105e-07 $layer=POLY_cond $X=0.94 $Y=1.325
+ $X2=1.04 $Y2=1.16
r37 7 9 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.94 $Y=1.325 $X2=0.94
+ $Y2=1.5
r38 6 10 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.91 $Y=2.09 $X2=0.91
+ $Y2=1.62
r39 1 14 64.1867 $w=3.1e-07 $l=3.89615e-07 $layer=POLY_cond $X=0.91 $Y=0.83
+ $X2=1.04 $Y2=1.16
r40 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.91 $Y=0.83 $X2=0.91
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%X 1 2 10 11 12 13 14 15
r28 14 15 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.22 $Y=1.87
+ $X2=0.22 $Y2=2.21
r29 11 14 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.22 $Y=1.695
+ $X2=0.22 $Y2=1.87
r30 11 12 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=1.695
+ $X2=0.22 $Y2=1.56
r31 10 12 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.17 $Y=0.76 $X2=0.17
+ $Y2=1.56
r32 9 13 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=0.215 $Y=0.63
+ $X2=0.215 $Y2=0.51
r33 9 10 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=0.63
+ $X2=0.215 $Y2=0.76
r34 2 14 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.695 $X2=0.26 $Y2=1.895
r35 1 13 182 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%KAPWR 1 8 10 12 15 21
c27 10 0 4.19985e-20 $X=0.55 $Y=2.21
r28 12 21 0.001875 $w=2e-07 $l=3e-09 $layer=MET1_cond $X=0.467 $Y=2.24 $X2=0.47
+ $Y2=2.24
r29 10 21 0.05 $w=2e-07 $l=8e-08 $layer=MET1_cond $X=0.55 $Y=2.24 $X2=0.47
+ $Y2=2.24
r30 9 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=2.21 $X2=0.69
+ $Y2=1.96
r31 8 10 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.695 $Y=2.21
+ $X2=0.55 $Y2=2.21
r32 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=2.21
+ $X2=0.695 $Y2=2.21
r33 1 15 300 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.695 $X2=0.69 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%VGND 1 6 8 10 17 21
r26 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r28 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.15
+ $Y2=0
r29 13 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r30 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r31 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r32 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.23
+ $Y2=0
r33 8 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r34 8 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r36 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r37 1 6 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%VPWR 1 8
r19 4 8 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=1.15
+ $Y2=2.72
r20 4 5 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r21 1 5 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72 $X2=0.23
+ $Y2=2.72
r22 1 8 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72 $X2=1.15
+ $Y2=2.72
.ends


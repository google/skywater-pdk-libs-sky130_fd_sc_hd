# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__sdfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.18000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.325000 4.025000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.415000 0.255000 14.665000 0.825000 ;
        RECT 14.415000 1.445000 14.665000 2.465000 ;
        RECT 14.460000 0.825000 14.665000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.580000 0.255000 12.830000 0.715000 ;
        RECT 12.580000 1.630000 12.830000 2.465000 ;
        RECT 12.660000 0.715000 12.830000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.590000 1.095000 12.070000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.025000 1.695000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.345000 2.145000 0.765000 ;
        RECT 1.935000 0.765000 2.335000 1.095000 ;
        RECT 1.935000 1.095000 2.155000 1.695000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.735000 6.295000 0.965000 ;
        RECT 5.885000 0.965000 6.215000 1.065000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 0.735000 10.130000 1.065000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065000 0.735000  6.355000 0.780000 ;
        RECT 6.065000 0.780000 10.035000 0.920000 ;
        RECT 6.065000 0.920000  6.355000 0.965000 ;
        RECT 9.745000 0.735000 10.035000 0.780000 ;
        RECT 9.745000 0.920000 10.035000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.180000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  1.430000  0.085000  1.705000 0.635000 ;
        RECT  3.370000  0.085000  3.700000 0.445000 ;
        RECT  5.885000  0.085000  6.055000 0.525000 ;
        RECT  7.645000  0.085000  7.975000 0.465000 ;
        RECT  9.560000  0.085000  9.820000 0.525000 ;
        RECT 12.080000  0.085000 12.410000 0.805000 ;
        RECT 13.000000  0.085000 13.235000 0.885000 ;
        RECT 13.950000  0.085000 14.245000 0.545000 ;
        RECT 14.835000  0.085000 15.075000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.180000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 15.180000 2.805000 ;
        RECT  0.515000 2.135000  0.845000 2.635000 ;
        RECT  1.430000 1.885000  1.785000 2.635000 ;
        RECT  3.295000 2.215000  3.640000 2.635000 ;
        RECT  5.705000 2.205000  6.085000 2.635000 ;
        RECT  7.175000 1.915000  7.505000 2.635000 ;
        RECT  9.620000 2.255000 10.000000 2.635000 ;
        RECT 10.940000 2.255000 12.410000 2.635000 ;
        RECT 13.000000 1.495000 13.235000 2.635000 ;
        RECT 13.950000 1.765000 14.245000 2.635000 ;
        RECT 14.835000 1.495000 15.075000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.180000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.170000 0.345000  0.345000 0.635000 ;
      RECT  0.170000 0.635000  0.835000 0.805000 ;
      RECT  0.170000 1.795000  0.835000 1.965000 ;
      RECT  0.170000 1.965000  0.345000 2.465000 ;
      RECT  0.605000 0.805000  0.835000 1.795000 ;
      RECT  1.015000 0.345000  1.235000 2.465000 ;
      RECT  2.215000 1.875000  2.575000 2.385000 ;
      RECT  2.315000 0.265000  2.730000 0.595000 ;
      RECT  2.405000 1.250000  3.075000 1.405000 ;
      RECT  2.405000 1.405000  2.575000 1.875000 ;
      RECT  2.435000 1.235000  3.075000 1.250000 ;
      RECT  2.560000 0.595000  2.730000 1.075000 ;
      RECT  2.560000 1.075000  3.075000 1.235000 ;
      RECT  2.745000 1.575000  3.645000 1.745000 ;
      RECT  2.745000 1.745000  3.065000 1.905000 ;
      RECT  2.895000 1.905000  3.065000 2.465000 ;
      RECT  2.955000 0.305000  3.125000 0.625000 ;
      RECT  2.955000 0.625000  3.645000 0.765000 ;
      RECT  2.955000 0.765000  3.770000 0.795000 ;
      RECT  3.475000 0.795000  3.770000 1.095000 ;
      RECT  3.475000 1.095000  3.645000 1.575000 ;
      RECT  4.230000 0.305000  4.455000 2.465000 ;
      RECT  4.625000 0.705000  4.845000 1.575000 ;
      RECT  4.625000 1.575000  5.125000 1.955000 ;
      RECT  4.635000 2.250000  5.465000 2.420000 ;
      RECT  4.700000 0.265000  5.715000 0.465000 ;
      RECT  5.025000 0.645000  5.375000 1.015000 ;
      RECT  5.295000 1.195000  5.715000 1.235000 ;
      RECT  5.295000 1.235000  6.645000 1.405000 ;
      RECT  5.295000 1.405000  5.465000 2.250000 ;
      RECT  5.545000 0.465000  5.715000 1.195000 ;
      RECT  5.635000 1.575000  5.885000 1.785000 ;
      RECT  5.635000 1.785000  6.985000 2.035000 ;
      RECT  6.225000 0.255000  7.375000 0.425000 ;
      RECT  6.225000 0.425000  6.555000 0.505000 ;
      RECT  6.385000 2.035000  6.555000 2.375000 ;
      RECT  6.395000 1.405000  6.645000 1.485000 ;
      RECT  6.425000 1.155000  6.645000 1.235000 ;
      RECT  6.705000 0.595000  7.035000 0.765000 ;
      RECT  6.815000 0.765000  7.035000 0.895000 ;
      RECT  6.815000 0.895000  8.125000 1.065000 ;
      RECT  6.815000 1.065000  6.985000 1.785000 ;
      RECT  7.155000 1.235000  7.485000 1.415000 ;
      RECT  7.155000 1.415000  8.160000 1.655000 ;
      RECT  7.205000 0.425000  7.375000 0.715000 ;
      RECT  7.795000 1.065000  8.125000 1.235000 ;
      RECT  8.360000 1.575000  8.595000 1.985000 ;
      RECT  8.420000 0.705000  8.705000 1.125000 ;
      RECT  8.420000 1.125000  9.040000 1.305000 ;
      RECT  8.550000 2.250000  9.380000 2.420000 ;
      RECT  8.615000 0.265000  9.380000 0.465000 ;
      RECT  8.835000 1.305000  9.040000 1.905000 ;
      RECT  9.210000 0.465000  9.380000 1.235000 ;
      RECT  9.210000 1.235000 10.560000 1.405000 ;
      RECT  9.210000 1.405000  9.380000 2.250000 ;
      RECT  9.550000 1.575000  9.800000 1.915000 ;
      RECT  9.550000 1.915000 12.410000 2.085000 ;
      RECT 10.080000 0.255000 11.250000 0.425000 ;
      RECT 10.080000 0.425000 10.410000 0.545000 ;
      RECT 10.240000 2.085000 10.410000 2.375000 ;
      RECT 10.340000 1.075000 10.560000 1.235000 ;
      RECT 10.580000 0.595000 10.910000 0.780000 ;
      RECT 10.730000 0.780000 10.910000 1.915000 ;
      RECT 11.080000 0.425000 11.250000 0.585000 ;
      RECT 11.080000 0.755000 11.845000 0.925000 ;
      RECT 11.080000 0.925000 11.355000 1.575000 ;
      RECT 11.080000 1.575000 11.925000 1.745000 ;
      RECT 11.620000 0.265000 11.845000 0.755000 ;
      RECT 12.240000 0.995000 12.480000 1.325000 ;
      RECT 12.240000 1.325000 12.410000 1.915000 ;
      RECT 13.455000 0.255000 13.770000 0.995000 ;
      RECT 13.455000 0.995000 14.290000 1.325000 ;
      RECT 13.455000 1.325000 13.770000 2.415000 ;
    LAYER mcon ;
      RECT  0.605000 0.765000  0.775000 0.935000 ;
      RECT  1.065000 1.785000  1.235000 1.955000 ;
      RECT  2.905000 1.105000  3.075000 1.275000 ;
      RECT  4.285000 1.105000  4.455000 1.275000 ;
      RECT  4.745000 1.785000  4.915000 1.955000 ;
      RECT  5.205000 0.765000  5.375000 0.935000 ;
      RECT  7.965000 1.445000  8.135000 1.615000 ;
      RECT  8.425000 1.105000  8.595000 1.275000 ;
      RECT  8.425000 1.785000  8.595000 1.955000 ;
      RECT 11.185000 1.445000 11.355000 1.615000 ;
    LAYER met1 ;
      RECT  0.545000 0.735000  0.835000 0.780000 ;
      RECT  0.545000 0.780000  5.435000 0.920000 ;
      RECT  0.545000 0.920000  0.835000 0.965000 ;
      RECT  1.005000 1.755000  1.295000 1.800000 ;
      RECT  1.005000 1.800000  8.655000 1.940000 ;
      RECT  1.005000 1.940000  1.295000 1.985000 ;
      RECT  2.845000 1.075000  3.135000 1.120000 ;
      RECT  2.845000 1.120000  4.515000 1.260000 ;
      RECT  2.845000 1.260000  3.135000 1.305000 ;
      RECT  4.225000 1.075000  4.515000 1.120000 ;
      RECT  4.225000 1.260000  4.515000 1.305000 ;
      RECT  4.685000 1.755000  4.975000 1.800000 ;
      RECT  4.685000 1.940000  4.975000 1.985000 ;
      RECT  5.145000 0.735000  5.435000 0.780000 ;
      RECT  5.145000 0.920000  5.435000 0.965000 ;
      RECT  5.220000 0.965000  5.435000 1.120000 ;
      RECT  5.220000 1.120000  8.655000 1.260000 ;
      RECT  7.905000 1.415000  8.195000 1.460000 ;
      RECT  7.905000 1.460000 11.415000 1.600000 ;
      RECT  7.905000 1.600000  8.195000 1.645000 ;
      RECT  8.365000 1.075000  8.655000 1.120000 ;
      RECT  8.365000 1.260000  8.655000 1.305000 ;
      RECT  8.365000 1.755000  8.655000 1.800000 ;
      RECT  8.365000 1.940000  8.655000 1.985000 ;
      RECT 11.125000 1.415000 11.415000 1.460000 ;
      RECT 11.125000 1.600000 11.415000 1.645000 ;
  END
END sky130_fd_sc_hd__sdfbbn_2
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_1269_47# A3 a_911_47# VNB nshort w=650000u l=150000u
+  ad=8.84e+11p pd=9.22e+06u as=7.02e+11p ps=7.36e+06u
M1001 VGND A4 a_1269_47# VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=9.16e+06u as=0p ps=0u
M1002 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.405e+12p pd=2.881e+07u as=2.905e+12p ps=2.181e+07u
M1003 Y A1 a_493_47# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=8.645e+11p ps=9.16e+06u
M1004 a_493_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1006 a_493_47# A2 a_911_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A4 a_1269_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A1 a_493_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_493_47# A2 a_911_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_911_47# A2 a_493_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_493_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_297# A4 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1269_47# A4 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A4 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_297# A4 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_911_47# A3 a_1269_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR A4 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1269_47# A3 a_911_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_911_47# A3 a_1269_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_27_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1269_47# A4 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_911_47# A2 a_493_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

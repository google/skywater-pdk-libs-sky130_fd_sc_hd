* File: sky130_fd_sc_hd__o211ai_1.spice
* Created: Thu Aug 27 14:34:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o211ai_1.spice.pex"
.subckt sky130_fd_sc_hd__o211ai_1  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A1_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.17225 PD=1.04 PS=1.83 NRD=12.912 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1004_d N_A2_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.12675 PD=1.04 PS=1.04 NRD=11.076 NRS=7.38 M=1 R=4.33333
+ SA=75000.7 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1006 A_326_47# N_B1_M1006_g N_A_27_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.12675 PD=0.86 PS=1.04 NRD=9.228 NRS=9.228 M=1 R=4.33333
+ SA=75001.3 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g A_326_47# VNB NSHORT L=0.15 W=0.65 AD=0.39325
+ AS=0.06825 PD=2.51 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.6 SB=75000.5
+ A=0.0975 P=1.6 MULT=1
MM1003 A_110_297# N_A1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.265 PD=1.21 PS=2.53 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A2_M1001_g A_110_297# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.105 PD=1.39 PS=1.21 NRD=11.8003 NRS=9.8303 M=1 R=6.66667 SA=75000.5
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.195 PD=1.39 PS=1.39 NRD=3.9203 NRS=9.8303 M=1 R=6.66667 SA=75001.1
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_C1_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.635
+ AS=0.195 PD=3.27 PS=1.39 NRD=1.9503 NRS=17.73 M=1 R=6.66667 SA=75001.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__o211ai_1.spice.SKY130_FD_SC_HD__O211AI_1.pxi"
*
.ends
*
*

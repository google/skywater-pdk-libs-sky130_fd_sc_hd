# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.100000 1.075000 3.595000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.075000 2.930000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.325000 ;
        RECT 0.595000 1.325000 0.775000 1.695000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.255000 1.240000 0.595000 ;
        RECT 0.945000 0.595000 1.115000 1.495000 ;
        RECT 0.945000 1.495000 1.350000 1.695000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.430000 0.345000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 0.395000 1.865000 ;
      RECT 0.085000  1.865000 1.935000 2.035000 ;
      RECT 0.520000  2.205000 0.910000 2.635000 ;
      RECT 0.595000  0.085000 0.775000 0.825000 ;
      RECT 1.285000  0.890000 1.595000 1.060000 ;
      RECT 1.285000  1.060000 1.455000 1.325000 ;
      RECT 1.410000  0.085000 1.770000 0.485000 ;
      RECT 1.415000  2.205000 2.230000 2.635000 ;
      RECT 1.425000  0.655000 2.275000 0.825000 ;
      RECT 1.425000  0.825000 1.595000 0.890000 ;
      RECT 1.765000  0.995000 1.935000 1.865000 ;
      RECT 1.940000  0.255000 2.275000 0.655000 ;
      RECT 2.105000  0.825000 2.275000 1.455000 ;
      RECT 2.105000  1.455000 2.725000 2.035000 ;
      RECT 2.400000  2.035000 2.725000 2.465000 ;
      RECT 2.445000  0.365000 2.745000 0.735000 ;
      RECT 2.445000  0.735000 3.590000 0.905000 ;
      RECT 2.915000  0.085000 3.085000 0.555000 ;
      RECT 3.200000  1.875000 3.530000 2.635000 ;
      RECT 3.255000  0.270000 3.590000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ba_2
END LIBRARY

* File: sky130_fd_sc_hd__a2111oi_4.spice.pex
* Created: Thu Aug 27 13:59:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2111OI_4%D1 3 5 7 8 10 13 15 17 20 22 24 27 29 41
+ 42
r76 40 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.68 $Y=1.16 $X2=1.77
+ $Y2=1.16
r77 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.16 $X2=1.68 $Y2=1.16
r78 38 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.34 $Y=1.16
+ $X2=1.68 $Y2=1.16
r79 37 38 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.34 $Y2=1.16
r80 35 37 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.66 $Y=1.16
+ $X2=0.91 $Y2=1.16
r81 33 35 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.66 $Y2=1.16
r82 31 33 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.48 $Y=1.16 $X2=0.49
+ $Y2=1.16
r83 29 41 46.0977 $w=2.53e-07 $l=1.02e-06 $layer=LI1_cond $X=0.66 $Y=1.147
+ $X2=1.68 $Y2=1.147
r84 29 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.66
+ $Y=1.16 $X2=0.66 $Y2=1.16
r85 25 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=1.16
r86 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=1.985
r87 22 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=0.995
+ $X2=1.77 $Y2=1.16
r88 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.77 $Y=0.995
+ $X2=1.77 $Y2=0.56
r89 18 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=1.16
r90 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=1.985
r91 15 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=0.995
+ $X2=1.34 $Y2=1.16
r92 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.34 $Y=0.995
+ $X2=1.34 $Y2=0.56
r93 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r94 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r95 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r96 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r97 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r98 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
r99 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r100 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%C1 3 5 7 10 12 14 17 19 21 24 26 28 29 44
+ 45
r85 44 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.58
+ $Y=1.16 $X2=3.58 $Y2=1.16
r86 42 44 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=3.57 $Y=1.16 $X2=3.58
+ $Y2=1.16
r87 41 42 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.49 $Y=1.16 $X2=3.57
+ $Y2=1.16
r88 40 41 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.14 $Y=1.16
+ $X2=3.49 $Y2=1.16
r89 39 40 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.06 $Y=1.16 $X2=3.14
+ $Y2=1.16
r90 38 39 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=3.06 $Y2=1.16
r91 37 38 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.63 $Y=1.16 $X2=2.71
+ $Y2=1.16
r92 36 37 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=2.28 $Y=1.16
+ $X2=2.63 $Y2=1.16
r93 34 36 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.22 $Y=1.16 $X2=2.28
+ $Y2=1.16
r94 34 35 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.22
+ $Y=1.16 $X2=2.22 $Y2=1.16
r95 31 34 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.2 $Y=1.16 $X2=2.22
+ $Y2=1.16
r96 29 45 47.2276 $w=2.53e-07 $l=1.045e-06 $layer=LI1_cond $X=2.535 $Y=1.147
+ $X2=3.58 $Y2=1.147
r97 29 35 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=2.535 $Y=1.147
+ $X2=2.22 $Y2=1.147
r98 26 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=0.995
+ $X2=3.57 $Y2=1.16
r99 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.57 $Y=0.995
+ $X2=3.57 $Y2=0.56
r100 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.325
+ $X2=3.49 $Y2=1.16
r101 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.49 $Y=1.325
+ $X2=3.49 $Y2=1.985
r102 19 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=0.995
+ $X2=3.14 $Y2=1.16
r103 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.14 $Y=0.995
+ $X2=3.14 $Y2=0.56
r104 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.325
+ $X2=3.06 $Y2=1.16
r105 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.06 $Y=1.325
+ $X2=3.06 $Y2=1.985
r106 12 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=0.995
+ $X2=2.71 $Y2=1.16
r107 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.71 $Y=0.995
+ $X2=2.71 $Y2=0.56
r108 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.325
+ $X2=2.63 $Y2=1.16
r109 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.63 $Y=1.325
+ $X2=2.63 $Y2=1.985
r110 5 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=0.995
+ $X2=2.28 $Y2=1.16
r111 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.28 $Y=0.995
+ $X2=2.28 $Y2=0.56
r112 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.325
+ $X2=2.2 $Y2=1.16
r113 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.2 $Y=1.325 $X2=2.2
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 44
+ 45
r83 43 45 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.48 $Y=1.16
+ $X2=5.73 $Y2=1.16
r84 43 44 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.48
+ $Y=1.16 $X2=5.48 $Y2=1.16
r85 41 43 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.4 $Y=1.16 $X2=5.48
+ $Y2=1.16
r86 40 41 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=5.3 $Y=1.16 $X2=5.4
+ $Y2=1.16
r87 39 40 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.97 $Y=1.16 $X2=5.3
+ $Y2=1.16
r88 38 39 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.87 $Y=1.16 $X2=4.97
+ $Y2=1.16
r89 37 38 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.54 $Y=1.16
+ $X2=4.87 $Y2=1.16
r90 36 37 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.44 $Y=1.16 $X2=4.54
+ $Y2=1.16
r91 34 36 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=4.12 $Y=1.16
+ $X2=4.44 $Y2=1.16
r92 34 35 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.12
+ $Y=1.16 $X2=4.12 $Y2=1.16
r93 31 34 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.11 $Y=1.16 $X2=4.12
+ $Y2=1.16
r94 29 44 49.9392 $w=2.53e-07 $l=1.105e-06 $layer=LI1_cond $X=4.375 $Y=1.147
+ $X2=5.48 $Y2=1.147
r95 29 35 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=4.375 $Y=1.147
+ $X2=4.12 $Y2=1.147
r96 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=1.325
+ $X2=5.73 $Y2=1.16
r97 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.73 $Y=1.325
+ $X2=5.73 $Y2=1.985
r98 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=0.995
+ $X2=5.4 $Y2=1.16
r99 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.4 $Y=0.995 $X2=5.4
+ $Y2=0.56
r100 18 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.3 $Y=1.325
+ $X2=5.3 $Y2=1.16
r101 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.3 $Y=1.325
+ $X2=5.3 $Y2=1.985
r102 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=0.995
+ $X2=4.97 $Y2=1.16
r103 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.97 $Y=0.995
+ $X2=4.97 $Y2=0.56
r104 11 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.87 $Y=1.325
+ $X2=4.87 $Y2=1.16
r105 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.87 $Y=1.325
+ $X2=4.87 $Y2=1.985
r106 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=0.995
+ $X2=4.54 $Y2=1.16
r107 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.54 $Y=0.995
+ $X2=4.54 $Y2=0.56
r108 4 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.44 $Y=1.325
+ $X2=4.44 $Y2=1.16
r109 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.44 $Y=1.325
+ $X2=4.44 $Y2=1.985
r110 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.11 $Y=0.995
+ $X2=4.11 $Y2=1.16
r111 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.11 $Y=0.995
+ $X2=4.11 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 29 44
+ 45
c72 3 0 4.3865e-20 $X=6.17 $Y=1.985
r73 43 45 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=7.55 $Y=1.16
+ $X2=7.67 $Y2=1.16
r74 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.55
+ $Y=1.16 $X2=7.55 $Y2=1.16
r75 41 43 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.48 $Y=1.16 $X2=7.55
+ $Y2=1.16
r76 40 41 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=7.24 $Y=1.16
+ $X2=7.48 $Y2=1.16
r77 39 40 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.03 $Y=1.16
+ $X2=7.24 $Y2=1.16
r78 38 39 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=6.81 $Y=1.16
+ $X2=7.03 $Y2=1.16
r79 37 38 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.6 $Y=1.16 $X2=6.81
+ $Y2=1.16
r80 36 44 46.0977 $w=2.53e-07 $l=1.02e-06 $layer=LI1_cond $X=6.53 $Y=1.147
+ $X2=7.55 $Y2=1.147
r81 35 37 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.53 $Y=1.16 $X2=6.6
+ $Y2=1.16
r82 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.16 $X2=6.53 $Y2=1.16
r83 33 35 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.38 $Y=1.16
+ $X2=6.53 $Y2=1.16
r84 31 33 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.17 $Y=1.16
+ $X2=6.38 $Y2=1.16
r85 29 36 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=6.225 $Y=1.147
+ $X2=6.53 $Y2=1.147
r86 26 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=0.995
+ $X2=7.67 $Y2=1.16
r87 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.67 $Y=0.995
+ $X2=7.67 $Y2=0.56
r88 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.48 $Y=1.325
+ $X2=7.48 $Y2=1.16
r89 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.48 $Y=1.325
+ $X2=7.48 $Y2=1.985
r90 19 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.24 $Y=0.995
+ $X2=7.24 $Y2=1.16
r91 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.24 $Y=0.995
+ $X2=7.24 $Y2=0.56
r92 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.03 $Y=1.325
+ $X2=7.03 $Y2=1.16
r93 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.03 $Y=1.325
+ $X2=7.03 $Y2=1.985
r94 12 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.81 $Y=0.995
+ $X2=6.81 $Y2=1.16
r95 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.81 $Y=0.995
+ $X2=6.81 $Y2=0.56
r96 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.6 $Y=1.325 $X2=6.6
+ $Y2=1.16
r97 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.6 $Y=1.325 $X2=6.6
+ $Y2=1.985
r98 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.38 $Y=0.995
+ $X2=6.38 $Y2=1.16
r99 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.38 $Y=0.995 $X2=6.38
+ $Y2=0.56
r100 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.325
+ $X2=6.17 $Y2=1.16
r101 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.17 $Y=1.325
+ $X2=6.17 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 31
+ 33 40
c70 5 0 9.1669e-20 $X=8.195 $Y=0.995
r71 46 47 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.41 $Y=1.16
+ $X2=9.485 $Y2=1.16
r72 45 46 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=9.055 $Y=1.16
+ $X2=9.41 $Y2=1.16
r73 44 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.98 $Y=1.16
+ $X2=9.055 $Y2=1.16
r74 43 44 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.625 $Y=1.16
+ $X2=8.98 $Y2=1.16
r75 42 43 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.46 $Y=1.16
+ $X2=8.625 $Y2=1.16
r76 41 42 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=8.195 $Y=1.16
+ $X2=8.46 $Y2=1.16
r77 39 41 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.125 $Y=1.16
+ $X2=8.195 $Y2=1.16
r78 39 40 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=8.125
+ $Y=1.16 $X2=8.125 $Y2=1.16
r79 36 39 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=8.03 $Y=1.16
+ $X2=8.125 $Y2=1.16
r80 33 40 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=9.825
+ $Y=1.16 $X2=9.825 $Y2=1.16
r81 31 47 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.56 $Y=1.16
+ $X2=9.485 $Y2=1.16
r82 31 33 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=9.56 $Y=1.16
+ $X2=9.825 $Y2=1.16
r83 29 40 0.180296 $w=2.028e-06 $l=3e-08 $layer=LI1_cond $X=8.975 $Y=1.19
+ $X2=8.975 $Y2=1.16
r84 26 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.485 $Y=0.995
+ $X2=9.485 $Y2=1.16
r85 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.485 $Y=0.995
+ $X2=9.485 $Y2=0.56
r86 22 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.41 $Y=1.325
+ $X2=9.41 $Y2=1.16
r87 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.41 $Y=1.325
+ $X2=9.41 $Y2=1.985
r88 19 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.055 $Y=0.995
+ $X2=9.055 $Y2=1.16
r89 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.055 $Y=0.995
+ $X2=9.055 $Y2=0.56
r90 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.98 $Y=1.325
+ $X2=8.98 $Y2=1.16
r91 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.98 $Y=1.325
+ $X2=8.98 $Y2=1.985
r92 12 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=0.995
+ $X2=8.625 $Y2=1.16
r93 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.625 $Y=0.995
+ $X2=8.625 $Y2=0.56
r94 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.46 $Y=1.325
+ $X2=8.46 $Y2=1.16
r95 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.46 $Y=1.325
+ $X2=8.46 $Y2=1.985
r96 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=0.995
+ $X2=8.195 $Y2=1.16
r97 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.195 $Y=0.995
+ $X2=8.195 $Y2=0.56
r98 1 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.03 $Y=1.325
+ $X2=8.03 $Y2=1.16
r99 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.03 $Y=1.325 $X2=8.03
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%A_28_297# 1 2 3 4 5 16 18 20 24 26 30 32
+ 36 38 40 42 47 49 51
r63 40 53 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=3.74 $Y=2.255
+ $X2=3.74 $Y2=2.35
r64 40 42 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=3.74 $Y=2.255
+ $X2=3.74 $Y2=2
r65 39 51 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.94 $Y=2.35
+ $X2=2.845 $Y2=2.35
r66 38 53 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=3.61 $Y=2.35 $X2=3.74
+ $Y2=2.35
r67 38 39 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=3.61 $Y=2.35 $X2=2.94
+ $Y2=2.35
r68 34 51 1.34256 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.845 $Y=2.255
+ $X2=2.845 $Y2=2.35
r69 34 36 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=2.845 $Y=2.255
+ $X2=2.845 $Y2=2.02
r70 33 49 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.08 $Y=2.35
+ $X2=1.985 $Y2=2.35
r71 32 51 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.75 $Y=2.35
+ $X2=2.845 $Y2=2.35
r72 32 33 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=2.75 $Y=2.35 $X2=2.08
+ $Y2=2.35
r73 28 49 1.34256 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.985 $Y=2.255
+ $X2=1.985 $Y2=2.35
r74 28 30 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.985 $Y=2.255
+ $X2=1.985 $Y2=2.02
r75 27 47 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.22 $Y=2.35
+ $X2=1.125 $Y2=2.35
r76 26 49 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.89 $Y=2.35
+ $X2=1.985 $Y2=2.35
r77 26 27 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.89 $Y=2.35 $X2=1.22
+ $Y2=2.35
r78 22 47 1.34256 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.125 $Y=2.255
+ $X2=1.125 $Y2=2.35
r79 22 24 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.125 $Y=2.255
+ $X2=1.125 $Y2=2.02
r80 21 45 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=0.36 $Y=2.35 $X2=0.23
+ $Y2=2.35
r81 20 47 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.03 $Y=2.35
+ $X2=1.125 $Y2=2.35
r82 20 21 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.03 $Y=2.35 $X2=0.36
+ $Y2=2.35
r83 16 45 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=0.23 $Y=2.255
+ $X2=0.23 $Y2=2.35
r84 16 18 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.23 $Y=2.255
+ $X2=0.23 $Y2=2
r85 5 53 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.485 $X2=3.7 $Y2=2.34
r86 5 42 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.485 $X2=3.7 $Y2=2
r87 4 51 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.485 $X2=2.845 $Y2=2.36
r88 4 36 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.485 $X2=2.845 $Y2=2.02
r89 3 49 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.485 $X2=1.985 $Y2=2.36
r90 3 30 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.485 $X2=1.985 $Y2=2.02
r91 2 47 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.125 $Y2=2.36
r92 2 24 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.125 $Y2=2.02
r93 1 45 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=2.34
r94 1 18 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%Y 1 2 3 4 5 6 7 8 9 10 31 32 35 37 41 43
+ 45 47 53 57 59 64 66 71 76 81 86 90 94 96
c157 53 0 9.1669e-20 $X=7.455 $Y=0.7
r158 94 96 4.11948 $w=1.73e-07 $l=6.5e-08 $layer=LI1_cond $X=0.232 $Y=0.785
+ $X2=0.232 $Y2=0.85
r159 90 94 3.35006 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.232 $Y=0.7
+ $X2=0.232 $Y2=0.785
r160 90 96 0.633766 $w=1.73e-07 $l=1e-08 $layer=LI1_cond $X=0.232 $Y=0.86
+ $X2=0.232 $Y2=0.85
r161 81 83 3.84148 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=4.3 $Y=0.62 $X2=4.3
+ $Y2=0.7
r162 76 78 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.385 $Y=0.62
+ $X2=3.385 $Y2=0.7
r163 71 73 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=2.495 $Y=0.62
+ $X2=2.495 $Y2=0.7
r164 66 68 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=1.555 $Y=0.62
+ $X2=1.555 $Y2=0.7
r165 59 90 17.3683 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.615 $Y=0.7
+ $X2=0.32 $Y2=0.7
r166 55 90 38.9766 $w=1.73e-07 $l=6.15e-07 $layer=LI1_cond $X=0.232 $Y=1.475
+ $X2=0.232 $Y2=0.86
r167 51 53 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=6.595 $Y=0.7
+ $X2=7.455 $Y2=0.7
r168 49 51 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=5.275 $Y=0.7
+ $X2=6.595 $Y2=0.7
r169 48 83 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.42 $Y=0.7 $X2=4.3
+ $Y2=0.7
r170 47 49 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=5.182 $Y=0.7
+ $X2=5.275 $Y2=0.7
r171 47 86 4.79607 $w=1.83e-07 $l=8e-08 $layer=LI1_cond $X=5.182 $Y=0.7
+ $X2=5.182 $Y2=0.62
r172 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.09 $Y=0.7
+ $X2=4.42 $Y2=0.7
r173 46 78 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.51 $Y=0.7
+ $X2=3.385 $Y2=0.7
r174 45 83 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.18 $Y=0.7 $X2=4.3
+ $Y2=0.7
r175 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.18 $Y=0.7
+ $X2=3.51 $Y2=0.7
r176 44 73 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.59 $Y=0.7 $X2=2.495
+ $Y2=0.7
r177 43 78 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.26 $Y=0.7
+ $X2=3.385 $Y2=0.7
r178 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.26 $Y=0.7
+ $X2=2.59 $Y2=0.7
r179 42 68 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.65 $Y=0.7 $X2=1.555
+ $Y2=0.7
r180 41 73 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.4 $Y=0.7 $X2=2.495
+ $Y2=0.7
r181 41 42 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.4 $Y=0.7 $X2=1.65
+ $Y2=0.7
r182 38 57 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.58
+ $X2=0.695 $Y2=1.58
r183 37 64 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.58
+ $X2=1.555 $Y2=1.58
r184 37 38 27.9913 $w=2.08e-07 $l=5.3e-07 $layer=LI1_cond $X=1.39 $Y=1.58
+ $X2=0.86 $Y2=1.58
r185 36 59 0.89264 $w=1.7e-07 $l=1.21589e-07 $layer=LI1_cond $X=0.79 $Y=0.7
+ $X2=0.702 $Y2=0.62
r186 35 68 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.46 $Y=0.7 $X2=1.555
+ $Y2=0.7
r187 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.46 $Y=0.7
+ $X2=0.79 $Y2=0.7
r188 32 55 6.81825 $w=1.8e-07 $l=1.2657e-07 $layer=LI1_cond $X=0.32 $Y=1.565
+ $X2=0.232 $Y2=1.475
r189 31 57 7.80489 $w=1.95e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.53 $Y=1.565
+ $X2=0.695 $Y2=1.58
r190 31 32 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.53 $Y=1.565
+ $X2=0.32 $Y2=1.565
r191 10 64 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.485 $X2=1.555 $Y2=1.655
r192 9 57 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.695 $Y2=1.64
r193 8 53 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=7.315
+ $Y=0.235 $X2=7.455 $Y2=0.7
r194 7 51 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=6.455
+ $Y=0.235 $X2=6.595 $Y2=0.7
r195 6 86 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.185 $Y2=0.62
r196 5 81 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=4.185
+ $Y=0.235 $X2=4.325 $Y2=0.62
r197 4 76 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.235 $X2=3.355 $Y2=0.62
r198 3 71 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.495 $Y2=0.62
r199 2 66 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.62
r200 1 59 182 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%A_455_297# 1 2 3 4 15 19 23 28 30 32 34
c70 34 0 4.3865e-20 $X=5.515 $Y=1.655
r71 24 32 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=1.58
+ $X2=4.655 $Y2=1.58
r72 23 34 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=1.58
+ $X2=5.515 $Y2=1.58
r73 23 24 27.9913 $w=2.08e-07 $l=5.3e-07 $layer=LI1_cond $X=5.35 $Y=1.58
+ $X2=4.82 $Y2=1.58
r74 20 30 7.80489 $w=1.95e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.44 $Y=1.565
+ $X2=3.275 $Y2=1.58
r75 19 32 7.80489 $w=1.95e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.49 $Y=1.565
+ $X2=4.655 $Y2=1.58
r76 19 20 64.697 $w=1.78e-07 $l=1.05e-06 $layer=LI1_cond $X=4.49 $Y=1.565
+ $X2=3.44 $Y2=1.565
r77 16 28 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=1.58
+ $X2=2.415 $Y2=1.58
r78 15 30 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=1.58
+ $X2=3.275 $Y2=1.58
r79 15 16 27.9913 $w=2.08e-07 $l=5.3e-07 $layer=LI1_cond $X=3.11 $Y=1.58
+ $X2=2.58 $Y2=1.58
r80 4 34 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=5.375
+ $Y=1.485 $X2=5.515 $Y2=1.655
r81 3 32 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=4.515
+ $Y=1.485 $X2=4.655 $Y2=1.655
r82 2 30 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=3.135
+ $Y=1.485 $X2=3.275 $Y2=1.655
r83 1 28 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.485 $X2=2.415 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%A_821_297# 1 2 3 4 5 6 7 22 24 26 30 32 38
+ 39 42 44 48 52 54 58 63 64 66 67
r88 56 58 2.64102 $w=2.38e-07 $l=5.5e-08 $layer=LI1_cond $X=9.65 $Y=1.67
+ $X2=9.65 $Y2=1.725
r89 55 67 5.8691 $w=2.22e-07 $l=1.3e-07 $layer=LI1_cond $X=8.84 $Y=1.557
+ $X2=8.71 $Y2=1.557
r90 54 56 6.82572 $w=2.25e-07 $l=1.67212e-07 $layer=LI1_cond $X=9.53 $Y=1.557
+ $X2=9.65 $Y2=1.67
r91 54 55 35.3416 $w=2.23e-07 $l=6.9e-07 $layer=LI1_cond $X=9.53 $Y=1.557
+ $X2=8.84 $Y2=1.557
r92 50 67 0.788168 $w=2.6e-07 $l=1.13e-07 $layer=LI1_cond $X=8.71 $Y=1.67
+ $X2=8.71 $Y2=1.557
r93 50 52 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=8.71 $Y=1.67
+ $X2=8.71 $Y2=1.725
r94 49 66 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=7.91 $Y=1.555
+ $X2=7.745 $Y2=1.555
r95 48 67 5.8691 $w=2.22e-07 $l=1.30996e-07 $layer=LI1_cond $X=8.58 $Y=1.555
+ $X2=8.71 $Y2=1.557
r96 48 49 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=8.58 $Y=1.555
+ $X2=7.91 $Y2=1.555
r97 45 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.91 $Y=1.53
+ $X2=6.815 $Y2=1.53
r98 44 66 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=7.58 $Y=1.53
+ $X2=7.745 $Y2=1.555
r99 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.58 $Y=1.53
+ $X2=6.91 $Y2=1.53
r100 40 64 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=1.615
+ $X2=6.815 $Y2=1.53
r101 40 42 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=6.815 $Y=1.615
+ $X2=6.815 $Y2=1.63
r102 38 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.72 $Y=1.53
+ $X2=6.815 $Y2=1.53
r103 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.72 $Y=1.53
+ $X2=6.05 $Y2=1.53
r104 35 37 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=5.955 $Y=2.275
+ $X2=5.955 $Y2=1.63
r105 34 39 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.955 $Y=1.615
+ $X2=6.05 $Y2=1.53
r106 34 37 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=5.955 $Y=1.615
+ $X2=5.955 $Y2=1.63
r107 33 63 5.40251 $w=1.8e-07 $l=9.98749e-08 $layer=LI1_cond $X=5.18 $Y=2.36
+ $X2=5.085 $Y2=2.35
r108 32 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.86 $Y=2.36
+ $X2=5.955 $Y2=2.275
r109 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.86 $Y=2.36
+ $X2=5.18 $Y2=2.36
r110 28 63 1.14861 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=5.085 $Y=2.255
+ $X2=5.085 $Y2=2.35
r111 28 30 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=5.085 $Y=2.255
+ $X2=5.085 $Y2=2.02
r112 27 61 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=4.32 $Y=2.35
+ $X2=4.19 $Y2=2.35
r113 26 63 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.99 $Y=2.35
+ $X2=5.085 $Y2=2.35
r114 26 27 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=4.99 $Y=2.35 $X2=4.32
+ $Y2=2.35
r115 22 61 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=4.19 $Y=2.255
+ $X2=4.19 $Y2=2.35
r116 22 24 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=4.19 $Y=2.255
+ $X2=4.19 $Y2=2
r117 7 58 300 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=2 $X=9.485
+ $Y=1.485 $X2=9.625 $Y2=1.725
r118 6 52 300 $w=1.7e-07 $l=3.15595e-07 $layer=licon1_PDIFF $count=2 $X=8.535
+ $Y=1.485 $X2=8.71 $Y2=1.725
r119 5 66 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.555
+ $Y=1.485 $X2=7.695 $Y2=1.63
r120 4 42 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.675
+ $Y=1.485 $X2=6.815 $Y2=1.63
r121 3 37 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.485 $X2=5.955 $Y2=1.63
r122 2 63 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.485 $X2=5.085 $Y2=2.36
r123 2 30 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.485 $X2=5.085 $Y2=2.02
r124 1 61 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.485 $X2=4.23 $Y2=2.34
r125 1 24 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.485 $X2=4.23 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%VPWR 1 2 3 4 15 17 21 25 29 31 32 34 35 37
+ 38 39 56 57 60
r131 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r132 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r133 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r134 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r135 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r136 51 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.13 $Y2=2.72
r137 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r138 48 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=2.72
+ $X2=7.245 $Y2=2.72
r139 48 50 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=7.41 $Y=2.72
+ $X2=8.05 $Y2=2.72
r140 47 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r141 46 47 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r142 42 46 390.139 $w=1.68e-07 $l=5.98e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=6.21 $Y2=2.72
r143 39 47 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=6.21 $Y2=2.72
r144 39 42 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 37 53 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=9.03 $Y=2.72 $X2=8.97
+ $Y2=2.72
r146 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.03 $Y=2.72
+ $X2=9.195 $Y2=2.72
r147 36 56 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=9.36 $Y=2.72
+ $X2=9.89 $Y2=2.72
r148 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.36 $Y=2.72
+ $X2=9.195 $Y2=2.72
r149 34 50 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=8.08 $Y=2.72 $X2=8.05
+ $Y2=2.72
r150 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.08 $Y=2.72
+ $X2=8.245 $Y2=2.72
r151 33 53 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.41 $Y=2.72
+ $X2=8.97 $Y2=2.72
r152 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.41 $Y=2.72
+ $X2=8.245 $Y2=2.72
r153 31 46 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.22 $Y=2.72
+ $X2=6.21 $Y2=2.72
r154 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.22 $Y=2.72
+ $X2=6.385 $Y2=2.72
r155 27 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.195 $Y=2.635
+ $X2=9.195 $Y2=2.72
r156 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=9.195 $Y=2.635
+ $X2=9.195 $Y2=2
r157 23 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.245 $Y=2.635
+ $X2=8.245 $Y2=2.72
r158 23 25 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=8.245 $Y=2.635
+ $X2=8.245 $Y2=1.98
r159 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.245 $Y=2.635
+ $X2=7.245 $Y2=2.72
r160 19 21 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=7.245 $Y=2.635
+ $X2=7.245 $Y2=1.89
r161 18 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.55 $Y=2.72
+ $X2=6.385 $Y2=2.72
r162 17 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.08 $Y=2.72
+ $X2=7.245 $Y2=2.72
r163 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.08 $Y=2.72
+ $X2=6.55 $Y2=2.72
r164 13 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=2.635
+ $X2=6.385 $Y2=2.72
r165 13 15 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=6.385 $Y=2.635
+ $X2=6.385 $Y2=1.89
r166 4 29 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=9.055
+ $Y=1.485 $X2=9.195 $Y2=2
r167 3 25 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=8.105
+ $Y=1.485 $X2=8.245 $Y2=1.98
r168 2 21 300 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=2 $X=7.105
+ $Y=1.485 $X2=7.245 $Y2=1.89
r169 1 15 300 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=2 $X=6.245
+ $Y=1.485 $X2=6.385 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46
+ 50 54 58 61 62 64 65 66 68 73 78 83 88 93 106 107 113 117 123 126 129 132 136
r175 132 133 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r176 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r177 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r178 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r179 117 120 10.119 $w=4.08e-07 $l=3.6e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.025 $Y2=0.36
r180 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r181 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r182 110 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r183 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r184 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r185 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r186 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r187 101 133 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=5.75 $Y2=0
r188 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r189 98 132 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=5.78 $Y=0
+ $X2=5.612 $Y2=0
r190 98 100 148.096 $w=1.68e-07 $l=2.27e-06 $layer=LI1_cond $X=5.78 $Y=0
+ $X2=8.05 $Y2=0
r191 97 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r192 97 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r193 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r194 94 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=0
+ $X2=4.755 $Y2=0
r195 94 96 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=5.29
+ $Y2=0
r196 93 132 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=5.445 $Y=0
+ $X2=5.612 $Y2=0
r197 93 96 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.445 $Y=0
+ $X2=5.29 $Y2=0
r198 92 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r199 92 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r200 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r201 89 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=0
+ $X2=3.845 $Y2=0
r202 89 91 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.01 $Y=0 $X2=4.37
+ $Y2=0
r203 88 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=0
+ $X2=4.755 $Y2=0
r204 88 91 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.59 $Y=0 $X2=4.37
+ $Y2=0
r205 87 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r206 87 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.99 $Y2=0
r207 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r208 84 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=0
+ $X2=2.925 $Y2=0
r209 84 86 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=3.45
+ $Y2=0
r210 83 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.68 $Y=0
+ $X2=3.845 $Y2=0
r211 83 86 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.68 $Y=0 $X2=3.45
+ $Y2=0
r212 82 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.99 $Y2=0
r213 82 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r214 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r215 79 117 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.23 $Y=0
+ $X2=2.025 $Y2=0
r216 79 81 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.23 $Y=0 $X2=2.53
+ $Y2=0
r217 78 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=0
+ $X2=2.925 $Y2=0
r218 78 81 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.53
+ $Y2=0
r219 77 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r220 77 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r221 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r222 74 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0
+ $X2=1.125 $Y2=0
r223 74 76 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.61
+ $Y2=0
r224 73 117 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.82 $Y=0
+ $X2=2.025 $Y2=0
r225 73 76 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.61
+ $Y2=0
r226 72 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r227 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r228 69 110 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r229 69 71 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.69
+ $Y2=0
r230 68 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0
+ $X2=1.125 $Y2=0
r231 68 71 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.69
+ $Y2=0
r232 66 72 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r233 66 136 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r234 64 103 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.105 $Y=0
+ $X2=8.97 $Y2=0
r235 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=0 $X2=9.27
+ $Y2=0
r236 63 106 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=9.435 $Y=0
+ $X2=9.89 $Y2=0
r237 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=0 $X2=9.27
+ $Y2=0
r238 61 100 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.245 $Y=0
+ $X2=8.05 $Y2=0
r239 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=8.41
+ $Y2=0
r240 60 103 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.575 $Y=0
+ $X2=8.97 $Y2=0
r241 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.575 $Y=0 $X2=8.41
+ $Y2=0
r242 56 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.27 $Y=0.085
+ $X2=9.27 $Y2=0
r243 56 58 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.27 $Y=0.085
+ $X2=9.27 $Y2=0.36
r244 52 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0
r245 52 54 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0.36
r246 48 132 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.612 $Y=0.085
+ $X2=5.612 $Y2=0
r247 48 50 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=5.612 $Y=0.085
+ $X2=5.612 $Y2=0.36
r248 44 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=0.085
+ $X2=4.755 $Y2=0
r249 44 46 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.755 $Y=0.085
+ $X2=4.755 $Y2=0.36
r250 40 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=0.085
+ $X2=3.845 $Y2=0
r251 40 42 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.845 $Y=0.085
+ $X2=3.845 $Y2=0.36
r252 36 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.085
+ $X2=2.925 $Y2=0
r253 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.925 $Y=0.085
+ $X2=2.925 $Y2=0.36
r254 32 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0
r255 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0.36
r256 28 110 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r257 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.36
r258 9 58 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=9.13
+ $Y=0.235 $X2=9.27 $Y2=0.36
r259 8 54 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.235 $X2=8.41 $Y2=0.36
r260 7 50 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.475
+ $Y=0.235 $X2=5.61 $Y2=0.36
r261 6 46 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.235 $X2=4.755 $Y2=0.36
r262 5 42 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.235 $X2=3.845 $Y2=0.36
r263 4 38 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.235 $X2=2.925 $Y2=0.36
r264 3 120 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=2.065 $Y2=0.36
r265 2 34 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.125 $Y2=0.36
r266 1 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_4%A_1205_47# 1 2 3 4 5 16 25 26 27 30 32 36
+ 38
r53 34 36 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=9.735 $Y=0.615
+ $X2=9.735 $Y2=0.51
r54 33 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.935 $Y=0.7 $X2=8.84
+ $Y2=0.7
r55 32 34 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.605 $Y=0.7
+ $X2=9.735 $Y2=0.615
r56 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.605 $Y=0.7
+ $X2=8.935 $Y2=0.7
r57 28 38 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.84 $Y=0.615
+ $X2=8.84 $Y2=0.7
r58 28 30 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=8.84 $Y=0.615
+ $X2=8.84 $Y2=0.51
r59 26 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.745 $Y=0.7 $X2=8.84
+ $Y2=0.7
r60 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.745 $Y=0.7
+ $X2=8.075 $Y2=0.7
r61 23 27 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.98 $Y=0.615
+ $X2=8.075 $Y2=0.7
r62 23 25 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=7.98 $Y=0.615
+ $X2=7.98 $Y2=0.51
r63 22 25 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=7.98 $Y=0.445
+ $X2=7.98 $Y2=0.51
r64 18 21 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=6.17 $Y=0.36
+ $X2=7.025 $Y2=0.36
r65 16 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.885 $Y=0.36
+ $X2=7.98 $Y2=0.445
r66 16 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=7.885 $Y=0.36
+ $X2=7.025 $Y2=0.36
r67 5 36 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.56
+ $Y=0.235 $X2=9.7 $Y2=0.51
r68 4 30 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=8.7
+ $Y=0.235 $X2=8.84 $Y2=0.51
r69 3 25 182 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_NDIFF $count=1 $X=7.745
+ $Y=0.235 $X2=7.975 $Y2=0.51
r70 2 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=6.885
+ $Y=0.235 $X2=7.025 $Y2=0.36
r71 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.025
+ $Y=0.235 $X2=6.17 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__xor2_4.spice.SKY130_FD_SC_HD__XOR2_4.pxi
* Created: Thu Aug 27 14:49:57 2020
* 
x_PM_SKY130_FD_SC_HD__XOR2_4%A N_A_c_161_n N_A_M1012_g N_A_M1004_g N_A_c_162_n
+ N_A_M1017_g N_A_M1018_g N_A_c_163_n N_A_M1028_g N_A_M1025_g N_A_c_164_n
+ N_A_M1030_g N_A_M1038_g N_A_c_165_n N_A_M1005_g N_A_M1009_g N_A_c_166_n
+ N_A_M1011_g N_A_M1019_g N_A_c_167_n N_A_M1015_g N_A_M1033_g N_A_c_168_n
+ N_A_M1023_g N_A_M1039_g N_A_c_180_n N_A_c_181_n N_A_c_188_p N_A_c_182_n
+ N_A_c_206_p N_A_c_237_p N_A_c_169_n A N_A_c_170_n N_A_c_171_n
+ PM_SKY130_FD_SC_HD__XOR2_4%A
x_PM_SKY130_FD_SC_HD__XOR2_4%B N_B_c_390_n N_B_M1021_g N_B_M1003_g N_B_c_391_n
+ N_B_M1029_g N_B_M1006_g N_B_c_392_n N_B_M1034_g N_B_M1007_g N_B_c_393_n
+ N_B_M1036_g N_B_M1026_g N_B_c_394_n N_B_c_395_n N_B_c_396_n N_B_M1010_g
+ N_B_M1000_g N_B_c_397_n N_B_M1013_g N_B_M1002_g N_B_c_398_n N_B_M1014_g
+ N_B_M1008_g N_B_c_399_n N_B_M1020_g N_B_M1027_g B N_B_c_400_n N_B_c_401_n
+ PM_SKY130_FD_SC_HD__XOR2_4%B
x_PM_SKY130_FD_SC_HD__XOR2_4%A_112_47# N_A_112_47#_M1012_d N_A_112_47#_M1028_d
+ N_A_112_47#_M1021_s N_A_112_47#_M1034_s N_A_112_47#_M1003_s
+ N_A_112_47#_M1007_s N_A_112_47#_c_544_n N_A_112_47#_M1024_g
+ N_A_112_47#_M1001_g N_A_112_47#_c_545_n N_A_112_47#_M1031_g
+ N_A_112_47#_M1016_g N_A_112_47#_c_546_n N_A_112_47#_M1032_g
+ N_A_112_47#_M1022_g N_A_112_47#_c_547_n N_A_112_47#_M1037_g
+ N_A_112_47#_M1035_g N_A_112_47#_c_548_n N_A_112_47#_c_549_n
+ N_A_112_47#_c_550_n N_A_112_47#_c_579_n N_A_112_47#_c_551_n
+ N_A_112_47#_c_586_n N_A_112_47#_c_552_n N_A_112_47#_c_591_n
+ N_A_112_47#_c_592_n N_A_112_47#_c_553_n N_A_112_47#_c_646_n
+ N_A_112_47#_c_554_n N_A_112_47#_c_555_n N_A_112_47#_c_728_p
+ N_A_112_47#_c_732_p N_A_112_47#_c_567_n N_A_112_47#_c_556_n
+ N_A_112_47#_c_557_n N_A_112_47#_c_558_n N_A_112_47#_c_568_n
+ N_A_112_47#_c_616_n N_A_112_47#_c_655_n N_A_112_47#_c_617_n
+ N_A_112_47#_c_559_n N_A_112_47#_c_569_n N_A_112_47#_c_570_n
+ N_A_112_47#_c_571_n N_A_112_47#_c_572_n N_A_112_47#_c_560_n
+ PM_SKY130_FD_SC_HD__XOR2_4%A_112_47#
x_PM_SKY130_FD_SC_HD__XOR2_4%A_27_297# N_A_27_297#_M1004_s N_A_27_297#_M1018_s
+ N_A_27_297#_M1038_s N_A_27_297#_M1006_d N_A_27_297#_M1026_d
+ N_A_27_297#_c_820_n N_A_27_297#_c_822_n N_A_27_297#_c_837_n
+ N_A_27_297#_c_825_n N_A_27_297#_c_856_p N_A_27_297#_c_815_n
+ N_A_27_297#_c_824_n N_A_27_297#_c_816_n N_A_27_297#_c_848_n
+ N_A_27_297#_c_849_n PM_SKY130_FD_SC_HD__XOR2_4%A_27_297#
x_PM_SKY130_FD_SC_HD__XOR2_4%VPWR N_VPWR_M1004_d N_VPWR_M1025_d N_VPWR_M1000_s
+ N_VPWR_M1008_s N_VPWR_M1009_s N_VPWR_M1033_s N_VPWR_c_880_n N_VPWR_c_881_n
+ N_VPWR_c_882_n N_VPWR_c_883_n N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n
+ N_VPWR_c_887_n N_VPWR_c_888_n N_VPWR_c_889_n VPWR N_VPWR_c_890_n
+ N_VPWR_c_891_n N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_879_n N_VPWR_c_895_n
+ N_VPWR_c_896_n N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_899_n
+ PM_SKY130_FD_SC_HD__XOR2_4%VPWR
x_PM_SKY130_FD_SC_HD__XOR2_4%A_806_297# N_A_806_297#_M1000_d
+ N_A_806_297#_M1002_d N_A_806_297#_M1027_d N_A_806_297#_M1019_d
+ N_A_806_297#_M1039_d N_A_806_297#_M1001_s N_A_806_297#_M1022_s
+ N_A_806_297#_c_1043_n N_A_806_297#_c_1044_n N_A_806_297#_c_1045_n
+ N_A_806_297#_c_1036_n N_A_806_297#_c_1055_n N_A_806_297#_c_1037_n
+ N_A_806_297#_c_1080_n N_A_806_297#_c_1038_n N_A_806_297#_c_1118_n
+ N_A_806_297#_c_1139_p N_A_806_297#_c_1082_n N_A_806_297#_c_1143_p
+ N_A_806_297#_c_1039_n N_A_806_297#_c_1060_n N_A_806_297#_c_1061_n
+ N_A_806_297#_c_1128_n N_A_806_297#_c_1130_n
+ PM_SKY130_FD_SC_HD__XOR2_4%A_806_297#
x_PM_SKY130_FD_SC_HD__XOR2_4%X N_X_M1010_s N_X_M1014_s N_X_M1024_s N_X_M1032_s
+ N_X_M1001_d N_X_M1016_d N_X_M1035_d N_X_c_1156_n N_X_c_1157_n N_X_c_1158_n
+ N_X_c_1203_n N_X_c_1145_n N_X_c_1159_n N_X_c_1214_n N_X_c_1146_n N_X_c_1147_n
+ N_X_c_1148_n N_X_c_1149_n N_X_c_1161_n N_X_c_1150_n N_X_c_1162_n X
+ N_X_c_1151_n N_X_c_1152_n N_X_c_1153_n N_X_c_1154_n N_X_c_1155_n
+ PM_SKY130_FD_SC_HD__XOR2_4%X
x_PM_SKY130_FD_SC_HD__XOR2_4%VGND N_VGND_M1012_s N_VGND_M1017_s N_VGND_M1030_s
+ N_VGND_M1029_d N_VGND_M1036_d N_VGND_M1005_d N_VGND_M1015_d N_VGND_M1024_d
+ N_VGND_M1031_d N_VGND_M1037_d N_VGND_c_1307_n N_VGND_c_1308_n N_VGND_c_1309_n
+ N_VGND_c_1310_n N_VGND_c_1311_n N_VGND_c_1312_n N_VGND_c_1313_n
+ N_VGND_c_1314_n N_VGND_c_1315_n N_VGND_c_1316_n N_VGND_c_1317_n
+ N_VGND_c_1318_n N_VGND_c_1319_n N_VGND_c_1320_n N_VGND_c_1321_n
+ N_VGND_c_1322_n N_VGND_c_1323_n N_VGND_c_1324_n N_VGND_c_1325_n
+ N_VGND_c_1326_n N_VGND_c_1327_n N_VGND_c_1328_n N_VGND_c_1329_n
+ N_VGND_c_1330_n N_VGND_c_1331_n N_VGND_c_1332_n N_VGND_c_1333_n VGND
+ N_VGND_c_1334_n N_VGND_c_1335_n N_VGND_c_1336_n N_VGND_c_1337_n
+ PM_SKY130_FD_SC_HD__XOR2_4%VGND
x_PM_SKY130_FD_SC_HD__XOR2_4%A_806_47# N_A_806_47#_M1010_d N_A_806_47#_M1013_d
+ N_A_806_47#_M1020_d N_A_806_47#_M1011_s N_A_806_47#_M1023_s
+ N_A_806_47#_c_1488_n N_A_806_47#_c_1494_n N_A_806_47#_c_1489_n
+ N_A_806_47#_c_1490_n N_A_806_47#_c_1504_n N_A_806_47#_c_1491_n
+ N_A_806_47#_c_1492_n N_A_806_47#_c_1493_n PM_SKY130_FD_SC_HD__XOR2_4%A_806_47#
cc_1 VNB N_A_c_161_n 0.0192198f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_A_c_162_n 0.0157984f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_A_c_163_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=0.995
cc_4 VNB N_A_c_164_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=0.995
cc_5 VNB N_A_c_165_n 0.0158649f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=0.995
cc_6 VNB N_A_c_166_n 0.0156747f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=0.995
cc_7 VNB N_A_c_167_n 0.0156747f $X=-0.19 $Y=-0.24 $X2=6.885 $Y2=0.995
cc_8 VNB N_A_c_168_n 0.0205818f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=0.995
cc_9 VNB N_A_c_169_n 0.00467216f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=1.175
cc_10 VNB N_A_c_170_n 0.0654734f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=1.16
cc_11 VNB N_A_c_171_n 0.0700147f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=1.16
cc_12 VNB N_B_c_390_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_13 VNB N_B_c_391_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_14 VNB N_B_c_392_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=0.995
cc_15 VNB N_B_c_393_n 0.0214817f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=0.995
cc_16 VNB N_B_c_394_n 0.0462482f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=0.995
cc_17 VNB N_B_c_395_n 0.0574269f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=0.56
cc_18 VNB N_B_c_396_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=0.56
cc_19 VNB N_B_c_397_n 0.0157834f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=0.56
cc_20 VNB N_B_c_398_n 0.0155532f $X=-0.19 $Y=-0.24 $X2=6.885 $Y2=0.56
cc_21 VNB N_B_c_399_n 0.0158403f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=0.56
cc_22 VNB N_B_c_400_n 0.00199483f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_23 VNB N_B_c_401_n 0.0575844f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_24 VNB N_A_112_47#_c_544_n 0.020524f $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=1.985
cc_25 VNB N_A_112_47#_c_545_n 0.0157963f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=1.985
cc_26 VNB N_A_112_47#_c_546_n 0.0157983f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=1.985
cc_27 VNB N_A_112_47#_c_547_n 0.0192096f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=1.985
cc_28 VNB N_A_112_47#_c_548_n 0.0190232f $X=-0.19 $Y=-0.24 $X2=6.885 $Y2=1.985
cc_29 VNB N_A_112_47#_c_549_n 0.00203902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_112_47#_c_550_n 0.00773467f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=0.995
cc_31 VNB N_A_112_47#_c_551_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=1.985
cc_32 VNB N_A_112_47#_c_552_n 0.00238002f $X=-0.19 $Y=-0.24 $X2=6.08 $Y2=1.275
cc_33 VNB N_A_112_47#_c_553_n 0.00470005f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=1.175
cc_34 VNB N_A_112_47#_c_554_n 7.98352e-19 $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=1.16
cc_35 VNB N_A_112_47#_c_555_n 0.00353971f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.16
cc_36 VNB N_A_112_47#_c_556_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=1.16
cc_37 VNB N_A_112_47#_c_557_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_112_47#_c_558_n 0.00209731f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.175
cc_39 VNB N_A_112_47#_c_559_n 0.0137744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_112_47#_c_560_n 0.0725826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_879_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_42 VNB N_X_c_1145_n 0.00217862f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=0.995
cc_43 VNB N_X_c_1146_n 0.0124013f $X=-0.19 $Y=-0.24 $X2=6.885 $Y2=1.325
cc_44 VNB N_X_c_1147_n 0.0219841f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_1148_n 0.00434087f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=0.56
cc_46 VNB N_X_c_1149_n 0.00231911f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=1.325
cc_47 VNB N_X_c_1150_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_1151_n 0.0112778f $X=-0.19 $Y=-0.24 $X2=6.08 $Y2=1.445
cc_49 VNB N_X_c_1152_n 0.00123766f $X=-0.19 $Y=-0.24 $X2=6.165 $Y2=1.175
cc_50 VNB N_X_c_1153_n 0.00144825f $X=-0.19 $Y=-0.24 $X2=6.17 $Y2=1.16
cc_51 VNB N_X_c_1154_n 0.00243579f $X=-0.19 $Y=-0.24 $X2=7.19 $Y2=1.16
cc_52 VNB N_X_c_1155_n 0.00542965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1307_n 0.0101714f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=0.56
cc_54 VNB N_VGND_c_1308_n 0.0177171f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=1.985
cc_55 VNB N_VGND_c_1309_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=0.56
cc_56 VNB N_VGND_c_1310_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=1.985
cc_57 VNB N_VGND_c_1311_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=6.885 $Y2=0.56
cc_58 VNB N_VGND_c_1312_n 0.014329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1313_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=7.305 $Y2=1.325
cc_60 VNB N_VGND_c_1314_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=2.715 $Y2=1.275
cc_61 VNB N_VGND_c_1315_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=6.08 $Y2=1.275
cc_62 VNB N_VGND_c_1316_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=6.17 $Y2=1.16
cc_63 VNB N_VGND_c_1317_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=7.19 $Y2=1.16
cc_64 VNB N_VGND_c_1318_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_65 VNB N_VGND_c_1319_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1320_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1321_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_68 VNB N_VGND_c_1322_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_69 VNB N_VGND_c_1323_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_70 VNB N_VGND_c_1324_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.16
cc_71 VNB N_VGND_c_1325_n 0.00519006f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.16
cc_72 VNB N_VGND_c_1326_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=1.16
cc_73 VNB N_VGND_c_1327_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1328_n 0.0205009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1329_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=6.17 $Y2=1.16
cc_76 VNB N_VGND_c_1330_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=6.885 $Y2=1.16
cc_77 VNB N_VGND_c_1331_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=7.19 $Y2=1.16
cc_78 VNB N_VGND_c_1332_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1333_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.175
cc_80 VNB N_VGND_c_1334_n 0.0545905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1335_n 0.0111912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1336_n 0.477585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1337_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_806_47#_c_1488_n 0.00266706f $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=0.56
cc_85 VNB N_A_806_47#_c_1489_n 0.00191802f $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=0.56
cc_86 VNB N_A_806_47#_c_1490_n 9.214e-19 $X=-0.19 $Y=-0.24 $X2=1.745 $Y2=0.56
cc_87 VNB N_A_806_47#_c_1491_n 0.00388751f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=0.56
cc_88 VNB N_A_806_47#_c_1492_n 0.00554991f $X=-0.19 $Y=-0.24 $X2=6.045 $Y2=1.985
cc_89 VNB N_A_806_47#_c_1493_n 9.22322e-19 $X=-0.19 $Y=-0.24 $X2=6.465 $Y2=1.985
cc_90 VPB N_A_M1004_g 0.022025f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_91 VPB N_A_M1018_g 0.0181185f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_92 VPB N_A_M1025_g 0.018138f $X=-0.19 $Y=1.305 $X2=1.325 $Y2=1.985
cc_93 VPB N_A_M1038_g 0.0184041f $X=-0.19 $Y=1.305 $X2=1.745 $Y2=1.985
cc_94 VPB N_A_M1009_g 0.0178886f $X=-0.19 $Y=1.305 $X2=6.045 $Y2=1.985
cc_95 VPB N_A_M1019_g 0.0182783f $X=-0.19 $Y=1.305 $X2=6.465 $Y2=1.985
cc_96 VPB N_A_M1033_g 0.0182798f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=1.985
cc_97 VPB N_A_M1039_g 0.0221099f $X=-0.19 $Y=1.305 $X2=7.305 $Y2=1.985
cc_98 VPB N_A_c_180_n 0.00111437f $X=-0.19 $Y=1.305 $X2=2.715 $Y2=1.445
cc_99 VPB N_A_c_181_n 0.0303803f $X=-0.19 $Y=1.305 $X2=5.995 $Y2=1.53
cc_100 VPB N_A_c_182_n 0.00118978f $X=-0.19 $Y=1.305 $X2=6.08 $Y2=1.445
cc_101 VPB N_A_c_170_n 0.0102666f $X=-0.19 $Y=1.305 $X2=1.745 $Y2=1.16
cc_102 VPB N_A_c_171_n 0.0113889f $X=-0.19 $Y=1.305 $X2=7.305 $Y2=1.16
cc_103 VPB N_B_M1003_g 0.0182124f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_104 VPB N_B_M1006_g 0.0177057f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_105 VPB N_B_M1007_g 0.0180908f $X=-0.19 $Y=1.305 $X2=1.325 $Y2=1.985
cc_106 VPB N_B_M1026_g 0.025024f $X=-0.19 $Y=1.305 $X2=1.745 $Y2=1.985
cc_107 VPB N_B_c_394_n 0.0160453f $X=-0.19 $Y=1.305 $X2=6.045 $Y2=0.995
cc_108 VPB N_B_c_395_n 0.0099693f $X=-0.19 $Y=1.305 $X2=6.045 $Y2=0.56
cc_109 VPB N_B_M1000_g 0.025044f $X=-0.19 $Y=1.305 $X2=6.465 $Y2=0.995
cc_110 VPB N_B_M1002_g 0.018138f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=0.995
cc_111 VPB N_B_M1008_g 0.018138f $X=-0.19 $Y=1.305 $X2=7.305 $Y2=0.995
cc_112 VPB N_B_M1027_g 0.0183686f $X=-0.19 $Y=1.305 $X2=2.715 $Y2=1.275
cc_113 VPB N_B_c_401_n 0.00974451f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_114 VPB N_A_112_47#_M1001_g 0.0226826f $X=-0.19 $Y=1.305 $X2=1.745 $Y2=0.56
cc_115 VPB N_A_112_47#_M1016_g 0.018138f $X=-0.19 $Y=1.305 $X2=6.045 $Y2=0.56
cc_116 VPB N_A_112_47#_M1022_g 0.0181184f $X=-0.19 $Y=1.305 $X2=6.465 $Y2=0.56
cc_117 VPB N_A_112_47#_M1035_g 0.0220113f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=0.56
cc_118 VPB N_A_112_47#_c_548_n 0.00683654f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=1.985
cc_119 VPB N_A_112_47#_c_554_n 0.00603241f $X=-0.19 $Y=1.305 $X2=1.325 $Y2=1.16
cc_120 VPB N_A_112_47#_c_567_n 0.00783783f $X=-0.19 $Y=1.305 $X2=7.19 $Y2=1.16
cc_121 VPB N_A_112_47#_c_568_n 0.0116758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_112_47#_c_569_n 0.00341908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_112_47#_c_570_n 0.0016129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_112_47#_c_571_n 0.00685751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_112_47#_c_572_n 0.00165362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_112_47#_c_560_n 0.0105189f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_297#_c_815_n 0.00148118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_297#_c_816_n 0.0280239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_880_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_881_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.745 $Y2=1.325
cc_131 VPB N_VPWR_c_882_n 0.00454762f $X=-0.19 $Y=1.305 $X2=6.045 $Y2=0.995
cc_132 VPB N_VPWR_c_883_n 0.0150723f $X=-0.19 $Y=1.305 $X2=6.045 $Y2=0.56
cc_133 VPB N_VPWR_c_884_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_885_n 0.0150723f $X=-0.19 $Y=1.305 $X2=6.465 $Y2=0.56
cc_135 VPB N_VPWR_c_886_n 0.00393015f $X=-0.19 $Y=1.305 $X2=6.465 $Y2=1.985
cc_136 VPB N_VPWR_c_887_n 0.00454762f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=0.56
cc_137 VPB N_VPWR_c_888_n 0.0664284f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=1.985
cc_138 VPB N_VPWR_c_889_n 0.00478085f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=1.985
cc_139 VPB N_VPWR_c_890_n 0.0166842f $X=-0.19 $Y=1.305 $X2=7.305 $Y2=0.56
cc_140 VPB N_VPWR_c_891_n 0.0150723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_892_n 0.0150723f $X=-0.19 $Y=1.305 $X2=6.17 $Y2=1.16
cc_142 VPB N_VPWR_c_893_n 0.0701463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_879_n 0.0594487f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_144 VPB N_VPWR_c_895_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_145 VPB N_VPWR_c_896_n 0.00478085f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.16
cc_146 VPB N_VPWR_c_897_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_898_n 0.00478085f $X=-0.19 $Y=1.305 $X2=6.17 $Y2=1.16
cc_148 VPB N_VPWR_c_899_n 0.00478085f $X=-0.19 $Y=1.305 $X2=7.19 $Y2=1.16
cc_149 VPB N_A_806_297#_c_1036_n 0.00262696f $X=-0.19 $Y=1.305 $X2=6.465
+ $Y2=0.995
cc_150 VPB N_A_806_297#_c_1037_n 0.001919f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_806_297#_c_1038_n 0.012098f $X=-0.19 $Y=1.305 $X2=6.885 $Y2=0.56
cc_152 VPB N_A_806_297#_c_1039_n 0.00198578f $X=-0.19 $Y=1.305 $X2=2.715
+ $Y2=1.275
cc_153 VPB N_X_c_1156_n 0.00424523f $X=-0.19 $Y=1.305 $X2=1.745 $Y2=1.985
cc_154 VPB N_X_c_1157_n 0.0050778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_X_c_1158_n 0.00235314f $X=-0.19 $Y=1.305 $X2=6.045 $Y2=0.56
cc_156 VPB N_X_c_1159_n 0.00238764f $X=-0.19 $Y=1.305 $X2=6.465 $Y2=1.985
cc_157 VPB N_X_c_1147_n 0.00788529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_X_c_1161_n 0.00202537f $X=-0.19 $Y=1.305 $X2=7.305 $Y2=1.985
cc_159 VPB N_X_c_1162_n 0.0103627f $X=-0.19 $Y=1.305 $X2=5.995 $Y2=1.53
cc_160 VPB X 0.0386269f $X=-0.19 $Y=1.305 $X2=2.8 $Y2=1.53
cc_161 N_A_c_164_n N_B_c_390_n 0.0240976f $X=1.745 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_162 N_A_M1038_g N_B_M1003_g 0.0240976f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_c_180_n N_B_M1003_g 5.91037e-19 $X=2.715 $Y=1.445 $X2=0 $Y2=0
cc_164 N_A_c_188_p N_B_M1003_g 2.10088e-19 $X=2.8 $Y=1.53 $X2=0 $Y2=0
cc_165 N_A_c_180_n N_B_M1006_g 0.00263969f $X=2.715 $Y=1.445 $X2=0 $Y2=0
cc_166 N_A_c_188_p N_B_M1006_g 0.00382121f $X=2.8 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A_c_180_n N_B_M1007_g 0.0025712f $X=2.715 $Y=1.445 $X2=0 $Y2=0
cc_168 N_A_c_181_n N_B_M1007_g 0.0108527f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_169 N_A_c_181_n N_B_M1026_g 0.0170519f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_170 N_A_c_181_n N_B_c_394_n 0.0145065f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_171 N_A_c_180_n N_B_c_395_n 0.00598194f $X=2.715 $Y=1.445 $X2=0 $Y2=0
cc_172 N_A_c_181_n N_B_c_395_n 0.00325236f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_173 N_A_c_169_n N_B_c_395_n 0.0358208f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_174 N_A_c_170_n N_B_c_395_n 0.0240976f $X=1.745 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_c_181_n N_B_M1000_g 0.0124706f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_176 N_A_c_181_n N_B_M1002_g 0.0103677f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_177 N_A_c_181_n N_B_M1008_g 0.0103557f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_178 N_A_c_165_n N_B_c_399_n 0.0196357f $X=6.045 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_M1009_g N_B_M1027_g 0.0196357f $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_c_181_n N_B_M1027_g 0.0103139f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_181 N_A_c_181_n N_B_c_400_n 0.177613f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_182 N_A_c_206_p N_B_c_400_n 0.0110392f $X=6.165 $Y=1.175 $X2=0 $Y2=0
cc_183 N_A_c_169_n N_B_c_400_n 0.0167609f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_184 N_A_c_171_n N_B_c_400_n 0.00135129f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_c_181_n N_B_c_401_n 0.00642092f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_186 N_A_c_182_n N_B_c_401_n 0.00106864f $X=6.08 $Y=1.445 $X2=0 $Y2=0
cc_187 N_A_c_206_p N_B_c_401_n 4.0849e-19 $X=6.165 $Y=1.175 $X2=0 $Y2=0
cc_188 N_A_c_171_n N_B_c_401_n 0.0196357f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_c_181_n N_A_112_47#_M1007_s 0.00165831f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_190 N_A_c_161_n N_A_112_47#_c_548_n 0.0181146f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_169_n N_A_112_47#_c_548_n 0.015823f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_192 N_A_c_161_n N_A_112_47#_c_549_n 0.0101732f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_169_n N_A_112_47#_c_549_n 0.00717314f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_194 N_A_c_161_n N_A_112_47#_c_579_n 0.0106039f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_162_n N_A_112_47#_c_579_n 0.00630972f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_163_n N_A_112_47#_c_579_n 5.22228e-19 $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_162_n N_A_112_47#_c_551_n 0.00870364f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_c_163_n N_A_112_47#_c_551_n 0.00870364f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_c_169_n N_A_112_47#_c_551_n 0.036111f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_200 N_A_c_170_n N_A_112_47#_c_551_n 0.00222133f $X=1.745 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_c_162_n N_A_112_47#_c_586_n 5.22228e-19 $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_163_n N_A_112_47#_c_586_n 0.00630972f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_164_n N_A_112_47#_c_586_n 0.00630972f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_164_n N_A_112_47#_c_552_n 0.00865686f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_c_169_n N_A_112_47#_c_552_n 0.0364455f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_206 N_A_c_164_n N_A_112_47#_c_591_n 5.22228e-19 $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_c_181_n N_A_112_47#_c_592_n 0.0139853f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_208 N_A_c_188_p N_A_112_47#_c_592_n 0.00809252f $X=2.8 $Y=1.53 $X2=0 $Y2=0
cc_209 N_A_c_169_n N_A_112_47#_c_592_n 0.00150764f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_210 N_A_c_181_n N_A_112_47#_c_553_n 0.00432883f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_211 N_A_c_169_n N_A_112_47#_c_553_n 0.0188803f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_212 N_A_c_171_n N_A_112_47#_c_554_n 0.00609322f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_c_237_p N_A_112_47#_c_555_n 0.0150669f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_c_171_n N_A_112_47#_c_555_n 0.00470444f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_c_161_n N_A_112_47#_c_556_n 0.00158032f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_c_162_n N_A_112_47#_c_556_n 0.00113286f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_c_169_n N_A_112_47#_c_556_n 0.0265405f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_218 N_A_c_170_n N_A_112_47#_c_556_n 0.00230339f $X=1.745 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_c_163_n N_A_112_47#_c_557_n 0.00113286f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_164_n N_A_112_47#_c_557_n 0.00113286f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_c_169_n N_A_112_47#_c_557_n 0.0265405f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_222 N_A_c_170_n N_A_112_47#_c_557_n 0.00230339f $X=1.745 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_c_169_n N_A_112_47#_c_558_n 0.0256811f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_224 N_A_M1004_g N_A_112_47#_c_568_n 0.012039f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_M1018_g N_A_112_47#_c_568_n 0.0103677f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A_M1025_g N_A_112_47#_c_568_n 0.0103677f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_M1038_g N_A_112_47#_c_568_n 0.0103235f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_c_188_p N_A_112_47#_c_568_n 0.00983136f $X=2.8 $Y=1.53 $X2=0 $Y2=0
cc_229 N_A_c_169_n N_A_112_47#_c_568_n 0.140206f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_230 N_A_c_170_n N_A_112_47#_c_568_n 0.00642092f $X=1.745 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_c_169_n N_A_112_47#_c_616_n 7.43958e-19 $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_232 N_A_c_181_n N_A_112_47#_c_617_n 0.0108571f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_233 N_A_M1019_g N_A_112_47#_c_569_n 0.00410596f $X=6.465 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_M1033_g N_A_112_47#_c_569_n 0.00410596f $X=6.885 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_M1039_g N_A_112_47#_c_569_n 0.00137956f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A_c_181_n N_A_112_47#_c_569_n 0.14787f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_237 N_A_c_188_p N_A_112_47#_c_569_n 0.00925036f $X=2.8 $Y=1.53 $X2=0 $Y2=0
cc_238 N_A_c_237_p N_A_112_47#_c_569_n 0.012924f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_c_169_n N_A_112_47#_c_569_n 0.00698296f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_240 N_A_c_171_n N_A_112_47#_c_569_n 0.00319534f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_M1038_g N_A_112_47#_c_570_n 9.85556e-19 $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A_c_180_n N_A_112_47#_c_570_n 9.2125e-19 $X=2.715 $Y=1.445 $X2=0 $Y2=0
cc_243 N_A_c_169_n N_A_112_47#_c_570_n 0.0077295f $X=2.63 $Y=1.175 $X2=0 $Y2=0
cc_244 N_A_M1039_g N_A_112_47#_c_571_n 0.00157208f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_M1033_g N_A_112_47#_c_572_n 6.78268e-19 $X=6.885 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A_M1039_g N_A_112_47#_c_572_n 0.0100813f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_c_237_p N_A_112_47#_c_572_n 0.00660761f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_c_181_n N_A_27_297#_M1006_d 7.6724e-19 $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_249 N_A_c_188_p N_A_27_297#_M1006_d 9.14305e-19 $X=2.8 $Y=1.53 $X2=0 $Y2=0
cc_250 N_A_c_181_n N_A_27_297#_M1026_d 0.00277065f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_251 N_A_M1004_g N_A_27_297#_c_820_n 0.0113824f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_M1018_g N_A_27_297#_c_820_n 0.0113824f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_M1025_g N_A_27_297#_c_822_n 0.0113251f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A_M1038_g N_A_27_297#_c_822_n 0.0113824f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A_c_181_n N_A_27_297#_c_824_n 0.0140276f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_256 N_A_c_181_n N_VPWR_M1000_s 0.00166235f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_257 N_A_c_181_n N_VPWR_M1008_s 0.00166235f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_258 N_A_M1004_g N_VPWR_c_880_n 0.00302074f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A_M1018_g N_VPWR_c_880_n 0.00157837f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_M1025_g N_VPWR_c_881_n 0.00157837f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A_M1038_g N_VPWR_c_881_n 0.00302074f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A_M1009_g N_VPWR_c_885_n 0.00436487f $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_M1009_g N_VPWR_c_886_n 0.00157837f $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A_M1019_g N_VPWR_c_886_n 0.00157837f $X=6.465 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A_M1033_g N_VPWR_c_887_n 0.00157837f $X=6.885 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A_M1039_g N_VPWR_c_887_n 0.00302074f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A_M1038_g N_VPWR_c_888_n 0.00436487f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A_M1004_g N_VPWR_c_890_n 0.00436487f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A_M1018_g N_VPWR_c_891_n 0.00436487f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_M1025_g N_VPWR_c_891_n 0.00436487f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_M1019_g N_VPWR_c_892_n 0.00436487f $X=6.465 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_M1033_g N_VPWR_c_892_n 0.00436487f $X=6.885 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_M1039_g N_VPWR_c_893_n 0.00436487f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A_M1004_g N_VPWR_c_879_n 0.00673011f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A_M1018_g N_VPWR_c_879_n 0.00576179f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A_M1025_g N_VPWR_c_879_n 0.00576179f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_M1038_g N_VPWR_c_879_n 0.00578899f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A_M1009_g N_VPWR_c_879_n 0.00578899f $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A_M1019_g N_VPWR_c_879_n 0.00576179f $X=6.465 $Y=1.985 $X2=0 $Y2=0
cc_280 N_A_M1033_g N_VPWR_c_879_n 0.00576179f $X=6.885 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_M1039_g N_VPWR_c_879_n 0.00708786f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A_c_181_n N_A_806_297#_M1000_d 0.00272914f $X=5.995 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_283 N_A_c_181_n N_A_806_297#_M1002_d 0.00165831f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_284 N_A_c_181_n N_A_806_297#_M1027_d 0.00165831f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_285 N_A_c_181_n N_A_806_297#_c_1043_n 0.0292185f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_286 N_A_c_181_n N_A_806_297#_c_1044_n 0.0292185f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_287 N_A_M1009_g N_A_806_297#_c_1045_n 0.0112896f $X=6.045 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_M1019_g N_A_806_297#_c_1045_n 0.0127541f $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_A_c_181_n N_A_806_297#_c_1045_n 0.0101711f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_290 N_A_c_237_p N_A_806_297#_c_1045_n 0.00442469f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A_c_171_n N_A_806_297#_c_1045_n 0.00167017f $X=7.305 $Y=1.16 $X2=0
+ $Y2=0
cc_292 N_A_M1019_g N_A_806_297#_c_1036_n 6.25986e-19 $X=6.465 $Y=1.985 $X2=0
+ $Y2=0
cc_293 N_A_M1033_g N_A_806_297#_c_1036_n 7.04624e-19 $X=6.885 $Y=1.985 $X2=0
+ $Y2=0
cc_294 N_A_c_181_n N_A_806_297#_c_1036_n 0.00285531f $X=5.995 $Y=1.53 $X2=0
+ $Y2=0
cc_295 N_A_c_237_p N_A_806_297#_c_1036_n 0.0169277f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_c_171_n N_A_806_297#_c_1036_n 0.00221654f $X=7.305 $Y=1.16 $X2=0
+ $Y2=0
cc_297 N_A_M1033_g N_A_806_297#_c_1055_n 0.0126968f $X=6.885 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_M1039_g N_A_806_297#_c_1055_n 0.0115989f $X=7.305 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A_c_237_p N_A_806_297#_c_1055_n 0.00507953f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_c_171_n N_A_806_297#_c_1055_n 0.00167017f $X=7.305 $Y=1.16 $X2=0
+ $Y2=0
cc_301 N_A_c_181_n N_A_806_297#_c_1039_n 0.0148561f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_302 N_A_c_181_n N_A_806_297#_c_1060_n 0.0114165f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_303 N_A_c_181_n N_A_806_297#_c_1061_n 0.0114165f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_304 N_A_M1039_g N_X_c_1156_n 0.00213556f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A_M1039_g N_X_c_1157_n 0.00284818f $X=7.305 $Y=1.985 $X2=0 $Y2=0
cc_306 N_A_c_168_n N_X_c_1148_n 9.12162e-19 $X=7.305 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_c_165_n N_X_c_1151_n 0.00162479f $X=6.045 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_c_166_n N_X_c_1151_n 0.00154513f $X=6.465 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_c_167_n N_X_c_1151_n 0.00154513f $X=6.885 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A_c_168_n N_X_c_1151_n 0.00172908f $X=7.305 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A_c_181_n N_X_c_1151_n 0.00251758f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_312 N_A_c_206_p N_X_c_1151_n 0.00174064f $X=6.165 $Y=1.175 $X2=0 $Y2=0
cc_313 N_A_c_237_p N_X_c_1151_n 0.0121354f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_c_171_n N_X_c_1151_n 0.00502053f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_c_165_n N_X_c_1153_n 3.27985e-19 $X=6.045 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A_c_168_n N_X_c_1154_n 5.99935e-19 $X=7.305 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_c_161_n N_VGND_c_1308_n 0.00322518f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A_c_162_n N_VGND_c_1309_n 0.00146448f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_c_163_n N_VGND_c_1309_n 0.00146448f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_c_164_n N_VGND_c_1310_n 0.00146448f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_c_165_n N_VGND_c_1313_n 0.00268723f $X=6.045 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_c_166_n N_VGND_c_1313_n 0.00146448f $X=6.465 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_c_167_n N_VGND_c_1314_n 0.00146448f $X=6.885 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_c_168_n N_VGND_c_1314_n 0.00268723f $X=7.305 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_c_168_n N_VGND_c_1315_n 0.00191367f $X=7.305 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_c_161_n N_VGND_c_1318_n 0.00424416f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_c_162_n N_VGND_c_1318_n 0.00423334f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_c_163_n N_VGND_c_1320_n 0.00423334f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A_c_164_n N_VGND_c_1320_n 0.00423334f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_c_166_n N_VGND_c_1326_n 0.00423334f $X=6.465 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_c_167_n N_VGND_c_1326_n 0.00423334f $X=6.885 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_c_168_n N_VGND_c_1328_n 0.00423334f $X=7.305 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_c_165_n N_VGND_c_1334_n 0.00421816f $X=6.045 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_c_161_n N_VGND_c_1336_n 0.00670439f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_c_162_n N_VGND_c_1336_n 0.0057163f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A_c_163_n N_VGND_c_1336_n 0.0057163f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A_c_164_n N_VGND_c_1336_n 0.0057435f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_c_165_n N_VGND_c_1336_n 0.00544403f $X=6.045 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_c_166_n N_VGND_c_1336_n 0.0054081f $X=6.465 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_c_167_n N_VGND_c_1336_n 0.0054081f $X=6.885 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A_c_168_n N_VGND_c_1336_n 0.00673417f $X=7.305 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A_c_165_n N_A_806_47#_c_1494_n 0.00255288f $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A_c_165_n N_A_806_47#_c_1489_n 0.00491819f $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A_c_166_n N_A_806_47#_c_1489_n 4.58193e-19 $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A_c_181_n N_A_806_47#_c_1489_n 0.00482919f $X=5.995 $Y=1.53 $X2=0 $Y2=0
cc_346 N_A_c_206_p N_A_806_47#_c_1489_n 3.31463e-19 $X=6.165 $Y=1.175 $X2=0
+ $Y2=0
cc_347 N_A_c_165_n N_A_806_47#_c_1490_n 0.00796409f $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_348 N_A_c_166_n N_A_806_47#_c_1490_n 0.00792293f $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_c_206_p N_A_806_47#_c_1490_n 0.0109022f $X=6.165 $Y=1.175 $X2=0 $Y2=0
cc_350 N_A_c_237_p N_A_806_47#_c_1490_n 0.0214391f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A_c_171_n N_A_806_47#_c_1490_n 0.00218025f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A_c_165_n N_A_806_47#_c_1504_n 5.22228e-19 $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_353 N_A_c_166_n N_A_806_47#_c_1504_n 0.00630972f $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_354 N_A_c_167_n N_A_806_47#_c_1504_n 0.00630972f $X=6.885 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A_c_168_n N_A_806_47#_c_1504_n 5.22228e-19 $X=7.305 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_c_167_n N_A_806_47#_c_1491_n 0.00796971f $X=6.885 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_c_168_n N_A_806_47#_c_1491_n 0.00917009f $X=7.305 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A_c_237_p N_A_806_47#_c_1491_n 0.0327612f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A_c_171_n N_A_806_47#_c_1491_n 0.00218025f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A_c_167_n N_A_806_47#_c_1492_n 5.22228e-19 $X=6.885 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_c_168_n N_A_806_47#_c_1492_n 0.00630972f $X=7.305 $Y=0.995 $X2=0
+ $Y2=0
cc_362 N_A_c_166_n N_A_806_47#_c_1493_n 9.29836e-19 $X=6.465 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_c_167_n N_A_806_47#_c_1493_n 9.29836e-19 $X=6.885 $Y=0.995 $X2=0
+ $Y2=0
cc_364 N_A_c_237_p N_A_806_47#_c_1493_n 0.0212739f $X=7.19 $Y=1.16 $X2=0 $Y2=0
cc_365 N_A_c_171_n N_A_806_47#_c_1493_n 0.00221535f $X=7.305 $Y=1.16 $X2=0 $Y2=0
cc_366 N_B_c_390_n N_A_112_47#_c_586_n 5.22228e-19 $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_367 N_B_c_390_n N_A_112_47#_c_552_n 0.00864834f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_368 N_B_c_390_n N_A_112_47#_c_591_n 0.00630972f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_369 N_B_c_391_n N_A_112_47#_c_591_n 0.00630972f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_370 N_B_c_392_n N_A_112_47#_c_591_n 5.22228e-19 $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_371 N_B_M1006_g N_A_112_47#_c_592_n 0.0102928f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_372 N_B_M1007_g N_A_112_47#_c_592_n 0.00916638f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_373 N_B_c_395_n N_A_112_47#_c_592_n 2.49536e-19 $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_374 N_B_c_391_n N_A_112_47#_c_553_n 0.00869626f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_375 N_B_c_392_n N_A_112_47#_c_553_n 0.0102974f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_376 N_B_c_393_n N_A_112_47#_c_553_n 0.00299088f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_377 N_B_c_395_n N_A_112_47#_c_553_n 0.00470323f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_378 N_B_c_400_n N_A_112_47#_c_553_n 0.0310079f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_379 N_B_c_391_n N_A_112_47#_c_646_n 5.22228e-19 $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_380 N_B_c_392_n N_A_112_47#_c_646_n 0.00630972f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_381 N_B_c_393_n N_A_112_47#_c_646_n 0.00538815f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_382 N_B_c_390_n N_A_112_47#_c_558_n 0.00107362f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_383 N_B_c_391_n N_A_112_47#_c_558_n 0.00113127f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_384 N_B_c_395_n N_A_112_47#_c_558_n 0.00230339f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_385 N_B_M1003_g N_A_112_47#_c_568_n 0.010997f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_386 N_B_M1006_g N_A_112_47#_c_568_n 0.00112412f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_387 N_B_c_395_n N_A_112_47#_c_568_n 0.00222344f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_388 N_B_M1006_g N_A_112_47#_c_655_n 0.00374677f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_389 N_B_M1006_g N_A_112_47#_c_569_n 0.00310092f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_390 N_B_c_400_n N_A_112_47#_c_569_n 0.0178034f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_391 N_B_M1003_g N_A_112_47#_c_570_n 0.00717649f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_392 N_B_M1003_g N_A_27_297#_c_825_n 0.0121306f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_393 N_B_M1006_g N_A_27_297#_c_825_n 0.00851673f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_394 N_B_M1007_g N_A_27_297#_c_815_n 0.00851673f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_395 N_B_M1026_g N_A_27_297#_c_815_n 0.0121306f $X=3.425 $Y=1.985 $X2=0 $Y2=0
cc_396 N_B_M1000_g N_VPWR_c_882_n 0.00302074f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_397 N_B_M1002_g N_VPWR_c_882_n 0.00157837f $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_398 N_B_M1002_g N_VPWR_c_883_n 0.00436487f $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_399 N_B_M1008_g N_VPWR_c_883_n 0.00436487f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_400 N_B_M1008_g N_VPWR_c_884_n 0.00157837f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_401 N_B_M1027_g N_VPWR_c_884_n 0.00157837f $X=5.625 $Y=1.985 $X2=0 $Y2=0
cc_402 N_B_M1027_g N_VPWR_c_885_n 0.00436487f $X=5.625 $Y=1.985 $X2=0 $Y2=0
cc_403 N_B_M1003_g N_VPWR_c_888_n 0.00357877f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_404 N_B_M1006_g N_VPWR_c_888_n 0.00357877f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_405 N_B_M1007_g N_VPWR_c_888_n 0.00357877f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_406 N_B_M1026_g N_VPWR_c_888_n 0.00357877f $X=3.425 $Y=1.985 $X2=0 $Y2=0
cc_407 N_B_M1000_g N_VPWR_c_888_n 0.00436487f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_408 N_B_M1003_g N_VPWR_c_879_n 0.00525237f $X=2.165 $Y=1.985 $X2=0 $Y2=0
cc_409 N_B_M1006_g N_VPWR_c_879_n 0.00522516f $X=2.585 $Y=1.985 $X2=0 $Y2=0
cc_410 N_B_M1007_g N_VPWR_c_879_n 0.00522516f $X=3.005 $Y=1.985 $X2=0 $Y2=0
cc_411 N_B_M1026_g N_VPWR_c_879_n 0.00655123f $X=3.425 $Y=1.985 $X2=0 $Y2=0
cc_412 N_B_M1000_g N_VPWR_c_879_n 0.00708786f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_413 N_B_M1002_g N_VPWR_c_879_n 0.00576179f $X=4.785 $Y=1.985 $X2=0 $Y2=0
cc_414 N_B_M1008_g N_VPWR_c_879_n 0.00576179f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_415 N_B_M1027_g N_VPWR_c_879_n 0.00578899f $X=5.625 $Y=1.985 $X2=0 $Y2=0
cc_416 N_B_M1000_g N_A_806_297#_c_1043_n 0.0113077f $X=4.365 $Y=1.985 $X2=0
+ $Y2=0
cc_417 N_B_M1002_g N_A_806_297#_c_1043_n 0.0112504f $X=4.785 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_B_M1008_g N_A_806_297#_c_1044_n 0.0113077f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_419 N_B_M1027_g N_A_806_297#_c_1044_n 0.0113077f $X=5.625 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_B_c_399_n N_X_c_1151_n 0.00255345f $X=5.625 $Y=0.995 $X2=0 $Y2=0
cc_421 N_B_c_400_n N_X_c_1151_n 0.00286238f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_422 N_B_c_397_n N_X_c_1152_n 3.17759e-19 $X=4.785 $Y=0.995 $X2=0 $Y2=0
cc_423 N_B_c_398_n N_X_c_1152_n 0.00226352f $X=5.205 $Y=0.995 $X2=0 $Y2=0
cc_424 N_B_c_399_n N_X_c_1152_n 4.89226e-19 $X=5.625 $Y=0.995 $X2=0 $Y2=0
cc_425 N_B_c_400_n N_X_c_1152_n 0.00301398f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_426 N_B_c_401_n N_X_c_1152_n 0.00127791f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_427 N_B_c_397_n N_X_c_1153_n 3.04965e-19 $X=4.785 $Y=0.995 $X2=0 $Y2=0
cc_428 N_B_c_398_n N_X_c_1153_n 0.0073213f $X=5.205 $Y=0.995 $X2=0 $Y2=0
cc_429 N_B_c_399_n N_X_c_1153_n 0.00428123f $X=5.625 $Y=0.995 $X2=0 $Y2=0
cc_430 N_B_c_400_n N_X_c_1153_n 0.0269599f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_431 N_B_c_401_n N_X_c_1153_n 0.00229185f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_432 N_B_c_393_n N_X_c_1155_n 8.28316e-19 $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_433 N_B_c_394_n N_X_c_1155_n 8.71943e-19 $X=4.29 $Y=1.16 $X2=0 $Y2=0
cc_434 N_B_c_396_n N_X_c_1155_n 0.0123073f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_435 N_B_c_397_n N_X_c_1155_n 0.0109499f $X=4.785 $Y=0.995 $X2=0 $Y2=0
cc_436 N_B_c_398_n N_X_c_1155_n 0.00393598f $X=5.205 $Y=0.995 $X2=0 $Y2=0
cc_437 N_B_c_400_n N_X_c_1155_n 0.0685937f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_438 N_B_c_401_n N_X_c_1155_n 0.00450248f $X=5.625 $Y=1.16 $X2=0 $Y2=0
cc_439 N_B_c_390_n N_VGND_c_1310_n 0.00146448f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_440 N_B_c_391_n N_VGND_c_1311_n 0.00146448f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_441 N_B_c_392_n N_VGND_c_1311_n 0.00146448f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_442 N_B_c_393_n N_VGND_c_1312_n 0.00344333f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_443 N_B_c_394_n N_VGND_c_1312_n 0.00585142f $X=4.29 $Y=1.16 $X2=0 $Y2=0
cc_444 N_B_c_396_n N_VGND_c_1312_n 0.00685325f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_445 N_B_c_400_n N_VGND_c_1312_n 0.02016f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_446 N_B_c_390_n N_VGND_c_1322_n 0.00423334f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_447 N_B_c_391_n N_VGND_c_1322_n 0.00423334f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_448 N_B_c_392_n N_VGND_c_1324_n 0.00423334f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_449 N_B_c_393_n N_VGND_c_1324_n 0.00541359f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_450 N_B_c_396_n N_VGND_c_1334_n 0.00357877f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_451 N_B_c_397_n N_VGND_c_1334_n 0.00357877f $X=4.785 $Y=0.995 $X2=0 $Y2=0
cc_452 N_B_c_398_n N_VGND_c_1334_n 0.00357877f $X=5.205 $Y=0.995 $X2=0 $Y2=0
cc_453 N_B_c_399_n N_VGND_c_1334_n 0.00357877f $X=5.625 $Y=0.995 $X2=0 $Y2=0
cc_454 N_B_c_390_n N_VGND_c_1336_n 0.0057435f $X=2.165 $Y=0.995 $X2=0 $Y2=0
cc_455 N_B_c_391_n N_VGND_c_1336_n 0.0057163f $X=2.585 $Y=0.995 $X2=0 $Y2=0
cc_456 N_B_c_392_n N_VGND_c_1336_n 0.0057163f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_457 N_B_c_393_n N_VGND_c_1336_n 0.0108276f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_458 N_B_c_396_n N_VGND_c_1336_n 0.00655123f $X=4.365 $Y=0.995 $X2=0 $Y2=0
cc_459 N_B_c_397_n N_VGND_c_1336_n 0.00522516f $X=4.785 $Y=0.995 $X2=0 $Y2=0
cc_460 N_B_c_398_n N_VGND_c_1336_n 0.00513402f $X=5.205 $Y=0.995 $X2=0 $Y2=0
cc_461 N_B_c_399_n N_VGND_c_1336_n 0.00519981f $X=5.625 $Y=0.995 $X2=0 $Y2=0
cc_462 N_B_c_394_n N_A_806_47#_c_1488_n 0.00316065f $X=4.29 $Y=1.16 $X2=0 $Y2=0
cc_463 N_B_c_396_n N_A_806_47#_c_1488_n 0.00892725f $X=4.365 $Y=0.995 $X2=0
+ $Y2=0
cc_464 N_B_c_397_n N_A_806_47#_c_1488_n 0.00892725f $X=4.785 $Y=0.995 $X2=0
+ $Y2=0
cc_465 N_B_c_398_n N_A_806_47#_c_1488_n 0.00887963f $X=5.205 $Y=0.995 $X2=0
+ $Y2=0
cc_466 N_B_c_399_n N_A_806_47#_c_1488_n 0.0103901f $X=5.625 $Y=0.995 $X2=0 $Y2=0
cc_467 N_B_c_400_n N_A_806_47#_c_1488_n 0.00610045f $X=4.835 $Y=1.16 $X2=0 $Y2=0
cc_468 N_B_c_399_n N_A_806_47#_c_1489_n 2.75855e-19 $X=5.625 $Y=0.995 $X2=0
+ $Y2=0
cc_469 N_A_112_47#_c_567_n N_A_27_297#_M1004_s 0.00201153f $X=0.255 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_470 N_A_112_47#_c_568_n N_A_27_297#_M1004_s 0.00103113f $X=2.25 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_471 N_A_112_47#_c_568_n N_A_27_297#_M1018_s 0.00165831f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_472 N_A_112_47#_c_568_n N_A_27_297#_M1038_s 0.00101922f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_473 N_A_112_47#_c_570_n N_A_27_297#_M1038_s 0.00216671f $X=2.215 $Y=1.53
+ $X2=0 $Y2=0
cc_474 N_A_112_47#_c_592_n N_A_27_297#_M1006_d 0.00302367f $X=3.09 $Y=1.87 $X2=0
+ $Y2=0
cc_475 N_A_112_47#_c_568_n N_A_27_297#_c_820_n 0.0322288f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_476 N_A_112_47#_c_568_n N_A_27_297#_c_822_n 0.0322288f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_477 N_A_112_47#_c_568_n N_A_27_297#_c_837_n 0.0123683f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_478 N_A_112_47#_c_570_n N_A_27_297#_c_837_n 0.0045571f $X=2.215 $Y=1.53 $X2=0
+ $Y2=0
cc_479 N_A_112_47#_M1003_s N_A_27_297#_c_825_n 0.00312348f $X=2.24 $Y=1.485
+ $X2=0 $Y2=0
cc_480 N_A_112_47#_c_592_n N_A_27_297#_c_825_n 0.00506389f $X=3.09 $Y=1.87 $X2=0
+ $Y2=0
cc_481 N_A_112_47#_c_616_n N_A_27_297#_c_825_n 0.0117584f $X=2.375 $Y=1.87 $X2=0
+ $Y2=0
cc_482 N_A_112_47#_M1007_s N_A_27_297#_c_815_n 0.00312348f $X=3.08 $Y=1.485
+ $X2=0 $Y2=0
cc_483 N_A_112_47#_c_592_n N_A_27_297#_c_815_n 0.00506389f $X=3.09 $Y=1.87 $X2=0
+ $Y2=0
cc_484 N_A_112_47#_c_617_n N_A_27_297#_c_815_n 0.0112811f $X=3.215 $Y=1.87 $X2=0
+ $Y2=0
cc_485 N_A_112_47#_c_569_n N_A_27_297#_c_824_n 0.00206914f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_486 N_A_112_47#_c_567_n N_A_27_297#_c_816_n 0.0154106f $X=0.255 $Y=1.53 $X2=0
+ $Y2=0
cc_487 N_A_112_47#_c_568_n N_A_27_297#_c_816_n 0.00793666f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_488 N_A_112_47#_c_568_n N_A_27_297#_c_848_n 0.0126919f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_489 N_A_112_47#_c_592_n N_A_27_297#_c_849_n 0.0112429f $X=3.09 $Y=1.87 $X2=0
+ $Y2=0
cc_490 N_A_112_47#_c_568_n N_VPWR_M1004_d 0.00166235f $X=2.25 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_491 N_A_112_47#_c_568_n N_VPWR_M1025_d 0.00166235f $X=2.25 $Y=1.53 $X2=0
+ $Y2=0
cc_492 N_A_112_47#_c_569_n N_VPWR_M1009_s 0.00179738f $X=7.445 $Y=1.53 $X2=0
+ $Y2=0
cc_493 N_A_112_47#_c_569_n N_VPWR_M1033_s 0.00224381f $X=7.445 $Y=1.53 $X2=0
+ $Y2=0
cc_494 N_A_112_47#_M1001_g N_VPWR_c_893_n 0.00357877f $X=8.255 $Y=1.985 $X2=0
+ $Y2=0
cc_495 N_A_112_47#_M1016_g N_VPWR_c_893_n 0.00357877f $X=8.675 $Y=1.985 $X2=0
+ $Y2=0
cc_496 N_A_112_47#_M1022_g N_VPWR_c_893_n 0.00357877f $X=9.095 $Y=1.985 $X2=0
+ $Y2=0
cc_497 N_A_112_47#_M1035_g N_VPWR_c_893_n 0.00585385f $X=9.515 $Y=1.985 $X2=0
+ $Y2=0
cc_498 N_A_112_47#_M1003_s N_VPWR_c_879_n 0.0021603f $X=2.24 $Y=1.485 $X2=0
+ $Y2=0
cc_499 N_A_112_47#_M1007_s N_VPWR_c_879_n 0.0021603f $X=3.08 $Y=1.485 $X2=0
+ $Y2=0
cc_500 N_A_112_47#_M1001_g N_VPWR_c_879_n 0.00660224f $X=8.255 $Y=1.985 $X2=0
+ $Y2=0
cc_501 N_A_112_47#_M1016_g N_VPWR_c_879_n 0.00522516f $X=8.675 $Y=1.985 $X2=0
+ $Y2=0
cc_502 N_A_112_47#_M1022_g N_VPWR_c_879_n 0.00522516f $X=9.095 $Y=1.985 $X2=0
+ $Y2=0
cc_503 N_A_112_47#_M1035_g N_VPWR_c_879_n 0.0117207f $X=9.515 $Y=1.985 $X2=0
+ $Y2=0
cc_504 N_A_112_47#_c_592_n N_VPWR_c_879_n 0.00127799f $X=3.09 $Y=1.87 $X2=0
+ $Y2=0
cc_505 N_A_112_47#_c_554_n N_A_806_297#_M1039_d 9.21756e-19 $X=7.625 $Y=1.445
+ $X2=0 $Y2=0
cc_506 N_A_112_47#_c_571_n N_A_806_297#_M1039_d 0.00200707f $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_507 N_A_112_47#_c_572_n N_A_806_297#_M1039_d 5.28034e-19 $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_508 N_A_112_47#_c_569_n N_A_806_297#_c_1043_n 0.00434997f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_509 N_A_112_47#_c_569_n N_A_806_297#_c_1044_n 0.00434997f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_510 N_A_112_47#_c_569_n N_A_806_297#_c_1045_n 0.0121139f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_511 N_A_112_47#_c_569_n N_A_806_297#_c_1036_n 0.0259796f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_512 N_A_112_47#_c_572_n N_A_806_297#_c_1036_n 0.00274272f $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_513 N_A_112_47#_c_569_n N_A_806_297#_c_1055_n 0.0136724f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_514 N_A_112_47#_c_572_n N_A_806_297#_c_1055_n 0.0074925f $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_515 N_A_112_47#_c_554_n N_A_806_297#_c_1037_n 0.00721577f $X=7.625 $Y=1.445
+ $X2=0 $Y2=0
cc_516 N_A_112_47#_c_569_n N_A_806_297#_c_1037_n 4.56591e-19 $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_517 N_A_112_47#_c_571_n N_A_806_297#_c_1037_n 0.00573091f $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_518 N_A_112_47#_c_572_n N_A_806_297#_c_1037_n 0.00726173f $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_519 N_A_112_47#_M1001_g N_A_806_297#_c_1080_n 0.00398343f $X=8.255 $Y=1.985
+ $X2=0 $Y2=0
cc_520 N_A_112_47#_M1001_g N_A_806_297#_c_1038_n 0.011858f $X=8.255 $Y=1.985
+ $X2=0 $Y2=0
cc_521 N_A_112_47#_M1016_g N_A_806_297#_c_1082_n 0.00971087f $X=8.675 $Y=1.985
+ $X2=0 $Y2=0
cc_522 N_A_112_47#_M1022_g N_A_806_297#_c_1082_n 0.00988743f $X=9.095 $Y=1.985
+ $X2=0 $Y2=0
cc_523 N_A_112_47#_c_569_n N_A_806_297#_c_1039_n 0.00209664f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_524 N_A_112_47#_c_569_n N_A_806_297#_c_1060_n 0.00209664f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_525 N_A_112_47#_c_569_n N_A_806_297#_c_1061_n 0.00209664f $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_526 N_A_112_47#_c_554_n N_X_c_1156_n 0.0126709f $X=7.625 $Y=1.445 $X2=0 $Y2=0
cc_527 N_A_112_47#_c_559_n N_X_c_1156_n 0.0234895f $X=8.54 $Y=1.175 $X2=0 $Y2=0
cc_528 N_A_112_47#_c_571_n N_X_c_1156_n 0.00755503f $X=7.59 $Y=1.53 $X2=0 $Y2=0
cc_529 N_A_112_47#_M1001_g N_X_c_1158_n 0.0126358f $X=8.255 $Y=1.985 $X2=0 $Y2=0
cc_530 N_A_112_47#_M1016_g N_X_c_1158_n 0.0123223f $X=8.675 $Y=1.985 $X2=0 $Y2=0
cc_531 N_A_112_47#_c_559_n N_X_c_1158_n 0.0419387f $X=8.54 $Y=1.175 $X2=0 $Y2=0
cc_532 N_A_112_47#_c_560_n N_X_c_1158_n 0.00215368f $X=9.515 $Y=1.16 $X2=0 $Y2=0
cc_533 N_A_112_47#_c_544_n N_X_c_1203_n 0.00717371f $X=8.255 $Y=0.995 $X2=0
+ $Y2=0
cc_534 N_A_112_47#_c_545_n N_X_c_1203_n 0.00630972f $X=8.675 $Y=0.995 $X2=0
+ $Y2=0
cc_535 N_A_112_47#_c_546_n N_X_c_1203_n 5.22228e-19 $X=9.095 $Y=0.995 $X2=0
+ $Y2=0
cc_536 N_A_112_47#_c_545_n N_X_c_1145_n 0.00850187f $X=8.675 $Y=0.995 $X2=0
+ $Y2=0
cc_537 N_A_112_47#_c_546_n N_X_c_1145_n 0.00850187f $X=9.095 $Y=0.995 $X2=0
+ $Y2=0
cc_538 N_A_112_47#_c_728_p N_X_c_1145_n 0.0359162f $X=8.64 $Y=1.175 $X2=0 $Y2=0
cc_539 N_A_112_47#_c_560_n N_X_c_1145_n 0.00221825f $X=9.515 $Y=1.16 $X2=0 $Y2=0
cc_540 N_A_112_47#_M1022_g N_X_c_1159_n 0.0113735f $X=9.095 $Y=1.985 $X2=0 $Y2=0
cc_541 N_A_112_47#_M1035_g N_X_c_1159_n 0.0143734f $X=9.515 $Y=1.985 $X2=0 $Y2=0
cc_542 N_A_112_47#_c_732_p N_X_c_1159_n 0.0392817f $X=9.385 $Y=1.16 $X2=0 $Y2=0
cc_543 N_A_112_47#_c_560_n N_X_c_1159_n 0.00214321f $X=9.515 $Y=1.16 $X2=0 $Y2=0
cc_544 N_A_112_47#_c_545_n N_X_c_1214_n 5.51569e-19 $X=8.675 $Y=0.995 $X2=0
+ $Y2=0
cc_545 N_A_112_47#_c_546_n N_X_c_1214_n 0.0064836f $X=9.095 $Y=0.995 $X2=0 $Y2=0
cc_546 N_A_112_47#_c_547_n N_X_c_1214_n 0.0113689f $X=9.515 $Y=0.995 $X2=0 $Y2=0
cc_547 N_A_112_47#_c_547_n N_X_c_1146_n 0.0105378f $X=9.515 $Y=0.995 $X2=0 $Y2=0
cc_548 N_A_112_47#_c_732_p N_X_c_1146_n 0.00648676f $X=9.385 $Y=1.16 $X2=0 $Y2=0
cc_549 N_A_112_47#_c_547_n N_X_c_1147_n 0.0192258f $X=9.515 $Y=0.995 $X2=0 $Y2=0
cc_550 N_A_112_47#_c_732_p N_X_c_1147_n 0.0164962f $X=9.385 $Y=1.16 $X2=0 $Y2=0
cc_551 N_A_112_47#_c_544_n N_X_c_1148_n 0.0111764f $X=8.255 $Y=0.995 $X2=0 $Y2=0
cc_552 N_A_112_47#_c_559_n N_X_c_1148_n 0.0299713f $X=8.54 $Y=1.175 $X2=0 $Y2=0
cc_553 N_A_112_47#_c_544_n N_X_c_1149_n 0.00161854f $X=8.255 $Y=0.995 $X2=0
+ $Y2=0
cc_554 N_A_112_47#_c_545_n N_X_c_1149_n 0.00145906f $X=8.675 $Y=0.995 $X2=0
+ $Y2=0
cc_555 N_A_112_47#_c_728_p N_X_c_1149_n 0.00717779f $X=8.64 $Y=1.175 $X2=0 $Y2=0
cc_556 N_A_112_47#_c_559_n N_X_c_1149_n 0.0169619f $X=8.54 $Y=1.175 $X2=0 $Y2=0
cc_557 N_A_112_47#_c_560_n N_X_c_1149_n 0.00235411f $X=9.515 $Y=1.16 $X2=0 $Y2=0
cc_558 N_A_112_47#_c_732_p N_X_c_1161_n 0.0203891f $X=9.385 $Y=1.16 $X2=0 $Y2=0
cc_559 N_A_112_47#_c_560_n N_X_c_1161_n 0.00222344f $X=9.515 $Y=1.16 $X2=0 $Y2=0
cc_560 N_A_112_47#_c_546_n N_X_c_1150_n 0.00110555f $X=9.095 $Y=0.995 $X2=0
+ $Y2=0
cc_561 N_A_112_47#_c_547_n N_X_c_1150_n 0.00110555f $X=9.515 $Y=0.995 $X2=0
+ $Y2=0
cc_562 N_A_112_47#_c_732_p N_X_c_1150_n 0.0265405f $X=9.385 $Y=1.16 $X2=0 $Y2=0
cc_563 N_A_112_47#_c_560_n N_X_c_1150_n 0.00230339f $X=9.515 $Y=1.16 $X2=0 $Y2=0
cc_564 N_A_112_47#_c_555_n N_X_c_1151_n 0.00260969f $X=7.71 $Y=1.19 $X2=0 $Y2=0
cc_565 N_A_112_47#_c_559_n N_X_c_1151_n 0.00627324f $X=8.54 $Y=1.175 $X2=0 $Y2=0
cc_566 N_A_112_47#_c_569_n N_X_c_1151_n 0.0880549f $X=7.445 $Y=1.53 $X2=0 $Y2=0
cc_567 N_A_112_47#_c_571_n N_X_c_1151_n 0.0143979f $X=7.59 $Y=1.53 $X2=0 $Y2=0
cc_568 N_A_112_47#_c_572_n N_X_c_1151_n 0.00120991f $X=7.59 $Y=1.53 $X2=0 $Y2=0
cc_569 N_A_112_47#_c_569_n N_X_c_1152_n 0.0135076f $X=7.445 $Y=1.53 $X2=0 $Y2=0
cc_570 N_A_112_47#_c_544_n N_X_c_1154_n 0.00105713f $X=8.255 $Y=0.995 $X2=0
+ $Y2=0
cc_571 N_A_112_47#_c_559_n N_X_c_1154_n 0.00817708f $X=8.54 $Y=1.175 $X2=0 $Y2=0
cc_572 N_A_112_47#_c_549_n N_VGND_M1012_s 0.00100734f $X=0.53 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_573 N_A_112_47#_c_550_n N_VGND_M1012_s 0.002086f $X=0.255 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_574 N_A_112_47#_c_551_n N_VGND_M1017_s 0.00162089f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_575 N_A_112_47#_c_552_n N_VGND_M1030_s 0.00162089f $X=2.21 $Y=0.815 $X2=0
+ $Y2=0
cc_576 N_A_112_47#_c_553_n N_VGND_M1029_d 0.00162089f $X=3.05 $Y=0.815 $X2=0
+ $Y2=0
cc_577 N_A_112_47#_c_549_n N_VGND_c_1308_n 0.00765622f $X=0.53 $Y=0.82 $X2=0
+ $Y2=0
cc_578 N_A_112_47#_c_550_n N_VGND_c_1308_n 0.0148186f $X=0.255 $Y=0.82 $X2=0
+ $Y2=0
cc_579 N_A_112_47#_c_551_n N_VGND_c_1309_n 0.0122559f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_580 N_A_112_47#_c_552_n N_VGND_c_1310_n 0.0122559f $X=2.21 $Y=0.815 $X2=0
+ $Y2=0
cc_581 N_A_112_47#_c_553_n N_VGND_c_1311_n 0.0122559f $X=3.05 $Y=0.815 $X2=0
+ $Y2=0
cc_582 N_A_112_47#_c_553_n N_VGND_c_1312_n 0.00752587f $X=3.05 $Y=0.815 $X2=0
+ $Y2=0
cc_583 N_A_112_47#_c_544_n N_VGND_c_1315_n 0.00316354f $X=8.255 $Y=0.995 $X2=0
+ $Y2=0
cc_584 N_A_112_47#_c_545_n N_VGND_c_1316_n 0.00146448f $X=8.675 $Y=0.995 $X2=0
+ $Y2=0
cc_585 N_A_112_47#_c_546_n N_VGND_c_1316_n 0.00146448f $X=9.095 $Y=0.995 $X2=0
+ $Y2=0
cc_586 N_A_112_47#_c_547_n N_VGND_c_1317_n 0.00316354f $X=9.515 $Y=0.995 $X2=0
+ $Y2=0
cc_587 N_A_112_47#_c_549_n N_VGND_c_1318_n 0.00193763f $X=0.53 $Y=0.82 $X2=0
+ $Y2=0
cc_588 N_A_112_47#_c_579_n N_VGND_c_1318_n 0.0188551f $X=0.695 $Y=0.39 $X2=0
+ $Y2=0
cc_589 N_A_112_47#_c_551_n N_VGND_c_1318_n 0.00198695f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_590 N_A_112_47#_c_551_n N_VGND_c_1320_n 0.00198695f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_591 N_A_112_47#_c_586_n N_VGND_c_1320_n 0.0188551f $X=1.535 $Y=0.39 $X2=0
+ $Y2=0
cc_592 N_A_112_47#_c_552_n N_VGND_c_1320_n 0.00198695f $X=2.21 $Y=0.815 $X2=0
+ $Y2=0
cc_593 N_A_112_47#_c_552_n N_VGND_c_1322_n 0.00198695f $X=2.21 $Y=0.815 $X2=0
+ $Y2=0
cc_594 N_A_112_47#_c_591_n N_VGND_c_1322_n 0.0188551f $X=2.375 $Y=0.39 $X2=0
+ $Y2=0
cc_595 N_A_112_47#_c_553_n N_VGND_c_1322_n 0.00198695f $X=3.05 $Y=0.815 $X2=0
+ $Y2=0
cc_596 N_A_112_47#_c_553_n N_VGND_c_1324_n 0.00198695f $X=3.05 $Y=0.815 $X2=0
+ $Y2=0
cc_597 N_A_112_47#_c_646_n N_VGND_c_1324_n 0.0188551f $X=3.215 $Y=0.39 $X2=0
+ $Y2=0
cc_598 N_A_112_47#_c_544_n N_VGND_c_1330_n 0.00423334f $X=8.255 $Y=0.995 $X2=0
+ $Y2=0
cc_599 N_A_112_47#_c_545_n N_VGND_c_1330_n 0.00424416f $X=8.675 $Y=0.995 $X2=0
+ $Y2=0
cc_600 N_A_112_47#_c_546_n N_VGND_c_1332_n 0.00424416f $X=9.095 $Y=0.995 $X2=0
+ $Y2=0
cc_601 N_A_112_47#_c_547_n N_VGND_c_1332_n 0.00424416f $X=9.515 $Y=0.995 $X2=0
+ $Y2=0
cc_602 N_A_112_47#_M1012_d N_VGND_c_1336_n 0.00215201f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_603 N_A_112_47#_M1028_d N_VGND_c_1336_n 0.00215201f $X=1.4 $Y=0.235 $X2=0
+ $Y2=0
cc_604 N_A_112_47#_M1021_s N_VGND_c_1336_n 0.00215201f $X=2.24 $Y=0.235 $X2=0
+ $Y2=0
cc_605 N_A_112_47#_M1034_s N_VGND_c_1336_n 0.00215201f $X=3.08 $Y=0.235 $X2=0
+ $Y2=0
cc_606 N_A_112_47#_c_544_n N_VGND_c_1336_n 0.00700051f $X=8.255 $Y=0.995 $X2=0
+ $Y2=0
cc_607 N_A_112_47#_c_545_n N_VGND_c_1336_n 0.00573607f $X=8.675 $Y=0.995 $X2=0
+ $Y2=0
cc_608 N_A_112_47#_c_546_n N_VGND_c_1336_n 0.00573607f $X=9.095 $Y=0.995 $X2=0
+ $Y2=0
cc_609 N_A_112_47#_c_547_n N_VGND_c_1336_n 0.00679692f $X=9.515 $Y=0.995 $X2=0
+ $Y2=0
cc_610 N_A_112_47#_c_549_n N_VGND_c_1336_n 0.004202f $X=0.53 $Y=0.82 $X2=0 $Y2=0
cc_611 N_A_112_47#_c_550_n N_VGND_c_1336_n 7.18354e-19 $X=0.255 $Y=0.82 $X2=0
+ $Y2=0
cc_612 N_A_112_47#_c_579_n N_VGND_c_1336_n 0.0122069f $X=0.695 $Y=0.39 $X2=0
+ $Y2=0
cc_613 N_A_112_47#_c_551_n N_VGND_c_1336_n 0.00835832f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_614 N_A_112_47#_c_586_n N_VGND_c_1336_n 0.0122069f $X=1.535 $Y=0.39 $X2=0
+ $Y2=0
cc_615 N_A_112_47#_c_552_n N_VGND_c_1336_n 0.00835832f $X=2.21 $Y=0.815 $X2=0
+ $Y2=0
cc_616 N_A_112_47#_c_591_n N_VGND_c_1336_n 0.0122069f $X=2.375 $Y=0.39 $X2=0
+ $Y2=0
cc_617 N_A_112_47#_c_553_n N_VGND_c_1336_n 0.00835832f $X=3.05 $Y=0.815 $X2=0
+ $Y2=0
cc_618 N_A_112_47#_c_646_n N_VGND_c_1336_n 0.0122069f $X=3.215 $Y=0.39 $X2=0
+ $Y2=0
cc_619 N_A_112_47#_c_569_n N_A_806_47#_c_1489_n 3.15059e-19 $X=7.445 $Y=1.53
+ $X2=0 $Y2=0
cc_620 N_A_112_47#_c_544_n N_A_806_47#_c_1491_n 6.15638e-19 $X=8.255 $Y=0.995
+ $X2=0 $Y2=0
cc_621 N_A_112_47#_c_555_n N_A_806_47#_c_1491_n 0.00872176f $X=7.71 $Y=1.19
+ $X2=0 $Y2=0
cc_622 N_A_112_47#_c_571_n N_A_806_47#_c_1491_n 5.92311e-19 $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_623 N_A_112_47#_c_572_n N_A_806_47#_c_1491_n 0.00341172f $X=7.59 $Y=1.53
+ $X2=0 $Y2=0
cc_624 N_A_112_47#_c_544_n N_A_806_47#_c_1492_n 0.00308231f $X=8.255 $Y=0.995
+ $X2=0 $Y2=0
cc_625 N_A_27_297#_c_820_n N_VPWR_M1004_d 0.00318567f $X=0.99 $Y=1.895 $X2=-0.19
+ $Y2=1.305
cc_626 N_A_27_297#_c_822_n N_VPWR_M1025_d 0.00318567f $X=1.83 $Y=1.895 $X2=0
+ $Y2=0
cc_627 N_A_27_297#_c_820_n N_VPWR_c_880_n 0.0123861f $X=0.99 $Y=1.895 $X2=0
+ $Y2=0
cc_628 N_A_27_297#_c_822_n N_VPWR_c_881_n 0.0123861f $X=1.83 $Y=1.895 $X2=0
+ $Y2=0
cc_629 N_A_27_297#_c_822_n N_VPWR_c_888_n 0.00223194f $X=1.83 $Y=1.895 $X2=0
+ $Y2=0
cc_630 N_A_27_297#_c_825_n N_VPWR_c_888_n 0.0330174f $X=2.67 $Y=2.38 $X2=0 $Y2=0
cc_631 N_A_27_297#_c_856_p N_VPWR_c_888_n 0.0143053f $X=2.08 $Y=2.38 $X2=0 $Y2=0
cc_632 N_A_27_297#_c_815_n N_VPWR_c_888_n 0.0489446f $X=3.51 $Y=2.38 $X2=0 $Y2=0
cc_633 N_A_27_297#_c_849_n N_VPWR_c_888_n 0.0137033f $X=2.795 $Y=2.3 $X2=0 $Y2=0
cc_634 N_A_27_297#_c_820_n N_VPWR_c_890_n 0.00223194f $X=0.99 $Y=1.895 $X2=0
+ $Y2=0
cc_635 N_A_27_297#_c_816_n N_VPWR_c_890_n 0.0204751f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_636 N_A_27_297#_c_820_n N_VPWR_c_891_n 0.00223194f $X=0.99 $Y=1.895 $X2=0
+ $Y2=0
cc_637 N_A_27_297#_c_822_n N_VPWR_c_891_n 0.00223194f $X=1.83 $Y=1.895 $X2=0
+ $Y2=0
cc_638 N_A_27_297#_c_848_n N_VPWR_c_891_n 0.0142343f $X=1.115 $Y=1.96 $X2=0
+ $Y2=0
cc_639 N_A_27_297#_M1004_s N_VPWR_c_879_n 0.00225153f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_640 N_A_27_297#_M1018_s N_VPWR_c_879_n 0.00222276f $X=0.98 $Y=1.485 $X2=0
+ $Y2=0
cc_641 N_A_27_297#_M1038_s N_VPWR_c_879_n 0.00219542f $X=1.82 $Y=1.485 $X2=0
+ $Y2=0
cc_642 N_A_27_297#_M1006_d N_VPWR_c_879_n 0.00213597f $X=2.66 $Y=1.485 $X2=0
+ $Y2=0
cc_643 N_A_27_297#_M1026_d N_VPWR_c_879_n 0.0020932f $X=3.5 $Y=1.485 $X2=0 $Y2=0
cc_644 N_A_27_297#_c_820_n N_VPWR_c_879_n 0.00843576f $X=0.99 $Y=1.895 $X2=0
+ $Y2=0
cc_645 N_A_27_297#_c_822_n N_VPWR_c_879_n 0.00843576f $X=1.83 $Y=1.895 $X2=0
+ $Y2=0
cc_646 N_A_27_297#_c_825_n N_VPWR_c_879_n 0.0204667f $X=2.67 $Y=2.38 $X2=0 $Y2=0
cc_647 N_A_27_297#_c_856_p N_VPWR_c_879_n 0.00962794f $X=2.08 $Y=2.38 $X2=0
+ $Y2=0
cc_648 N_A_27_297#_c_815_n N_VPWR_c_879_n 0.0300909f $X=3.51 $Y=2.38 $X2=0 $Y2=0
cc_649 N_A_27_297#_c_816_n N_VPWR_c_879_n 0.0120542f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_650 N_A_27_297#_c_848_n N_VPWR_c_879_n 0.00955092f $X=1.115 $Y=1.96 $X2=0
+ $Y2=0
cc_651 N_A_27_297#_c_849_n N_VPWR_c_879_n 0.00938745f $X=2.795 $Y=2.3 $X2=0
+ $Y2=0
cc_652 N_A_27_297#_c_815_n N_A_806_297#_c_1039_n 0.0100846f $X=3.51 $Y=2.38
+ $X2=0 $Y2=0
cc_653 N_A_27_297#_c_824_n N_A_806_297#_c_1039_n 0.0282783f $X=3.635 $Y=1.96
+ $X2=0 $Y2=0
cc_654 N_VPWR_c_879_n N_A_806_297#_M1000_d 0.00212053f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_655 N_VPWR_c_879_n N_A_806_297#_M1002_d 0.00222276f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_879_n N_A_806_297#_M1027_d 0.00222276f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_879_n N_A_806_297#_M1019_d 0.00222276f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_879_n N_A_806_297#_M1039_d 0.00213659f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_879_n N_A_806_297#_M1001_s 0.00215203f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_879_n N_A_806_297#_M1022_s 0.00246446f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_661 N_VPWR_M1000_s N_A_806_297#_c_1043_n 0.00304824f $X=4.44 $Y=1.485 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_882_n N_A_806_297#_c_1043_n 0.0120197f $X=4.575 $Y=2.34 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_883_n N_A_806_297#_c_1043_n 0.00223194f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_888_n N_A_806_297#_c_1043_n 0.00223194f $X=4.45 $Y=2.72 $X2=0
+ $Y2=0
cc_665 N_VPWR_c_879_n N_A_806_297#_c_1043_n 0.00843576f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_666 N_VPWR_M1008_s N_A_806_297#_c_1044_n 0.00304824f $X=5.28 $Y=1.485 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_883_n N_A_806_297#_c_1044_n 0.00223194f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_884_n N_A_806_297#_c_1044_n 0.0120197f $X=5.415 $Y=2.34 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_885_n N_A_806_297#_c_1044_n 0.00223194f $X=6.13 $Y=2.72 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_879_n N_A_806_297#_c_1044_n 0.00843576f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_671 N_VPWR_M1009_s N_A_806_297#_c_1045_n 0.00383085f $X=6.12 $Y=1.485 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_885_n N_A_806_297#_c_1045_n 0.00223194f $X=6.13 $Y=2.72 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_886_n N_A_806_297#_c_1045_n 0.0120197f $X=6.255 $Y=2.34 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_892_n N_A_806_297#_c_1045_n 0.00223194f $X=6.97 $Y=2.72 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_879_n N_A_806_297#_c_1045_n 0.00843576f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_676 N_VPWR_M1033_s N_A_806_297#_c_1055_n 0.00383085f $X=6.96 $Y=1.485 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_887_n N_A_806_297#_c_1055_n 0.0120197f $X=7.095 $Y=2.34 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_892_n N_A_806_297#_c_1055_n 0.00223194f $X=6.97 $Y=2.72 $X2=0
+ $Y2=0
cc_679 N_VPWR_c_893_n N_A_806_297#_c_1055_n 0.00223194f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_680 N_VPWR_c_879_n N_A_806_297#_c_1055_n 0.00843576f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_681 N_VPWR_c_893_n N_A_806_297#_c_1038_n 0.0424325f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_682 N_VPWR_c_879_n N_A_806_297#_c_1038_n 0.0253118f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_683 N_VPWR_c_893_n N_A_806_297#_c_1118_n 0.0159427f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_684 N_VPWR_c_879_n N_A_806_297#_c_1118_n 0.00962794f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_685 N_VPWR_c_893_n N_A_806_297#_c_1082_n 0.0473107f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_686 N_VPWR_c_879_n N_A_806_297#_c_1082_n 0.0300869f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_687 N_VPWR_c_888_n N_A_806_297#_c_1039_n 0.0158369f $X=4.45 $Y=2.72 $X2=0
+ $Y2=0
cc_688 N_VPWR_c_879_n N_A_806_297#_c_1039_n 0.00955092f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_689 N_VPWR_c_883_n N_A_806_297#_c_1060_n 0.0142343f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_879_n N_A_806_297#_c_1060_n 0.00955092f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_885_n N_A_806_297#_c_1061_n 0.0142343f $X=6.13 $Y=2.72 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_879_n N_A_806_297#_c_1061_n 0.00955092f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_892_n N_A_806_297#_c_1128_n 0.0142343f $X=6.97 $Y=2.72 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_879_n N_A_806_297#_c_1128_n 0.00955092f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_893_n N_A_806_297#_c_1130_n 0.014244f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_879_n N_A_806_297#_c_1130_n 0.00960883f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_697 N_VPWR_c_879_n N_X_M1001_d 0.00218346f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_698 N_VPWR_c_879_n N_X_M1016_d 0.00216833f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_699 N_VPWR_c_879_n N_X_M1035_d 0.00260431f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_700 N_VPWR_c_893_n X 0.0290717f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_701 N_VPWR_c_879_n X 0.0166756f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_702 N_A_806_297#_c_1038_n N_X_M1001_d 0.00510164f $X=8.34 $Y=2.38 $X2=0 $Y2=0
cc_703 N_A_806_297#_c_1082_n N_X_M1016_d 0.00312348f $X=9.18 $Y=2.38 $X2=0 $Y2=0
cc_704 N_A_806_297#_c_1037_n N_X_c_1157_n 0.0147657f $X=7.515 $Y=2.005 $X2=0
+ $Y2=0
cc_705 N_A_806_297#_c_1080_n N_X_c_1157_n 0.00740213f $X=7.515 $Y=2.295 $X2=0
+ $Y2=0
cc_706 N_A_806_297#_c_1038_n N_X_c_1157_n 0.0185233f $X=8.34 $Y=2.38 $X2=0 $Y2=0
cc_707 N_A_806_297#_M1001_s N_X_c_1158_n 0.00167154f $X=8.33 $Y=1.485 $X2=0
+ $Y2=0
cc_708 N_A_806_297#_c_1038_n N_X_c_1158_n 0.00347015f $X=8.34 $Y=2.38 $X2=0
+ $Y2=0
cc_709 N_A_806_297#_c_1139_p N_X_c_1158_n 0.0128373f $X=8.465 $Y=2 $X2=0 $Y2=0
cc_710 N_A_806_297#_c_1082_n N_X_c_1158_n 0.00347015f $X=9.18 $Y=2.38 $X2=0
+ $Y2=0
cc_711 N_A_806_297#_M1022_s N_X_c_1159_n 0.00166124f $X=9.17 $Y=1.485 $X2=0
+ $Y2=0
cc_712 N_A_806_297#_c_1082_n N_X_c_1159_n 0.00322336f $X=9.18 $Y=2.38 $X2=0
+ $Y2=0
cc_713 N_A_806_297#_c_1143_p N_X_c_1159_n 0.0127256f $X=9.305 $Y=1.96 $X2=0
+ $Y2=0
cc_714 N_A_806_297#_c_1082_n N_X_c_1161_n 0.0118865f $X=9.18 $Y=2.38 $X2=0 $Y2=0
cc_715 N_X_c_1148_n N_VGND_M1024_d 0.00316909f $X=8.3 $Y=0.83 $X2=0 $Y2=0
cc_716 N_X_c_1145_n N_VGND_M1031_d 0.00165819f $X=9.14 $Y=0.82 $X2=0 $Y2=0
cc_717 N_X_c_1146_n N_VGND_M1037_d 0.00379521f $X=9.735 $Y=0.82 $X2=0 $Y2=0
cc_718 N_X_c_1155_n N_VGND_c_1312_n 0.0128219f $X=5.15 $Y=0.79 $X2=0 $Y2=0
cc_719 N_X_c_1151_n N_VGND_c_1313_n 8.00522e-19 $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_720 N_X_c_1151_n N_VGND_c_1314_n 8.00522e-19 $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_721 N_X_c_1148_n N_VGND_c_1315_n 0.01153f $X=8.3 $Y=0.83 $X2=0 $Y2=0
cc_722 N_X_c_1154_n N_VGND_c_1315_n 8.69875e-19 $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_723 N_X_c_1145_n N_VGND_c_1316_n 0.0116528f $X=9.14 $Y=0.82 $X2=0 $Y2=0
cc_724 N_X_c_1146_n N_VGND_c_1317_n 0.012644f $X=9.735 $Y=0.82 $X2=0 $Y2=0
cc_725 N_X_c_1148_n N_VGND_c_1328_n 0.00166406f $X=8.3 $Y=0.83 $X2=0 $Y2=0
cc_726 N_X_c_1203_n N_VGND_c_1330_n 0.018856f $X=8.465 $Y=0.39 $X2=0 $Y2=0
cc_727 N_X_c_1145_n N_VGND_c_1330_n 0.00193763f $X=9.14 $Y=0.82 $X2=0 $Y2=0
cc_728 N_X_c_1148_n N_VGND_c_1330_n 0.00200317f $X=8.3 $Y=0.83 $X2=0 $Y2=0
cc_729 N_X_c_1145_n N_VGND_c_1332_n 0.00193763f $X=9.14 $Y=0.82 $X2=0 $Y2=0
cc_730 N_X_c_1214_n N_VGND_c_1332_n 0.0188551f $X=9.305 $Y=0.39 $X2=0 $Y2=0
cc_731 N_X_c_1146_n N_VGND_c_1332_n 0.00193763f $X=9.735 $Y=0.82 $X2=0 $Y2=0
cc_732 N_X_c_1146_n N_VGND_c_1335_n 0.00369499f $X=9.735 $Y=0.82 $X2=0 $Y2=0
cc_733 N_X_M1010_s N_VGND_c_1336_n 0.00216833f $X=4.44 $Y=0.235 $X2=0 $Y2=0
cc_734 N_X_M1014_s N_VGND_c_1336_n 0.00174764f $X=5.28 $Y=0.235 $X2=0 $Y2=0
cc_735 N_X_M1024_s N_VGND_c_1336_n 0.00215201f $X=8.33 $Y=0.235 $X2=0 $Y2=0
cc_736 N_X_M1032_s N_VGND_c_1336_n 0.00215201f $X=9.17 $Y=0.235 $X2=0 $Y2=0
cc_737 N_X_c_1203_n N_VGND_c_1336_n 0.0122071f $X=8.465 $Y=0.39 $X2=0 $Y2=0
cc_738 N_X_c_1145_n N_VGND_c_1336_n 0.00827287f $X=9.14 $Y=0.82 $X2=0 $Y2=0
cc_739 N_X_c_1214_n N_VGND_c_1336_n 0.0122069f $X=9.305 $Y=0.39 $X2=0 $Y2=0
cc_740 N_X_c_1146_n N_VGND_c_1336_n 0.0108275f $X=9.735 $Y=0.82 $X2=0 $Y2=0
cc_741 N_X_c_1148_n N_VGND_c_1336_n 0.00461222f $X=8.3 $Y=0.83 $X2=0 $Y2=0
cc_742 N_X_c_1151_n N_VGND_c_1336_n 0.11241f $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_743 N_X_c_1152_n N_VGND_c_1336_n 0.0144123f $X=5.435 $Y=0.85 $X2=0 $Y2=0
cc_744 N_X_c_1154_n N_VGND_c_1336_n 0.0137327f $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_745 N_X_c_1155_n N_A_806_47#_M1010_d 0.0040802f $X=5.15 $Y=0.79 $X2=-0.19
+ $Y2=-0.24
cc_746 N_X_c_1155_n N_A_806_47#_M1013_d 0.00162317f $X=5.15 $Y=0.79 $X2=0 $Y2=0
cc_747 N_X_c_1151_n N_A_806_47#_M1020_d 3.83093e-19 $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_748 N_X_M1010_s N_A_806_47#_c_1488_n 0.00305026f $X=4.44 $Y=0.235 $X2=0 $Y2=0
cc_749 N_X_M1014_s N_A_806_47#_c_1488_n 0.00294958f $X=5.28 $Y=0.235 $X2=0 $Y2=0
cc_750 N_X_c_1151_n N_A_806_47#_c_1488_n 0.00259909f $X=7.905 $Y=0.85 $X2=0
+ $Y2=0
cc_751 N_X_c_1152_n N_A_806_47#_c_1488_n 0.00100468f $X=5.435 $Y=0.85 $X2=0
+ $Y2=0
cc_752 N_X_c_1155_n N_A_806_47#_c_1488_n 0.0696782f $X=5.15 $Y=0.79 $X2=0 $Y2=0
cc_753 N_X_c_1151_n N_A_806_47#_c_1489_n 0.014335f $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_754 N_X_c_1152_n N_A_806_47#_c_1489_n 2.69214e-19 $X=5.435 $Y=0.85 $X2=0
+ $Y2=0
cc_755 N_X_c_1153_n N_A_806_47#_c_1489_n 0.00916987f $X=5.29 $Y=0.85 $X2=0 $Y2=0
cc_756 N_X_c_1151_n N_A_806_47#_c_1490_n 0.0163519f $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_757 N_X_c_1148_n N_A_806_47#_c_1491_n 0.014034f $X=8.3 $Y=0.83 $X2=0 $Y2=0
cc_758 N_X_c_1151_n N_A_806_47#_c_1491_n 0.0336415f $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_759 N_X_c_1154_n N_A_806_47#_c_1491_n 3.29239e-19 $X=8.05 $Y=0.85 $X2=0 $Y2=0
cc_760 N_X_c_1203_n N_A_806_47#_c_1492_n 0.00502037f $X=8.465 $Y=0.39 $X2=0
+ $Y2=0
cc_761 N_X_c_1151_n N_A_806_47#_c_1493_n 0.0144518f $X=7.905 $Y=0.85 $X2=0 $Y2=0
cc_762 N_VGND_c_1336_n N_A_806_47#_M1010_d 0.00209344f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_763 N_VGND_c_1336_n N_A_806_47#_M1013_d 0.00215227f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_764 N_VGND_c_1336_n N_A_806_47#_M1020_d 0.00177027f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_765 N_VGND_c_1336_n N_A_806_47#_M1011_s 0.00177024f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_766 N_VGND_c_1336_n N_A_806_47#_M1023_s 0.00172424f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_767 N_VGND_c_1312_n N_A_806_47#_c_1488_n 0.0190115f $X=3.635 $Y=0.39 $X2=0
+ $Y2=0
cc_768 N_VGND_c_1334_n N_A_806_47#_c_1488_n 0.0991765f $X=6.17 $Y=0 $X2=0 $Y2=0
cc_769 N_VGND_c_1336_n N_A_806_47#_c_1488_n 0.0511951f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_770 N_VGND_c_1334_n N_A_806_47#_c_1494_n 0.0152108f $X=6.17 $Y=0 $X2=0 $Y2=0
cc_771 N_VGND_c_1336_n N_A_806_47#_c_1494_n 0.00447564f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_772 N_VGND_M1005_d N_A_806_47#_c_1490_n 0.00162089f $X=6.12 $Y=0.235 $X2=0
+ $Y2=0
cc_773 N_VGND_c_1313_n N_A_806_47#_c_1490_n 0.0111016f $X=6.255 $Y=0.39 $X2=0
+ $Y2=0
cc_774 N_VGND_c_1326_n N_A_806_47#_c_1490_n 0.00198695f $X=7.01 $Y=0 $X2=0 $Y2=0
cc_775 N_VGND_c_1334_n N_A_806_47#_c_1490_n 0.00198695f $X=6.17 $Y=0 $X2=0 $Y2=0
cc_776 N_VGND_c_1336_n N_A_806_47#_c_1490_n 0.00370618f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_777 N_VGND_c_1326_n N_A_806_47#_c_1504_n 0.0188551f $X=7.01 $Y=0 $X2=0 $Y2=0
cc_778 N_VGND_c_1336_n N_A_806_47#_c_1504_n 0.00580811f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_779 N_VGND_M1015_d N_A_806_47#_c_1491_n 0.00162089f $X=6.96 $Y=0.235 $X2=0
+ $Y2=0
cc_780 N_VGND_c_1314_n N_A_806_47#_c_1491_n 0.0111016f $X=7.095 $Y=0.39 $X2=0
+ $Y2=0
cc_781 N_VGND_c_1326_n N_A_806_47#_c_1491_n 0.00198695f $X=7.01 $Y=0 $X2=0 $Y2=0
cc_782 N_VGND_c_1328_n N_A_806_47#_c_1491_n 0.00198695f $X=7.96 $Y=0 $X2=0 $Y2=0
cc_783 N_VGND_c_1336_n N_A_806_47#_c_1491_n 0.00370618f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_784 N_VGND_c_1315_n N_A_806_47#_c_1492_n 0.016379f $X=8.045 $Y=0.39 $X2=0
+ $Y2=0
cc_785 N_VGND_c_1328_n N_A_806_47#_c_1492_n 0.0209752f $X=7.96 $Y=0 $X2=0 $Y2=0
cc_786 N_VGND_c_1336_n N_A_806_47#_c_1492_n 0.00590515f $X=9.89 $Y=0 $X2=0 $Y2=0

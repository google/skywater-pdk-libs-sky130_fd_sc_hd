* File: sky130_fd_sc_hd__o21bai_2.spice.pex
* Created: Thu Aug 27 14:36:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21BAI_2%B1_N 3 6 8 11 12 13
r30 11 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.16
+ $X2=0.362 $Y2=1.325
r31 11 13 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.16
+ $X2=0.362 $Y2=0.995
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.355
+ $Y=1.16 $X2=0.355 $Y2=1.16
r33 8 12 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.23 $Y=1.16
+ $X2=0.355 $Y2=1.16
r34 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.475 $Y=1.695
+ $X2=0.475 $Y2=1.325
r35 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.675
+ $X2=0.475 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%A_28_297# 1 2 9 13 15 17 18 20 21 24 26 29
+ 32 40 42 48
c74 26 0 1.5158e-19 $X=0.78 $Y=1.495
c75 18 0 1.56657e-19 $X=1.9 $Y=0.995
r76 47 48 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.48 $Y=1.16 $X2=1.9
+ $Y2=1.16
r77 46 47 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.38 $Y=1.16 $X2=1.48
+ $Y2=1.16
r78 38 40 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=0.685 $Y=0.635
+ $X2=0.78 $Y2=0.635
r79 32 35 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.265 $Y=1.58
+ $X2=0.265 $Y2=1.725
r80 30 46 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.38 $Y2=1.16
r81 30 43 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=0.96 $Y2=1.16
r82 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r83 27 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=1.16
+ $X2=0.78 $Y2=1.16
r84 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.865 $Y=1.16
+ $X2=1.17 $Y2=1.16
r85 25 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.245
+ $X2=0.78 $Y2=1.16
r86 25 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.78 $Y=1.245
+ $X2=0.78 $Y2=1.495
r87 24 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.075
+ $X2=0.78 $Y2=1.16
r88 23 40 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.78 $Y=0.825
+ $X2=0.78 $Y2=0.635
r89 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.78 $Y=0.825
+ $X2=0.78 $Y2=1.075
r90 22 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.58
+ $X2=0.265 $Y2=1.58
r91 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.695 $Y=1.58
+ $X2=0.78 $Y2=1.495
r92 21 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.695 $Y=1.58
+ $X2=0.35 $Y2=1.58
r93 18 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=1.16
r94 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995 $X2=1.9
+ $Y2=0.56
r95 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.16
r96 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=0.56
r97 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.325
+ $X2=1.38 $Y2=1.16
r98 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.38 $Y=1.325
+ $X2=1.38 $Y2=1.985
r99 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.325
+ $X2=0.96 $Y2=1.16
r100 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.96 $Y=1.325
+ $X2=0.96 $Y2=1.985
r101 2 35 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.725
r102 1 38 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.465 $X2=0.685 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%A2 1 3 6 8 10 13 15 22
c52 22 0 1.26413e-19 $X=2.74 $Y=1.16
c53 1 0 8.54869e-20 $X=2.32 $Y=0.995
r54 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.53 $Y=1.16
+ $X2=2.74 $Y2=1.16
r55 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.32 $Y=1.16
+ $X2=2.53 $Y2=1.16
r56 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.16 $X2=2.53 $Y2=1.16
r57 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.325
+ $X2=2.74 $Y2=1.16
r58 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.74 $Y=1.325
+ $X2=2.74 $Y2=1.985
r59 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=0.995
+ $X2=2.74 $Y2=1.16
r60 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.74 $Y=0.995
+ $X2=2.74 $Y2=0.56
r61 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.325
+ $X2=2.32 $Y2=1.16
r62 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.32 $Y=1.325 $X2=2.32
+ $Y2=1.985
r63 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=0.995
+ $X2=2.32 $Y2=1.16
r64 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.32 $Y=0.995 $X2=2.32
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%A1 1 3 6 8 10 13 15 22
c38 15 0 1.26413e-19 $X=3.45 $Y=1.19
r39 20 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=3.425 $Y=1.16
+ $X2=3.58 $Y2=1.16
r40 17 20 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=3.16 $Y=1.16
+ $X2=3.425 $Y2=1.16
r41 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.16 $X2=3.425 $Y2=1.16
r42 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.325
+ $X2=3.58 $Y2=1.16
r43 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.58 $Y=1.325
+ $X2=3.58 $Y2=1.985
r44 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=0.995
+ $X2=3.58 $Y2=1.16
r45 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.58 $Y=0.995
+ $X2=3.58 $Y2=0.56
r46 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=1.325
+ $X2=3.16 $Y2=1.16
r47 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.16 $Y=1.325 $X2=3.16
+ $Y2=1.985
r48 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=0.995
+ $X2=3.16 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.16 $Y=0.995 $X2=3.16
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%VPWR 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
c61 2 0 1.3066e-19 $X=1.455 $Y=1.485
c62 1 0 1.5158e-19 $X=0.55 $Y=1.485
r63 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r64 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r65 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 45 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.37 $Y2=2.72
r69 42 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 41 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r71 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r72 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 37 40 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r76 35 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.72 $Y=2.72
+ $X2=1.595 $Y2=2.72
r77 35 37 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.72 $Y=2.72
+ $X2=2.07 $Y2=2.72
r78 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=3.37 $Y2=2.72
r79 34 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=2.99 $Y2=2.72
r80 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.75 $Y2=2.72
r84 30 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 29 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.595 $Y2=2.72
r86 29 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.47 $Y=2.72 $X2=1.15
+ $Y2=2.72
r87 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=2.72
+ $X2=0.75 $Y2=2.72
r88 24 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.585 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=2.635
+ $X2=3.37 $Y2=2.72
r92 18 20 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.37 $Y=2.635
+ $X2=3.37 $Y2=2
r93 14 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=2.635
+ $X2=1.595 $Y2=2.72
r94 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.595 $Y=2.635
+ $X2=1.595 $Y2=1.96
r95 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r96 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r97 3 20 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.235
+ $Y=1.485 $X2=3.37 $Y2=2
r98 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.455
+ $Y=1.485 $X2=1.59 $Y2=1.96
r99 1 12 300 $w=1.7e-07 $l=5.66238e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%Y 1 2 3 12 16 20 22 25 28
c43 28 0 1.3066e-19 $X=1.61 $Y=1.53
c44 25 0 8.54869e-20 $X=1.69 $Y=0.73
r45 27 28 15.8578 $w=4.23e-07 $l=5.4e-07 $layer=LI1_cond $X=1.652 $Y=0.905
+ $X2=1.652 $Y2=1.445
r46 25 27 6.73672 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.69 $Y=0.73
+ $X2=1.69 $Y2=0.905
r47 22 28 10.5913 $w=3.38e-07 $l=2.7e-07 $layer=LI1_cond $X=1.255 $Y=1.53
+ $X2=1.525 $Y2=1.53
r48 18 20 0.235192 $w=2.43e-07 $l=5e-09 $layer=LI1_cond $X=2.527 $Y=1.615
+ $X2=2.527 $Y2=1.62
r49 17 28 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.78 $Y=1.53
+ $X2=1.652 $Y2=1.53
r50 16 18 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.405 $Y=1.53
+ $X2=2.527 $Y2=1.615
r51 16 17 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.405 $Y=1.53
+ $X2=1.78 $Y2=1.53
r52 12 14 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=1.62
+ $X2=1.17 $Y2=2.3
r53 10 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.17 $Y=1.615
+ $X2=1.255 $Y2=1.53
r54 10 12 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.62
r55 3 20 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.395
+ $Y=1.485 $X2=2.53 $Y2=1.62
r56 2 14 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.485 $X2=1.17 $Y2=2.3
r57 2 12 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.485 $X2=1.17 $Y2=1.62
r58 1 25 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%A_397_297# 1 2 3 12 14 15 16 17 18 20 22
r38 20 29 3.02719 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=3.842 $Y=1.665
+ $X2=3.842 $Y2=1.56
r39 20 22 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=3.842 $Y=1.665
+ $X2=3.842 $Y2=2.3
r40 19 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=1.56
+ $X2=2.95 $Y2=1.56
r41 18 29 3.94976 $w=2.1e-07 $l=1.37e-07 $layer=LI1_cond $X=3.705 $Y=1.56
+ $X2=3.842 $Y2=1.56
r42 18 19 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=3.705 $Y=1.56
+ $X2=3.035 $Y2=1.56
r43 17 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=2.295
+ $X2=2.95 $Y2=2.38
r44 16 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.95 $Y=1.665
+ $X2=2.95 $Y2=1.56
r45 16 17 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.95 $Y=1.665
+ $X2=2.95 $Y2=2.295
r46 14 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=2.38
+ $X2=2.95 $Y2=2.38
r47 14 15 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.865 $Y=2.38
+ $X2=2.235 $Y2=2.38
r48 10 15 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.095 $Y=2.295
+ $X2=2.235 $Y2=2.38
r49 10 12 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.095 $Y=2.295
+ $X2=2.095 $Y2=1.96
r50 3 29 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.655
+ $Y=1.485 $X2=3.79 $Y2=1.62
r51 3 22 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.655
+ $Y=1.485 $X2=3.79 $Y2=2.3
r52 2 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.485 $X2=2.95 $Y2=2.3
r53 2 25 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.485 $X2=2.95 $Y2=1.62
r54 1 12 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=1.985
+ $Y=1.485 $X2=2.11 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%VGND 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r59 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r60 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r61 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r62 38 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r63 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r64 35 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.53
+ $Y2=0
r65 35 37 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.99
+ $Y2=0
r66 34 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r67 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r68 31 34 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r69 30 33 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r70 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r71 28 44 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.175
+ $Y2=0
r72 28 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.69
+ $Y2=0
r73 27 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.53
+ $Y2=0
r74 27 33 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.07
+ $Y2=0
r75 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r76 25 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r77 23 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.285 $Y=0 $X2=2.99
+ $Y2=0
r78 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.37
+ $Y2=0
r79 22 40 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.91
+ $Y2=0
r80 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.37
+ $Y2=0
r81 18 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=0.085
+ $X2=3.37 $Y2=0
r82 18 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.37 $Y=0.085
+ $X2=3.37 $Y2=0.39
r83 14 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0
r84 14 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0.39
r85 10 44 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.175 $Y2=0
r86 10 12 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.66
r87 3 20 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.235 $X2=3.37 $Y2=0.39
r88 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.53 $Y2=0.39
r89 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.465 $X2=0.265 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BAI_2%A_229_47# 1 2 3 4 13 15 17 19 20 21 25 27
+ 31 39
c70 20 0 1.56657e-19 $X=2.15 $Y=0.725
r71 29 31 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=3.802 $Y=0.725
+ $X2=3.802 $Y2=0.39
r72 28 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0.815
+ $X2=2.95 $Y2=0.815
r73 27 29 7.81092 $w=1.8e-07 $l=2.17391e-07 $layer=LI1_cond $X=3.625 $Y=0.815
+ $X2=3.802 $Y2=0.725
r74 27 28 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.625 $Y=0.815
+ $X2=3.115 $Y2=0.815
r75 23 39 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.95 $Y=0.725 $X2=2.95
+ $Y2=0.815
r76 23 25 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.95 $Y=0.725
+ $X2=2.95 $Y2=0.39
r77 22 38 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.275 $Y=0.815
+ $X2=2.15 $Y2=0.815
r78 21 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.785 $Y=0.815
+ $X2=2.95 $Y2=0.815
r79 21 22 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.785 $Y=0.815
+ $X2=2.275 $Y2=0.815
r80 20 38 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.15 $Y=0.725 $X2=2.15
+ $Y2=0.815
r81 19 36 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2.15 $Y=0.475
+ $X2=2.15 $Y2=0.365
r82 19 20 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.15 $Y=0.475
+ $X2=2.15 $Y2=0.725
r83 18 34 3.88917 $w=2.2e-07 $l=1.4e-07 $layer=LI1_cond $X=1.355 $Y=0.365
+ $X2=1.215 $Y2=0.365
r84 17 36 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=0.365
+ $X2=2.15 $Y2=0.365
r85 17 18 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=0.365
+ $X2=1.355 $Y2=0.365
r86 13 34 3.05577 $w=2.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.215 $Y=0.475
+ $X2=1.215 $Y2=0.365
r87 13 15 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=1.215 $Y=0.475
+ $X2=1.215 $Y2=0.73
r88 4 31 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.655
+ $Y=0.235 $X2=3.79 $Y2=0.39
r89 3 25 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.815
+ $Y=0.235 $X2=2.95 $Y2=0.39
r90 2 38 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.73
r91 2 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.39
r92 1 34 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.235 $X2=1.27 $Y2=0.39
r93 1 15 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.235 $X2=1.27 $Y2=0.73
.ends


* File: sky130_fd_sc_hd__dlrbn_2.pex.spice
* Created: Thu Aug 27 14:16:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRBN_2%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.35704e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%A_27_47# 1 2 9 13 17 20 24 28 29 30 38 42 45
+ 47 52 54 56 57 60 63 64 68 71 75 79
c168 20 0 1.41946e-19 $X=3.335 $Y=2.275
c169 13 0 2.67852e-20 $X=0.89 $Y=2.135
c170 9 0 2.67852e-20 $X=0.89 $Y=0.445
r171 64 79 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.095 $Y=1.53
+ $X2=3.095 $Y2=1.415
r172 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.53
+ $X2=3.015 $Y2=1.53
r173 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r175 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=3.015 $Y2=1.53
r176 56 57 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=0.84 $Y2=1.53
r177 52 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=0.87
+ $X2=2.8 $Y2=0.705
r178 51 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=0.87
+ $X2=3.01 $Y2=0.87
r179 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=0.87 $X2=2.8 $Y2=0.87
r180 49 60 16.7948 $w=1.73e-07 $l=2.65e-07 $layer=LI1_cond $X=0.692 $Y=1.795
+ $X2=0.692 $Y2=1.53
r181 48 60 8.23896 $w=1.73e-07 $l=1.3e-07 $layer=LI1_cond $X=0.692 $Y=1.4
+ $X2=0.692 $Y2=1.53
r182 46 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r183 45 48 8.86758 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.722 $Y=1.235
+ $X2=0.722 $Y2=1.4
r184 45 47 8.86758 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.722 $Y=1.235
+ $X2=0.722 $Y2=1.07
r185 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r186 39 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.335 $Y2=1.74
r187 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r188 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.53
r189 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.74
r190 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=0.87
r191 34 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=1.415
r192 32 47 16.7948 $w=1.73e-07 $l=2.65e-07 $layer=LI1_cond $X=0.692 $Y=0.805
+ $X2=0.692 $Y2=1.07
r193 31 42 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r194 30 49 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.692 $Y2=1.795
r195 30 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.345 $Y2=1.88
r196 28 32 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.692 $Y2=0.805
r197 28 29 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.345 $Y2=0.72
r198 22 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r199 22 24 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r200 18 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=1.74
r201 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=2.275
r202 17 71 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.79 $Y=0.415
+ $X2=2.79 $Y2=0.705
r203 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r204 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r205 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r206 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r207 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r208 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%A_299_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c83 32 0 1.12109e-19 $X=2.255 $Y=0.93
c84 18 0 7.13094e-20 $X=1.97 $Y=0.7
r85 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=1.095
r86 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=0.765
r87 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r88 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r89 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.155 $Y2=0.93
r90 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.055 $Y2=1.495
r91 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=2.055 $Y2=1.495
r92 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=1.785 $Y2=1.58
r93 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r94 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=2.155 $Y2=0.93
r95 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=1.705 $Y2=0.7
r96 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r97 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r98 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=2.165
+ $X2=2.25 $Y2=1.095
r99 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.765
r100 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r101 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%A_193_47# 1 2 9 11 12 15 19 22 24 26 27 30
+ 33 37 38
c112 38 0 1.41946e-19 $X=2.67 $Y=1.52
r113 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r114 34 38 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.612 $Y=1.87
+ $X2=2.612 $Y2=1.52
r115 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.87
+ $X2=2.555 $Y2=1.87
r116 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r117 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r118 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=2.555 $Y2=1.87
r119 26 27 1.37376 $w=1.4e-07 $l=1.11e-06 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=1.3 $Y2=1.87
r120 24 30 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r121 24 25 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r122 22 25 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r123 18 37 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r124 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r125 17 37 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r126 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.22 $Y=1.245
+ $X2=3.22 $Y2=0.415
r127 12 17 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r128 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=3.22 $Y2=1.245
r129 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=2.805 $Y2=1.32
r130 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.73 $Y=2.275
+ $X2=2.73 $Y2=1.685
r131 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r132 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%A_724_21# 1 2 9 13 15 17 20 22 24 27 29 30
+ 31 32 33 35 36 38 42 44 47 49 53 55 60 62 67 69 71
c147 69 0 1.12853e-19 $X=5.535 $Y=1.16
c148 60 0 1.05093e-19 $X=5.395 $Y=1.495
c149 31 0 9.0697e-20 $X=6.77 $Y=1.325
c150 9 0 1.27208e-19 $X=3.695 $Y=0.445
r151 70 80 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=5.535 $Y=1.16
+ $X2=5.95 $Y2=1.16
r152 70 77 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.535 $Y=1.16
+ $X2=5.475 $Y2=1.16
r153 69 72 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=1.16
+ $X2=5.465 $Y2=1.325
r154 69 71 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=1.16
+ $X2=5.465 $Y2=0.995
r155 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.535
+ $Y=1.16 $X2=5.535 $Y2=1.16
r156 62 64 8.3814 $w=2.18e-07 $l=1.6e-07 $layer=LI1_cond $X=4.45 $Y=0.58
+ $X2=4.45 $Y2=0.74
r157 60 72 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.395 $Y=1.495
+ $X2=5.395 $Y2=1.325
r158 57 71 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.395 $Y=0.825
+ $X2=5.395 $Y2=0.995
r159 56 67 3.46198 $w=2.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.93 $Y=1.58
+ $X2=4.845 $Y2=1.68
r160 55 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.31 $Y=1.58
+ $X2=5.395 $Y2=1.495
r161 55 56 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.31 $Y=1.58
+ $X2=4.93 $Y2=1.58
r162 51 67 3.05049 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.845 $Y=1.865
+ $X2=4.845 $Y2=1.68
r163 51 53 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.845 $Y=1.865
+ $X2=4.845 $Y2=2.27
r164 50 64 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.56 $Y=0.74 $X2=4.45
+ $Y2=0.74
r165 49 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.31 $Y=0.74
+ $X2=5.395 $Y2=0.825
r166 49 50 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.31 $Y=0.74
+ $X2=4.56 $Y2=0.74
r167 47 73 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.695 $Y2=1.7
r168 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r169 44 67 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=1.68
+ $X2=4.845 $Y2=1.68
r170 44 46 26.0078 $w=3.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.76 $Y=1.68
+ $X2=3.925 $Y2=1.68
r171 40 42 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=6.77 $Y=1.695
+ $X2=6.9 $Y2=1.695
r172 36 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.9 $Y=1.77 $X2=6.9
+ $Y2=1.695
r173 36 38 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.9 $Y=1.77
+ $X2=6.9 $Y2=2.165
r174 33 35 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.9 $Y=0.73 $X2=6.9
+ $Y2=0.445
r175 32 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.77 $Y=1.62
+ $X2=6.77 $Y2=1.695
r176 31 32 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=6.77 $Y=1.325
+ $X2=6.77 $Y2=1.62
r177 30 80 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.025 $Y=1.16
+ $X2=5.95 $Y2=1.16
r178 29 31 45.3305 $w=1.82e-07 $l=1.94808e-07 $layer=POLY_cond $X=6.835 $Y=1.16
+ $X2=6.77 $Y2=1.325
r179 29 33 115.512 $w=1.82e-07 $l=4.61357e-07 $layer=POLY_cond $X=6.835 $Y=1.16
+ $X2=6.9 $Y2=0.73
r180 29 30 117.157 $w=3.3e-07 $l=6.7e-07 $layer=POLY_cond $X=6.695 $Y=1.16
+ $X2=6.025 $Y2=1.16
r181 25 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.325
+ $X2=5.95 $Y2=1.16
r182 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.95 $Y=1.325
+ $X2=5.95 $Y2=1.985
r183 22 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=0.995
+ $X2=5.95 $Y2=1.16
r184 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.95 $Y=0.995
+ $X2=5.95 $Y2=0.56
r185 18 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.325
+ $X2=5.475 $Y2=1.16
r186 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.475 $Y=1.325
+ $X2=5.475 $Y2=1.985
r187 15 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=0.995
+ $X2=5.475 $Y2=1.16
r188 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.475 $Y=0.995
+ $X2=5.475 $Y2=0.56
r189 11 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=1.7
r190 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=2.275
r191 7 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=1.7
r192 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=0.445
r193 2 67 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.845 $Y2=1.755
r194 2 53 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.845 $Y2=2.27
r195 1 62 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.235 $X2=4.425 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%A_561_413# 1 2 7 9 12 14 15 16 20 25 26 27
+ 30
c81 26 0 1.57048e-19 $X=3.565 $Y=1.325
r82 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.16 $X2=4.115 $Y2=1.16
r83 28 30 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.65 $Y=1.16
+ $X2=4.115 $Y2=1.16
r84 26 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.49 $Y2=1.16
r85 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=2.255
r86 25 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.415 $Y=0.995
+ $X2=3.49 $Y2=1.16
r87 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=0.995
r88 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.565 $Y2=2.255
r89 20 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.065 $Y2=2.34
r90 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r91 16 18 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.005 $Y2=0.45
r92 14 31 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.115 $Y2=1.16
r93 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.635 $Y2=1.16
r94 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=1.325
+ $X2=4.635 $Y2=1.16
r95 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.635 $Y=1.325
+ $X2=4.635 $Y2=1.985
r96 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=0.995
+ $X2=4.635 $Y2=1.16
r97 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.635 $Y=0.995
+ $X2=4.635 $Y2=0.56
r98 2 22 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.065 $X2=3.065 $Y2=2.34
r99 1 18 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3.005 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%RESET_B 1 3 6 8 11 12
c37 12 0 1.27208e-19 $X=5.055 $Y=1.16
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.16 $X2=5.055 $Y2=1.16
r39 8 12 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.875 $Y=1.16
+ $X2=5.055 $Y2=1.16
r40 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.325
+ $X2=5.055 $Y2=1.16
r41 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.055 $Y=1.325
+ $X2=5.055 $Y2=1.985
r42 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=0.995
+ $X2=5.055 $Y2=1.16
r43 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.055 $Y=0.995
+ $X2=5.055 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%A_1313_47# 1 2 7 9 12 14 15 18 22 24 27 31
+ 35 38
c77 14 0 1.35563e-19 $X=7.725 $Y=1.16
r78 36 41 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=7.29 $Y=1.16
+ $X2=7.375 $Y2=1.16
r79 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.29
+ $Y=1.16 $X2=7.29 $Y2=1.16
r80 33 38 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.855 $Y=1.16
+ $X2=6.69 $Y2=1.16
r81 33 35 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.855 $Y=1.16
+ $X2=7.29 $Y2=1.16
r82 29 38 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=1.325
+ $X2=6.69 $Y2=1.16
r83 29 31 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.69 $Y=1.325
+ $X2=6.69 $Y2=2
r84 25 38 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=0.995
+ $X2=6.69 $Y2=1.16
r85 25 27 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=6.69 $Y=0.995
+ $X2=6.69 $Y2=0.51
r86 20 24 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.8 $Y=1.295
+ $X2=7.8 $Y2=1.16
r87 20 22 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.8 $Y=1.295 $X2=7.8
+ $Y2=1.985
r88 16 24 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.8 $Y=1.025
+ $X2=7.8 $Y2=1.16
r89 16 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.8 $Y=1.025
+ $X2=7.8 $Y2=0.56
r90 15 41 15.1926 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.45 $Y=1.16
+ $X2=7.375 $Y2=1.16
r91 14 24 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=7.725 $Y=1.16
+ $X2=7.8 $Y2=1.16
r92 14 15 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=7.725 $Y=1.16
+ $X2=7.45 $Y2=1.16
r93 10 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.375 $Y=1.325
+ $X2=7.375 $Y2=1.16
r94 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.375 $Y=1.325
+ $X2=7.375 $Y2=1.985
r95 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.375 $Y=0.995
+ $X2=7.375 $Y2=1.16
r96 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.375 $Y=0.995
+ $X2=7.375 $Y2=0.56
r97 2 31 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=6.565
+ $Y=1.845 $X2=6.69 $Y2=2
r98 1 27 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.69 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 45 47 52
+ 53 54 56 61 78 82 87 93 96 100 106 108 111 115
c126 5 0 1.05093e-19 $X=5.13 $Y=1.485
r127 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r128 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r129 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r130 105 106 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=2.47
+ $X2=4.59 $Y2=2.47
r131 102 105 0.981855 $w=6.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.37 $Y=2.47
+ $X2=4.425 $Y2=2.47
r132 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 99 102 8.30114 $w=6.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.905 $Y=2.47
+ $X2=4.37 $Y2=2.47
r134 99 100 9.18355 $w=6.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=2.47
+ $X2=3.82 $Y2=2.47
r135 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r137 91 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r138 91 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r139 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r140 88 111 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.33 $Y=2.72
+ $X2=7.182 $Y2=2.72
r141 88 90 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.33 $Y=2.72
+ $X2=7.59 $Y2=2.72
r142 87 114 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.925 $Y=2.72
+ $X2=8.102 $Y2=2.72
r143 87 90 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.925 $Y=2.72
+ $X2=7.59 $Y2=2.72
r144 86 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r145 86 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r146 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r147 83 108 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.355 $Y=2.72
+ $X2=6.22 $Y2=2.72
r148 83 85 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.355 $Y=2.72
+ $X2=6.67 $Y2=2.72
r149 82 111 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=7.182 $Y2=2.72
r150 82 85 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=6.67 $Y2=2.72
r151 81 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r152 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r153 78 108 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=6.22 $Y2=2.72
r154 78 80 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=5.75 $Y2=2.72
r155 77 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r156 77 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r157 76 106 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=4.59 $Y2=2.72
r158 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r159 73 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r160 72 100 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.82 $Y2=2.72
r161 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r162 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r163 70 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r164 69 72 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r165 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r166 67 96 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r167 67 69 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r168 65 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r169 65 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r170 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r171 62 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r172 62 64 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r173 61 96 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r174 61 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r175 56 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r176 56 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r177 54 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r178 54 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r179 52 76 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.1 $Y=2.72 $X2=4.83
+ $Y2=2.72
r180 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=2.72
+ $X2=5.225 $Y2=2.72
r181 51 80 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.35 $Y=2.72 $X2=5.75
+ $Y2=2.72
r182 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.35 $Y=2.72
+ $X2=5.225 $Y2=2.72
r183 47 50 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.06 $Y=1.66
+ $X2=8.06 $Y2=2.34
r184 45 114 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=8.06 $Y=2.635
+ $X2=8.102 $Y2=2.72
r185 45 50 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.06 $Y=2.635
+ $X2=8.06 $Y2=2.34
r186 41 111 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.182 $Y=2.635
+ $X2=7.182 $Y2=2.72
r187 41 43 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=7.182 $Y=2.635
+ $X2=7.182 $Y2=2
r188 37 108 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2.72
r189 37 39 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2
r190 33 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=2.635
+ $X2=5.225 $Y2=2.72
r191 33 35 28.3501 $w=2.48e-07 $l=6.15e-07 $layer=LI1_cond $X=5.225 $Y=2.635
+ $X2=5.225 $Y2=2.02
r192 29 96 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r193 29 31 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r194 25 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r195 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r196 8 50 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.485 $X2=8.01 $Y2=2.34
r197 8 47 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.485 $X2=8.01 $Y2=1.66
r198 7 43 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=6.975
+ $Y=1.845 $X2=7.165 $Y2=2
r199 6 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.025
+ $Y=1.485 $X2=6.17 $Y2=2
r200 5 35 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=5.13
+ $Y=1.485 $X2=5.265 $Y2=2.02
r201 4 105 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.485 $X2=4.425 $Y2=2.34
r202 3 99 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.77
+ $Y=2.065 $X2=3.905 $Y2=2.3
r203 2 31 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r204 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%Q 1 2 7 10 11 12 13 14 19
r34 13 19 10.8721 $w=2.63e-07 $l=2.5e-07 $layer=LI1_cond $X=5.782 $Y=2.21
+ $X2=5.782 $Y2=1.96
r35 12 14 19.9904 $w=4.15e-07 $l=8.44985e-07 $layer=LI1_cond $X=5.795 $Y=0.51
+ $X2=6.165 $Y2=1.19
r36 11 19 13.0465 $w=2.63e-07 $l=3e-07 $layer=LI1_cond $X=5.782 $Y=1.66
+ $X2=5.782 $Y2=1.96
r37 10 11 8.23835 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.812 $Y=1.495
+ $X2=5.812 $Y2=1.66
r38 7 14 7.7687 $w=4.15e-07 $l=3.43939e-07 $layer=LI1_cond $X=5.882 $Y=1.325
+ $X2=6.165 $Y2=1.19
r39 7 10 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=5.882 $Y=1.325
+ $X2=5.882 $Y2=1.495
r40 2 19 300 $w=1.7e-07 $l=5.59911e-07 $layer=licon1_PDIFF $count=2 $X=5.55
+ $Y=1.485 $X2=5.735 $Y2=1.96
r41 1 12 182 $w=1.7e-07 $l=4.2761e-07 $layer=licon1_NDIFF $count=1 $X=5.55
+ $Y=0.235 $X2=5.735 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%Q_N 1 2 8 10 11 14 15 16 17 33
c29 11 0 1.50259e-19 $X=7.627 $Y=1.572
c30 10 0 1.35563e-19 $X=7.627 $Y=0.825
r31 17 33 0.853661 $w=2.68e-07 $l=2e-08 $layer=LI1_cond $X=8.07 $Y=1.19 $X2=8.05
+ $Y2=1.19
r32 15 16 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=7.627 $Y=1.82
+ $X2=7.627 $Y2=2.21
r33 13 33 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.755 $Y=1.19
+ $X2=8.05 $Y2=1.19
r34 11 15 11.2081 $w=2.53e-07 $l=2.48e-07 $layer=LI1_cond $X=7.627 $Y=1.572
+ $X2=7.627 $Y2=1.82
r35 11 13 18.526 $w=2.55e-07 $l=3.82e-07 $layer=LI1_cond $X=7.627 $Y=1.572
+ $X2=7.627 $Y2=1.19
r36 9 14 8.49644 $w=2.53e-07 $l=1.88e-07 $layer=LI1_cond $X=7.627 $Y=0.698
+ $X2=7.627 $Y2=0.51
r37 9 10 6.13261 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=7.627 $Y=0.698
+ $X2=7.627 $Y2=0.825
r38 8 13 7.49469 $w=2.21e-07 $l=1.46048e-07 $layer=LI1_cond $X=7.65 $Y=1.055
+ $X2=7.627 $Y2=1.19
r39 8 10 12.1472 $w=2.08e-07 $l=2.3e-07 $layer=LI1_cond $X=7.65 $Y=1.055
+ $X2=7.65 $Y2=0.825
r40 2 15 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=7.45
+ $Y=1.485 $X2=7.585 $Y2=1.82
r41 1 14 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=7.45
+ $Y=0.235 $X2=7.585 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 50 52 57 62 70 75 80 85 91 94 97 100 103 106 110
c136 110 0 2.71124e-20 $X=8.05 $Y=0
c137 2 0 7.13094e-20 $X=1.905 $Y=0.235
r138 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r139 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r140 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r141 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r142 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r143 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r144 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r145 89 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r146 89 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r147 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r148 86 106 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.33 $Y=0
+ $X2=7.177 $Y2=0
r149 86 88 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.33 $Y=0 $X2=7.59
+ $Y2=0
r150 85 109 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.925 $Y=0
+ $X2=8.102 $Y2=0
r151 85 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.925 $Y=0
+ $X2=7.59 $Y2=0
r152 84 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r153 84 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r154 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r155 81 103 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.355 $Y=0
+ $X2=6.22 $Y2=0
r156 81 83 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.355 $Y=0
+ $X2=6.67 $Y2=0
r157 80 106 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.025 $Y=0
+ $X2=7.177 $Y2=0
r158 80 83 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.025 $Y=0
+ $X2=6.67 $Y2=0
r159 79 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r160 79 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r161 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r162 76 100 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.48 $Y=0 $X2=5.29
+ $Y2=0
r163 76 78 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.48 $Y=0 $X2=5.75
+ $Y2=0
r164 75 103 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=6.22 $Y2=0
r165 75 78 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=5.75 $Y2=0
r166 74 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r167 74 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r168 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r169 71 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.905
+ $Y2=0
r170 71 73 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.83
+ $Y2=0
r171 70 100 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=5.29
+ $Y2=0
r172 70 73 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.1 $Y=0 $X2=4.83
+ $Y2=0
r173 69 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r174 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r175 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r176 66 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r177 65 68 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r178 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r179 63 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r180 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r181 62 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.905
+ $Y2=0
r182 62 68 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.45
+ $Y2=0
r183 61 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r184 61 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r185 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r186 58 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r187 58 60 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r188 57 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r189 57 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r190 52 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r191 52 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r192 50 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r193 50 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r194 46 109 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=8.06 $Y=0.085
+ $X2=8.102 $Y2=0
r195 46 48 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.06 $Y=0.085
+ $X2=8.06 $Y2=0.38
r196 42 106 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.177 $Y=0.085
+ $X2=7.177 $Y2=0
r197 42 44 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=7.177 $Y=0.085
+ $X2=7.177 $Y2=0.38
r198 38 103 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=0.085
+ $X2=6.22 $Y2=0
r199 38 40 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.22 $Y=0.085
+ $X2=6.22 $Y2=0.38
r200 34 100 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0
r201 34 36 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0.36
r202 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0
r203 30 32 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0.445
r204 26 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r205 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r206 22 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r207 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r208 7 48 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.875
+ $Y=0.235 $X2=8.01 $Y2=0.38
r209 6 44 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=6.975
+ $Y=0.235 $X2=7.165 $Y2=0.38
r210 5 40 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.025
+ $Y=0.235 $X2=6.17 $Y2=0.38
r211 4 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.13
+ $Y=0.235 $X2=5.265 $Y2=0.36
r212 3 32 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.235 $X2=3.905 $Y2=0.445
r213 2 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r214 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


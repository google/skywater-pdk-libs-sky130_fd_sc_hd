* File: sky130_fd_sc_hd__o32ai_2.spice.SKY130_FD_SC_HD__O32AI_2.pxi
* Created: Thu Aug 27 14:41:24 2020
* 
x_PM_SKY130_FD_SC_HD__O32AI_2%B2 N_B2_c_87_n N_B2_M1009_g N_B2_M1003_g
+ N_B2_c_88_n N_B2_M1018_g N_B2_M1015_g B2 B2 N_B2_c_90_n
+ PM_SKY130_FD_SC_HD__O32AI_2%B2
x_PM_SKY130_FD_SC_HD__O32AI_2%B1 N_B1_c_125_n N_B1_M1013_g N_B1_M1000_g
+ N_B1_c_126_n N_B1_M1014_g N_B1_M1017_g B1 B1 N_B1_c_128_n
+ PM_SKY130_FD_SC_HD__O32AI_2%B1
x_PM_SKY130_FD_SC_HD__O32AI_2%A3 N_A3_M1010_g N_A3_c_174_n N_A3_M1001_g
+ N_A3_c_175_n N_A3_M1016_g N_A3_M1004_g A3 N_A3_c_176_n N_A3_c_177_n
+ N_A3_c_178_n PM_SKY130_FD_SC_HD__O32AI_2%A3
x_PM_SKY130_FD_SC_HD__O32AI_2%A2 N_A2_c_227_n N_A2_M1005_g N_A2_M1008_g
+ N_A2_c_228_n N_A2_M1006_g N_A2_M1011_g A2 A2 N_A2_c_230_n
+ PM_SKY130_FD_SC_HD__O32AI_2%A2
x_PM_SKY130_FD_SC_HD__O32AI_2%A1 N_A1_c_273_n N_A1_M1002_g N_A1_M1007_g
+ N_A1_c_274_n N_A1_M1019_g N_A1_M1012_g A1 A1 A1 N_A1_c_276_n
+ PM_SKY130_FD_SC_HD__O32AI_2%A1
x_PM_SKY130_FD_SC_HD__O32AI_2%A_27_297# N_A_27_297#_M1003_d N_A_27_297#_M1015_d
+ N_A_27_297#_M1017_s N_A_27_297#_c_312_n N_A_27_297#_c_313_n
+ N_A_27_297#_c_316_n N_A_27_297#_c_319_n N_A_27_297#_c_320_n
+ N_A_27_297#_c_322_n N_A_27_297#_c_314_n PM_SKY130_FD_SC_HD__O32AI_2%A_27_297#
x_PM_SKY130_FD_SC_HD__O32AI_2%Y N_Y_M1009_s N_Y_M1013_s N_Y_M1003_s N_Y_M1001_s
+ N_Y_c_352_n N_Y_c_361_n N_Y_c_354_n N_Y_c_362_n N_Y_c_384_n Y Y Y
+ PM_SKY130_FD_SC_HD__O32AI_2%Y
x_PM_SKY130_FD_SC_HD__O32AI_2%VPWR N_VPWR_M1000_d N_VPWR_M1007_d N_VPWR_M1012_d
+ N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n
+ N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n VPWR N_VPWR_c_432_n
+ N_VPWR_c_423_n PM_SKY130_FD_SC_HD__O32AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O32AI_2%A_475_297# N_A_475_297#_M1001_d
+ N_A_475_297#_M1004_d N_A_475_297#_M1011_d N_A_475_297#_c_498_n
+ N_A_475_297#_c_499_n N_A_475_297#_c_502_n N_A_475_297#_c_504_n
+ N_A_475_297#_c_506_n N_A_475_297#_c_500_n N_A_475_297#_c_501_n
+ N_A_475_297#_c_529_n PM_SKY130_FD_SC_HD__O32AI_2%A_475_297#
x_PM_SKY130_FD_SC_HD__O32AI_2%A_729_297# N_A_729_297#_M1008_s
+ N_A_729_297#_M1007_s N_A_729_297#_c_538_n N_A_729_297#_c_548_n
+ N_A_729_297#_c_552_n N_A_729_297#_c_541_n
+ PM_SKY130_FD_SC_HD__O32AI_2%A_729_297#
x_PM_SKY130_FD_SC_HD__O32AI_2%A_27_47# N_A_27_47#_M1009_d N_A_27_47#_M1018_d
+ N_A_27_47#_M1014_d N_A_27_47#_M1016_d N_A_27_47#_M1006_d N_A_27_47#_M1019_s
+ N_A_27_47#_c_567_n N_A_27_47#_c_568_n N_A_27_47#_c_578_n N_A_27_47#_c_584_n
+ N_A_27_47#_c_569_n N_A_27_47#_c_570_n N_A_27_47#_c_591_n N_A_27_47#_c_571_n
+ N_A_27_47#_c_572_n N_A_27_47#_c_573_n N_A_27_47#_c_574_n N_A_27_47#_c_575_n
+ PM_SKY130_FD_SC_HD__O32AI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__O32AI_2%VGND N_VGND_M1010_s N_VGND_M1005_s N_VGND_M1002_d
+ N_VGND_c_659_n N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n
+ N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n VGND
+ N_VGND_c_668_n N_VGND_c_669_n PM_SKY130_FD_SC_HD__O32AI_2%VGND
cc_1 VNB N_B2_c_87_n 0.0213689f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B2_c_88_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB B2 0.0135148f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_4 VNB N_B2_c_90_n 0.0377314f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_B1_c_125_n 0.0159967f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B1_c_126_n 0.0159701f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_7 VNB B1 0.00363163f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_B1_c_128_n 0.0315417f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_9 VNB N_A3_M1010_g 0.0285182f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A3_c_174_n 0.0084854f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_11 VNB N_A3_c_175_n 0.0217006f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_12 VNB N_A3_c_176_n 0.0293787f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_13 VNB N_A3_c_177_n 0.00295465f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_14 VNB N_A3_c_178_n 0.0381424f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_15 VNB N_A2_c_227_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_A2_c_228_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_17 VNB A2 0.00989386f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_18 VNB N_A2_c_230_n 0.0391114f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_19 VNB N_A1_c_273_n 0.0212108f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_A1_c_274_n 0.0213225f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_21 VNB A1 0.0207295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_276_n 0.0475875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_352_n 0.00824807f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_24 VNB Y 0.0055537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_423_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_567_n 0.0100703f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_27 VNB N_A_27_47#_c_568_n 0.0183982f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_28 VNB N_A_27_47#_c_569_n 0.003827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_570_n 0.00191967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_571_n 0.0144518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_572_n 0.0180521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_573_n 0.00484878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_574_n 0.00246923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_575_n 0.00822315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_659_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_36 VNB N_VGND_c_660_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_37 VNB N_VGND_c_661_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_662_n 0.0623145f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.16
cc_39 VNB N_VGND_c_663_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_40 VNB N_VGND_c_664_n 0.0170602f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_41 VNB N_VGND_c_665_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_666_n 0.0259816f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=1.2
cc_43 VNB N_VGND_c_667_n 0.00436611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_668_n 0.0209894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_669_n 0.301374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_B2_M1003_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_47 VPB N_B2_M1015_g 0.0188371f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_48 VPB B2 0.00503392f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_49 VPB N_B2_c_90_n 0.00429053f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_50 VPB N_B1_M1000_g 0.0188311f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_51 VPB N_B1_M1017_g 0.0218926f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_52 VPB B1 0.00215893f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_53 VPB N_B1_c_128_n 0.00409488f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_54 VPB N_A3_M1001_g 0.0229395f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_55 VPB N_A3_M1004_g 0.0188371f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_56 VPB N_A3_c_177_n 0.00247431f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_57 VPB N_A3_c_178_n 0.00424573f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_58 VPB N_A2_M1008_g 0.0188371f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_59 VPB N_A2_M1011_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_60 VPB A2 0.00489054f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_61 VPB N_A2_c_230_n 0.00742087f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_62 VPB N_A1_M1007_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_63 VPB N_A1_M1012_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_64 VPB A1 0.0108238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A1_c_276_n 0.00689228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_297#_c_312_n 0.00753428f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_67 VPB N_A_27_297#_c_313_n 0.0305647f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_A_27_297#_c_314_n 0.00663738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_Y_c_354_n 0.00929876f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_70 VPB Y 0.0044334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB Y 0.00357952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_424_n 0.00462218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_73 VPB N_VPWR_c_425_n 0.004361f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_74 VPB N_VPWR_c_426_n 0.0148582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_427_n 0.00444474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_428_n 0.0357516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_429_n 0.003239f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_78 VPB N_VPWR_c_430_n 0.0736785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_431_n 0.00391557f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.2
cc_80 VPB N_VPWR_c_432_n 0.0181025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_423_n 0.0707433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_475_297#_c_498_n 0.00213564f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_83 VPB N_A_475_297#_c_499_n 0.00428417f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_84 VPB N_A_475_297#_c_500_n 0.00211678f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_85 VPB N_A_475_297#_c_501_n 0.00431617f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_86 VPB N_A_729_297#_c_538_n 0.0133368f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_87 N_B2_c_88_n N_B1_c_125_n 0.024858f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_88 N_B2_M1015_g N_B1_M1000_g 0.024858f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_89 B2 B1 0.0221327f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B2_c_90_n B1 0.00234073f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B2_c_90_n N_B1_c_128_n 0.024858f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_92 B2 N_A_27_297#_c_313_n 0.021306f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B2_M1003_g N_A_27_297#_c_316_n 0.011323f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_94 N_B2_M1015_g N_A_27_297#_c_316_n 0.00934626f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_95 N_B2_c_87_n N_Y_c_352_n 0.00376463f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B2_c_88_n N_Y_c_352_n 0.0121388f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_97 B2 N_Y_c_352_n 0.0248006f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B2_c_90_n N_Y_c_352_n 0.00223984f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B2_M1015_g N_Y_c_361_n 0.0102605f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B2_M1003_g N_Y_c_362_n 0.0074304f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B2_M1015_g N_Y_c_362_n 0.00713556f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_102 B2 N_Y_c_362_n 0.0211943f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B2_c_90_n N_Y_c_362_n 0.00208544f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B2_M1003_g N_VPWR_c_428_n 0.00357877f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B2_M1015_g N_VPWR_c_428_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B2_M1003_g N_VPWR_c_423_n 0.00617937f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B2_M1015_g N_VPWR_c_423_n 0.00525237f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B2_c_87_n N_A_27_47#_c_568_n 4.62114e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_109 B2 N_A_27_47#_c_568_n 0.0218655f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_110 N_B2_c_87_n N_A_27_47#_c_578_n 0.0108017f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B2_c_88_n N_A_27_47#_c_578_n 0.00918728f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_112 B2 N_A_27_47#_c_578_n 0.00389697f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_113 N_B2_c_87_n N_VGND_c_662_n 0.00357877f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B2_c_88_n N_VGND_c_662_n 0.00357877f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B2_c_87_n N_VGND_c_669_n 0.00617937f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B2_c_88_n N_VGND_c_669_n 0.00525237f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B1_c_126_n N_A3_M1010_g 0.0181595f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_c_128_n N_A3_c_174_n 0.0181595f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B1_M1000_g N_A_27_297#_c_316_n 0.00202914f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B1_M1000_g N_A_27_297#_c_319_n 8.8323e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B1_M1000_g N_A_27_297#_c_320_n 0.00418215f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_M1017_g N_A_27_297#_c_320_n 4.70065e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_M1000_g N_A_27_297#_c_322_n 0.00844123f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_M1017_g N_A_27_297#_c_322_n 0.00839707f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_125 N_B1_M1000_g N_A_27_297#_c_314_n 5.16334e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B1_M1017_g N_A_27_297#_c_314_n 0.0069824f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B1_c_125_n N_Y_c_352_n 0.010631f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_c_126_n N_Y_c_352_n 0.0113463f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_129 B1 N_Y_c_352_n 0.0524345f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_130 N_B1_c_128_n N_Y_c_352_n 0.00223984f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B1_M1000_g N_Y_c_361_n 0.0103223f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_132 N_B1_M1017_g N_Y_c_361_n 0.0137453f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_133 B1 N_Y_c_361_n 0.0437923f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B1_c_128_n N_Y_c_361_n 0.00201785f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B1_M1000_g N_Y_c_362_n 7.7319e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B1_c_126_n Y 0.00475726f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_M1017_g Y 0.00475726f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_138 B1 Y 0.020483f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_139 N_B1_c_128_n Y 0.00475726f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B1_M1000_g N_VPWR_c_424_n 0.00268723f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B1_M1017_g N_VPWR_c_424_n 0.00268723f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B1_M1000_g N_VPWR_c_428_n 0.00420723f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B1_M1017_g N_VPWR_c_430_n 0.00422645f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B1_M1000_g N_VPWR_c_423_n 0.00573284f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B1_M1017_g N_VPWR_c_423_n 0.00702302f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_146 N_B1_c_125_n N_A_27_47#_c_578_n 0.00918728f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B1_c_126_n N_A_27_47#_c_578_n 0.00918728f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_148 N_B1_c_125_n N_VGND_c_662_n 0.00357877f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_149 N_B1_c_126_n N_VGND_c_662_n 0.00357877f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B1_c_125_n N_VGND_c_669_n 0.00525237f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B1_c_126_n N_VGND_c_669_n 0.00525237f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A3_c_175_n N_A2_c_227_n 0.0124239f $X=3.09 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_153 N_A3_M1004_g N_A2_M1008_g 0.0151563f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A3_c_177_n A2 0.0142213f $X=2.9 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A3_c_178_n A2 0.00228619f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A3_c_177_n N_A2_c_230_n 2.2138e-19 $X=2.9 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A3_c_178_n N_A2_c_230_n 0.0229806f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A3_M1010_g N_Y_c_352_n 0.00116103f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A3_c_174_n N_Y_c_354_n 0.00610428f $X=2.225 $Y=1.19 $X2=0 $Y2=0
cc_160 N_A3_M1001_g N_Y_c_354_n 0.010778f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A3_c_176_n N_Y_c_354_n 0.00140486f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A3_c_177_n N_Y_c_354_n 0.0253373f $X=2.9 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A3_M1001_g N_Y_c_384_n 0.0115378f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A3_M1004_g N_Y_c_384_n 0.00735116f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A3_c_177_n N_Y_c_384_n 0.0185297f $X=2.9 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A3_c_178_n N_Y_c_384_n 0.00208443f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A3_M1010_g Y 0.00743278f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A3_c_174_n Y 0.00705208f $X=2.225 $Y=1.19 $X2=0 $Y2=0
cc_169 N_A3_c_177_n Y 0.0152726f $X=2.9 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A3_c_178_n Y 0.00471841f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A3_M1001_g N_VPWR_c_430_n 0.00362032f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A3_M1004_g N_VPWR_c_430_n 0.00362032f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A3_M1001_g N_VPWR_c_423_n 0.00655665f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A3_M1004_g N_VPWR_c_423_n 0.00525778f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A3_M1001_g N_A_475_297#_c_502_n 0.00986542f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A3_M1004_g N_A_475_297#_c_502_n 0.0120057f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A3_M1010_g N_A_27_47#_c_578_n 0.0137645f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A3_c_175_n N_A_27_47#_c_584_n 0.00374992f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A3_c_175_n N_A_27_47#_c_569_n 0.0126951f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A3_c_176_n N_A_27_47#_c_569_n 0.00160685f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A3_c_177_n N_A_27_47#_c_569_n 0.0497557f $X=2.9 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A3_c_178_n N_A_27_47#_c_569_n 0.0100576f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A3_M1010_g N_A_27_47#_c_570_n 0.00391811f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A3_c_176_n N_A_27_47#_c_570_n 0.0041434f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A3_c_175_n N_A_27_47#_c_591_n 0.010934f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A3_c_175_n N_A_27_47#_c_573_n 0.00223339f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A3_c_178_n N_A_27_47#_c_573_n 0.00313057f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A3_M1010_g N_VGND_c_659_n 0.00427695f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A3_c_175_n N_VGND_c_659_n 0.011703f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A3_M1010_g N_VGND_c_662_n 0.00357877f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A3_c_175_n N_VGND_c_664_n 0.00422241f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A3_M1010_g N_VGND_c_669_n 0.00662944f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A3_c_175_n N_VGND_c_669_n 0.00718253f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_194 A2 A1 0.0167879f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_195 N_A2_c_230_n A1 8.78255e-19 $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_196 A2 N_A1_c_276_n 0.00167412f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_197 N_A2_M1011_g N_VPWR_c_425_n 0.00227006f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A2_M1008_g N_VPWR_c_430_n 0.00362032f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A2_M1011_g N_VPWR_c_430_n 0.00362032f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A2_M1008_g N_VPWR_c_423_n 0.00525778f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A2_M1011_g N_VPWR_c_423_n 0.00655665f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_202 A2 N_A_475_297#_c_504_n 0.00598284f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A2_c_230_n N_A_475_297#_c_504_n 2.26876e-19 $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A2_M1008_g N_A_475_297#_c_506_n 0.0120057f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A2_M1011_g N_A_475_297#_c_506_n 0.00986542f $X=3.99 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A2_M1011_g N_A_729_297#_c_538_n 0.010778f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_207 A2 N_A_729_297#_c_538_n 0.0380967f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_208 N_A2_M1008_g N_A_729_297#_c_541_n 0.00695277f $X=3.57 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A2_M1011_g N_A_729_297#_c_541_n 0.0115378f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_210 A2 N_A_729_297#_c_541_n 0.0211713f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_211 N_A2_c_230_n N_A_729_297#_c_541_n 0.00232108f $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A2_c_227_n N_A_27_47#_c_591_n 0.00641078f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A2_c_228_n N_A_27_47#_c_591_n 5.362e-19 $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A2_c_227_n N_A_27_47#_c_573_n 0.00115517f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_215 A2 N_A_27_47#_c_573_n 0.0079569f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A2_c_227_n N_A_27_47#_c_574_n 0.00890471f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A2_c_228_n N_A_27_47#_c_574_n 0.0151866f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_218 A2 N_A_27_47#_c_574_n 0.0792307f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_219 N_A2_c_230_n N_A_27_47#_c_574_n 0.00422891f $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A2_c_227_n N_VGND_c_660_n 0.00268723f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A2_c_228_n N_VGND_c_660_n 0.00268723f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_227_n N_VGND_c_664_n 0.00422241f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A2_c_228_n N_VGND_c_666_n 0.00436487f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A2_c_227_n N_VGND_c_669_n 0.00572376f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A2_c_228_n N_VGND_c_669_n 0.00728351f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A1_M1007_g N_VPWR_c_425_n 0.00318713f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A1_M1012_g N_VPWR_c_427_n 0.00319616f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_228 A1 N_VPWR_c_427_n 0.0182541f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_229 N_A1_M1007_g N_VPWR_c_432_n 0.00541562f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A1_M1012_g N_VPWR_c_432_n 0.00541562f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_M1007_g N_VPWR_c_423_n 0.0108278f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A1_M1012_g N_VPWR_c_423_n 0.0105657f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_M1007_g N_A_729_297#_c_538_n 0.0128219f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_234 A1 N_A_729_297#_c_538_n 0.0154908f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_235 N_A1_c_276_n N_A_729_297#_c_538_n 0.00198379f $X=5.37 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A1_M1007_g N_A_729_297#_c_548_n 8.84614e-19 $X=4.95 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A1_M1012_g N_A_729_297#_c_548_n 0.00229676f $X=5.37 $Y=1.985 $X2=0
+ $Y2=0
cc_238 A1 N_A_729_297#_c_548_n 0.0213676f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A1_c_276_n N_A_729_297#_c_548_n 0.00241214f $X=5.37 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A1_M1007_g N_A_729_297#_c_552_n 0.0145112f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A1_M1012_g N_A_729_297#_c_552_n 0.00897627f $X=5.37 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A1_c_273_n N_A_27_47#_c_571_n 0.0147143f $X=4.87 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A1_c_274_n N_A_27_47#_c_571_n 0.0144325f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_244 A1 N_A_27_47#_c_571_n 0.0775525f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_245 N_A1_c_276_n N_A_27_47#_c_571_n 0.00490423f $X=5.37 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A1_c_274_n N_A_27_47#_c_572_n 0.0136394f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A1_c_273_n N_A_27_47#_c_575_n 0.0142899f $X=4.87 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A1_c_273_n N_VGND_c_661_n 0.00996796f $X=4.87 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A1_c_274_n N_VGND_c_661_n 0.00873867f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A1_c_273_n N_VGND_c_666_n 0.00319306f $X=4.87 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_274_n N_VGND_c_668_n 0.00377504f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_273_n N_VGND_c_669_n 0.00522424f $X=4.87 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_274_n N_VGND_c_669_n 0.0055953f $X=5.29 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_27_297#_c_316_n N_Y_M1003_s 0.00324321f $X=1.015 $Y=2.38 $X2=0 $Y2=0
cc_255 N_A_27_297#_M1015_d N_Y_c_361_n 0.00332066f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_256 N_A_27_297#_M1017_s N_Y_c_361_n 3.49698e-19 $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_257 N_A_27_297#_c_316_n N_Y_c_361_n 0.00271653f $X=1.015 $Y=2.38 $X2=0 $Y2=0
cc_258 N_A_27_297#_c_319_n N_Y_c_361_n 0.0148421f $X=1.14 $Y=2.005 $X2=0 $Y2=0
cc_259 N_A_27_297#_c_322_n N_Y_c_361_n 0.0275303f $X=1.775 $Y=1.92 $X2=0 $Y2=0
cc_260 N_A_27_297#_c_314_n N_Y_c_361_n 0.00323992f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_261 N_A_27_297#_c_316_n N_Y_c_362_n 0.0137059f $X=1.015 $Y=2.38 $X2=0 $Y2=0
cc_262 N_A_27_297#_M1017_s Y 0.00284298f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_263 N_A_27_297#_c_314_n Y 0.0206123f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_264 N_A_27_297#_c_322_n N_VPWR_M1000_d 0.00317424f $X=1.775 $Y=1.92 $X2=-0.19
+ $Y2=1.305
cc_265 N_A_27_297#_c_322_n N_VPWR_c_424_n 0.012179f $X=1.775 $Y=1.92 $X2=0 $Y2=0
cc_266 N_A_27_297#_c_312_n N_VPWR_c_428_n 0.0177497f $X=0.217 $Y=2.295 $X2=0
+ $Y2=0
cc_267 N_A_27_297#_c_316_n N_VPWR_c_428_n 0.0510205f $X=1.015 $Y=2.38 $X2=0
+ $Y2=0
cc_268 N_A_27_297#_c_322_n N_VPWR_c_428_n 0.0020257f $X=1.775 $Y=1.92 $X2=0
+ $Y2=0
cc_269 N_A_27_297#_c_322_n N_VPWR_c_430_n 0.0020257f $X=1.775 $Y=1.92 $X2=0
+ $Y2=0
cc_270 N_A_27_297#_c_314_n N_VPWR_c_430_n 0.0196584f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_271 N_A_27_297#_M1003_d N_VPWR_c_423_n 0.00209324f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_272 N_A_27_297#_M1015_d N_VPWR_c_423_n 0.00215206f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_273 N_A_27_297#_M1017_s N_VPWR_c_423_n 0.00209642f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_274 N_A_27_297#_c_312_n N_VPWR_c_423_n 0.00981527f $X=0.217 $Y=2.295 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_c_316_n N_VPWR_c_423_n 0.0328416f $X=1.015 $Y=2.38 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_c_322_n N_VPWR_c_423_n 0.00841425f $X=1.775 $Y=1.92 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_c_314_n N_VPWR_c_423_n 0.0123353f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_278 N_A_27_297#_c_314_n N_A_475_297#_c_498_n 0.0135924f $X=1.94 $Y=2 $X2=0
+ $Y2=0
cc_279 N_A_27_297#_c_314_n N_A_475_297#_c_499_n 0.0283667f $X=1.94 $Y=2 $X2=0
+ $Y2=0
cc_280 N_Y_c_361_n N_VPWR_M1000_d 0.00311888f $X=1.875 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_281 N_Y_M1003_s N_VPWR_c_423_n 0.00216833f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_282 N_Y_M1001_s N_VPWR_c_423_n 0.00217706f $X=2.805 $Y=1.485 $X2=0 $Y2=0
cc_283 N_Y_c_354_n N_A_475_297#_M1001_d 0.00549184f $X=2.775 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_284 N_Y_c_354_n N_A_475_297#_c_499_n 0.0201185f $X=2.775 $Y=1.58 $X2=0 $Y2=0
cc_285 N_Y_c_384_n N_A_475_297#_c_499_n 0.0174368f $X=2.94 $Y=1.66 $X2=0 $Y2=0
cc_286 N_Y_M1001_s N_A_475_297#_c_502_n 0.0031999f $X=2.805 $Y=1.485 $X2=0 $Y2=0
cc_287 N_Y_c_354_n N_A_475_297#_c_502_n 0.00327285f $X=2.775 $Y=1.58 $X2=0 $Y2=0
cc_288 N_Y_c_384_n N_A_475_297#_c_502_n 0.0160339f $X=2.94 $Y=1.66 $X2=0 $Y2=0
cc_289 N_Y_c_352_n N_A_27_47#_M1018_d 0.00162409f $X=1.875 $Y=0.78 $X2=0 $Y2=0
cc_290 N_Y_c_352_n N_A_27_47#_M1014_d 0.00206002f $X=1.875 $Y=0.78 $X2=0 $Y2=0
cc_291 N_Y_c_352_n N_A_27_47#_c_568_n 0.01117f $X=1.875 $Y=0.78 $X2=0 $Y2=0
cc_292 N_Y_M1009_s N_A_27_47#_c_578_n 0.00305179f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_293 N_Y_M1013_s N_A_27_47#_c_578_n 0.00305179f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_294 N_Y_c_352_n N_A_27_47#_c_578_n 0.0786734f $X=1.875 $Y=0.78 $X2=0 $Y2=0
cc_295 Y N_A_27_47#_c_578_n 0.00299102f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_296 N_Y_c_384_n N_A_27_47#_c_569_n 9.21061e-19 $X=2.94 $Y=1.66 $X2=0 $Y2=0
cc_297 N_Y_c_352_n N_A_27_47#_c_570_n 0.00164322f $X=1.875 $Y=0.78 $X2=0 $Y2=0
cc_298 N_Y_c_354_n N_A_27_47#_c_570_n 0.00590606f $X=2.775 $Y=1.58 $X2=0 $Y2=0
cc_299 N_Y_M1009_s N_VGND_c_669_n 0.00216833f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_300 N_Y_M1013_s N_VGND_c_669_n 0.00216833f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_301 N_VPWR_c_423_n N_A_475_297#_M1001_d 0.00226598f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_302 N_VPWR_c_423_n N_A_475_297#_M1004_d 0.00216056f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_423_n N_A_475_297#_M1011_d 0.00226598f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_430_n N_A_475_297#_c_498_n 0.0155085f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_423_n N_A_475_297#_c_498_n 0.00950669f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_430_n N_A_475_297#_c_502_n 0.0329469f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_423_n N_A_475_297#_c_502_n 0.0239272f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_430_n N_A_475_297#_c_506_n 0.0329469f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_423_n N_A_475_297#_c_506_n 0.0239272f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_425_n N_A_475_297#_c_500_n 0.0126677f $X=4.74 $Y=2 $X2=0 $Y2=0
cc_311 N_VPWR_c_430_n N_A_475_297#_c_500_n 0.0155085f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_423_n N_A_475_297#_c_500_n 0.00950669f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_425_n N_A_475_297#_c_501_n 0.0256956f $X=4.74 $Y=2 $X2=0 $Y2=0
cc_314 N_VPWR_c_430_n N_A_475_297#_c_529_n 0.0101645f $X=4.62 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_423_n N_A_475_297#_c_529_n 0.00648411f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_423_n N_A_729_297#_M1008_s 0.00217706f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_317 N_VPWR_c_423_n N_A_729_297#_M1007_s 0.00215347f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_318 N_VPWR_M1007_d N_A_729_297#_c_538_n 0.00636722f $X=4.615 $Y=1.485 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_425_n N_A_729_297#_c_538_n 0.0160276f $X=4.74 $Y=2 $X2=0 $Y2=0
cc_320 N_VPWR_c_432_n N_A_729_297#_c_552_n 0.0183232f $X=5.495 $Y=2.72 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_423_n N_A_729_297#_c_552_n 0.0121916f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_322 N_A_475_297#_c_506_n N_A_729_297#_M1008_s 0.0031999f $X=4.135 $Y=2.35
+ $X2=-0.19 $Y2=1.305
cc_323 N_A_475_297#_M1011_d N_A_729_297#_c_538_n 0.00578441f $X=4.065 $Y=1.485
+ $X2=0 $Y2=0
cc_324 N_A_475_297#_c_506_n N_A_729_297#_c_538_n 0.00327285f $X=4.135 $Y=2.35
+ $X2=0 $Y2=0
cc_325 N_A_475_297#_c_501_n N_A_729_297#_c_538_n 0.0201185f $X=4.22 $Y=2 $X2=0
+ $Y2=0
cc_326 N_A_475_297#_c_506_n N_A_729_297#_c_541_n 0.0160339f $X=4.135 $Y=2.35
+ $X2=0 $Y2=0
cc_327 N_A_475_297#_c_501_n N_A_729_297#_c_541_n 0.0174368f $X=4.22 $Y=2 $X2=0
+ $Y2=0
cc_328 N_A_475_297#_c_504_n N_A_27_47#_c_573_n 0.00338865f $X=3.36 $Y=1.66 $X2=0
+ $Y2=0
cc_329 N_A_729_297#_c_538_n N_A_27_47#_c_575_n 0.0092242f $X=4.995 $Y=1.58 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_578_n N_VGND_M1010_s 0.00377834f $X=2.235 $Y=0.37 $X2=-0.19
+ $Y2=-0.24
cc_331 N_A_27_47#_c_584_n N_VGND_M1010_s 0.00382853f $X=2.32 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_332 N_A_27_47#_c_569_n N_VGND_M1010_s 0.0116591f $X=3.135 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_333 N_A_27_47#_c_570_n N_VGND_M1010_s 0.00115737f $X=2.405 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_334 N_A_27_47#_c_574_n N_VGND_M1005_s 0.00162148f $X=4.055 $Y=0.58 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_571_n N_VGND_M1002_d 0.00162148f $X=5.425 $Y=0.81 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_578_n N_VGND_c_659_n 0.0164488f $X=2.235 $Y=0.37 $X2=0 $Y2=0
cc_337 N_A_27_47#_c_584_n N_VGND_c_659_n 0.00382373f $X=2.32 $Y=0.715 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_569_n N_VGND_c_659_n 0.0257931f $X=3.135 $Y=0.81 $X2=0 $Y2=0
cc_339 N_A_27_47#_c_591_n N_VGND_c_659_n 0.0210898f $X=3.3 $Y=0.38 $X2=0 $Y2=0
cc_340 N_A_27_47#_c_574_n N_VGND_c_660_n 0.0122675f $X=4.055 $Y=0.58 $X2=0 $Y2=0
cc_341 N_A_27_47#_c_571_n N_VGND_c_661_n 0.016455f $X=5.425 $Y=0.81 $X2=0 $Y2=0
cc_342 N_A_27_47#_c_572_n N_VGND_c_661_n 0.0206616f $X=5.59 $Y=0.38 $X2=0 $Y2=0
cc_343 N_A_27_47#_c_575_n N_VGND_c_661_n 0.0228041f $X=4.725 $Y=0.58 $X2=0 $Y2=0
cc_344 N_A_27_47#_c_567_n N_VGND_c_662_n 0.0176918f $X=0.217 $Y=0.485 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_578_n N_VGND_c_662_n 0.115793f $X=2.235 $Y=0.37 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_569_n N_VGND_c_662_n 0.00318662f $X=3.135 $Y=0.81 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_569_n N_VGND_c_664_n 0.00221227f $X=3.135 $Y=0.81 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_591_n N_VGND_c_664_n 0.0188551f $X=3.3 $Y=0.38 $X2=0 $Y2=0
cc_349 N_A_27_47#_c_574_n N_VGND_c_664_n 0.00203746f $X=4.055 $Y=0.58 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_571_n N_VGND_c_666_n 0.00214783f $X=5.425 $Y=0.81 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_574_n N_VGND_c_666_n 0.00285442f $X=4.055 $Y=0.58 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_575_n N_VGND_c_666_n 0.0464092f $X=4.725 $Y=0.58 $X2=0 $Y2=0
cc_353 N_A_27_47#_c_571_n N_VGND_c_668_n 0.00226063f $X=5.425 $Y=0.81 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_572_n N_VGND_c_668_n 0.0230421f $X=5.59 $Y=0.38 $X2=0 $Y2=0
cc_355 N_A_27_47#_M1009_d N_VGND_c_669_n 0.00209324f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_M1018_d N_VGND_c_669_n 0.00215227f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_M1014_d N_VGND_c_669_n 0.00215227f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_M1016_d N_VGND_c_669_n 0.00215201f $X=3.165 $Y=0.235 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_M1006_d N_VGND_c_669_n 0.00699525f $X=4.005 $Y=0.235 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_M1019_s N_VGND_c_669_n 0.00312036f $X=5.365 $Y=0.235 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_567_n N_VGND_c_669_n 0.00980895f $X=0.217 $Y=0.485 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_578_n N_VGND_c_669_n 0.0736174f $X=2.235 $Y=0.37 $X2=0 $Y2=0
cc_363 N_A_27_47#_c_569_n N_VGND_c_669_n 0.0114487f $X=3.135 $Y=0.81 $X2=0 $Y2=0
cc_364 N_A_27_47#_c_591_n N_VGND_c_669_n 0.0122069f $X=3.3 $Y=0.38 $X2=0 $Y2=0
cc_365 N_A_27_47#_c_571_n N_VGND_c_669_n 0.00999938f $X=5.425 $Y=0.81 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_572_n N_VGND_c_669_n 0.0126169f $X=5.59 $Y=0.38 $X2=0 $Y2=0
cc_367 N_A_27_47#_c_574_n N_VGND_c_669_n 0.0104483f $X=4.055 $Y=0.58 $X2=0 $Y2=0
cc_368 N_A_27_47#_c_575_n N_VGND_c_669_n 0.0257581f $X=4.725 $Y=0.58 $X2=0 $Y2=0

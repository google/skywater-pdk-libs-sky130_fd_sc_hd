* File: sky130_fd_sc_hd__o31a_2.spice.SKY130_FD_SC_HD__O31A_2.pxi
* Created: Thu Aug 27 14:39:57 2020
* 
x_PM_SKY130_FD_SC_HD__O31A_2%A_108_21# N_A_108_21#_M1010_d N_A_108_21#_M1005_d
+ N_A_108_21#_c_65_n N_A_108_21#_M1002_g N_A_108_21#_M1000_g N_A_108_21#_c_66_n
+ N_A_108_21#_c_67_n N_A_108_21#_M1003_g N_A_108_21#_M1011_g N_A_108_21#_c_68_n
+ N_A_108_21#_c_76_n N_A_108_21#_c_69_n N_A_108_21#_c_78_n N_A_108_21#_c_79_n
+ N_A_108_21#_c_85_p N_A_108_21#_c_96_p N_A_108_21#_c_86_p N_A_108_21#_c_100_p
+ N_A_108_21#_c_101_p N_A_108_21#_c_80_n N_A_108_21#_c_70_n N_A_108_21#_c_71_n
+ PM_SKY130_FD_SC_HD__O31A_2%A_108_21#
x_PM_SKY130_FD_SC_HD__O31A_2%A1 N_A1_M1009_g N_A1_M1004_g A1 N_A1_c_174_n
+ N_A1_c_175_n PM_SKY130_FD_SC_HD__O31A_2%A1
x_PM_SKY130_FD_SC_HD__O31A_2%A2 N_A2_c_206_n N_A2_M1007_g N_A2_M1001_g A2 A2 A2
+ N_A2_c_208_n PM_SKY130_FD_SC_HD__O31A_2%A2
x_PM_SKY130_FD_SC_HD__O31A_2%A3 N_A3_c_242_n N_A3_M1008_g N_A3_M1005_g A3
+ N_A3_c_244_n PM_SKY130_FD_SC_HD__O31A_2%A3
x_PM_SKY130_FD_SC_HD__O31A_2%B1 N_B1_M1010_g N_B1_M1006_g B1 N_B1_c_278_n
+ N_B1_c_279_n PM_SKY130_FD_SC_HD__O31A_2%B1
x_PM_SKY130_FD_SC_HD__O31A_2%VPWR N_VPWR_M1000_d N_VPWR_M1011_d N_VPWR_M1006_d
+ N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n
+ N_VPWR_c_316_n N_VPWR_c_317_n VPWR N_VPWR_c_318_n N_VPWR_c_310_n
+ PM_SKY130_FD_SC_HD__O31A_2%VPWR
x_PM_SKY130_FD_SC_HD__O31A_2%X N_X_M1002_s N_X_M1000_s X X X X X X X N_X_c_357_n
+ X N_X_c_375_n X PM_SKY130_FD_SC_HD__O31A_2%X
x_PM_SKY130_FD_SC_HD__O31A_2%VGND N_VGND_M1002_d N_VGND_M1003_d N_VGND_M1007_d
+ N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n
+ VGND N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n N_VGND_c_406_n
+ PM_SKY130_FD_SC_HD__O31A_2%VGND
x_PM_SKY130_FD_SC_HD__O31A_2%A_346_47# N_A_346_47#_M1009_d N_A_346_47#_M1008_d
+ N_A_346_47#_c_466_n N_A_346_47#_c_453_n N_A_346_47#_c_454_n
+ N_A_346_47#_c_461_n PM_SKY130_FD_SC_HD__O31A_2%A_346_47#
cc_1 VNB N_A_108_21#_c_65_n 0.021741f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.995
cc_2 VNB N_A_108_21#_c_66_n 0.0158815f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=1.16
cc_3 VNB N_A_108_21#_c_67_n 0.0177204f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=0.995
cc_4 VNB N_A_108_21#_c_68_n 0.0162344f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.16
cc_5 VNB N_A_108_21#_c_69_n 0.0136458f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_6 VNB N_A_108_21#_c_70_n 0.0231573f $X=-0.19 $Y=-0.24 $X2=3.51 $Y2=1.495
cc_7 VNB N_A_108_21#_c_71_n 0.0272789f $X=-0.19 $Y=-0.24 $X2=3.275 $Y2=0.36
cc_8 VNB A1 0.00751177f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.56
cc_9 VNB N_A1_c_174_n 0.0190063f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.985
cc_10 VNB N_A1_c_175_n 0.017251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_206_n 0.0167675f $X=-0.19 $Y=-0.24 $X2=3.11 $Y2=0.235
cc_12 VNB A2 8.31138e-19 $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.56
cc_13 VNB N_A2_c_208_n 0.0222913f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_14 VNB N_A3_c_242_n 0.0171433f $X=-0.19 $Y=-0.24 $X2=3.11 $Y2=0.235
cc_15 VNB A3 0.00290055f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.56
cc_16 VNB N_A3_c_244_n 0.0203366f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.985
cc_17 VNB B1 0.00577659f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.56
cc_18 VNB N_B1_c_278_n 0.0264604f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.985
cc_19 VNB N_B1_c_279_n 0.0203196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_310_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_357_n 0.027911f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.16
cc_22 VNB X 0.00114446f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=1.53
cc_23 VNB N_VGND_c_398_n 0.0105866f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.325
cc_24 VNB N_VGND_c_399_n 0.0341703f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.985
cc_25 VNB N_VGND_c_400_n 5.61383e-19 $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=0.995
cc_26 VNB N_VGND_c_401_n 0.0196699f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.325
cc_27 VNB N_VGND_c_402_n 0.00617014f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.985
cc_28 VNB N_VGND_c_403_n 0.0117788f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=1.16
cc_29 VNB N_VGND_c_404_n 0.0299592f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=2.38
cc_30 VNB N_VGND_c_405_n 0.200107f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=2.38
cc_31 VNB N_VGND_c_406_n 0.00598854f $X=-0.19 $Y=-0.24 $X2=2.955 $Y2=1.58
cc_32 VPB N_A_108_21#_M1000_g 0.0256894f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_33 VPB N_A_108_21#_c_66_n 0.00576892f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.16
cc_34 VPB N_A_108_21#_M1011_g 0.0190672f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.985
cc_35 VPB N_A_108_21#_c_68_n 0.00142224f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.16
cc_36 VPB N_A_108_21#_c_76_n 0.00214903f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_37 VPB N_A_108_21#_c_69_n 0.002223f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_38 VPB N_A_108_21#_c_78_n 0.00599705f $X=-0.19 $Y=1.305 $X2=1.65 $Y2=1.53
cc_39 VPB N_A_108_21#_c_79_n 2.62111e-19 $X=-0.19 $Y=1.305 $X2=1.2 $Y2=1.53
cc_40 VPB N_A_108_21#_c_80_n 0.00785406f $X=-0.19 $Y=1.305 $X2=3.425 $Y2=1.58
cc_41 VPB N_A_108_21#_c_70_n 0.00934765f $X=-0.19 $Y=1.305 $X2=3.51 $Y2=1.495
cc_42 VPB N_A1_M1004_g 0.019844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A1_c_174_n 0.00406143f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_44 VPB N_A2_M1001_g 0.0179385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB A2 0.00164103f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=0.56
cc_46 VPB A2 0.00256075f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=0.56
cc_47 VPB N_A2_c_208_n 0.00525592f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_48 VPB N_A3_M1005_g 0.0194949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB A3 0.00315937f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=0.56
cc_50 VPB N_A3_c_244_n 0.00566534f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_51 VPB N_B1_M1006_g 0.0240229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB B1 0.00118297f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=0.56
cc_53 VPB N_B1_c_278_n 0.00531816f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_54 VPB N_VPWR_c_311_n 0.0105574f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.325
cc_55 VPB N_VPWR_c_312_n 0.0476707f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_56 VPB N_VPWR_c_313_n 0.00271285f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=0.56
cc_57 VPB N_VPWR_c_314_n 0.0113853f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.985
cc_58 VPB N_VPWR_c_315_n 0.0312537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_316_n 0.0195868f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_60 VPB N_VPWR_c_317_n 0.0048162f $X=-0.19 $Y=1.305 $X2=1.115 $Y2=1.16
cc_61 VPB N_VPWR_c_318_n 0.0424511f $X=-0.19 $Y=1.305 $X2=2.83 $Y2=2.38
cc_62 VPB N_VPWR_c_310_n 0.0425769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB X 9.753e-19 $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.985
cc_64 N_A_108_21#_M1011_g N_A1_M1004_g 0.0170252f $X=1.115 $Y=1.985 $X2=0 $Y2=0
cc_65 N_A_108_21#_c_76_n N_A1_M1004_g 0.00201299f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_108_21#_c_78_n N_A1_M1004_g 0.0109966f $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_67 N_A_108_21#_c_85_p N_A1_M1004_g 0.0147648f $X=1.735 $Y=2.295 $X2=0 $Y2=0
cc_68 N_A_108_21#_c_86_p N_A1_M1004_g 0.00500312f $X=1.82 $Y=2.38 $X2=0 $Y2=0
cc_69 N_A_108_21#_c_76_n A1 0.0214385f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_108_21#_c_69_n A1 0.00195764f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_108_21#_c_78_n A1 0.029767f $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_72 N_A_108_21#_c_76_n N_A1_c_174_n 5.86485e-19 $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_108_21#_c_69_n N_A1_c_174_n 0.0218666f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_108_21#_c_78_n N_A1_c_174_n 0.00285216f $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_75 N_A_108_21#_c_67_n N_A1_c_175_n 0.00783657f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_108_21#_c_78_n N_A2_M1001_g 6.63228e-19 $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_77 N_A_108_21#_c_85_p N_A2_M1001_g 0.00499689f $X=1.735 $Y=2.295 $X2=0 $Y2=0
cc_78 N_A_108_21#_c_96_p N_A2_M1001_g 0.00984966f $X=2.83 $Y=2.38 $X2=0 $Y2=0
cc_79 N_A_108_21#_c_78_n A2 0.00921084f $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_80 N_A_108_21#_c_96_p A2 0.0106994f $X=2.83 $Y=2.38 $X2=0 $Y2=0
cc_81 N_A_108_21#_c_96_p N_A3_M1005_g 0.010625f $X=2.83 $Y=2.38 $X2=0 $Y2=0
cc_82 N_A_108_21#_c_100_p N_A3_M1005_g 7.54408e-19 $X=2.955 $Y=1.665 $X2=0 $Y2=0
cc_83 N_A_108_21#_c_101_p N_A3_M1005_g 0.00559579f $X=2.955 $Y=2.295 $X2=0 $Y2=0
cc_84 N_A_108_21#_c_96_p A3 0.0131377f $X=2.83 $Y=2.38 $X2=0 $Y2=0
cc_85 N_A_108_21#_c_96_p N_B1_M1006_g 0.00204575f $X=2.83 $Y=2.38 $X2=0 $Y2=0
cc_86 N_A_108_21#_c_100_p N_B1_M1006_g 7.32094e-19 $X=2.955 $Y=1.665 $X2=0 $Y2=0
cc_87 N_A_108_21#_c_101_p N_B1_M1006_g 0.0150705f $X=2.955 $Y=2.295 $X2=0 $Y2=0
cc_88 N_A_108_21#_c_80_n N_B1_M1006_g 0.0127201f $X=3.425 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_108_21#_c_100_p B1 0.0160964f $X=2.955 $Y=1.665 $X2=0 $Y2=0
cc_90 N_A_108_21#_c_80_n B1 0.0109744f $X=3.425 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_108_21#_c_70_n B1 0.0265259f $X=3.51 $Y=1.495 $X2=0 $Y2=0
cc_92 N_A_108_21#_c_71_n B1 0.00948181f $X=3.275 $Y=0.36 $X2=0 $Y2=0
cc_93 N_A_108_21#_c_100_p N_B1_c_278_n 0.00381184f $X=2.955 $Y=1.665 $X2=0 $Y2=0
cc_94 N_A_108_21#_c_70_n N_B1_c_278_n 0.00753568f $X=3.51 $Y=1.495 $X2=0 $Y2=0
cc_95 N_A_108_21#_c_71_n N_B1_c_278_n 0.0023839f $X=3.275 $Y=0.36 $X2=0 $Y2=0
cc_96 N_A_108_21#_c_70_n N_B1_c_279_n 0.00408814f $X=3.51 $Y=1.495 $X2=0 $Y2=0
cc_97 N_A_108_21#_c_78_n N_VPWR_M1011_d 0.00434929f $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_98 N_A_108_21#_c_80_n N_VPWR_M1006_d 0.00777396f $X=3.425 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A_108_21#_M1000_g N_VPWR_c_312_n 0.0240327f $X=0.615 $Y=1.985 $X2=0
+ $Y2=0
cc_100 N_A_108_21#_M1000_g N_VPWR_c_313_n 9.72969e-19 $X=0.615 $Y=1.985 $X2=0
+ $Y2=0
cc_101 N_A_108_21#_M1011_g N_VPWR_c_313_n 0.0127611f $X=1.115 $Y=1.985 $X2=0
+ $Y2=0
cc_102 N_A_108_21#_c_78_n N_VPWR_c_313_n 0.0188752f $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_103 N_A_108_21#_c_79_n N_VPWR_c_313_n 0.00197512f $X=1.2 $Y=1.53 $X2=0 $Y2=0
cc_104 N_A_108_21#_c_85_p N_VPWR_c_313_n 0.0375609f $X=1.735 $Y=2.295 $X2=0
+ $Y2=0
cc_105 N_A_108_21#_c_86_p N_VPWR_c_313_n 0.0139612f $X=1.82 $Y=2.38 $X2=0 $Y2=0
cc_106 N_A_108_21#_c_80_n N_VPWR_c_315_n 0.028122f $X=3.425 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A_108_21#_M1000_g N_VPWR_c_316_n 0.00374367f $X=0.615 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_108_21#_M1011_g N_VPWR_c_316_n 0.00486043f $X=1.115 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_108_21#_c_96_p N_VPWR_c_318_n 0.0725033f $X=2.83 $Y=2.38 $X2=0 $Y2=0
cc_110 N_A_108_21#_c_86_p N_VPWR_c_318_n 0.00979741f $X=1.82 $Y=2.38 $X2=0 $Y2=0
cc_111 N_A_108_21#_M1005_d N_VPWR_c_310_n 0.00341579f $X=2.63 $Y=1.485 $X2=0
+ $Y2=0
cc_112 N_A_108_21#_M1000_g N_VPWR_c_310_n 0.00693752f $X=0.615 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_108_21#_M1011_g N_VPWR_c_310_n 0.00847989f $X=1.115 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_108_21#_c_96_p N_VPWR_c_310_n 0.0456869f $X=2.83 $Y=2.38 $X2=0 $Y2=0
cc_115 N_A_108_21#_c_86_p N_VPWR_c_310_n 0.00618115f $X=1.82 $Y=2.38 $X2=0 $Y2=0
cc_116 N_A_108_21#_c_66_n X 0.00658616f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_108_21#_c_68_n X 0.00290026f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_108_21#_c_76_n X 0.0167586f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_108_21#_M1000_g X 0.0181119f $X=0.615 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_108_21#_c_66_n X 0.00279725f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_108_21#_M1011_g X 0.005479f $X=1.115 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_108_21#_c_68_n X 0.00151846f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_108_21#_c_76_n X 0.0115216f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_108_21#_c_79_n X 0.00866303f $X=1.2 $Y=1.53 $X2=0 $Y2=0
cc_125 N_A_108_21#_c_68_n N_X_c_357_n 0.00582195f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_108_21#_c_65_n X 0.00710709f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_108_21#_c_66_n X 0.0042679f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_108_21#_c_67_n X 0.00400284f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_108_21#_c_68_n X 0.0041365f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_108_21#_c_76_n X 0.00564724f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_108_21#_c_65_n N_X_c_375_n 0.0113819f $X=0.615 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_108_21#_c_66_n N_X_c_375_n 0.0038784f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_108_21#_M1000_g X 0.0125862f $X=0.615 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_108_21#_c_66_n X 0.00275532f $X=1.04 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_108_21#_c_78_n A_346_297# 0.00113639f $X=1.65 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_108_21#_c_85_p A_346_297# 0.00624788f $X=1.735 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_137 N_A_108_21#_c_96_p A_346_297# 0.00580081f $X=2.83 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_138 N_A_108_21#_c_86_p A_346_297# 3.22723e-19 $X=1.82 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_139 N_A_108_21#_c_96_p A_430_297# 0.00938948f $X=2.83 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_140 N_A_108_21#_c_65_n N_VGND_c_399_n 0.0173387f $X=0.615 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_108_21#_c_65_n N_VGND_c_400_n 0.00103077f $X=0.615 $Y=0.995 $X2=0
+ $Y2=0
cc_142 N_A_108_21#_c_67_n N_VGND_c_400_n 0.0122541f $X=1.115 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_108_21#_c_76_n N_VGND_c_400_n 0.00277103f $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A_108_21#_c_69_n N_VGND_c_400_n 0.00106074f $X=1.115 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_108_21#_c_78_n N_VGND_c_400_n 0.00469622f $X=1.65 $Y=1.53 $X2=0 $Y2=0
cc_146 N_A_108_21#_c_65_n N_VGND_c_401_n 0.00376303f $X=0.615 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A_108_21#_c_67_n N_VGND_c_401_n 0.0046653f $X=1.115 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_108_21#_c_71_n N_VGND_c_404_n 0.0320206f $X=3.275 $Y=0.36 $X2=0 $Y2=0
cc_149 N_A_108_21#_M1010_d N_VGND_c_405_n 0.00250309f $X=3.11 $Y=0.235 $X2=0
+ $Y2=0
cc_150 N_A_108_21#_c_65_n N_VGND_c_405_n 0.00693946f $X=0.615 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_A_108_21#_c_67_n N_VGND_c_405_n 0.00817276f $X=1.115 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_108_21#_c_71_n N_VGND_c_405_n 0.0185458f $X=3.275 $Y=0.36 $X2=0 $Y2=0
cc_153 N_A_108_21#_c_100_p N_A_346_47#_c_453_n 7.86906e-19 $X=2.955 $Y=1.665
+ $X2=0 $Y2=0
cc_154 N_A_108_21#_c_78_n N_A_346_47#_c_454_n 0.00130321f $X=1.65 $Y=1.53 $X2=0
+ $Y2=0
cc_155 N_A1_c_175_n N_A2_c_206_n 0.0235606f $X=1.595 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A1_M1004_g N_A2_M1001_g 0.0602645f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_157 A1 A2 0.0206392f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A1_c_174_n A2 6.78235e-19 $X=1.595 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A1_M1004_g A2 0.00280499f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_160 A1 N_A2_c_208_n 0.00159548f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A1_c_174_n N_A2_c_208_n 0.020542f $X=1.595 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A1_M1004_g N_VPWR_c_313_n 0.00510722f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A1_M1004_g N_VPWR_c_318_n 0.00463936f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A1_M1004_g N_VPWR_c_310_n 0.00809909f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_165 A1 N_VGND_c_400_n 0.017196f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A1_c_174_n N_VGND_c_400_n 7.77033e-19 $X=1.595 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A1_c_175_n N_VGND_c_400_n 0.0108291f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A1_c_175_n N_VGND_c_403_n 0.0046653f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_175_n N_VGND_c_405_n 0.00799591f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_c_175_n N_VGND_c_406_n 5.59196e-19 $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A2_c_206_n N_A3_c_242_n 0.0218007f $X=2.075 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_172 N_A2_M1001_g N_A3_M1005_g 0.0477842f $X=2.075 $Y=1.985 $X2=0 $Y2=0
cc_173 A2 N_A3_M1005_g 9.18397e-19 $X=1.99 $Y=1.445 $X2=0 $Y2=0
cc_174 N_A2_M1001_g A3 0.00263562f $X=2.075 $Y=1.985 $X2=0 $Y2=0
cc_175 A2 A3 0.0550984f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A2_c_208_n A3 0.00185237f $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_177 A2 N_A3_c_244_n 3.8169e-19 $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A2_c_208_n N_A3_c_244_n 0.0203414f $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A2_M1001_g N_VPWR_c_318_n 0.00357877f $X=2.075 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_VPWR_c_310_n 0.00546655f $X=2.075 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A2_c_206_n N_VGND_c_400_n 6.91082e-19 $X=2.075 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_c_206_n N_VGND_c_403_n 0.00342417f $X=2.075 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_c_206_n N_VGND_c_405_n 0.00405449f $X=2.075 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_c_206_n N_VGND_c_406_n 0.00707893f $X=2.075 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A2_c_206_n N_A_346_47#_c_453_n 0.0104349f $X=2.075 $Y=0.995 $X2=0 $Y2=0
cc_186 A2 N_A_346_47#_c_453_n 0.0149998f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A2_c_208_n N_A_346_47#_c_453_n 4.76779e-19 $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A3_M1005_g N_B1_M1006_g 0.0231582f $X=2.555 $Y=1.985 $X2=0 $Y2=0
cc_189 A3 N_B1_M1006_g 0.00281575f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_190 A3 B1 0.0217777f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A3_c_244_n B1 0.00207233f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_192 A3 N_B1_c_278_n 3.51722e-19 $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_193 N_A3_c_244_n N_B1_c_278_n 0.0203288f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A3_c_242_n N_B1_c_279_n 0.0188926f $X=2.555 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A3_M1005_g N_VPWR_c_318_n 0.00357877f $X=2.555 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A3_M1005_g N_VPWR_c_310_n 0.00581352f $X=2.555 $Y=1.985 $X2=0 $Y2=0
cc_197 A3 A_430_297# 0.0062622f $X=2.45 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_198 N_A3_c_242_n N_VGND_c_404_n 0.00256813f $X=2.555 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A3_c_242_n N_VGND_c_405_n 0.00335748f $X=2.555 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A3_c_242_n N_VGND_c_406_n 0.0101098f $X=2.555 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A3_c_242_n N_A_346_47#_c_453_n 0.0103396f $X=2.555 $Y=0.995 $X2=0 $Y2=0
cc_202 A3 N_A_346_47#_c_453_n 0.016853f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A3_c_244_n N_A_346_47#_c_453_n 0.00138218f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A3_c_242_n N_A_346_47#_c_461_n 0.00462294f $X=2.555 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_B1_M1006_g N_VPWR_c_315_n 0.0170878f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B1_M1006_g N_VPWR_c_318_n 0.00547432f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1006_g N_VPWR_c_310_n 0.0111484f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_c_279_n N_VGND_c_404_n 0.00585385f $X=3.052 $Y=0.995 $X2=0 $Y2=0
cc_209 N_B1_c_279_n N_VGND_c_405_n 0.0119949f $X=3.052 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B1_c_279_n N_VGND_c_406_n 0.00119839f $X=3.052 $Y=0.995 $X2=0 $Y2=0
cc_211 B1 N_A_346_47#_c_453_n 0.0054881f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_212 N_B1_c_278_n N_A_346_47#_c_453_n 8.18609e-19 $X=3.035 $Y=1.16 $X2=0 $Y2=0
cc_213 N_VPWR_c_310_n N_X_M1000_s 0.00457293f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_312_n X 0.0778839f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_215 N_VPWR_c_313_n X 0.00243345f $X=1.385 $Y=1.96 $X2=0 $Y2=0
cc_216 N_VPWR_c_312_n N_X_c_357_n 0.0251894f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_217 N_VPWR_c_316_n X 0.028227f $X=1.165 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_310_n X 0.0161501f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_310_n A_346_297# 0.00216824f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_220 N_VPWR_c_310_n A_430_297# 0.00265018f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_221 N_X_c_357_n N_VGND_c_399_n 0.0251894f $X=0.55 $Y=1.185 $X2=0 $Y2=0
cc_222 N_X_c_375_n N_VGND_c_399_n 0.0501637f $X=0.825 $Y=0.36 $X2=0 $Y2=0
cc_223 N_X_c_375_n N_VGND_c_401_n 0.0264535f $X=0.825 $Y=0.36 $X2=0 $Y2=0
cc_224 N_X_M1002_s N_VGND_c_405_n 0.00457664f $X=0.69 $Y=0.235 $X2=0 $Y2=0
cc_225 N_X_c_375_n N_VGND_c_405_n 0.0160507f $X=0.825 $Y=0.36 $X2=0 $Y2=0
cc_226 N_VGND_c_405_n N_A_346_47#_M1009_d 0.00412745f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_227 N_VGND_c_405_n N_A_346_47#_M1008_d 0.00370961f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_403_n N_A_346_47#_c_466_n 0.0112554f $X=2.12 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_405_n N_A_346_47#_c_466_n 0.00644035f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_M1007_d N_A_346_47#_c_453_n 0.00943141f $X=2.15 $Y=0.235 $X2=0
+ $Y2=0
cc_231 N_VGND_c_403_n N_A_346_47#_c_453_n 0.00233324f $X=2.12 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_404_n N_A_346_47#_c_453_n 0.00230733f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_405_n N_A_346_47#_c_453_n 0.0102298f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_406_n N_A_346_47#_c_453_n 0.022823f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_404_n N_A_346_47#_c_461_n 0.0146061f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_c_405_n N_A_346_47#_c_461_n 0.00874048f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_406_n N_A_346_47#_c_461_n 0.0176937f $X=2.53 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nor2_4.spice.SKY130_FD_SC_HD__NOR2_4.pxi
* Created: Thu Aug 27 14:31:24 2020
* 
x_PM_SKY130_FD_SC_HD__NOR2_4%A N_A_c_68_n N_A_M1002_g N_A_M1001_g N_A_c_69_n
+ N_A_M1003_g N_A_M1010_g N_A_c_70_n N_A_M1007_g N_A_M1012_g N_A_c_71_n
+ N_A_M1008_g N_A_M1015_g A A N_A_c_72_n N_A_c_73_n PM_SKY130_FD_SC_HD__NOR2_4%A
x_PM_SKY130_FD_SC_HD__NOR2_4%B N_B_c_148_n N_B_M1004_g N_B_M1000_g N_B_c_149_n
+ N_B_M1009_g N_B_M1005_g N_B_c_150_n N_B_M1011_g N_B_M1006_g N_B_c_151_n
+ N_B_M1014_g N_B_M1013_g B N_B_c_160_n N_B_c_152_n PM_SKY130_FD_SC_HD__NOR2_4%B
x_PM_SKY130_FD_SC_HD__NOR2_4%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1010_s
+ N_A_27_297#_M1015_s N_A_27_297#_M1005_d N_A_27_297#_M1013_d
+ N_A_27_297#_c_236_n N_A_27_297#_c_237_n N_A_27_297#_c_238_n
+ N_A_27_297#_c_279_p N_A_27_297#_c_239_n N_A_27_297#_c_240_n
+ N_A_27_297#_c_254_n N_A_27_297#_c_262_n N_A_27_297#_c_264_n
+ N_A_27_297#_c_268_n N_A_27_297#_c_241_n N_A_27_297#_c_270_n
+ N_A_27_297#_c_242_n PM_SKY130_FD_SC_HD__NOR2_4%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR2_4%VPWR N_VPWR_M1001_d N_VPWR_M1012_d N_VPWR_c_314_n
+ N_VPWR_c_315_n VPWR N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n
+ N_VPWR_c_313_n N_VPWR_c_320_n N_VPWR_c_321_n PM_SKY130_FD_SC_HD__NOR2_4%VPWR
x_PM_SKY130_FD_SC_HD__NOR2_4%Y N_Y_M1002_d N_Y_M1007_d N_Y_M1004_s N_Y_M1011_s
+ N_Y_M1000_s N_Y_M1006_s N_Y_c_383_n N_Y_c_369_n N_Y_c_370_n N_Y_c_394_n
+ N_Y_c_371_n N_Y_c_399_n N_Y_c_378_n N_Y_c_444_n N_Y_c_379_n N_Y_c_372_n
+ N_Y_c_421_n N_Y_c_449_n N_Y_c_380_n N_Y_c_373_n N_Y_c_374_n N_Y_c_375_n
+ N_Y_c_376_n N_Y_c_381_n Y PM_SKY130_FD_SC_HD__NOR2_4%Y
x_PM_SKY130_FD_SC_HD__NOR2_4%VGND N_VGND_M1002_s N_VGND_M1003_s N_VGND_M1008_s
+ N_VGND_M1009_d N_VGND_M1014_d N_VGND_c_490_n N_VGND_c_491_n N_VGND_c_492_n
+ N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n
+ N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ N_VGND_c_503_n VGND N_VGND_c_504_n N_VGND_c_505_n
+ PM_SKY130_FD_SC_HD__NOR2_4%VGND
cc_1 VNB N_A_c_68_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_69_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_A_c_70_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_A_c_71_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB N_A_c_72_n 0.0151855f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_6 VNB N_A_c_73_n 0.0705772f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_7 VNB N_B_c_148_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B_c_149_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_9 VNB N_B_c_150_n 0.0157984f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_10 VNB N_B_c_151_n 0.0192147f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_11 VNB N_B_c_152_n 0.0667613f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_12 VNB N_VPWR_c_313_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_13 VNB N_Y_c_369_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_14 VNB N_Y_c_370_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_15 VNB N_Y_c_371_n 0.00410518f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_16 VNB N_Y_c_372_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_17 VNB N_Y_c_373_n 0.0151086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_374_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_375_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_376_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB Y 0.0241147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_490_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_23 VNB N_VGND_c_491_n 0.0332455f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.325
cc_24 VNB N_VGND_c_492_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_25 VNB N_VGND_c_493_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_26 VNB N_VGND_c_494_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_27 VNB N_VGND_c_495_n 0.0179705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_496_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_29 VNB N_VGND_c_497_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_30 VNB N_VGND_c_498_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_31 VNB N_VGND_c_499_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_32 VNB N_VGND_c_500_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_33 VNB N_VGND_c_501_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_502_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_503_n 0.00545092f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_36 VNB N_VGND_c_504_n 0.0108937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_505_n 0.220103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_A_M1001_g 0.0250431f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_39 VPB N_A_M1010_g 0.0179946f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_40 VPB N_A_M1012_g 0.0179946f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_41 VPB N_A_M1015_g 0.0184982f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_42 VPB N_A_c_73_n 0.0108808f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_43 VPB N_B_M1000_g 0.0186339f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_44 VPB N_B_M1005_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_45 VPB N_B_M1006_g 0.0181185f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_46 VPB N_B_M1013_g 0.022018f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_47 VPB N_B_c_152_n 0.0102634f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_48 VPB N_A_27_297#_c_236_n 0.0119249f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_49 VPB N_A_27_297#_c_237_n 0.0307403f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.325
cc_50 VPB N_A_27_297#_c_238_n 0.00315624f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_51 VPB N_A_27_297#_c_239_n 0.00269564f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_52 VPB N_A_27_297#_c_240_n 0.00422862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_297#_c_241_n 0.00131915f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_54 VPB N_A_27_297#_c_242_n 0.0252915f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_55 VPB N_VPWR_c_314_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_56 VPB N_VPWR_c_315_n 0.00221708f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_57 VPB N_VPWR_c_316_n 0.015553f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_58 VPB N_VPWR_c_317_n 0.0124915f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.995
cc_59 VPB N_VPWR_c_318_n 0.0618174f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_60 VPB N_VPWR_c_313_n 0.0512465f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_61 VPB N_VPWR_c_320_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_62 VPB N_VPWR_c_321_n 0.00353635f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_63 VPB N_Y_c_378_n 0.00158719f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_64 VPB N_Y_c_379_n 0.00311424f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.16
cc_65 VPB N_Y_c_380_n 0.0024274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_Y_c_381_n 0.00127413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB Y 0.0319103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 N_A_c_71_n N_B_c_148_n 0.0199001f $X=1.75 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_69 N_A_M1015_g N_B_M1000_g 0.0199001f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A_c_72_n N_B_c_160_n 0.0100567f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_73_n N_B_c_160_n 8.57456e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_72_n N_B_c_152_n 8.57456e-19 $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_c_73_n N_B_c_152_n 0.0199001f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_c_72_n N_A_27_297#_c_236_n 0.018453f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_M1001_g N_A_27_297#_c_238_n 0.0138748f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1010_g N_A_27_297#_c_238_n 0.0136248f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_c_72_n N_A_27_297#_c_238_n 0.046205f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_c_73_n N_A_27_297#_c_238_n 0.00213789f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_M1012_g N_A_27_297#_c_239_n 0.0136248f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_M1015_g N_A_27_297#_c_239_n 0.0118246f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_c_72_n N_A_27_297#_c_239_n 0.0404893f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_c_73_n N_A_27_297#_c_239_n 0.00213789f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1015_g N_A_27_297#_c_240_n 0.00167295f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_c_72_n N_A_27_297#_c_240_n 3.67829e-19 $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_M1012_g N_A_27_297#_c_254_n 4.50937e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1015_g N_A_27_297#_c_254_n 0.00997294f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_c_72_n N_A_27_297#_c_241_n 0.0132812f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_c_73_n N_A_27_297#_c_241_n 0.00221654f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_M1001_g N_VPWR_c_314_n 0.0129691f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_M1010_g N_VPWR_c_314_n 0.0110282f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_M1012_g N_VPWR_c_314_n 6.32588e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_M1010_g N_VPWR_c_315_n 6.27883e-19 $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_M1012_g N_VPWR_c_315_n 0.0106598f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_M1015_g N_VPWR_c_315_n 0.00279634f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_M1001_g N_VPWR_c_316_n 0.0046653f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_M1010_g N_VPWR_c_317_n 0.0046653f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_M1012_g N_VPWR_c_317_n 0.0046653f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_M1015_g N_VPWR_c_318_n 0.00539841f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_M1001_g N_VPWR_c_313_n 0.00886468f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_M1010_g N_VPWR_c_313_n 0.00789179f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_M1012_g N_VPWR_c_313_n 0.00789179f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_M1015_g N_VPWR_c_313_n 0.00949176f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_c_68_n N_Y_c_383_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_69_n N_Y_c_383_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_c_70_n N_Y_c_383_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_c_69_n N_Y_c_369_n 0.00870364f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_c_70_n N_Y_c_369_n 0.00870364f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_c_72_n N_Y_c_369_n 0.036111f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_c_73_n N_Y_c_369_n 0.00222133f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_c_68_n N_Y_c_370_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_c_69_n N_Y_c_370_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_c_72_n N_Y_c_370_n 0.0265405f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_c_73_n N_Y_c_370_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_c_69_n N_Y_c_394_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_c_70_n N_Y_c_394_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_c_71_n N_Y_c_394_n 0.00630972f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_c_71_n N_Y_c_371_n 0.00896662f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_72_n N_Y_c_371_n 0.00651491f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_c_71_n N_Y_c_399_n 5.22228e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_70_n N_Y_c_374_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_c_71_n N_Y_c_374_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_72_n N_Y_c_374_n 0.0265405f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_c_73_n N_Y_c_374_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_c_68_n N_VGND_c_491_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_72_n N_VGND_c_491_n 0.019131f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_c_69_n N_VGND_c_492_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_70_n N_VGND_c_492_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_71_n N_VGND_c_493_n 0.00146448f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_68_n N_VGND_c_496_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_69_n N_VGND_c_496_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_70_n N_VGND_c_498_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_71_n N_VGND_c_498_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_68_n N_VGND_c_505_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_69_n N_VGND_c_505_n 0.0057163f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_70_n N_VGND_c_505_n 0.0057163f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_71_n N_VGND_c_505_n 0.0057435f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B_M1000_g N_A_27_297#_c_240_n 0.00329439f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B_c_160_n N_A_27_297#_c_240_n 3.67829e-19 $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B_M1000_g N_A_27_297#_c_254_n 0.00843121f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B_M1005_g N_A_27_297#_c_254_n 5.461e-19 $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B_M1000_g N_A_27_297#_c_262_n 0.0101149f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B_M1005_g N_A_27_297#_c_262_n 0.00795376f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B_M1000_g N_A_27_297#_c_264_n 4.89808e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B_M1005_g N_A_27_297#_c_264_n 0.00534818f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B_M1006_g N_A_27_297#_c_264_n 0.00534818f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_146 N_B_M1013_g N_A_27_297#_c_264_n 4.89808e-19 $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_147 N_B_M1006_g N_A_27_297#_c_268_n 0.00795376f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B_M1013_g N_A_27_297#_c_268_n 0.00853389f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B_M1005_g N_A_27_297#_c_270_n 7.04098e-19 $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B_M1006_g N_A_27_297#_c_270_n 7.04098e-19 $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B_M1006_g N_A_27_297#_c_242_n 5.77441e-19 $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B_M1013_g N_A_27_297#_c_242_n 0.00674479f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B_M1000_g N_VPWR_c_318_n 0.00357835f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B_M1005_g N_VPWR_c_318_n 0.00357835f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_155 N_B_M1006_g N_VPWR_c_318_n 0.00357835f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_156 N_B_M1013_g N_VPWR_c_318_n 0.00359354f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_157 N_B_M1000_g N_VPWR_c_313_n 0.00525234f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_158 N_B_M1005_g N_VPWR_c_313_n 0.00522513f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B_M1006_g N_VPWR_c_313_n 0.00522513f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B_M1013_g N_VPWR_c_313_n 0.00633431f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_161 N_B_c_148_n N_Y_c_394_n 5.22228e-19 $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B_c_148_n N_Y_c_371_n 0.00896662f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B_c_160_n N_Y_c_371_n 0.00651491f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B_c_148_n N_Y_c_399_n 0.00630972f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_165 N_B_c_149_n N_Y_c_399_n 0.00630972f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_166 N_B_c_150_n N_Y_c_399_n 5.22228e-19 $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B_M1000_g N_Y_c_378_n 5.53367e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_168 N_B_c_160_n N_Y_c_378_n 0.0138639f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B_c_152_n N_Y_c_378_n 0.00222344f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B_M1005_g N_Y_c_379_n 0.0136843f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B_M1006_g N_Y_c_379_n 0.0137138f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_172 N_B_c_160_n N_Y_c_379_n 0.0494751f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B_c_152_n N_Y_c_379_n 0.00217081f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B_c_149_n N_Y_c_372_n 0.00870364f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B_c_150_n N_Y_c_372_n 0.00870364f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B_c_160_n N_Y_c_372_n 0.036111f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B_c_152_n N_Y_c_372_n 0.00222133f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B_c_149_n N_Y_c_421_n 5.22228e-19 $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B_c_150_n N_Y_c_421_n 0.00630972f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B_c_151_n N_Y_c_421_n 0.0109314f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B_M1013_g N_Y_c_380_n 0.0173729f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B_c_160_n N_Y_c_380_n 0.0130728f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B_c_151_n N_Y_c_373_n 0.0109523f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_160_n N_Y_c_373_n 0.0068596f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_185 N_B_c_148_n N_Y_c_375_n 0.00113286f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B_c_149_n N_Y_c_375_n 0.00113286f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B_c_160_n N_Y_c_375_n 0.0265405f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B_c_152_n N_Y_c_375_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B_c_150_n N_Y_c_376_n 0.00113286f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B_c_151_n N_Y_c_376_n 0.00113286f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B_c_160_n N_Y_c_376_n 0.0265405f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B_c_152_n N_Y_c_376_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B_c_160_n N_Y_c_381_n 0.0138639f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B_c_152_n N_Y_c_381_n 0.00222344f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_195 N_B_c_151_n Y 0.0196229f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B_c_160_n Y 0.016859f $X=3.315 $Y=1.16 $X2=0 $Y2=0
cc_197 N_B_c_148_n N_VGND_c_493_n 0.00146448f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B_c_149_n N_VGND_c_494_n 0.00146448f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B_c_150_n N_VGND_c_494_n 0.00146448f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B_c_151_n N_VGND_c_495_n 0.00322989f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B_c_148_n N_VGND_c_500_n 0.00423334f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B_c_149_n N_VGND_c_500_n 0.00423334f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B_c_150_n N_VGND_c_502_n 0.00423334f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B_c_151_n N_VGND_c_502_n 0.00423334f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B_c_148_n N_VGND_c_505_n 0.0057435f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B_c_149_n N_VGND_c_505_n 0.0057163f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B_c_150_n N_VGND_c_505_n 0.0057163f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_208 N_B_c_151_n N_VGND_c_505_n 0.00683455f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_27_297#_c_238_n N_VPWR_M1001_d 0.00166915f $X=1.035 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_210 N_A_27_297#_c_239_n N_VPWR_M1012_d 0.00166915f $X=1.795 $Y=1.56 $X2=0
+ $Y2=0
cc_211 N_A_27_297#_c_238_n N_VPWR_c_314_n 0.0172742f $X=1.035 $Y=1.56 $X2=0
+ $Y2=0
cc_212 N_A_27_297#_c_239_n N_VPWR_c_315_n 0.0150746f $X=1.795 $Y=1.56 $X2=0
+ $Y2=0
cc_213 N_A_27_297#_c_237_n N_VPWR_c_316_n 0.019049f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_214 N_A_27_297#_c_279_p N_VPWR_c_317_n 0.0113958f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_215 N_A_27_297#_c_254_n N_VPWR_c_318_n 0.0190403f $X=1.96 $Y=2.295 $X2=0
+ $Y2=0
cc_216 N_A_27_297#_c_262_n N_VPWR_c_318_n 0.0286211f $X=2.635 $Y=2.38 $X2=0
+ $Y2=0
cc_217 N_A_27_297#_c_268_n N_VPWR_c_318_n 0.0286474f $X=3.475 $Y=2.38 $X2=0
+ $Y2=0
cc_218 N_A_27_297#_c_270_n N_VPWR_c_318_n 0.0187749f $X=2.8 $Y=2.38 $X2=0 $Y2=0
cc_219 N_A_27_297#_c_242_n N_VPWR_c_318_n 0.0267299f $X=3.64 $Y=2 $X2=0 $Y2=0
cc_220 N_A_27_297#_M1001_s N_VPWR_c_313_n 0.00399293f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_221 N_A_27_297#_M1010_s N_VPWR_c_313_n 0.00562358f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_222 N_A_27_297#_M1015_s N_VPWR_c_313_n 0.00215201f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_223 N_A_27_297#_M1005_d N_VPWR_c_313_n 0.00215201f $X=2.665 $Y=1.485 $X2=0
+ $Y2=0
cc_224 N_A_27_297#_M1013_d N_VPWR_c_313_n 0.00217517f $X=3.505 $Y=1.485 $X2=0
+ $Y2=0
cc_225 N_A_27_297#_c_237_n N_VPWR_c_313_n 0.0105137f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_226 N_A_27_297#_c_279_p N_VPWR_c_313_n 0.00646998f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_227 N_A_27_297#_c_254_n N_VPWR_c_313_n 0.0122896f $X=1.96 $Y=2.295 $X2=0
+ $Y2=0
cc_228 N_A_27_297#_c_262_n N_VPWR_c_313_n 0.0178969f $X=2.635 $Y=2.38 $X2=0
+ $Y2=0
cc_229 N_A_27_297#_c_268_n N_VPWR_c_313_n 0.0179004f $X=3.475 $Y=2.38 $X2=0
+ $Y2=0
cc_230 N_A_27_297#_c_270_n N_VPWR_c_313_n 0.0122096f $X=2.8 $Y=2.38 $X2=0 $Y2=0
cc_231 N_A_27_297#_c_242_n N_VPWR_c_313_n 0.0156135f $X=3.64 $Y=2 $X2=0 $Y2=0
cc_232 N_A_27_297#_c_262_n N_Y_M1000_s 0.00312348f $X=2.635 $Y=2.38 $X2=0 $Y2=0
cc_233 N_A_27_297#_c_268_n N_Y_M1006_s 0.00312348f $X=3.475 $Y=2.38 $X2=0 $Y2=0
cc_234 N_A_27_297#_c_240_n N_Y_c_371_n 0.0115682f $X=1.96 $Y=1.665 $X2=0 $Y2=0
cc_235 N_A_27_297#_c_240_n N_Y_c_378_n 0.010246f $X=1.96 $Y=1.665 $X2=0 $Y2=0
cc_236 N_A_27_297#_c_262_n N_Y_c_444_n 0.0118865f $X=2.635 $Y=2.38 $X2=0 $Y2=0
cc_237 N_A_27_297#_M1005_d N_Y_c_379_n 0.00176936f $X=2.665 $Y=1.485 $X2=0 $Y2=0
cc_238 N_A_27_297#_c_262_n N_Y_c_379_n 0.00321626f $X=2.635 $Y=2.38 $X2=0 $Y2=0
cc_239 N_A_27_297#_c_264_n N_Y_c_379_n 0.0159581f $X=2.8 $Y=2.02 $X2=0 $Y2=0
cc_240 N_A_27_297#_c_268_n N_Y_c_379_n 0.00321626f $X=3.475 $Y=2.38 $X2=0 $Y2=0
cc_241 N_A_27_297#_c_268_n N_Y_c_449_n 0.0118865f $X=3.475 $Y=2.38 $X2=0 $Y2=0
cc_242 N_A_27_297#_M1013_d N_Y_c_380_n 9.9523e-19 $X=3.505 $Y=1.485 $X2=0 $Y2=0
cc_243 N_A_27_297#_c_268_n N_Y_c_380_n 0.00322918f $X=3.475 $Y=2.38 $X2=0 $Y2=0
cc_244 N_A_27_297#_c_242_n N_Y_c_380_n 0.00991777f $X=3.64 $Y=2 $X2=0 $Y2=0
cc_245 N_A_27_297#_M1013_d Y 0.00262315f $X=3.505 $Y=1.485 $X2=0 $Y2=0
cc_246 N_A_27_297#_c_242_n Y 0.0211657f $X=3.64 $Y=2 $X2=0 $Y2=0
cc_247 N_A_27_297#_c_236_n N_VGND_c_491_n 0.00202255f $X=0.227 $Y=1.665 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_313_n N_Y_M1000_s 0.00216833f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_c_313_n N_Y_M1006_s 0.00216833f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_250 N_Y_c_369_n N_VGND_M1003_s 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_251 N_Y_c_371_n N_VGND_M1008_s 0.00162089f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_252 N_Y_c_372_n N_VGND_M1009_d 0.00162089f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_253 N_Y_c_373_n N_VGND_M1014_d 0.00285206f $X=3.655 $Y=0.815 $X2=0 $Y2=0
cc_254 N_Y_c_370_n N_VGND_c_491_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_255 N_Y_c_369_n N_VGND_c_492_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_256 N_Y_c_371_n N_VGND_c_493_n 0.0122559f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_257 N_Y_c_372_n N_VGND_c_494_n 0.0122559f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_258 N_Y_c_373_n N_VGND_c_495_n 0.0234351f $X=3.655 $Y=0.815 $X2=0 $Y2=0
cc_259 N_Y_c_383_n N_VGND_c_496_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_260 N_Y_c_369_n N_VGND_c_496_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_261 N_Y_c_369_n N_VGND_c_498_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_262 N_Y_c_394_n N_VGND_c_498_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_263 N_Y_c_371_n N_VGND_c_498_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_264 N_Y_c_371_n N_VGND_c_500_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_265 N_Y_c_399_n N_VGND_c_500_n 0.0188551f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_266 N_Y_c_372_n N_VGND_c_500_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_267 N_Y_c_372_n N_VGND_c_502_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_268 N_Y_c_421_n N_VGND_c_502_n 0.0188551f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_269 N_Y_c_373_n N_VGND_c_502_n 0.00198695f $X=3.655 $Y=0.815 $X2=0 $Y2=0
cc_270 N_Y_c_373_n N_VGND_c_504_n 0.00365233f $X=3.655 $Y=0.815 $X2=0 $Y2=0
cc_271 N_Y_M1002_d N_VGND_c_505_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_272 N_Y_M1007_d N_VGND_c_505_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_273 N_Y_M1004_s N_VGND_c_505_n 0.00215201f $X=2.245 $Y=0.235 $X2=0 $Y2=0
cc_274 N_Y_M1011_s N_VGND_c_505_n 0.00215201f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_275 N_Y_c_383_n N_VGND_c_505_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_276 N_Y_c_369_n N_VGND_c_505_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_277 N_Y_c_394_n N_VGND_c_505_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_278 N_Y_c_371_n N_VGND_c_505_n 0.00835832f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_279 N_Y_c_399_n N_VGND_c_505_n 0.0122069f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_280 N_Y_c_372_n N_VGND_c_505_n 0.00835832f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_281 N_Y_c_421_n N_VGND_c_505_n 0.0122069f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_282 N_Y_c_373_n N_VGND_c_505_n 0.0111264f $X=3.655 $Y=0.815 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dlrtp_2.pxi.spice
* Created: Thu Aug 27 14:17:35 2020
* 
x_PM_SKY130_FD_SC_HD__DLRTP_2%GATE N_GATE_c_147_n N_GATE_c_142_n N_GATE_M1020_g
+ N_GATE_c_148_n N_GATE_M1010_g N_GATE_c_143_n N_GATE_c_149_n GATE GATE
+ N_GATE_c_145_n N_GATE_c_146_n PM_SKY130_FD_SC_HD__DLRTP_2%GATE
x_PM_SKY130_FD_SC_HD__DLRTP_2%A_27_47# N_A_27_47#_M1020_s N_A_27_47#_M1010_s
+ N_A_27_47#_M1012_g N_A_27_47#_M1000_g N_A_27_47#_M1002_g N_A_27_47#_c_186_n
+ N_A_27_47#_c_187_n N_A_27_47#_M1018_g N_A_27_47#_c_199_n N_A_27_47#_c_189_n
+ N_A_27_47#_c_190_n N_A_27_47#_c_191_n N_A_27_47#_c_200_n N_A_27_47#_c_201_n
+ N_A_27_47#_c_192_n N_A_27_47#_c_193_n N_A_27_47#_c_203_n N_A_27_47#_c_204_n
+ N_A_27_47#_c_205_n N_A_27_47#_c_206_n N_A_27_47#_c_207_n N_A_27_47#_c_208_n
+ N_A_27_47#_c_194_n PM_SKY130_FD_SC_HD__DLRTP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRTP_2%D N_D_M1003_g N_D_M1016_g D N_D_c_338_n
+ N_D_c_339_n PM_SKY130_FD_SC_HD__DLRTP_2%D
x_PM_SKY130_FD_SC_HD__DLRTP_2%A_299_47# N_A_299_47#_M1003_s N_A_299_47#_M1016_s
+ N_A_299_47#_c_375_n N_A_299_47#_M1007_g N_A_299_47#_M1013_g
+ N_A_299_47#_c_383_n N_A_299_47#_c_377_n N_A_299_47#_c_378_n
+ N_A_299_47#_c_379_n N_A_299_47#_c_385_n N_A_299_47#_c_380_n
+ N_A_299_47#_c_381_n PM_SKY130_FD_SC_HD__DLRTP_2%A_299_47#
x_PM_SKY130_FD_SC_HD__DLRTP_2%A_193_47# N_A_193_47#_M1012_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1017_g N_A_193_47#_M1001_g N_A_193_47#_c_461_n
+ N_A_193_47#_c_462_n N_A_193_47#_c_463_n N_A_193_47#_c_464_n
+ N_A_193_47#_c_468_n N_A_193_47#_c_469_n N_A_193_47#_c_470_n
+ N_A_193_47#_c_471_n N_A_193_47#_c_472_n N_A_193_47#_c_473_n
+ N_A_193_47#_c_474_n PM_SKY130_FD_SC_HD__DLRTP_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRTP_2%A_711_307# N_A_711_307#_M1019_s
+ N_A_711_307#_M1006_d N_A_711_307#_M1011_g N_A_711_307#_M1005_g
+ N_A_711_307#_M1009_g N_A_711_307#_c_588_n N_A_711_307#_M1004_g
+ N_A_711_307#_c_589_n N_A_711_307#_M1008_g N_A_711_307#_M1014_g
+ N_A_711_307#_c_598_n N_A_711_307#_c_599_n N_A_711_307#_c_590_n
+ N_A_711_307#_c_591_n N_A_711_307#_c_612_p N_A_711_307#_c_630_p
+ N_A_711_307#_c_645_p N_A_711_307#_c_592_n N_A_711_307#_c_600_n
+ N_A_711_307#_c_633_p N_A_711_307#_c_608_p N_A_711_307#_c_609_p
+ N_A_711_307#_c_593_n PM_SKY130_FD_SC_HD__DLRTP_2%A_711_307#
x_PM_SKY130_FD_SC_HD__DLRTP_2%A_560_47# N_A_560_47#_M1017_d N_A_560_47#_M1002_d
+ N_A_560_47#_M1019_g N_A_560_47#_M1006_g N_A_560_47#_c_735_n
+ N_A_560_47#_c_736_n N_A_560_47#_c_744_n N_A_560_47#_c_745_n
+ N_A_560_47#_c_737_n N_A_560_47#_c_762_n N_A_560_47#_c_741_n
+ N_A_560_47#_c_738_n N_A_560_47#_c_739_n PM_SKY130_FD_SC_HD__DLRTP_2%A_560_47#
x_PM_SKY130_FD_SC_HD__DLRTP_2%RESET_B N_RESET_B_M1015_g N_RESET_B_M1021_g
+ RESET_B N_RESET_B_c_828_n N_RESET_B_c_829_n N_RESET_B_c_830_n
+ N_RESET_B_c_831_n RESET_B PM_SKY130_FD_SC_HD__DLRTP_2%RESET_B
x_PM_SKY130_FD_SC_HD__DLRTP_2%VPWR N_VPWR_M1010_d N_VPWR_M1016_d N_VPWR_M1011_d
+ N_VPWR_M1006_s N_VPWR_M1021_d N_VPWR_M1014_s N_VPWR_c_876_n N_VPWR_c_877_n
+ N_VPWR_c_878_n N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n
+ N_VPWR_c_883_n VPWR N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n
+ N_VPWR_c_887_n N_VPWR_c_888_n N_VPWR_c_889_n N_VPWR_c_890_n N_VPWR_c_891_n
+ N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_875_n PM_SKY130_FD_SC_HD__DLRTP_2%VPWR
x_PM_SKY130_FD_SC_HD__DLRTP_2%Q N_Q_M1004_d N_Q_M1009_d N_Q_c_992_n N_Q_c_996_n
+ N_Q_c_1000_n N_Q_c_1003_n N_Q_c_990_n Q Q Q N_Q_c_989_n Q
+ PM_SKY130_FD_SC_HD__DLRTP_2%Q
x_PM_SKY130_FD_SC_HD__DLRTP_2%VGND N_VGND_M1020_d N_VGND_M1003_d N_VGND_M1005_d
+ N_VGND_M1015_d N_VGND_M1008_s N_VGND_c_1035_n N_VGND_c_1036_n N_VGND_c_1037_n
+ N_VGND_c_1038_n N_VGND_c_1039_n N_VGND_c_1040_n VGND N_VGND_c_1041_n
+ N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n N_VGND_c_1045_n
+ N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n N_VGND_c_1049_n
+ N_VGND_c_1050_n PM_SKY130_FD_SC_HD__DLRTP_2%VGND
cc_1 VNB N_GATE_c_142_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_c_143_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE 0.0127963f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_c_145_n 0.0210048f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_c_146_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1012_g 0.0396846f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_186_n 0.0121234f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_c_187_n 0.00503399f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_9 VNB N_A_27_47#_M1018_g 0.0440053f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_10 VNB N_A_27_47#_c_189_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_190_n 0.00225297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_191_n 0.00809684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_192_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_193_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_194_n 0.0230161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1003_g 0.025882f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_17 VNB N_D_M1016_g 0.00623852f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_338_n 0.00396738f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_19 VNB N_D_c_339_n 0.0437054f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_20 VNB N_A_299_47#_c_375_n 0.0166791f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_21 VNB N_A_299_47#_M1013_g 0.0129633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_377_n 0.0021682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_47#_c_378_n 0.0053306f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_24 VNB N_A_299_47#_c_379_n 0.00331308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_299_47#_c_380_n 0.00282063f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_26 VNB N_A_299_47#_c_381_n 0.0266195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_M1017_g 0.0208902f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_28 VNB N_A_193_47#_c_461_n 0.0139557f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_29 VNB N_A_193_47#_c_462_n 0.0077229f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_30 VNB N_A_193_47#_c_463_n 0.0257799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_193_47#_c_464_n 0.00401932f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_32 VNB N_A_711_307#_M1005_g 0.0512645f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_33 VNB N_A_711_307#_c_588_n 0.0158942f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_34 VNB N_A_711_307#_c_589_n 0.019249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_711_307#_c_590_n 0.00478966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_711_307#_c_591_n 0.00340829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_711_307#_c_592_n 0.00111867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_711_307#_c_593_n 0.0401273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_560_47#_M1019_g 0.0243249f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_40 VNB N_A_560_47#_M1006_g 4.92816e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_41 VNB N_A_560_47#_c_735_n 0.0503735f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_42 VNB N_A_560_47#_c_736_n 0.0070289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_560_47#_c_737_n 0.00369082f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_44 VNB N_A_560_47#_c_738_n 0.00645421f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.53
cc_45 VNB N_A_560_47#_c_739_n 0.0105366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_828_n 0.0188248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_829_n 0.00310136f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_48 VNB N_RESET_B_c_830_n 0.0172478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_831_n 0.00251297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VPWR_c_875_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB Q 0.019138f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_52 VNB N_Q_c_989_n 0.00583f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.53
cc_53 VNB N_VGND_c_1035_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1036_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1037_n 0.00595133f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_56 VNB N_VGND_c_1038_n 0.00415973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1039_n 0.00988417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1040_n 0.0186875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1041_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1042_n 0.0270169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1043_n 0.040267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1044_n 0.0318162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1045_n 0.0173295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1046_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1047_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1048_n 0.00520851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1049_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1050_n 0.331845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VPB N_GATE_c_147_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_70 VPB N_GATE_c_148_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_71 VPB N_GATE_c_149_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_72 VPB GATE 0.0153801f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_73 VPB N_GATE_c_145_n 0.0106763f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_74 VPB N_A_27_47#_M1000_g 0.0394751f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_75 VPB N_A_27_47#_M1002_g 0.0300054f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_76 VPB N_A_27_47#_c_186_n 0.0171269f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_77 VPB N_A_27_47#_c_187_n 0.00734368f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_78 VPB N_A_27_47#_c_199_n 0.012166f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_79 VPB N_A_27_47#_c_200_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_201_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_192_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_203_n 0.0203003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_204_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_205_n 0.0054554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_206_n 0.00344459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_207_n 0.0062631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_47#_c_208_n 0.00916151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_47#_c_194_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_D_M1016_g 0.046254f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_90 VPB N_D_c_338_n 0.00249607f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_91 VPB N_A_299_47#_M1013_g 0.0366914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_299_47#_c_383_n 0.00820942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_299_47#_c_379_n 0.00343957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_299_47#_c_385_n 0.00734292f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_95 VPB N_A_193_47#_M1001_g 0.0203874f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_96 VPB N_A_193_47#_c_461_n 0.00798859f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_97 VPB N_A_193_47#_c_464_n 0.0023883f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_98 VPB N_A_193_47#_c_468_n 0.00290734f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_99 VPB N_A_193_47#_c_469_n 0.00816718f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.19
cc_100 VPB N_A_193_47#_c_470_n 0.00237364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_193_47#_c_471_n 0.00694487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_193_47#_c_472_n 0.00245022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_193_47#_c_473_n 0.0261435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_193_47#_c_474_n 0.00852821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_711_307#_M1011_g 0.0291391f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_106 VPB N_A_711_307#_M1005_g 0.0187255f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_107 VPB N_A_711_307#_M1009_g 0.0178942f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_108 VPB N_A_711_307#_M1014_g 0.0226986f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_109 VPB N_A_711_307#_c_598_n 0.00811709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_711_307#_c_599_n 0.0428181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_711_307#_c_600_n 0.00160584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_711_307#_c_593_n 0.00715816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_560_47#_M1006_g 0.0272227f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_114 VPB N_A_560_47#_c_741_n 0.00808746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_560_47#_c_738_n 0.00392171f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.53
cc_116 VPB N_A_560_47#_c_739_n 0.00401579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_RESET_B_M1021_g 0.0194172f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_118 VPB N_RESET_B_c_828_n 0.00406519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_RESET_B_c_829_n 0.00160346f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_120 VPB N_RESET_B_c_831_n 0.00205786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_876_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_877_n 0.00362994f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_123 VPB N_VPWR_c_878_n 0.00867107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_879_n 0.00598254f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.53
cc_125 VPB N_VPWR_c_880_n 0.00117743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_881_n 3.31047e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_882_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_883_n 0.0359186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_884_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_885_n 0.0292658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_886_n 0.039475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_887_n 0.014719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_888_n 0.0156539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_889_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_890_n 0.00413931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_891_n 0.00651127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_892_n 0.00423502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_893_n 0.00456844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_875_n 0.0572825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_Q_c_990_n 0.00642382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB Q 0.00390984f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_142 N_GATE_c_142_n N_A_27_47#_M1012_g 0.0187834f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_143 N_GATE_c_146_n N_A_27_47#_M1012_g 0.00419721f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_144 N_GATE_c_149_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_145 N_GATE_c_145_n N_A_27_47#_M1000_g 0.00527139f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_146 N_GATE_c_142_n N_A_27_47#_c_190_n 0.00674622f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_147 N_GATE_c_143_n N_A_27_47#_c_190_n 0.0105293f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_148 N_GATE_c_143_n N_A_27_47#_c_191_n 0.00672951f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_149 GATE N_A_27_47#_c_191_n 0.0198215f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_150 N_GATE_c_145_n N_A_27_47#_c_191_n 7.3212e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_151 N_GATE_c_148_n N_A_27_47#_c_200_n 0.0135489f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_152 N_GATE_c_149_n N_A_27_47#_c_200_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_153 N_GATE_c_148_n N_A_27_47#_c_201_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_154 N_GATE_c_149_n N_A_27_47#_c_201_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_155 GATE N_A_27_47#_c_201_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_156 N_GATE_c_145_n N_A_27_47#_c_201_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_157 N_GATE_c_145_n N_A_27_47#_c_192_n 0.00319349f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_158 N_GATE_c_143_n N_A_27_47#_c_193_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_159 GATE N_A_27_47#_c_193_n 0.0288278f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_160 N_GATE_c_146_n N_A_27_47#_c_193_n 0.00151818f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_161 N_GATE_c_147_n N_A_27_47#_c_204_n 0.0033897f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_162 N_GATE_c_149_n N_A_27_47#_c_204_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_163 GATE N_A_27_47#_c_204_n 0.00653562f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_164 N_GATE_c_147_n N_A_27_47#_c_205_n 7.602e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_165 N_GATE_c_149_n N_A_27_47#_c_205_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_166 GATE N_A_27_47#_c_194_n 9.06856e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_167 N_GATE_c_145_n N_A_27_47#_c_194_n 0.0165768f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_168 N_GATE_c_148_n N_VPWR_c_876_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_169 N_GATE_c_148_n N_VPWR_c_884_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_170 N_GATE_c_148_n N_VPWR_c_875_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_171 N_GATE_c_142_n N_VGND_c_1035_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_172 N_GATE_c_142_n N_VGND_c_1041_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_173 N_GATE_c_143_n N_VGND_c_1041_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_174 N_GATE_c_142_n N_VGND_c_1050_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_203_n N_D_M1016_g 0.00650345f $X=2.39 $Y=1.53 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_203_n N_D_c_338_n 0.00872077f $X=2.39 $Y=1.53 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1012_g N_D_c_339_n 0.00556424f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A_27_47#_M1002_g N_A_299_47#_M1013_g 0.0361306f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_187_n N_A_299_47#_M1013_g 0.0249798f $X=2.805 $Y=1.325 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_203_n N_A_299_47#_M1013_g 0.00512637f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_206_n N_A_299_47#_M1013_g 0.00142929f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_207_n N_A_299_47#_M1013_g 0.0023158f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_203_n N_A_299_47#_c_383_n 5.17324e-19 $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_207_n N_A_299_47#_c_383_n 5.26803e-19 $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_203_n N_A_299_47#_c_378_n 0.00730284f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_203_n N_A_299_47#_c_379_n 0.0112022f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_206_n N_A_299_47#_c_379_n 0.00124596f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_207_n N_A_299_47#_c_379_n 0.00574185f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_203_n N_A_299_47#_c_385_n 0.0201053f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_206_n N_A_299_47#_c_385_n 0.00130924f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_207_n N_A_299_47#_c_385_n 0.00667388f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_203_n N_A_299_47#_c_381_n 0.00107604f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1018_g N_A_193_47#_M1017_g 0.0193168f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1002_g N_A_193_47#_M1001_g 0.0194728f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1012_g N_A_193_47#_c_461_n 0.00777428f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_190_n N_A_193_47#_c_461_n 0.0100297f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_192_n N_A_193_47#_c_461_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_193_n N_A_193_47#_c_461_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_203_n N_A_193_47#_c_461_n 0.0183875f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_204_n N_A_193_47#_c_461_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_205_n N_A_193_47#_c_461_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_187_n N_A_193_47#_c_462_n 0.002062f $X=2.805 $Y=1.325 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1018_g N_A_193_47#_c_462_n 0.0022579f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_206_n N_A_193_47#_c_462_n 5.78162e-19 $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_207_n N_A_193_47#_c_462_n 0.00712428f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_187_n N_A_193_47#_c_463_n 0.0210448f $X=2.805 $Y=1.325 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1018_g N_A_193_47#_c_463_n 0.0157692f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_207_n N_A_193_47#_c_463_n 5.58275e-19 $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_186_n N_A_193_47#_c_464_n 0.0133783f $X=3.135 $Y=1.325 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_M1018_g N_A_193_47#_c_464_n 0.0046954f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_206_n N_A_193_47#_c_464_n 9.31908e-19 $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_207_n N_A_193_47#_c_464_n 0.0145048f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_208_n N_A_193_47#_c_464_n 0.00382314f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_200_n N_A_193_47#_c_468_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_203_n N_A_193_47#_c_468_n 0.00195186f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_194_n N_A_193_47#_c_468_n 0.00777428f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_M1002_g N_A_193_47#_c_469_n 0.00742914f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_218 N_A_27_47#_c_186_n N_A_193_47#_c_469_n 0.00109188f $X=3.135 $Y=1.325
+ $X2=0 $Y2=0
cc_219 N_A_27_47#_c_199_n N_A_193_47#_c_469_n 0.00192289f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_203_n N_A_193_47#_c_469_n 0.0854152f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_206_n N_A_193_47#_c_469_n 0.0266191f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_207_n N_A_193_47#_c_469_n 0.00975596f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_M1000_g N_A_193_47#_c_470_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_200_n N_A_193_47#_c_470_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_203_n N_A_193_47#_c_470_n 0.0259095f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_205_n N_A_193_47#_c_470_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_M1000_g N_A_193_47#_c_471_n 0.00777428f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1002_g N_A_193_47#_c_472_n 0.00145302f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_229 N_A_27_47#_c_186_n N_A_193_47#_c_472_n 0.00134584f $X=3.135 $Y=1.325
+ $X2=0 $Y2=0
cc_230 N_A_27_47#_M1002_g N_A_193_47#_c_473_n 0.0117523f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_186_n N_A_193_47#_c_473_n 0.0176547f $X=3.135 $Y=1.325 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_199_n N_A_193_47#_c_473_n 0.00459274f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_M1002_g N_A_193_47#_c_474_n 0.00486506f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_234 N_A_27_47#_c_186_n N_A_193_47#_c_474_n 0.00459229f $X=3.135 $Y=1.325
+ $X2=0 $Y2=0
cc_235 N_A_27_47#_c_199_n N_A_193_47#_c_474_n 0.00140206f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_206_n N_A_193_47#_c_474_n 4.84725e-19 $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_207_n N_A_193_47#_c_474_n 0.00836787f $X=2.535 $Y=1.53 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_M1018_g N_A_711_307#_M1005_g 0.0461684f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1018_g N_A_560_47#_c_744_n 0.0140034f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1002_g N_A_560_47#_c_745_n 0.00383536f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_241 N_A_27_47#_M1018_g N_A_560_47#_c_737_n 0.00990974f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_186_n N_A_560_47#_c_741_n 7.3591e-19 $X=3.135 $Y=1.325 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_186_n N_A_560_47#_c_738_n 0.00238788f $X=3.135 $Y=1.325
+ $X2=0 $Y2=0
cc_244 N_A_27_47#_M1018_g N_A_560_47#_c_738_n 0.00589168f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_200_n N_VPWR_M1010_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_246 N_A_27_47#_M1000_g N_VPWR_c_876_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_200_n N_VPWR_c_876_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_201_n N_VPWR_c_876_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_204_n N_VPWR_c_876_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_250 N_A_27_47#_M1002_g N_VPWR_c_877_n 0.00387673f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_203_n N_VPWR_c_877_n 0.00172226f $X=2.39 $Y=1.53 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_200_n N_VPWR_c_884_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_201_n N_VPWR_c_884_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_254 N_A_27_47#_M1000_g N_VPWR_c_885_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1002_g N_VPWR_c_886_n 0.0054153f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1000_g N_VPWR_c_875_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1002_g N_VPWR_c_875_n 0.00634589f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_200_n N_VPWR_c_875_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_201_n N_VPWR_c_875_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_190_n N_VGND_M1020_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_261 N_A_27_47#_M1012_g N_VGND_c_1035_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_190_n N_VGND_c_1035_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_192_n N_VGND_c_1035_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_194_n N_VGND_c_1035_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1018_g N_VGND_c_1037_n 0.00177134f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_189_n N_VGND_c_1041_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_190_n N_VGND_c_1041_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1012_g N_VGND_c_1042_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1018_g N_VGND_c_1043_n 0.00379791f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1020_s N_VGND_c_1050_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1012_g N_VGND_c_1050_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1018_g N_VGND_c_1050_n 0.00569125f $X=3.21 $Y=0.415 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_189_n N_VGND_c_1050_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_190_n N_VGND_c_1050_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_275 N_D_M1003_g N_A_299_47#_c_375_n 0.0152898f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_276 N_D_c_339_n N_A_299_47#_M1013_g 0.0386497f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_277 N_D_M1016_g N_A_299_47#_c_383_n 0.0130693f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_278 N_D_M1003_g N_A_299_47#_c_377_n 0.0149989f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_279 N_D_c_338_n N_A_299_47#_c_377_n 0.0048234f $X=1.605 $Y=1.04 $X2=0 $Y2=0
cc_280 N_D_c_339_n N_A_299_47#_c_377_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_281 N_D_M1003_g N_A_299_47#_c_378_n 0.00582093f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_282 N_D_c_338_n N_A_299_47#_c_378_n 0.0107934f $X=1.605 $Y=1.04 $X2=0 $Y2=0
cc_283 N_D_c_338_n N_A_299_47#_c_379_n 0.0164825f $X=1.605 $Y=1.04 $X2=0 $Y2=0
cc_284 N_D_c_339_n N_A_299_47#_c_379_n 0.00572971f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_285 N_D_M1016_g N_A_299_47#_c_385_n 0.0125532f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_286 N_D_c_338_n N_A_299_47#_c_385_n 0.0227226f $X=1.605 $Y=1.04 $X2=0 $Y2=0
cc_287 N_D_c_339_n N_A_299_47#_c_385_n 0.00134698f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_288 N_D_M1003_g N_A_299_47#_c_380_n 0.00120861f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_289 N_D_c_338_n N_A_299_47#_c_380_n 0.0154978f $X=1.605 $Y=1.04 $X2=0 $Y2=0
cc_290 N_D_c_339_n N_A_299_47#_c_380_n 0.00475215f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_291 N_D_M1003_g N_A_299_47#_c_381_n 0.0203485f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_292 N_D_M1003_g N_A_193_47#_c_461_n 0.00203363f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_293 N_D_M1016_g N_A_193_47#_c_461_n 0.00456749f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_294 N_D_c_338_n N_A_193_47#_c_461_n 0.0221156f $X=1.605 $Y=1.04 $X2=0 $Y2=0
cc_295 N_D_c_339_n N_A_193_47#_c_461_n 0.00258308f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_296 N_D_M1016_g N_A_193_47#_c_468_n 0.00126017f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_297 N_D_M1016_g N_A_193_47#_c_469_n 0.00297192f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_298 N_D_M1016_g N_VPWR_c_877_n 0.0030264f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_299 N_D_M1016_g N_VPWR_c_885_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_300 N_D_M1016_g N_VPWR_c_875_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_301 N_D_M1003_g N_VGND_c_1036_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_302 N_D_M1003_g N_VGND_c_1042_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_303 N_D_M1003_g N_VGND_c_1050_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_304 N_D_c_339_n N_VGND_c_1050_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_305 N_A_299_47#_c_375_n N_A_193_47#_M1017_g 0.026216f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_306 N_A_299_47#_c_381_n N_A_193_47#_M1017_g 2.04413e-19 $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_307 N_A_299_47#_c_383_n N_A_193_47#_c_461_n 0.00118895f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_308 N_A_299_47#_c_385_n N_A_193_47#_c_461_n 0.00908469f $X=2.035 $Y=1.58
+ $X2=0 $Y2=0
cc_309 N_A_299_47#_c_380_n N_A_193_47#_c_461_n 0.0201829f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_310 N_A_299_47#_c_375_n N_A_193_47#_c_462_n 2.58725e-19 $X=2.25 $Y=0.765
+ $X2=0 $Y2=0
cc_311 N_A_299_47#_c_378_n N_A_193_47#_c_462_n 0.0184755f $X=2.035 $Y=1.095
+ $X2=0 $Y2=0
cc_312 N_A_299_47#_c_381_n N_A_193_47#_c_462_n 0.00179935f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_313 N_A_299_47#_c_378_n N_A_193_47#_c_463_n 3.08309e-19 $X=2.035 $Y=1.095
+ $X2=0 $Y2=0
cc_314 N_A_299_47#_c_381_n N_A_193_47#_c_463_n 0.0167221f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_315 N_A_299_47#_M1013_g N_A_193_47#_c_464_n 0.00376144f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_316 N_A_299_47#_c_378_n N_A_193_47#_c_464_n 0.00160321f $X=2.035 $Y=1.095
+ $X2=0 $Y2=0
cc_317 N_A_299_47#_c_381_n N_A_193_47#_c_464_n 9.02285e-19 $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_318 N_A_299_47#_c_383_n N_A_193_47#_c_468_n 0.0510205f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_319 N_A_299_47#_M1013_g N_A_193_47#_c_469_n 0.00397068f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_320 N_A_299_47#_c_383_n N_A_193_47#_c_469_n 0.0217612f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_321 N_A_299_47#_c_385_n N_A_193_47#_c_469_n 0.00557533f $X=2.035 $Y=1.58
+ $X2=0 $Y2=0
cc_322 N_A_299_47#_c_383_n N_A_193_47#_c_470_n 0.0027642f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_323 N_A_299_47#_c_375_n N_A_560_47#_c_744_n 6.66585e-19 $X=2.25 $Y=0.765
+ $X2=0 $Y2=0
cc_324 N_A_299_47#_M1013_g N_A_560_47#_c_745_n 5.02989e-19 $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_325 N_A_299_47#_M1013_g N_VPWR_c_877_n 0.0215213f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_326 N_A_299_47#_c_383_n N_VPWR_c_877_n 0.0234575f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_327 N_A_299_47#_c_385_n N_VPWR_c_877_n 0.0110105f $X=2.035 $Y=1.58 $X2=0
+ $Y2=0
cc_328 N_A_299_47#_c_383_n N_VPWR_c_885_n 0.0170306f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_329 N_A_299_47#_M1013_g N_VPWR_c_886_n 0.00290915f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_330 N_A_299_47#_M1016_s N_VPWR_c_875_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_331 N_A_299_47#_M1013_g N_VPWR_c_875_n 0.00321027f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_332 N_A_299_47#_c_383_n N_VPWR_c_875_n 0.00612385f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_333 N_A_299_47#_c_378_n N_VGND_M1003_d 0.00165422f $X=2.035 $Y=1.095 $X2=0
+ $Y2=0
cc_334 N_A_299_47#_c_375_n N_VGND_c_1036_n 0.00941159f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_377_n N_VGND_c_1036_n 0.0020169f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_336 N_A_299_47#_c_378_n N_VGND_c_1036_n 0.0152179f $X=2.035 $Y=1.095 $X2=0
+ $Y2=0
cc_337 N_A_299_47#_c_377_n N_VGND_c_1042_n 0.00255672f $X=1.95 $Y=0.7 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_380_n N_VGND_c_1042_n 0.00797702f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_339 N_A_299_47#_c_375_n N_VGND_c_1043_n 0.0046653f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_340 N_A_299_47#_c_381_n N_VGND_c_1043_n 9.48611e-19 $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_341 N_A_299_47#_M1003_s N_VGND_c_1050_n 0.00258726f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_342 N_A_299_47#_c_375_n N_VGND_c_1050_n 0.00440683f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_343 N_A_299_47#_c_377_n N_VGND_c_1050_n 0.00463926f $X=1.95 $Y=0.7 $X2=0
+ $Y2=0
cc_344 N_A_299_47#_c_378_n N_VGND_c_1050_n 0.00543344f $X=2.035 $Y=1.095 $X2=0
+ $Y2=0
cc_345 N_A_299_47#_c_380_n N_VGND_c_1050_n 0.0068025f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_c_381_n N_VGND_c_1050_n 0.00117722f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_347 N_A_193_47#_M1001_g N_A_711_307#_M1011_g 0.0258097f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_348 N_A_193_47#_c_473_n N_A_711_307#_c_599_n 0.0167011f $X=3.18 $Y=1.745
+ $X2=0 $Y2=0
cc_349 N_A_193_47#_c_474_n N_A_711_307#_c_599_n 4.54087e-19 $X=3.18 $Y=1.745
+ $X2=0 $Y2=0
cc_350 N_A_193_47#_M1017_g N_A_560_47#_c_744_n 0.00414674f $X=2.725 $Y=0.415
+ $X2=0 $Y2=0
cc_351 N_A_193_47#_c_462_n N_A_560_47#_c_744_n 0.0194231f $X=2.93 $Y=0.887 $X2=0
+ $Y2=0
cc_352 N_A_193_47#_c_463_n N_A_560_47#_c_744_n 6.54407e-19 $X=2.76 $Y=0.905
+ $X2=0 $Y2=0
cc_353 N_A_193_47#_M1001_g N_A_560_47#_c_745_n 0.00881123f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_354 N_A_193_47#_c_469_n N_A_560_47#_c_745_n 0.0022889f $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_193_47#_c_472_n N_A_560_47#_c_745_n 0.00219471f $X=3.01 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_193_47#_c_473_n N_A_560_47#_c_745_n 0.00219212f $X=3.18 $Y=1.745
+ $X2=0 $Y2=0
cc_357 N_A_193_47#_c_474_n N_A_560_47#_c_745_n 0.0134954f $X=3.18 $Y=1.745 $X2=0
+ $Y2=0
cc_358 N_A_193_47#_M1017_g N_A_560_47#_c_737_n 8.29815e-19 $X=2.725 $Y=0.415
+ $X2=0 $Y2=0
cc_359 N_A_193_47#_c_462_n N_A_560_47#_c_737_n 0.0205197f $X=2.93 $Y=0.887 $X2=0
+ $Y2=0
cc_360 N_A_193_47#_M1001_g N_A_560_47#_c_762_n 0.00349107f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_361 N_A_193_47#_M1001_g N_A_560_47#_c_741_n 0.00256184f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_362 N_A_193_47#_c_464_n N_A_560_47#_c_741_n 0.0112187f $X=3.015 $Y=1.57 $X2=0
+ $Y2=0
cc_363 N_A_193_47#_c_472_n N_A_560_47#_c_741_n 0.00136609f $X=3.01 $Y=1.87 $X2=0
+ $Y2=0
cc_364 N_A_193_47#_c_473_n N_A_560_47#_c_741_n 0.00167058f $X=3.18 $Y=1.745
+ $X2=0 $Y2=0
cc_365 N_A_193_47#_c_474_n N_A_560_47#_c_741_n 0.0292265f $X=3.18 $Y=1.745 $X2=0
+ $Y2=0
cc_366 N_A_193_47#_c_462_n N_A_560_47#_c_738_n 0.00383982f $X=2.93 $Y=0.887
+ $X2=0 $Y2=0
cc_367 N_A_193_47#_c_464_n N_A_560_47#_c_738_n 0.0223371f $X=3.015 $Y=1.57 $X2=0
+ $Y2=0
cc_368 N_A_193_47#_c_473_n N_A_560_47#_c_738_n 0.00218481f $X=3.18 $Y=1.745
+ $X2=0 $Y2=0
cc_369 N_A_193_47#_c_469_n N_VPWR_M1016_d 6.81311e-19 $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_471_n N_VPWR_c_876_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_c_469_n N_VPWR_c_877_n 0.0177393f $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_372 N_A_193_47#_c_472_n N_VPWR_c_877_n 9.43467e-19 $X=3.01 $Y=1.87 $X2=0
+ $Y2=0
cc_373 N_A_193_47#_c_474_n N_VPWR_c_877_n 0.00218193f $X=3.18 $Y=1.745 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_471_n N_VPWR_c_885_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_375 N_A_193_47#_M1001_g N_VPWR_c_886_n 0.00366111f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_376 N_A_193_47#_M1001_g N_VPWR_c_875_n 0.00539375f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_c_469_n N_VPWR_c_875_n 0.0748399f $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_378 N_A_193_47#_c_470_n N_VPWR_c_875_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_379 N_A_193_47#_c_471_n N_VPWR_c_875_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_380 N_A_193_47#_c_472_n N_VPWR_c_875_n 0.0146567f $X=3.01 $Y=1.87 $X2=0 $Y2=0
cc_381 N_A_193_47#_c_469_n A_465_369# 0.00393496f $X=2.865 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_193_47#_M1017_g N_VGND_c_1036_n 0.0018389f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_c_461_n N_VGND_c_1042_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_384 N_A_193_47#_M1017_g N_VGND_c_1043_n 0.00427327f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_385 N_A_193_47#_c_462_n N_VGND_c_1043_n 0.00265165f $X=2.93 $Y=0.887 $X2=0
+ $Y2=0
cc_386 N_A_193_47#_M1012_d N_VGND_c_1050_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_387 N_A_193_47#_M1017_g N_VGND_c_1050_n 0.00631563f $X=2.725 $Y=0.415 $X2=0
+ $Y2=0
cc_388 N_A_193_47#_c_461_n N_VGND_c_1050_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_389 N_A_193_47#_c_462_n N_VGND_c_1050_n 0.00469826f $X=2.93 $Y=0.887 $X2=0
+ $Y2=0
cc_390 N_A_711_307#_c_590_n N_A_560_47#_M1019_g 0.00818164f $X=4.415 $Y=0.4
+ $X2=0 $Y2=0
cc_391 N_A_711_307#_c_591_n N_A_560_47#_M1019_g 8.65818e-19 $X=4.58 $Y=0.74
+ $X2=0 $Y2=0
cc_392 N_A_711_307#_c_608_p N_A_560_47#_M1019_g 0.00848342f $X=4.955 $Y=0.76
+ $X2=0 $Y2=0
cc_393 N_A_711_307#_c_609_p N_A_560_47#_M1019_g 9.60405e-19 $X=5.095 $Y=0.76
+ $X2=0 $Y2=0
cc_394 N_A_711_307#_c_598_n N_A_560_47#_M1006_g 0.0172268f $X=4.8 $Y=1.7 $X2=0
+ $Y2=0
cc_395 N_A_711_307#_c_599_n N_A_560_47#_M1006_g 0.00528335f $X=3.86 $Y=1.7 $X2=0
+ $Y2=0
cc_396 N_A_711_307#_c_612_p N_A_560_47#_M1006_g 0.00671349f $X=4.885 $Y=2.27
+ $X2=0 $Y2=0
cc_397 N_A_711_307#_M1005_g N_A_560_47#_c_735_n 0.0175191f $X=3.685 $Y=0.445
+ $X2=0 $Y2=0
cc_398 N_A_711_307#_c_598_n N_A_560_47#_c_735_n 0.0113699f $X=4.8 $Y=1.7 $X2=0
+ $Y2=0
cc_399 N_A_711_307#_c_599_n N_A_560_47#_c_735_n 0.00132537f $X=3.86 $Y=1.7 $X2=0
+ $Y2=0
cc_400 N_A_711_307#_c_591_n N_A_560_47#_c_735_n 0.010168f $X=4.58 $Y=0.74 $X2=0
+ $Y2=0
cc_401 N_A_711_307#_M1005_g N_A_560_47#_c_744_n 0.0015515f $X=3.685 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_711_307#_M1011_g N_A_560_47#_c_745_n 0.00438393f $X=3.63 $Y=2.275
+ $X2=0 $Y2=0
cc_403 N_A_711_307#_M1005_g N_A_560_47#_c_737_n 0.00982596f $X=3.685 $Y=0.445
+ $X2=0 $Y2=0
cc_404 N_A_711_307#_M1011_g N_A_560_47#_c_762_n 0.00586723f $X=3.63 $Y=2.275
+ $X2=0 $Y2=0
cc_405 N_A_711_307#_M1011_g N_A_560_47#_c_741_n 0.0115949f $X=3.63 $Y=2.275
+ $X2=0 $Y2=0
cc_406 N_A_711_307#_M1005_g N_A_560_47#_c_741_n 0.00747368f $X=3.685 $Y=0.445
+ $X2=0 $Y2=0
cc_407 N_A_711_307#_c_598_n N_A_560_47#_c_741_n 0.0247809f $X=4.8 $Y=1.7 $X2=0
+ $Y2=0
cc_408 N_A_711_307#_c_599_n N_A_560_47#_c_741_n 0.0094011f $X=3.86 $Y=1.7 $X2=0
+ $Y2=0
cc_409 N_A_711_307#_c_599_n N_A_560_47#_c_738_n 4.42372e-19 $X=3.86 $Y=1.7 $X2=0
+ $Y2=0
cc_410 N_A_711_307#_M1005_g N_A_560_47#_c_739_n 0.0259371f $X=3.685 $Y=0.445
+ $X2=0 $Y2=0
cc_411 N_A_711_307#_c_598_n N_A_560_47#_c_739_n 0.0310195f $X=4.8 $Y=1.7 $X2=0
+ $Y2=0
cc_412 N_A_711_307#_c_599_n N_A_560_47#_c_739_n 0.00507019f $X=3.86 $Y=1.7 $X2=0
+ $Y2=0
cc_413 N_A_711_307#_M1009_g N_RESET_B_M1021_g 0.0285211f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_414 N_A_711_307#_c_630_p N_RESET_B_M1021_g 0.0125688f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_415 N_A_711_307#_c_600_n N_RESET_B_M1021_g 0.00311258f $X=5.5 $Y=1.535 $X2=0
+ $Y2=0
cc_416 N_A_711_307#_c_592_n N_RESET_B_c_828_n 4.85636e-19 $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_417 N_A_711_307#_c_633_p N_RESET_B_c_828_n 0.00134512f $X=4.885 $Y=1.755
+ $X2=0 $Y2=0
cc_418 N_A_711_307#_c_608_p N_RESET_B_c_828_n 0.00102737f $X=4.955 $Y=0.76 $X2=0
+ $Y2=0
cc_419 N_A_711_307#_c_609_p N_RESET_B_c_828_n 0.00139297f $X=5.095 $Y=0.76 $X2=0
+ $Y2=0
cc_420 N_A_711_307#_c_593_n N_RESET_B_c_828_n 0.0217393f $X=5.97 $Y=1.16 $X2=0
+ $Y2=0
cc_421 N_A_711_307#_c_630_p N_RESET_B_c_829_n 0.0133125f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_422 N_A_711_307#_c_592_n N_RESET_B_c_829_n 0.0230924f $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_423 N_A_711_307#_c_633_p N_RESET_B_c_829_n 0.0108676f $X=4.885 $Y=1.755 $X2=0
+ $Y2=0
cc_424 N_A_711_307#_c_608_p N_RESET_B_c_829_n 0.00902483f $X=4.955 $Y=0.76 $X2=0
+ $Y2=0
cc_425 N_A_711_307#_c_609_p N_RESET_B_c_829_n 0.0166122f $X=5.095 $Y=0.76 $X2=0
+ $Y2=0
cc_426 N_A_711_307#_c_593_n N_RESET_B_c_829_n 0.00199264f $X=5.97 $Y=1.16 $X2=0
+ $Y2=0
cc_427 N_A_711_307#_c_588_n N_RESET_B_c_830_n 0.0233647f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A_711_307#_c_590_n N_RESET_B_c_830_n 0.00148099f $X=4.415 $Y=0.4 $X2=0
+ $Y2=0
cc_429 N_A_711_307#_c_645_p N_RESET_B_c_830_n 0.00610473f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_430 N_A_711_307#_c_592_n N_RESET_B_c_830_n 0.00249115f $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_431 N_A_711_307#_c_609_p N_RESET_B_c_830_n 0.00731779f $X=5.095 $Y=0.76 $X2=0
+ $Y2=0
cc_432 N_A_711_307#_c_598_n N_RESET_B_c_831_n 0.0175697f $X=4.8 $Y=1.7 $X2=0
+ $Y2=0
cc_433 N_A_711_307#_c_591_n N_RESET_B_c_831_n 0.00584602f $X=4.58 $Y=0.74 $X2=0
+ $Y2=0
cc_434 N_A_711_307#_c_592_n N_RESET_B_c_831_n 0.00117696f $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_435 N_A_711_307#_c_633_p N_RESET_B_c_831_n 0.00111997f $X=4.885 $Y=1.755
+ $X2=0 $Y2=0
cc_436 N_A_711_307#_c_608_p N_RESET_B_c_831_n 0.0155084f $X=4.955 $Y=0.76 $X2=0
+ $Y2=0
cc_437 N_A_711_307#_c_598_n N_VPWR_M1006_s 0.00719583f $X=4.8 $Y=1.7 $X2=0 $Y2=0
cc_438 N_A_711_307#_c_630_p N_VPWR_M1021_d 0.00467552f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_439 N_A_711_307#_M1011_g N_VPWR_c_878_n 0.00462652f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_440 N_A_711_307#_c_598_n N_VPWR_c_878_n 0.0154733f $X=4.8 $Y=1.7 $X2=0 $Y2=0
cc_441 N_A_711_307#_c_599_n N_VPWR_c_878_n 0.00540932f $X=3.86 $Y=1.7 $X2=0
+ $Y2=0
cc_442 N_A_711_307#_M1011_g N_VPWR_c_880_n 0.00111884f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_443 N_A_711_307#_c_598_n N_VPWR_c_880_n 0.0124093f $X=4.8 $Y=1.7 $X2=0 $Y2=0
cc_444 N_A_711_307#_c_612_p N_VPWR_c_880_n 0.0184572f $X=4.885 $Y=2.27 $X2=0
+ $Y2=0
cc_445 N_A_711_307#_M1009_g N_VPWR_c_881_n 0.0120946f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_446 N_A_711_307#_M1014_g N_VPWR_c_881_n 7.64344e-19 $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_447 N_A_711_307#_c_630_p N_VPWR_c_881_n 0.0185412f $X=5.415 $Y=1.62 $X2=0
+ $Y2=0
cc_448 N_A_711_307#_M1014_g N_VPWR_c_883_n 0.00439898f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_449 N_A_711_307#_M1011_g N_VPWR_c_886_n 0.00522066f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_450 N_A_711_307#_c_612_p N_VPWR_c_887_n 0.0116048f $X=4.885 $Y=2.27 $X2=0
+ $Y2=0
cc_451 N_A_711_307#_M1009_g N_VPWR_c_888_n 0.00407992f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_452 N_A_711_307#_M1014_g N_VPWR_c_888_n 0.00541359f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_453 N_A_711_307#_M1006_d N_VPWR_c_875_n 0.00502345f $X=4.7 $Y=1.485 $X2=0
+ $Y2=0
cc_454 N_A_711_307#_M1011_g N_VPWR_c_875_n 0.0103672f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_455 N_A_711_307#_M1009_g N_VPWR_c_875_n 0.00706053f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_456 N_A_711_307#_M1014_g N_VPWR_c_875_n 0.0105459f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_457 N_A_711_307#_c_598_n N_VPWR_c_875_n 0.0169079f $X=4.8 $Y=1.7 $X2=0 $Y2=0
cc_458 N_A_711_307#_c_599_n N_VPWR_c_875_n 0.00112448f $X=3.86 $Y=1.7 $X2=0
+ $Y2=0
cc_459 N_A_711_307#_c_612_p N_VPWR_c_875_n 0.00646998f $X=4.885 $Y=2.27 $X2=0
+ $Y2=0
cc_460 N_A_711_307#_c_588_n N_Q_c_992_n 0.0037375f $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_461 N_A_711_307#_c_589_n N_Q_c_992_n 0.00971895f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_462 N_A_711_307#_c_592_n N_Q_c_992_n 0.00546544f $X=5.5 $Y=1.325 $X2=0 $Y2=0
cc_463 N_A_711_307#_c_609_p N_Q_c_992_n 0.00103283f $X=5.095 $Y=0.76 $X2=0 $Y2=0
cc_464 N_A_711_307#_c_588_n N_Q_c_996_n 0.00357088f $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_465 N_A_711_307#_c_589_n N_Q_c_996_n 0.00285458f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_466 N_A_711_307#_c_592_n N_Q_c_996_n 5.96903e-19 $X=5.5 $Y=1.325 $X2=0 $Y2=0
cc_467 N_A_711_307#_c_593_n N_Q_c_996_n 0.00115756f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_468 N_A_711_307#_M1009_g N_Q_c_1000_n 0.00280459f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_469 N_A_711_307#_M1014_g N_Q_c_1000_n 0.00283598f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_470 N_A_711_307#_c_593_n N_Q_c_1000_n 0.00228063f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_471 N_A_711_307#_M1009_g N_Q_c_1003_n 0.00476088f $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_472 N_A_711_307#_M1014_g N_Q_c_1003_n 0.0120309f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_473 N_A_711_307#_c_630_p N_Q_c_1003_n 0.0133619f $X=5.415 $Y=1.62 $X2=0 $Y2=0
cc_474 N_A_711_307#_c_600_n N_Q_c_1003_n 0.00238698f $X=5.5 $Y=1.535 $X2=0 $Y2=0
cc_475 N_A_711_307#_M1009_g N_Q_c_990_n 7.59735e-19 $X=5.515 $Y=1.985 $X2=0
+ $Y2=0
cc_476 N_A_711_307#_M1014_g N_Q_c_990_n 0.0110611f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_477 N_A_711_307#_c_600_n N_Q_c_990_n 0.00895287f $X=5.5 $Y=1.535 $X2=0 $Y2=0
cc_478 N_A_711_307#_c_593_n N_Q_c_990_n 9.62648e-19 $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_479 N_A_711_307#_M1014_g Q 0.00617274f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_480 N_A_711_307#_M1009_g Q 3.91463e-19 $X=5.515 $Y=1.985 $X2=0 $Y2=0
cc_481 N_A_711_307#_c_588_n Q 6.98001e-19 $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_482 N_A_711_307#_c_589_n Q 0.00417216f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_483 N_A_711_307#_M1014_g Q 0.00239602f $X=5.97 $Y=1.985 $X2=0 $Y2=0
cc_484 N_A_711_307#_c_592_n Q 0.0323847f $X=5.5 $Y=1.325 $X2=0 $Y2=0
cc_485 N_A_711_307#_c_600_n Q 0.00413456f $X=5.5 $Y=1.535 $X2=0 $Y2=0
cc_486 N_A_711_307#_c_593_n Q 0.0202112f $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_487 N_A_711_307#_c_588_n N_Q_c_989_n 8.32935e-19 $X=5.55 $Y=0.995 $X2=0 $Y2=0
cc_488 N_A_711_307#_c_589_n N_Q_c_989_n 0.00811298f $X=5.97 $Y=0.995 $X2=0 $Y2=0
cc_489 N_A_711_307#_c_592_n N_Q_c_989_n 0.0104813f $X=5.5 $Y=1.325 $X2=0 $Y2=0
cc_490 N_A_711_307#_c_593_n N_Q_c_989_n 8.81346e-19 $X=5.97 $Y=1.16 $X2=0 $Y2=0
cc_491 N_A_711_307#_c_645_p N_VGND_M1015_d 0.00566049f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_492 N_A_711_307#_c_592_n N_VGND_M1015_d 2.45523e-19 $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_493 N_A_711_307#_M1005_g N_VGND_c_1037_n 0.012404f $X=3.685 $Y=0.445 $X2=0
+ $Y2=0
cc_494 N_A_711_307#_c_590_n N_VGND_c_1037_n 0.0220941f $X=4.415 $Y=0.4 $X2=0
+ $Y2=0
cc_495 N_A_711_307#_c_588_n N_VGND_c_1038_n 0.00151665f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_496 N_A_711_307#_c_590_n N_VGND_c_1038_n 0.00663311f $X=4.415 $Y=0.4 $X2=0
+ $Y2=0
cc_497 N_A_711_307#_c_645_p N_VGND_c_1038_n 0.0123135f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_498 N_A_711_307#_c_592_n N_VGND_c_1038_n 2.57371e-19 $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_499 N_A_711_307#_c_589_n N_VGND_c_1040_n 0.00360303f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_500 N_A_711_307#_M1005_g N_VGND_c_1043_n 0.00427505f $X=3.685 $Y=0.445 $X2=0
+ $Y2=0
cc_501 N_A_711_307#_c_590_n N_VGND_c_1044_n 0.0215017f $X=4.415 $Y=0.4 $X2=0
+ $Y2=0
cc_502 N_A_711_307#_c_645_p N_VGND_c_1044_n 0.00196578f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_503 N_A_711_307#_c_608_p N_VGND_c_1044_n 0.00756134f $X=4.955 $Y=0.76 $X2=0
+ $Y2=0
cc_504 N_A_711_307#_c_588_n N_VGND_c_1045_n 0.00428558f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_A_711_307#_c_589_n N_VGND_c_1045_n 0.00539883f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_711_307#_c_592_n N_VGND_c_1045_n 0.00214121f $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_507 N_A_711_307#_M1019_s N_VGND_c_1050_n 0.00209319f $X=4.29 $Y=0.235 $X2=0
+ $Y2=0
cc_508 N_A_711_307#_M1005_g N_VGND_c_1050_n 0.00751607f $X=3.685 $Y=0.445 $X2=0
+ $Y2=0
cc_509 N_A_711_307#_c_588_n N_VGND_c_1050_n 0.00609476f $X=5.55 $Y=0.995 $X2=0
+ $Y2=0
cc_510 N_A_711_307#_c_589_n N_VGND_c_1050_n 0.00674774f $X=5.97 $Y=0.995 $X2=0
+ $Y2=0
cc_511 N_A_711_307#_c_590_n N_VGND_c_1050_n 0.0127527f $X=4.415 $Y=0.4 $X2=0
+ $Y2=0
cc_512 N_A_711_307#_c_645_p N_VGND_c_1050_n 0.00458246f $X=5.415 $Y=0.78 $X2=0
+ $Y2=0
cc_513 N_A_711_307#_c_592_n N_VGND_c_1050_n 0.0040434f $X=5.5 $Y=1.325 $X2=0
+ $Y2=0
cc_514 N_A_711_307#_c_608_p N_VGND_c_1050_n 0.0134135f $X=4.955 $Y=0.76 $X2=0
+ $Y2=0
cc_515 N_A_711_307#_c_608_p A_940_47# 0.00564009f $X=4.955 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_516 N_A_711_307#_c_609_p A_940_47# 7.75098e-19 $X=5.095 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_517 N_A_560_47#_M1006_g N_RESET_B_M1021_g 0.0203794f $X=4.625 $Y=1.985 $X2=0
+ $Y2=0
cc_518 N_A_560_47#_M1019_g N_RESET_B_c_828_n 0.0212403f $X=4.625 $Y=0.56 $X2=0
+ $Y2=0
cc_519 N_A_560_47#_M1019_g N_RESET_B_c_830_n 0.0348688f $X=4.625 $Y=0.56 $X2=0
+ $Y2=0
cc_520 N_A_560_47#_M1019_g N_RESET_B_c_831_n 0.00308864f $X=4.625 $Y=0.56 $X2=0
+ $Y2=0
cc_521 N_A_560_47#_M1006_g N_RESET_B_c_831_n 0.00345126f $X=4.625 $Y=1.985 $X2=0
+ $Y2=0
cc_522 N_A_560_47#_c_735_n N_RESET_B_c_831_n 0.00866392f $X=4.55 $Y=1.16 $X2=0
+ $Y2=0
cc_523 N_A_560_47#_c_736_n N_RESET_B_c_831_n 0.00623852f $X=4.625 $Y=1.16 $X2=0
+ $Y2=0
cc_524 N_A_560_47#_c_739_n N_RESET_B_c_831_n 0.0201209f $X=4.135 $Y=1.16 $X2=0
+ $Y2=0
cc_525 N_A_560_47#_c_745_n N_VPWR_c_877_n 0.00531509f $X=3.41 $Y=2.34 $X2=0
+ $Y2=0
cc_526 N_A_560_47#_M1006_g N_VPWR_c_878_n 9.6561e-19 $X=4.625 $Y=1.985 $X2=0
+ $Y2=0
cc_527 N_A_560_47#_M1006_g N_VPWR_c_880_n 0.00859988f $X=4.625 $Y=1.985 $X2=0
+ $Y2=0
cc_528 N_A_560_47#_M1006_g N_VPWR_c_881_n 6.43646e-19 $X=4.625 $Y=1.985 $X2=0
+ $Y2=0
cc_529 N_A_560_47#_c_745_n N_VPWR_c_886_n 0.0361033f $X=3.41 $Y=2.34 $X2=0 $Y2=0
cc_530 N_A_560_47#_c_741_n N_VPWR_c_886_n 4.40954e-19 $X=3.52 $Y=1.985 $X2=0
+ $Y2=0
cc_531 N_A_560_47#_M1006_g N_VPWR_c_887_n 0.00544582f $X=4.625 $Y=1.985 $X2=0
+ $Y2=0
cc_532 N_A_560_47#_M1002_d N_VPWR_c_875_n 0.00173835f $X=2.8 $Y=2.065 $X2=0
+ $Y2=0
cc_533 N_A_560_47#_M1006_g N_VPWR_c_875_n 0.00522142f $X=4.625 $Y=1.985 $X2=0
+ $Y2=0
cc_534 N_A_560_47#_c_745_n N_VPWR_c_875_n 0.021096f $X=3.41 $Y=2.34 $X2=0 $Y2=0
cc_535 N_A_560_47#_c_741_n N_VPWR_c_875_n 6.17842e-19 $X=3.52 $Y=1.985 $X2=0
+ $Y2=0
cc_536 N_A_560_47#_c_745_n A_644_413# 0.0056626f $X=3.41 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_537 N_A_560_47#_c_762_n A_644_413# 0.00197555f $X=3.495 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_538 N_A_560_47#_c_741_n A_644_413# 2.3925e-19 $X=3.52 $Y=1.985 $X2=-0.19
+ $Y2=-0.24
cc_539 N_A_560_47#_c_744_n N_VGND_c_1036_n 0.00233775f $X=3.27 $Y=0.45 $X2=0
+ $Y2=0
cc_540 N_A_560_47#_M1019_g N_VGND_c_1037_n 0.00235562f $X=4.625 $Y=0.56 $X2=0
+ $Y2=0
cc_541 N_A_560_47#_c_735_n N_VGND_c_1037_n 5.64862e-19 $X=4.55 $Y=1.16 $X2=0
+ $Y2=0
cc_542 N_A_560_47#_c_744_n N_VGND_c_1037_n 0.00942912f $X=3.27 $Y=0.45 $X2=0
+ $Y2=0
cc_543 N_A_560_47#_c_739_n N_VGND_c_1037_n 0.0127094f $X=4.135 $Y=1.16 $X2=0
+ $Y2=0
cc_544 N_A_560_47#_c_744_n N_VGND_c_1043_n 0.0225727f $X=3.27 $Y=0.45 $X2=0
+ $Y2=0
cc_545 N_A_560_47#_M1019_g N_VGND_c_1044_n 0.00415469f $X=4.625 $Y=0.56 $X2=0
+ $Y2=0
cc_546 N_A_560_47#_M1017_d N_VGND_c_1050_n 0.00284725f $X=2.8 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_A_560_47#_M1019_g N_VGND_c_1050_n 0.00722231f $X=4.625 $Y=0.56 $X2=0
+ $Y2=0
cc_548 N_A_560_47#_c_744_n N_VGND_c_1050_n 0.0227907f $X=3.27 $Y=0.45 $X2=0
+ $Y2=0
cc_549 N_A_560_47#_c_744_n A_657_47# 0.00297704f $X=3.27 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_550 N_A_560_47#_c_737_n A_657_47# 0.00138052f $X=3.357 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_551 N_RESET_B_M1021_g N_VPWR_c_880_n 5.76295e-19 $X=5.095 $Y=1.985 $X2=0
+ $Y2=0
cc_552 N_RESET_B_M1021_g N_VPWR_c_881_n 0.010794f $X=5.095 $Y=1.985 $X2=0 $Y2=0
cc_553 N_RESET_B_M1021_g N_VPWR_c_887_n 0.0046653f $X=5.095 $Y=1.985 $X2=0 $Y2=0
cc_554 N_RESET_B_M1021_g N_VPWR_c_875_n 0.00811867f $X=5.095 $Y=1.985 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_830_n N_VGND_c_1038_n 0.00515466f $X=5.047 $Y=0.995 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_830_n N_VGND_c_1044_n 0.00430869f $X=5.047 $Y=0.995 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_830_n N_VGND_c_1050_n 0.00615788f $X=5.047 $Y=0.995 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_875_n A_465_369# 0.00469533f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_559 N_VPWR_c_875_n A_644_413# 0.0027197f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_560 N_VPWR_c_875_n N_Q_M1009_d 0.00468958f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_561 N_VPWR_c_881_n N_Q_c_1000_n 0.0452123f $X=5.305 $Y=2.02 $X2=0 $Y2=0
cc_562 N_VPWR_M1014_s N_Q_c_990_n 0.00231287f $X=6.045 $Y=1.485 $X2=0 $Y2=0
cc_563 N_VPWR_c_883_n N_Q_c_990_n 0.022894f $X=6.18 $Y=1.835 $X2=0 $Y2=0
cc_564 N_VPWR_c_888_n Q 0.0166934f $X=6.095 $Y=2.72 $X2=0 $Y2=0
cc_565 N_VPWR_c_875_n Q 0.010102f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_566 N_Q_c_989_n N_VGND_M1008_s 0.00273341f $X=6.07 $Y=0.89 $X2=0 $Y2=0
cc_567 N_Q_c_989_n N_VGND_c_1040_n 0.0221752f $X=6.07 $Y=0.89 $X2=0 $Y2=0
cc_568 N_Q_c_996_n N_VGND_c_1045_n 0.0178243f $X=5.84 $Y=0.37 $X2=0 $Y2=0
cc_569 N_Q_M1004_d N_VGND_c_1050_n 0.00215227f $X=5.625 $Y=0.235 $X2=0 $Y2=0
cc_570 N_Q_c_996_n N_VGND_c_1050_n 0.0119575f $X=5.84 $Y=0.37 $X2=0 $Y2=0
cc_571 N_Q_c_989_n N_VGND_c_1050_n 0.00719248f $X=6.07 $Y=0.89 $X2=0 $Y2=0
cc_572 N_VGND_c_1050_n A_465_47# 0.0105287f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_573 N_VGND_c_1050_n A_657_47# 0.00841175f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_574 N_VGND_c_1050_n A_940_47# 0.00382975f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__dlrtn_4.spice
* Created: Thu Aug 27 14:17:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlrtn_4.pex.spice"
.subckt sky130_fd_sc_hd__dlrtn_4  VNB VPB GATE_N D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE_N	GATE_N
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_GATE_N_M1024_g N_A_27_47#_M1024_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_193_47#_M1013_d N_A_27_47#_M1013_g N_VGND_M1024_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_D_M1022_g N_A_300_47#_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1005 A_466_47# N_A_300_47#_M1005_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0836769 AS=0.0567 PD=0.872308 PS=0.69 NRD=41.208 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1008 N_A_562_413#_M1008_d N_A_27_47#_M1008_g A_466_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0504 AS=0.0717231 PD=0.64 PS=0.747692 NRD=0 NRS=48.072 M=1 R=2.4
+ SA=75001.1 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1019 A_660_47# N_A_193_47#_M1019_g N_A_562_413#_M1008_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0504 PD=0.687692 PS=0.64 NRD=38.076 NRS=0 M=1 R=2.4
+ SA=75001.6 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1009 N_VGND_M1009_d N_A_725_21#_M1009_g A_660_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75001.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_943_47# N_A_562_413#_M1003_g N_A_725_21#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=14.76 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_RESET_B_M1021_g A_943_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1021_d N_A_725_21#_M1007_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.099125 PD=0.98 PS=0.955 NRD=9.228 NRS=3.684 M=1 R=4.33333
+ SA=75001.1 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_A_725_21#_M1017_g N_Q_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.099125 PD=0.935 PS=0.955 NRD=1.836 NRS=0.912 M=1 R=4.33333
+ SA=75001.5 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1017_d N_A_725_21#_M1018_g N_Q_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.10075 PD=0.935 PS=0.96 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75002
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A_725_21#_M1020_g N_Q_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10075 PD=1.82 PS=0.96 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_GATE_N_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_D_M1016_g N_A_300_47#_M1016_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1012 A_466_369# N_A_300_47#_M1012_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.116891 AS=0.0864 PD=1.17132 PS=0.91 NRD=39.2818 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1025 N_A_562_413#_M1025_d N_A_193_47#_M1025_g A_466_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09555 AS=0.0767094 PD=0.875 PS=0.768679 NRD=56.2829 NRS=59.8683
+ M=1 R=2.8 SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 A_683_413# N_A_27_47#_M1004_g N_A_562_413#_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.09555 PD=0.63 PS=0.875 NRD=23.443 NRS=25.7873 M=1 R=2.8
+ SA=75001.7 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_725_21#_M1006_g A_683_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_725_21#_M1001_d N_A_562_413#_M1001_g N_VPWR_M1001_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_RESET_B_M1010_g N_A_725_21#_M1001_d VPB PHIGHVT L=0.15
+ W=1 AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75002 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1010_d N_A_725_21#_M1002_g N_Q_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.1525 PD=1.33 PS=1.305 NRD=4.9053 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A_725_21#_M1014_g N_Q_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1425 AS=0.1525 PD=1.285 PS=1.305 NRD=1.9503 NRS=2.9353 M=1 R=6.66667
+ SA=75001.5 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1014_d N_A_725_21#_M1015_g N_Q_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1425 AS=0.155 PD=1.285 PS=1.31 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75002
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_A_725_21#_M1023_g N_Q_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.155 PD=2.52 PS=1.31 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=12.4227 P=18.69
c_151 VPB 0 1.65126e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__dlrtn_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a221o_2.pxi.spice
* Created: Thu Aug 27 14:01:45 2020
* 
x_PM_SKY130_FD_SC_HD__A221O_2%C1 N_C1_c_68_n N_C1_M1012_g N_C1_M1009_g C1
+ N_C1_c_70_n PM_SKY130_FD_SC_HD__A221O_2%C1
x_PM_SKY130_FD_SC_HD__A221O_2%B2 N_B2_M1002_g N_B2_M1007_g B2 N_B2_c_96_n
+ N_B2_c_97_n N_B2_c_98_n PM_SKY130_FD_SC_HD__A221O_2%B2
x_PM_SKY130_FD_SC_HD__A221O_2%B1 N_B1_M1008_g N_B1_M1000_g B1 B1 N_B1_c_130_n
+ N_B1_c_131_n PM_SKY130_FD_SC_HD__A221O_2%B1
x_PM_SKY130_FD_SC_HD__A221O_2%A1 N_A1_M1005_g N_A1_M1011_g A1 A1 N_A1_c_174_n
+ N_A1_c_175_n PM_SKY130_FD_SC_HD__A221O_2%A1
x_PM_SKY130_FD_SC_HD__A221O_2%A2 N_A2_M1006_g N_A2_M1004_g A2 N_A2_c_213_n
+ N_A2_c_214_n N_A2_c_215_n PM_SKY130_FD_SC_HD__A221O_2%A2
x_PM_SKY130_FD_SC_HD__A221O_2%A_27_47# N_A_27_47#_M1012_s N_A_27_47#_M1008_d
+ N_A_27_47#_M1005_s N_A_27_47#_M1009_s N_A_27_47#_c_249_n N_A_27_47#_M1010_g
+ N_A_27_47#_M1001_g N_A_27_47#_c_250_n N_A_27_47#_M1013_g N_A_27_47#_M1003_g
+ N_A_27_47#_c_361_p N_A_27_47#_c_335_p N_A_27_47#_c_251_n N_A_27_47#_c_252_n
+ N_A_27_47#_c_260_n N_A_27_47#_c_261_n N_A_27_47#_c_287_n N_A_27_47#_c_253_n
+ N_A_27_47#_c_292_n N_A_27_47#_c_301_n N_A_27_47#_c_254_n N_A_27_47#_c_255_n
+ N_A_27_47#_c_256_n N_A_27_47#_c_257_n PM_SKY130_FD_SC_HD__A221O_2%A_27_47#
x_PM_SKY130_FD_SC_HD__A221O_2%A_109_297# N_A_109_297#_M1009_d
+ N_A_109_297#_M1000_d N_A_109_297#_c_386_n N_A_109_297#_c_387_n
+ N_A_109_297#_c_385_n N_A_109_297#_c_390_n
+ PM_SKY130_FD_SC_HD__A221O_2%A_109_297#
x_PM_SKY130_FD_SC_HD__A221O_2%A_193_297# N_A_193_297#_M1002_d
+ N_A_193_297#_M1011_d N_A_193_297#_c_410_n N_A_193_297#_c_416_n
+ N_A_193_297#_c_425_p N_A_193_297#_c_412_n
+ PM_SKY130_FD_SC_HD__A221O_2%A_193_297#
x_PM_SKY130_FD_SC_HD__A221O_2%VPWR N_VPWR_M1011_s N_VPWR_M1004_d N_VPWR_M1003_d
+ N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n VPWR VPWR
+ N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n
+ N_VPWR_c_433_n PM_SKY130_FD_SC_HD__A221O_2%VPWR
x_PM_SKY130_FD_SC_HD__A221O_2%X N_X_M1010_d N_X_M1001_s N_X_c_495_n N_X_c_498_n
+ N_X_c_493_n X X N_X_c_508_n PM_SKY130_FD_SC_HD__A221O_2%X
x_PM_SKY130_FD_SC_HD__A221O_2%VGND N_VGND_M1012_d N_VGND_M1006_d N_VGND_M1013_s
+ N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n VGND VGND N_VGND_c_521_n
+ N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n
+ PM_SKY130_FD_SC_HD__A221O_2%VGND
cc_1 VNB N_C1_c_68_n 0.0219801f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB C1 0.0117053f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C1_c_70_n 0.0366682f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B2_c_96_n 0.0195311f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_5 VNB N_B2_c_97_n 0.00562927f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_6 VNB N_B2_c_98_n 0.016165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB B1 0.00548362f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB B1 0.0050594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_130_n 0.0237542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_c_131_n 0.0186691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A1 0.00161887f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB A1 0.00190698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A1_c_174_n 0.0270655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_175_n 0.0207121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_213_n 0.0194f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_16 VNB N_A2_c_214_n 0.00428746f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_17 VNB N_A2_c_215_n 0.016864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_249_n 0.015967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_250_n 0.0190558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_251_n 0.00582006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_252_n 0.00183184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_253_n 0.0126554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_254_n 0.00335714f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_255_n 0.00163224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_256_n 9.16142e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_257_n 0.0497212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_433_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_493_n 6.45185e-19 $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_29 VNB N_VGND_c_517_n 0.00224165f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_30 VNB N_VGND_c_518_n 0.0126443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_31 VNB N_VGND_c_519_n 0.0109111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB VGND 0.00507731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_521_n 0.0152765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_522_n 0.0441421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_523_n 0.0173056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_524_n 0.00507731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_525_n 0.225294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_526_n 0.00280453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VPB N_C1_M1009_g 0.0255531f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_40 VPB N_C1_c_70_n 0.0092301f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_41 VPB N_B2_M1002_g 0.0187873f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_42 VPB N_B2_c_96_n 0.00419673f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_43 VPB N_B1_M1000_g 0.0255531f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_B1_c_130_n 0.00478812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A1_M1011_g 0.0251751f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_46 VPB N_A1_c_174_n 0.0056937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A2_M1004_g 0.0198907f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_48 VPB N_A2_c_213_n 0.00407683f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_49 VPB N_A_27_47#_M1001_g 0.018071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_M1003_g 0.0242689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_260_n 0.0319812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_261_n 0.00227971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_256_n 0.00132789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_257_n 0.00820462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_109_297#_c_385_n 0.00256417f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_56 VPB N_A_193_297#_c_410_n 0.00819467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_434_n 0.0059122f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_58 VPB N_VPWR_c_435_n 0.00210326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_436_n 0.0126188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_437_n 0.00833018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_438_n 0.0480882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_439_n 0.0146389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_440_n 0.015316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_441_n 0.0054066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_442_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_433_n 0.0507932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_X_c_493_n 9.41128e-19 $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_68 N_C1_M1009_g N_B2_M1002_g 0.0283323f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 C1 N_B2_c_96_n 2.15083e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_70 N_C1_c_70_n N_B2_c_96_n 0.0221625f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_71 C1 N_B2_c_97_n 0.0162885f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_72 N_C1_c_70_n N_B2_c_97_n 0.00145945f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_73 N_C1_c_68_n N_B2_c_98_n 0.0189859f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_74 N_C1_c_68_n N_A_27_47#_c_251_n 0.0141248f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_75 C1 N_A_27_47#_c_251_n 0.00669468f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_76 N_C1_c_70_n N_A_27_47#_c_251_n 0.00122978f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_77 C1 N_A_27_47#_c_252_n 0.0138529f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_78 N_C1_c_70_n N_A_27_47#_c_252_n 0.00435101f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C1_M1009_g N_A_27_47#_c_260_n 0.0137688f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_80 C1 N_A_27_47#_c_260_n 0.00669486f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_81 N_C1_c_70_n N_A_27_47#_c_260_n 0.00117267f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_82 C1 N_A_27_47#_c_261_n 0.0139066f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_83 N_C1_c_70_n N_A_27_47#_c_261_n 0.00415632f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_84 N_C1_M1009_g N_A_109_297#_c_386_n 0.00589212f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_85 N_C1_M1009_g N_A_109_297#_c_387_n 0.00211624f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_86 N_C1_M1009_g N_VPWR_c_438_n 0.00539841f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_87 N_C1_M1009_g N_VPWR_c_433_n 0.0105687f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_88 N_C1_c_68_n N_VGND_c_521_n 0.00350562f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_89 N_C1_c_68_n N_VGND_c_525_n 0.00517665f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C1_c_68_n N_VGND_c_526_n 0.00956923f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B2_M1002_g N_B1_M1000_g 0.0444451f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B2_c_96_n B1 3.76715e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B2_c_96_n B1 6.45094e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B2_c_97_n B1 0.0174856f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B2_c_96_n N_B1_c_130_n 0.038331f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B2_c_97_n N_B1_c_130_n 6.68726e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B2_c_98_n N_B1_c_131_n 0.038331f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B2_c_96_n N_A_27_47#_c_251_n 0.00321555f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B2_c_97_n N_A_27_47#_c_251_n 0.0323232f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B2_c_98_n N_A_27_47#_c_251_n 0.0120087f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B2_M1002_g N_A_27_47#_c_260_n 0.0121487f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B2_c_96_n N_A_27_47#_c_260_n 0.00308238f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B2_c_97_n N_A_27_47#_c_260_n 0.0309701f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B2_M1002_g N_A_109_297#_c_386_n 0.00692418f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_105 N_B2_M1002_g N_A_109_297#_c_387_n 7.04098e-19 $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_106 N_B2_M1002_g N_A_109_297#_c_390_n 0.00824396f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_107 N_B2_M1002_g N_VPWR_c_438_n 0.00357835f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B2_M1002_g N_VPWR_c_433_n 0.00528059f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_109 N_B2_c_98_n N_VGND_c_522_n 0.00439206f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B2_c_98_n N_VGND_c_525_n 0.00598982f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B2_c_98_n N_VGND_c_526_n 0.00313179f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_112 B1 A1 0.0232166f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_113 N_B1_c_130_n A1 2.30657e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_114 B1 A1 0.0123226f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_115 N_B1_c_130_n A1 5.90294e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_116 B1 N_A1_c_174_n 3.14731e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_117 B1 N_A1_c_174_n 8.44e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B1_c_130_n N_A1_c_174_n 0.00768957f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_119 B1 N_A1_c_175_n 0.00146136f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_120 B1 N_A_27_47#_M1008_d 0.0036585f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_121 B1 N_A_27_47#_c_251_n 0.00758188f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_122 B1 N_A_27_47#_c_251_n 0.00123465f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B1_c_131_n N_A_27_47#_c_251_n 0.00323811f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B1_M1000_g N_A_27_47#_c_260_n 0.0124878f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_125 B1 N_A_27_47#_c_260_n 0.0330891f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B1_c_130_n N_A_27_47#_c_260_n 0.00330809f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B1_c_131_n N_A_27_47#_c_287_n 0.00847781f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_128 B1 N_A_27_47#_c_253_n 0.0198101f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_129 B1 N_A_27_47#_c_253_n 0.00425548f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_130 N_B1_c_130_n N_A_27_47#_c_253_n 3.50679e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B1_c_131_n N_A_27_47#_c_253_n 0.00843864f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_c_131_n N_A_27_47#_c_292_n 0.00166393f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B1_M1000_g N_A_109_297#_c_386_n 6.99628e-19 $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_B1_M1000_g N_A_109_297#_c_385_n 0.00185095f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_B1_M1000_g N_A_109_297#_c_390_n 0.00681763f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_B1_M1000_g N_A_193_297#_c_410_n 0.0131306f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B1_M1000_g N_A_193_297#_c_412_n 0.00406201f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_B1_M1000_g N_VPWR_c_434_n 0.00237859f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_139 N_B1_M1000_g N_VPWR_c_438_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B1_M1000_g N_VPWR_c_433_n 0.00657948f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B1_c_131_n N_VGND_c_522_n 0.0035787f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_c_131_n N_VGND_c_525_n 0.00641667f $X=1.38 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_M1011_g N_A2_M1004_g 0.0229849f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_144 A1 N_A2_c_213_n 4.72548e-19 $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_145 A1 N_A2_c_213_n 2.08304e-19 $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A1_c_174_n N_A2_c_213_n 0.0214975f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_147 A1 N_A2_c_214_n 0.0158728f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A1_c_174_n N_A2_c_214_n 0.0011832f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_149 A1 N_A2_c_215_n 6.34434e-19 $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_150 N_A1_c_175_n N_A2_c_215_n 0.0294157f $X=2.162 $Y=0.995 $X2=0 $Y2=0
cc_151 A1 N_A_27_47#_M1005_s 0.00427953f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_152 N_A1_M1011_g N_A_27_47#_c_260_n 0.0136041f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_153 A1 N_A_27_47#_c_260_n 0.0242436f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A1_c_174_n N_A_27_47#_c_260_n 0.00413287f $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_155 A1 N_A_27_47#_c_253_n 0.0173818f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_156 A1 N_A_27_47#_c_253_n 0.0011516f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A1_c_174_n N_A_27_47#_c_253_n 5.61513e-19 $X=2.135 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A1_c_175_n N_A_27_47#_c_253_n 0.0110135f $X=2.162 $Y=0.995 $X2=0 $Y2=0
cc_159 A1 N_A_27_47#_c_301_n 0.0041561f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_160 N_A1_c_175_n N_A_27_47#_c_301_n 0.00428119f $X=2.162 $Y=0.995 $X2=0 $Y2=0
cc_161 A1 N_A_27_47#_c_255_n 0.0133298f $X=2.01 $Y=0.765 $X2=0 $Y2=0
cc_162 N_A1_c_175_n N_A_27_47#_c_255_n 0.00135688f $X=2.162 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_M1011_g N_A_193_297#_c_410_n 0.0141907f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A1_M1011_g N_VPWR_c_434_n 0.00990552f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A1_M1011_g N_VPWR_c_439_n 0.00273041f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A1_M1011_g N_VPWR_c_433_n 0.00348631f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A1_c_175_n N_VGND_c_517_n 0.00125396f $X=2.162 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A1_c_175_n N_VGND_c_522_n 0.00357877f $X=2.162 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_175_n N_VGND_c_525_n 0.00672549f $X=2.162 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A2_c_215_n N_A_27_47#_c_249_n 0.0202981f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A2_M1004_g N_A_27_47#_M1001_g 0.0223617f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A2_M1004_g N_A_27_47#_c_260_n 0.015518f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A2_c_213_n N_A_27_47#_c_260_n 0.0028355f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A2_c_214_n N_A_27_47#_c_260_n 0.0251115f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A2_c_213_n N_A_27_47#_c_254_n 0.00122978f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A2_c_214_n N_A_27_47#_c_254_n 0.0161642f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A2_c_215_n N_A_27_47#_c_254_n 0.0117449f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A2_c_213_n N_A_27_47#_c_255_n 0.00179152f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A2_c_214_n N_A_27_47#_c_255_n 0.0112164f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A2_M1004_g N_A_27_47#_c_256_n 0.00243411f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A2_c_213_n N_A_27_47#_c_256_n 0.0010489f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A2_c_214_n N_A_27_47#_c_256_n 0.0120858f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A2_c_215_n N_A_27_47#_c_256_n 0.00167934f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_c_213_n N_A_27_47#_c_257_n 0.0225009f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A2_c_214_n N_A_27_47#_c_257_n 0.00137404f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_M1004_g N_VPWR_c_434_n 5.43585e-19 $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A2_M1004_g N_VPWR_c_435_n 0.00166715f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A2_M1004_g N_VPWR_c_439_n 0.00585385f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A2_M1004_g N_VPWR_c_433_n 0.0107512f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A2_c_215_n N_VGND_c_517_n 0.0088683f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_c_215_n N_VGND_c_522_n 0.00350562f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_215_n N_VGND_c_525_n 0.00436f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_260_n N_A_109_297#_M1009_d 0.00165831f $X=3.065 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_194 N_A_27_47#_c_260_n N_A_109_297#_M1000_d 0.00277869f $X=3.065 $Y=1.54
+ $X2=0 $Y2=0
cc_195 N_A_27_47#_c_260_n N_A_109_297#_c_386_n 0.0170052f $X=3.065 $Y=1.54 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_260_n N_A_109_297#_c_390_n 0.0025738f $X=3.065 $Y=1.54 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_260_n N_A_193_297#_M1002_d 0.00166235f $X=3.065 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_198 N_A_27_47#_c_260_n N_A_193_297#_M1011_d 0.00229659f $X=3.065 $Y=1.54
+ $X2=0 $Y2=0
cc_199 N_A_27_47#_c_260_n N_A_193_297#_c_416_n 0.0160896f $X=3.065 $Y=1.54 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_260_n N_A_193_297#_c_412_n 0.0851707f $X=3.065 $Y=1.54 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_260_n N_VPWR_M1011_s 0.00277869f $X=3.065 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_202 N_A_27_47#_c_260_n N_VPWR_M1004_d 0.00253908f $X=3.065 $Y=1.54 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1001_g N_VPWR_c_435_n 0.0108499f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_M1003_g N_VPWR_c_435_n 4.81859e-19 $X=3.615 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_260_n N_VPWR_c_435_n 0.0140564f $X=3.065 $Y=1.54 $X2=0 $Y2=0
cc_206 N_A_27_47#_M1003_g N_VPWR_c_437_n 0.0039228f $X=3.615 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_335_p N_VPWR_c_438_n 0.0116048f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1001_g N_VPWR_c_440_n 0.0046653f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_M1003_g N_VPWR_c_440_n 0.00533769f $X=3.615 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_M1009_s N_VPWR_c_433_n 0.00525232f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_M1001_g N_VPWR_c_433_n 0.00789179f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_M1003_g N_VPWR_c_433_n 0.0103321f $X=3.615 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_335_p N_VPWR_c_433_n 0.00646998f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_249_n N_X_c_495_n 0.00167752f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_250_n N_X_c_495_n 0.00532021f $X=3.615 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_257_n N_X_c_495_n 0.00146773f $X=3.615 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_27_47#_M1003_g N_X_c_498_n 0.00143964f $X=3.615 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_257_n N_X_c_498_n 0.00144574f $X=3.615 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_249_n N_X_c_493_n 0.00299217f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_27_47#_M1001_g N_X_c_493_n 0.00526836f $X=3.195 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_250_n N_X_c_493_n 0.0063906f $X=3.615 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_27_47#_M1003_g N_X_c_493_n 0.0118648f $X=3.615 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_260_n N_X_c_493_n 0.0134012f $X=3.065 $Y=1.54 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_254_n N_X_c_493_n 0.0133881f $X=3.065 $Y=0.82 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_256_n N_X_c_493_n 0.0379666f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_257_n N_X_c_493_n 0.024289f $X=3.615 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1003_g N_X_c_508_n 0.00642666f $X=3.615 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_251_n N_VGND_M1012_d 0.00224316f $X=1.07 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_229 N_A_27_47#_c_254_n N_VGND_M1006_d 0.00208738f $X=3.065 $Y=0.82 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_249_n N_VGND_c_517_n 0.00173437f $X=3.195 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_254_n N_VGND_c_517_n 0.0178614f $X=3.065 $Y=0.82 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_250_n N_VGND_c_519_n 0.00517995f $X=3.615 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_361_p N_VGND_c_521_n 0.0115672f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_251_n N_VGND_c_521_n 0.00193763f $X=1.07 $Y=0.82 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_251_n N_VGND_c_522_n 0.00252537f $X=1.07 $Y=0.82 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_253_n N_VGND_c_522_n 0.0839447f $X=2.435 $Y=0.38 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_292_n N_VGND_c_522_n 0.00951646f $X=1.24 $Y=0.38 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_254_n N_VGND_c_522_n 0.00194318f $X=3.065 $Y=0.82 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_249_n N_VGND_c_523_n 0.00473211f $X=3.195 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_250_n N_VGND_c_523_n 0.00532251f $X=3.615 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_254_n N_VGND_c_523_n 0.00176795f $X=3.065 $Y=0.82 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1012_s N_VGND_c_525_n 0.00377256f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_M1008_d N_VGND_c_525_n 0.00209344f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1005_s N_VGND_c_525_n 0.00209344f $X=1.915 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_249_n N_VGND_c_525_n 0.00701835f $X=3.195 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_250_n N_VGND_c_525_n 0.0102951f $X=3.615 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_361_p N_VGND_c_525_n 0.0064623f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_251_n N_VGND_c_525_n 0.0102369f $X=1.07 $Y=0.82 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_253_n N_VGND_c_525_n 0.0499293f $X=2.435 $Y=0.38 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_292_n N_VGND_c_525_n 0.00651637f $X=1.24 $Y=0.38 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_254_n N_VGND_c_525_n 0.00812503f $X=3.065 $Y=0.82 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_251_n N_VGND_c_526_n 0.0190384f $X=1.07 $Y=0.82 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_292_n A_205_47# 9.37539e-19 $X=1.24 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_254 N_A_27_47#_c_253_n A_465_47# 0.00542414f $X=2.435 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_255 N_A_27_47#_c_301_n A_465_47# 0.00274948f $X=2.52 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_256 N_A_27_47#_c_255_n A_465_47# 0.00164429f $X=2.605 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_257 N_A_109_297#_c_390_n N_A_193_297#_M1002_d 0.00312752f $X=1.355 $Y=2.36
+ $X2=-0.19 $Y2=1.305
cc_258 N_A_109_297#_M1000_d N_A_193_297#_c_410_n 0.00549596f $X=1.385 $Y=1.485
+ $X2=0 $Y2=0
cc_259 N_A_109_297#_c_385_n N_A_193_297#_c_410_n 0.0157397f $X=1.52 $Y=2.34
+ $X2=0 $Y2=0
cc_260 N_A_109_297#_c_390_n N_A_193_297#_c_410_n 0.0048504f $X=1.355 $Y=2.36
+ $X2=0 $Y2=0
cc_261 N_A_109_297#_c_390_n N_A_193_297#_c_412_n 0.0118327f $X=1.355 $Y=2.36
+ $X2=0 $Y2=0
cc_262 N_A_109_297#_c_385_n N_VPWR_c_434_n 0.0169231f $X=1.52 $Y=2.34 $X2=0
+ $Y2=0
cc_263 N_A_109_297#_c_387_n N_VPWR_c_438_n 0.0189915f $X=0.845 $Y=2.38 $X2=0
+ $Y2=0
cc_264 N_A_109_297#_c_390_n N_VPWR_c_438_n 0.0481435f $X=1.355 $Y=2.36 $X2=0
+ $Y2=0
cc_265 N_A_109_297#_M1009_d N_VPWR_c_433_n 0.00215201f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_266 N_A_109_297#_M1000_d N_VPWR_c_433_n 0.00209344f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_267 N_A_109_297#_c_387_n N_VPWR_c_433_n 0.0122801f $X=0.845 $Y=2.38 $X2=0
+ $Y2=0
cc_268 N_A_109_297#_c_390_n N_VPWR_c_433_n 0.030037f $X=1.355 $Y=2.36 $X2=0
+ $Y2=0
cc_269 N_A_193_297#_c_410_n N_VPWR_M1011_s 0.00525348f $X=2.4 $Y=1.915 $X2=-0.19
+ $Y2=1.305
cc_270 N_A_193_297#_c_410_n N_VPWR_c_434_n 0.0221078f $X=2.4 $Y=1.915 $X2=0
+ $Y2=0
cc_271 N_A_193_297#_c_425_p N_VPWR_c_434_n 0.0191044f $X=2.485 $Y=2.3 $X2=0
+ $Y2=0
cc_272 N_A_193_297#_c_410_n N_VPWR_c_438_n 0.00320421f $X=2.4 $Y=1.915 $X2=0
+ $Y2=0
cc_273 N_A_193_297#_c_410_n N_VPWR_c_439_n 0.00217595f $X=2.4 $Y=1.915 $X2=0
+ $Y2=0
cc_274 N_A_193_297#_c_425_p N_VPWR_c_439_n 0.0156476f $X=2.485 $Y=2.3 $X2=0
+ $Y2=0
cc_275 N_A_193_297#_M1002_d N_VPWR_c_433_n 0.00216833f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_276 N_A_193_297#_M1011_d N_VPWR_c_433_n 0.00314787f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_277 N_A_193_297#_c_410_n N_VPWR_c_433_n 0.0120275f $X=2.4 $Y=1.915 $X2=0
+ $Y2=0
cc_278 N_A_193_297#_c_425_p N_VPWR_c_433_n 0.00954719f $X=2.485 $Y=2.3 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_433_n N_X_M1001_s 0.0038878f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_437_n N_X_c_493_n 0.0374251f $X=3.83 $Y=1.62 $X2=0 $Y2=0
cc_281 N_VPWR_c_440_n N_X_c_508_n 0.0154848f $X=3.745 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_433_n N_X_c_508_n 0.00951427f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_c_437_n N_VGND_c_519_n 0.00781039f $X=3.83 $Y=1.62 $X2=0 $Y2=0
cc_284 N_X_c_493_n N_VGND_c_519_n 0.0141782f $X=3.447 $Y=1.795 $X2=0 $Y2=0
cc_285 N_X_c_495_n N_VGND_c_523_n 0.0153335f $X=3.49 $Y=0.665 $X2=0 $Y2=0
cc_286 N_X_M1010_d N_VGND_c_525_n 0.00385308f $X=3.27 $Y=0.235 $X2=0 $Y2=0
cc_287 N_X_c_495_n N_VGND_c_525_n 0.00953265f $X=3.49 $Y=0.665 $X2=0 $Y2=0
cc_288 N_VGND_c_525_n A_205_47# 0.0019167f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_289 N_VGND_c_525_n A_465_47# 0.002906f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a2bb2oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.310000 1.075000 4.205000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.455000 1.075000 5.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.710000 1.445000 ;
        RECT 0.085000 1.445000 2.030000 1.615000 ;
        RECT 1.700000 1.075000 2.030000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.075000 1.480000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 0.645000 1.400000 0.725000 ;
        RECT 1.070000 0.725000 2.660000 0.905000 ;
        RECT 2.330000 0.255000 2.660000 0.725000 ;
        RECT 2.370000 0.905000 2.660000 1.660000 ;
        RECT 2.370000 1.660000 2.620000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 0.310000  0.085000 0.480000 0.895000 ;
        RECT 1.990000  0.085000 2.160000 0.555000 ;
        RECT 2.830000  0.085000 3.520000 0.555000 ;
        RECT 4.190000  0.085000 4.360000 0.555000 ;
        RECT 5.030000  0.085000 5.200000 0.905000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.690000 2.135000 0.940000 2.635000 ;
        RECT 1.530000 2.135000 1.780000 2.635000 ;
        RECT 3.730000 2.135000 3.980000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.270000 1.785000 2.200000 1.955000 ;
      RECT 0.270000 1.955000 0.520000 2.465000 ;
      RECT 0.650000 0.255000 1.820000 0.475000 ;
      RECT 0.650000 0.475000 0.900000 0.895000 ;
      RECT 1.110000 1.955000 1.360000 2.465000 ;
      RECT 1.950000 1.955000 2.200000 2.295000 ;
      RECT 1.950000 2.295000 3.040000 2.465000 ;
      RECT 2.790000 1.795000 3.040000 2.295000 ;
      RECT 2.830000 0.995000 3.120000 1.325000 ;
      RECT 2.950000 0.725000 4.860000 0.905000 ;
      RECT 2.950000 0.905000 3.120000 0.995000 ;
      RECT 2.950000 1.325000 3.120000 1.445000 ;
      RECT 2.950000 1.445000 4.820000 1.615000 ;
      RECT 3.310000 1.785000 4.400000 1.965000 ;
      RECT 3.310000 1.965000 3.560000 2.465000 ;
      RECT 3.690000 0.255000 4.020000 0.725000 ;
      RECT 4.150000 1.965000 4.400000 2.295000 ;
      RECT 4.150000 2.295000 5.240000 2.465000 ;
      RECT 4.530000 0.255000 4.860000 0.725000 ;
      RECT 4.570000 1.615000 4.820000 2.125000 ;
      RECT 4.990000 1.455000 5.240000 2.295000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_2

* File: sky130_fd_sc_hd__and4bb_1.spice
* Created: Tue Sep  1 18:58:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and4bb_1.pex.spice"
.subckt sky130_fd_sc_hd__and4bb_1  VNB VPB A_N B_N C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_N_M1007_g N_A_27_47#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.168 PD=0.7 PS=1.64 NRD=0 NRS=38.568 M=1 R=2.8 SA=75000.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_223_47#_M1009_d N_B_N_M1009_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1386 AS=0.0588 PD=1.5 PS=0.7 NRD=18.564 NRS=1.428 M=1 R=2.8 SA=75000.8
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 A_429_93# N_A_27_47#_M1011_g N_A_343_93#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=24.276 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1001 A_515_93# N_A_223_47#_M1001_g A_429_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=34.284 NRS=24.276 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 A_615_93# N_C_M1000_g A_515_93# VNB NSHORT L=0.15 W=0.42 AD=0.0777
+ AS=0.0735 PD=0.79 PS=0.77 NRD=37.14 NRS=34.284 M=1 R=2.8 SA=75001.1 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_D_M1010_g A_615_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.0993084 AS=0.0777 PD=0.871402 PS=0.79 NRD=51.84 NRS=37.14 M=1 R=2.8
+ SA=75001.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_343_93#_M1005_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1654 AS=0.153692 PD=1.82 PS=1.3486 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_N_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.168 PD=0.7 PS=1.64 NRD=0 NRS=63.3158 M=1 R=2.8 SA=75000.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_A_223_47#_M1012_d N_B_N_M1012_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1344 AS=0.0588 PD=1.48 PS=0.7 NRD=25.7873 NRS=2.3443 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_343_93#_M1008_d N_A_27_47#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1218 PD=0.7 PS=1.42 NRD=2.3443 NRS=11.7215 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_223_47#_M1002_g N_A_343_93#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_343_93#_M1004_d N_C_M1004_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0777 AS=0.0735 PD=0.79 PS=0.77 NRD=14.0658 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_D_M1003_g N_A_343_93#_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.101746 AS=0.0777 PD=0.863662 PS=0.79 NRD=86.7588 NRS=28.1316 M=1 R=2.8
+ SA=75001.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_X_M1013_d N_A_343_93#_M1013_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.242254 PD=2.52 PS=2.05634 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__and4bb_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nor2_1.pex.spice
* Created: Tue Sep  1 19:17:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR2_1%B 1 3 6 8 14
c26 8 0 1.17796e-19 $X=0.23 $Y=1.19
r27 11 14 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.27 $Y=1.16 $X2=0.47
+ $Y2=1.16
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r29 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r31 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_1%A 3 5 7 8 11
c28 11 0 1.17796e-19 $X=0.89 $Y=1.16
r29 11 13 34.3172 $w=3.09e-07 $l=2.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.11 $Y2=1.16
r30 10 11 9.35922 $w=3.09e-07 $l=6e-08 $layer=POLY_cond $X=0.83 $Y=1.16 $X2=0.89
+ $Y2=1.16
r31 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.16 $X2=1.11 $Y2=1.16
r32 5 11 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r33 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
r34 1 10 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.83 $Y=1.325
+ $X2=0.83 $Y2=1.16
r35 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.83 $Y=1.325 $X2=0.83
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_1%Y 1 2 7 11 14 15 18 19
c33 14 0 9.89984e-20 $X=0.69 $Y=1.495
r34 19 24 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.21
+ $X2=0.26 $Y2=2.34
r35 15 19 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.21
r36 15 17 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.665 $X2=0.26
+ $Y2=1.58
r37 14 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.69 $Y=1.495 $X2=0.69
+ $Y2=0.895
r38 9 18 7.20219 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.73
+ $X2=0.68 $Y2=0.895
r39 9 11 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.73 $X2=0.68
+ $Y2=0.39
r40 8 17 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=1.58
+ $X2=0.26 $Y2=1.58
r41 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=1.58
+ $X2=0.69 $Y2=1.495
r42 7 8 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.605 $Y=1.58
+ $X2=0.425 $Y2=1.58
r43 2 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r44 2 17 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r45 1 11 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_1%VPWR 1 4 6 10 12 19 21
r16 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r17 15 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r18 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r19 12 18 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=1.167 $Y2=2.72
r20 12 14 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=0.69 $Y2=2.72
r21 10 15 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r22 10 21 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r23 6 9 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=1.66 $X2=1.12
+ $Y2=2.34
r24 4 18 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.167 $Y2=2.72
r25 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.34
r26 1 9 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.485 $X2=1.04 $Y2=2.34
r27 1 6 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.485 $X2=1.04 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_1%VGND 1 2 7 9 11 13 15 17 27
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r22 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r23 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r24 18 23 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r25 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r26 17 26 4.22234 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.197
+ $Y2=0
r27 17 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.69
+ $Y2=0
r28 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r29 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r30 11 26 3.06235 $w=2.7e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.197 $Y2=0
r31 11 13 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.39
r32 7 23 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r33 7 9 14.6456 $w=2.38e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.39
r34 2 13 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r35 1 9 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends


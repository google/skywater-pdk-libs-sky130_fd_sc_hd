* File: sky130_fd_sc_hd__nor3_1.pex.spice
* Created: Thu Aug 27 14:31:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR3_1%C 1 3 6 8 14
r27 11 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r29 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r31 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_1%B 1 3 6 12 13 15 16
c39 15 0 5.10403e-20 $X=0.695 $Y=1.53
r40 15 16 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.712 $Y=1.53
+ $X2=0.712 $Y2=1.87
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r42 9 15 10.0532 $w=2.33e-07 $l=2.05e-07 $layer=LI1_cond $X=0.712 $Y=1.325
+ $X2=0.712 $Y2=1.53
r43 8 12 6.21621 $w=3.28e-07 $l=1.78e-07 $layer=LI1_cond $X=0.712 $Y=1.16
+ $X2=0.89 $Y2=1.16
r44 8 9 2.74472 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=1.16
+ $X2=0.712 $Y2=1.325
r45 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r46 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r47 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_1%A 1 3 6 8 9 10 17
c36 8 0 5.10403e-20 $X=1.615 $Y=0.85
r37 14 17 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.57 $Y2=1.16
r38 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.62 $Y=1.16 $X2=1.62
+ $Y2=1.53
r39 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.16 $X2=1.57 $Y2=1.16
r40 8 9 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.62 $Y=0.85 $X2=1.62
+ $Y2=1.16
r41 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r42 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r43 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_1%Y 1 2 3 10 12 15 16 17 19 25 30 33 35 39
r58 33 39 2.40809 $w=3.33e-07 $l=7e-08 $layer=LI1_cond $X=0.257 $Y=2.28
+ $X2=0.257 $Y2=2.21
r59 30 33 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=2.365
+ $X2=0.257 $Y2=2.28
r60 30 39 0.27521 $w=3.33e-07 $l=8e-09 $layer=LI1_cond $X=0.257 $Y=2.202
+ $X2=0.257 $Y2=2.21
r61 30 35 18.6455 $w=3.33e-07 $l=5.42e-07 $layer=LI1_cond $X=0.257 $Y=2.202
+ $X2=0.257 $Y2=1.66
r62 28 29 10.5364 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.165 $Y=0.55
+ $X2=1.165 $Y2=0.74
r63 23 25 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.085 $Y=1.58
+ $X2=1.23 $Y2=1.58
r64 19 21 8.58683 $w=2.53e-07 $l=1.9e-07 $layer=LI1_cond $X=0.217 $Y=0.55
+ $X2=0.217 $Y2=0.74
r65 17 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=1.495
+ $X2=1.23 $Y2=1.58
r66 16 29 5.37557 $w=2.2e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.23 $Y=0.825
+ $X2=1.165 $Y2=0.74
r67 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.23 $Y=0.825
+ $X2=1.23 $Y2=1.495
r68 14 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=1.665
+ $X2=1.085 $Y2=1.58
r69 14 15 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.085 $Y=1.665
+ $X2=1.085 $Y2=2.28
r70 13 30 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=2.365
+ $X2=0.257 $Y2=2.365
r71 12 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1 $Y=2.365
+ $X2=1.085 $Y2=2.28
r72 12 13 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1 $Y=2.365
+ $X2=0.425 $Y2=2.365
r73 11 21 3.11056 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.217 $Y2=0.74
r74 10 29 2.2496 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.015 $Y=0.74
+ $X2=1.165 $Y2=0.74
r75 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.74
+ $X2=0.345 $Y2=0.74
r76 3 30 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r77 3 35 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r78 2 28 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.55
r79 1 19 182 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_1%VPWR 1 4 6 8 10 20
r22 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r23 17 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r24 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 12 16 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r26 10 19 4.64874 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.637 $Y2=2.72
r27 10 16 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r28 8 17 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 8 12 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r30 4 19 2.99176 $w=3.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.592 $Y=2.635
+ $X2=1.637 $Y2=2.72
r31 4 6 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=1.592 $Y=2.635
+ $X2=1.592 $Y2=2
r32 1 6 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_1%VGND 1 2 9 11 13 15 17 22 28 32
r34 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r35 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r36 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r37 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r38 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r39 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r40 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r41 22 31 4.65202 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.597
+ $Y2=0
r42 22 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.15
+ $Y2=0
r43 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r44 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r45 15 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r46 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r47 11 31 3.11416 $w=3.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.597 $Y2=0
r48 11 13 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.39
r49 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r50 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.39
r51 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r52 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__or4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 0.995000 2.010000 1.445000 ;
        RECT 1.840000 1.445000 2.275000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.280000 0.995000 1.610000 1.450000 ;
        RECT 1.400000 1.450000 1.610000 1.785000 ;
        RECT 1.400000 1.785000 1.720000 2.375000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.880000 0.995000 1.050000 1.620000 ;
        RECT 0.880000 1.620000 1.230000 2.375000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.370000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 1.455000 4.055000 1.625000 ;
        RECT 2.480000 1.625000 2.730000 2.465000 ;
        RECT 2.520000 0.255000 2.770000 0.725000 ;
        RECT 2.520000 0.725000 4.055000 0.905000 ;
        RECT 3.280000 0.255000 3.610000 0.725000 ;
        RECT 3.320000 1.625000 3.570000 2.465000 ;
        RECT 3.810000 0.905000 4.055000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.115000  1.495000 0.710000 1.665000 ;
      RECT 0.115000  1.665000 0.450000 2.450000 ;
      RECT 0.120000  0.085000 0.370000 0.585000 ;
      RECT 0.540000  0.655000 2.350000 0.825000 ;
      RECT 0.540000  0.825000 0.710000 1.495000 ;
      RECT 0.700000  0.305000 0.870000 0.655000 ;
      RECT 1.070000  0.085000 1.400000 0.485000 ;
      RECT 1.570000  0.305000 1.740000 0.655000 ;
      RECT 1.960000  0.085000 2.340000 0.485000 ;
      RECT 2.005000  1.795000 2.255000 2.635000 ;
      RECT 2.180000  0.825000 2.350000 1.075000 ;
      RECT 2.180000  1.075000 3.640000 1.245000 ;
      RECT 2.900000  1.795000 3.150000 2.635000 ;
      RECT 2.940000  0.085000 3.110000 0.555000 ;
      RECT 3.740000  1.795000 3.990000 2.635000 ;
      RECT 3.780000  0.085000 3.950000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or4_4
END LIBRARY

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 1.005000 2.160000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615000 0.255000 11.875000 0.825000 ;
        RECT 11.615000 1.445000 11.875000 2.465000 ;
        RECT 11.660000 0.825000 11.875000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.200000 0.255000 10.485000 0.715000 ;
        RECT 10.200000 1.630000 10.485000 2.465000 ;
        RECT 10.280000 0.715000 10.485000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315000 1.095000 9.690000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.590000 0.735000 4.000000 0.965000 ;
        RECT 3.590000 0.965000 3.920000 1.065000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.460000 0.735000 7.835000 1.065000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.770000 0.735000 4.060000 0.780000 ;
        RECT 3.770000 0.780000 7.740000 0.920000 ;
        RECT 3.770000 0.920000 4.060000 0.965000 ;
        RECT 7.450000 0.735000 7.740000 0.780000 ;
        RECT 7.450000 0.920000 7.740000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.960000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  1.435000  0.085000  1.785000 0.465000 ;
        RECT  3.570000  0.085000  3.740000 0.525000 ;
        RECT  5.350000  0.085000  5.680000 0.465000 ;
        RECT  7.265000  0.085000  7.525000 0.525000 ;
        RECT  9.700000  0.085000 10.030000 0.805000 ;
        RECT 11.150000  0.085000 11.445000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.960000 2.805000 ;
        RECT  0.515000 2.135000  0.845000 2.635000 ;
        RECT  1.435000 2.135000  1.785000 2.635000 ;
        RECT  3.410000 2.205000  3.790000 2.635000 ;
        RECT  4.880000 1.915000  5.210000 2.635000 ;
        RECT  7.325000 2.255000  7.705000 2.635000 ;
        RECT  8.645000 2.255000 10.030000 2.635000 ;
        RECT 11.150000 1.765000 11.445000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.345000  0.345000 0.635000 ;
      RECT  0.085000 0.635000  0.840000 0.805000 ;
      RECT  0.085000 1.795000  0.840000 1.965000 ;
      RECT  0.085000 1.965000  0.345000 2.465000 ;
      RECT  0.610000 0.805000  0.840000 1.795000 ;
      RECT  1.015000 0.345000  1.240000 2.465000 ;
      RECT  1.410000 0.635000  2.125000 0.825000 ;
      RECT  1.410000 0.825000  1.580000 1.795000 ;
      RECT  1.410000 1.795000  2.125000 1.965000 ;
      RECT  1.955000 0.305000  2.125000 0.635000 ;
      RECT  1.955000 1.965000  2.125000 2.465000 ;
      RECT  2.330000 0.705000  2.550000 1.575000 ;
      RECT  2.330000 1.575000  2.830000 1.955000 ;
      RECT  2.340000 2.250000  3.170000 2.420000 ;
      RECT  2.405000 0.265000  3.400000 0.465000 ;
      RECT  2.730000 0.645000  3.060000 1.015000 ;
      RECT  3.000000 1.195000  3.400000 1.235000 ;
      RECT  3.000000 1.235000  4.350000 1.405000 ;
      RECT  3.000000 1.405000  3.170000 2.250000 ;
      RECT  3.230000 0.465000  3.400000 1.195000 ;
      RECT  3.340000 1.575000  3.590000 1.785000 ;
      RECT  3.340000 1.785000  4.690000 2.035000 ;
      RECT  3.910000 0.255000  5.080000 0.425000 ;
      RECT  3.910000 0.425000  4.240000 0.545000 ;
      RECT  4.090000 2.035000  4.260000 2.375000 ;
      RECT  4.100000 1.405000  4.350000 1.485000 ;
      RECT  4.130000 1.155000  4.350000 1.235000 ;
      RECT  4.410000 0.595000  4.740000 0.765000 ;
      RECT  4.520000 0.765000  4.740000 0.895000 ;
      RECT  4.520000 0.895000  5.830000 1.065000 ;
      RECT  4.520000 1.065000  4.690000 1.785000 ;
      RECT  4.860000 1.235000  5.190000 1.415000 ;
      RECT  4.860000 1.415000  5.865000 1.655000 ;
      RECT  4.910000 0.425000  5.080000 0.715000 ;
      RECT  5.500000 1.065000  5.830000 1.235000 ;
      RECT  6.065000 1.575000  6.300000 1.985000 ;
      RECT  6.125000 0.705000  6.410000 1.125000 ;
      RECT  6.125000 1.125000  6.745000 1.305000 ;
      RECT  6.255000 2.250000  7.085000 2.420000 ;
      RECT  6.320000 0.265000  7.085000 0.465000 ;
      RECT  6.540000 1.305000  6.745000 1.905000 ;
      RECT  6.915000 0.465000  7.085000 1.235000 ;
      RECT  6.915000 1.235000  8.265000 1.405000 ;
      RECT  6.915000 1.405000  7.085000 2.250000 ;
      RECT  7.255000 1.575000  7.505000 1.915000 ;
      RECT  7.255000 1.915000 10.030000 2.085000 ;
      RECT  7.785000 0.255000  8.955000 0.425000 ;
      RECT  7.785000 0.425000  8.115000 0.545000 ;
      RECT  7.945000 2.085000  8.115000 2.375000 ;
      RECT  8.045000 1.075000  8.265000 1.235000 ;
      RECT  8.285000 0.595000  8.615000 0.780000 ;
      RECT  8.435000 0.780000  8.615000 1.915000 ;
      RECT  8.785000 0.425000  8.955000 0.585000 ;
      RECT  8.785000 0.755000  9.475000 0.925000 ;
      RECT  8.785000 0.925000  9.060000 1.575000 ;
      RECT  8.785000 1.575000  9.545000 1.745000 ;
      RECT  9.240000 0.265000  9.475000 0.755000 ;
      RECT  9.860000 0.995000 10.110000 1.325000 ;
      RECT  9.860000 1.325000 10.030000 1.915000 ;
      RECT 10.655000 0.255000 10.970000 0.995000 ;
      RECT 10.655000 0.995000 11.490000 1.325000 ;
      RECT 10.655000 1.325000 10.970000 2.415000 ;
    LAYER mcon ;
      RECT 0.610000 1.785000 0.780000 1.955000 ;
      RECT 1.070000 0.765000 1.240000 0.935000 ;
      RECT 2.450000 1.785000 2.620000 1.955000 ;
      RECT 2.890000 0.765000 3.060000 0.935000 ;
      RECT 5.670000 1.445000 5.840000 1.615000 ;
      RECT 6.130000 1.105000 6.300000 1.275000 ;
      RECT 6.130000 1.785000 6.300000 1.955000 ;
      RECT 8.890000 1.445000 9.060000 1.615000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 6.360000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 3.120000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.390000 1.755000 2.680000 1.800000 ;
      RECT 2.390000 1.940000 2.680000 1.985000 ;
      RECT 2.830000 0.735000 3.120000 0.780000 ;
      RECT 2.830000 0.920000 3.120000 0.965000 ;
      RECT 2.925000 0.965000 3.120000 1.120000 ;
      RECT 2.925000 1.120000 6.360000 1.260000 ;
      RECT 5.610000 1.415000 5.900000 1.460000 ;
      RECT 5.610000 1.460000 9.120000 1.600000 ;
      RECT 5.610000 1.600000 5.900000 1.645000 ;
      RECT 6.070000 1.075000 6.360000 1.120000 ;
      RECT 6.070000 1.260000 6.360000 1.305000 ;
      RECT 6.070000 1.755000 6.360000 1.800000 ;
      RECT 6.070000 1.940000 6.360000 1.985000 ;
      RECT 8.830000 1.415000 9.120000 1.460000 ;
      RECT 8.830000 1.600000 9.120000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbp_1
END LIBRARY

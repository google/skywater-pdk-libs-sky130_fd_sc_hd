* File: sky130_fd_sc_hd__clkdlybuf4s25_1.pex.spice
* Created: Tue Sep  1 19:00:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A 3 7 9 15
c33 9 0 2.11583e-19 $X=0.235 $Y=1.19
r34 12 15 33.0962 $w=2.9e-07 $l=1.6e-07 $layer=POLY_cond $X=0.32 $Y=1.16
+ $X2=0.48 $Y2=1.16
r35 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.16 $X2=0.32 $Y2=1.16
r36 5 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.48 $Y=1.305
+ $X2=0.48 $Y2=1.16
r37 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.48 $Y=1.305 $X2=0.48
+ $Y2=1.985
r38 1 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.48 $Y=1.015
+ $X2=0.48 $Y2=1.16
r39 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.48 $Y=1.015 $X2=0.48
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_27_47# 1 2 9 13 17 21 23 24 25 26
+ 27 28 35
c69 35 0 1.94337e-19 $X=1.095 $Y=1.16
c70 28 0 5.32225e-20 $X=0.83 $Y=1.49
c71 27 0 1.68905e-19 $X=0.83 $Y=1.295
c72 13 0 1.72457e-20 $X=1.095 $Y=2.075
r73 32 35 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=1.095 $Y2=1.16
r74 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r75 29 31 10.4221 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.88 $Y=0.82
+ $X2=0.88 $Y2=1.16
r76 27 31 4.34663 $w=3.98e-07 $l=1.58035e-07 $layer=LI1_cond $X=0.83 $Y=1.295
+ $X2=0.88 $Y2=1.16
r77 27 28 6.42075 $w=3.48e-07 $l=1.95e-07 $layer=LI1_cond $X=0.83 $Y=1.295
+ $X2=0.83 $Y2=1.49
r78 25 28 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.655 $Y=1.575
+ $X2=0.83 $Y2=1.49
r79 25 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.655 $Y=1.575
+ $X2=0.43 $Y2=1.575
r80 23 29 5.74796 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.655 $Y=0.82
+ $X2=0.88 $Y2=0.82
r81 23 24 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.655 $Y=0.82
+ $X2=0.41 $Y2=0.82
r82 19 26 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.257 $Y=1.66
+ $X2=0.43 $Y2=1.575
r83 19 21 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=1.66
+ $X2=0.257 $Y2=1.995
r84 15 24 7.72402 $w=1.7e-07 $l=2.01057e-07 $layer=LI1_cond $X=0.247 $Y=0.735
+ $X2=0.41 $Y2=0.82
r85 15 17 11.1698 $w=3.23e-07 $l=3.15e-07 $layer=LI1_cond $X=0.247 $Y=0.735
+ $X2=0.247 $Y2=0.42
r86 11 35 4.66776 $w=2.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=1.16
r87 11 13 193.794 $w=2.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=2.075
r88 7 35 4.66776 $w=2.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.095 $Y=1.025
+ $X2=1.095 $Y2=1.16
r89 7 9 115.531 $w=2.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.095 $Y=1.025
+ $X2=1.095 $Y2=0.56
r90 2 21 300 $w=1.7e-07 $l=5.71314e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.265 $Y2=1.995
r91 1 17 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_244_47# 1 2 11 15 18 23 24 27 31
+ 32 34
c66 24 0 1.68905e-19 $X=2.255 $Y=1.16
c67 23 0 1.65571e-19 $X=2.255 $Y=1.16
r68 31 32 10.0889 $w=4.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.42 $Y=1.995
+ $X2=1.42 $Y2=1.79
r69 27 29 16.5173 $w=4.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.41 $Y=0.4
+ $X2=1.41 $Y2=0.855
r70 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.255
+ $Y=1.16 $X2=2.255 $Y2=1.16
r71 21 34 1.34256 $w=1.75e-07 $l=8.8e-08 $layer=LI1_cond $X=1.645 $Y=1.162
+ $X2=1.557 $Y2=1.162
r72 21 23 38.6597 $w=1.73e-07 $l=6.1e-07 $layer=LI1_cond $X=1.645 $Y=1.162
+ $X2=2.255 $Y2=1.162
r73 19 34 5.16603 $w=1.75e-07 $l=8.8e-08 $layer=LI1_cond $X=1.557 $Y=1.25
+ $X2=1.557 $Y2=1.162
r74 19 32 34.2234 $w=1.73e-07 $l=5.4e-07 $layer=LI1_cond $X=1.557 $Y=1.25
+ $X2=1.557 $Y2=1.79
r75 18 34 5.16603 $w=1.75e-07 $l=8.7e-08 $layer=LI1_cond $X=1.557 $Y=1.075
+ $X2=1.557 $Y2=1.162
r76 18 29 13.9429 $w=1.73e-07 $l=2.2e-07 $layer=LI1_cond $X=1.557 $Y=1.075
+ $X2=1.557 $Y2=0.855
r77 13 24 21.7495 $w=2.5e-07 $l=1.64317e-07 $layer=POLY_cond $X=2.165 $Y=1.295
+ $X2=2.23 $Y2=1.16
r78 13 15 193.794 $w=2.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.165 $Y=1.295
+ $X2=2.165 $Y2=2.075
r79 9 24 21.7495 $w=2.5e-07 $l=1.64317e-07 $layer=POLY_cond $X=2.165 $Y=1.025
+ $X2=2.23 $Y2=1.16
r80 9 11 115.531 $w=2.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.165 $Y=1.025
+ $X2=2.165 $Y2=0.56
r81 2 31 300 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.665 $X2=1.36 $Y2=1.995
r82 1 27 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.22
+ $Y=0.235 $X2=1.36 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_355_47# 1 2 9 13 17 21 23 24 25 26
+ 27 28 32
c79 32 0 1.65571e-19 $X=2.915 $Y=1.16
c80 28 0 1.13255e-19 $X=2.68 $Y=1.495
r81 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.16
+ $X2=2.915 $Y2=1.325
r82 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.16
+ $X2=2.915 $Y2=0.995
r83 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.16 $X2=2.915 $Y2=1.16
r84 27 31 8.95891 $w=3.31e-07 $l=2.25067e-07 $layer=LI1_cond $X=2.68 $Y=1.325
+ $X2=2.822 $Y2=1.16
r85 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.68 $Y=1.325
+ $X2=2.68 $Y2=1.495
r86 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.595 $Y=1.58
+ $X2=2.68 $Y2=1.495
r87 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.595 $Y=1.58
+ $X2=2.065 $Y2=1.58
r88 23 31 12.5317 $w=3.31e-07 $l=4.39067e-07 $layer=LI1_cond $X=2.595 $Y=0.82
+ $X2=2.822 $Y2=1.16
r89 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.595 $Y=0.82
+ $X2=2.065 $Y2=0.82
r90 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.94 $Y=1.665
+ $X2=2.065 $Y2=1.58
r91 19 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=1.665
+ $X2=1.94 $Y2=1.96
r92 15 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=2.065 $Y2=0.82
r93 15 17 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.42
r94 13 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.975 $Y=1.985
+ $X2=2.975 $Y2=1.325
r95 9 34 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.975 $Y=0.445
+ $X2=2.975 $Y2=0.995
r96 2 21 300 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=2 $X=1.775
+ $Y=1.665 $X2=1.9 $Y2=1.96
r97 1 17 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.235 $X2=1.9 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%VPWR 1 2 9 13 15 17 22 32 33 36 39
c41 2 0 1.13255e-19 $X=2.29 $Y=1.665
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 33 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 30 39 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.54 $Y2=2.72
r47 30 32 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=3.45 $Y2=2.72
r48 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 25 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 23 36 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.762 $Y2=2.72
r55 23 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 22 39 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.54 $Y2=2.72
r57 22 28 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 17 36 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.762
+ $Y2=2.72
r59 17 19 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r60 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r62 11 39 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=2.635
+ $X2=2.54 $Y2=2.72
r63 11 13 12.549 $w=6.08e-07 $l=6.4e-07 $layer=LI1_cond $X=2.54 $Y=2.635
+ $X2=2.54 $Y2=1.995
r64 7 36 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.762 $Y=2.635
+ $X2=0.762 $Y2=2.72
r65 7 9 22.6943 $w=3.23e-07 $l=6.4e-07 $layer=LI1_cond $X=0.762 $Y=2.635
+ $X2=0.762 $Y2=1.995
r66 2 13 300 $w=1.7e-07 $l=5.29906e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.665 $X2=2.68 $Y2=1.995
r67 1 9 300 $w=1.7e-07 $l=6.03863e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.76 $Y2=1.995
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%X 1 2 7 8 9 10 11 12 29 32
r22 40 42 6.64526 $w=3.83e-07 $l=2.22e-07 $layer=LI1_cond $X=3.19 $Y=0.447
+ $X2=3.412 $Y2=0.447
r23 30 32 0.533964 $w=5.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.315 $Y=1.845
+ $X2=3.315 $Y2=1.87
r24 29 47 1.10508 $w=3.63e-07 $l=3.5e-08 $layer=LI1_cond $X=3.412 $Y=1.53
+ $X2=3.412 $Y2=1.565
r25 21 42 1.05553 $w=3.65e-07 $l=1.93e-07 $layer=LI1_cond $X=3.412 $Y=0.64
+ $X2=3.412 $Y2=0.447
r26 12 35 5.33964 $w=5.58e-07 $l=2.5e-07 $layer=LI1_cond $X=3.315 $Y=2.21
+ $X2=3.315 $Y2=1.96
r27 11 30 0.640756 $w=5.58e-07 $l=3e-08 $layer=LI1_cond $X=3.315 $Y=1.815
+ $X2=3.315 $Y2=1.845
r28 11 35 1.28151 $w=5.58e-07 $l=6e-08 $layer=LI1_cond $X=3.315 $Y=1.9 $X2=3.315
+ $Y2=1.96
r29 11 32 0.640756 $w=5.58e-07 $l=3e-08 $layer=LI1_cond $X=3.315 $Y=1.9
+ $X2=3.315 $Y2=1.87
r30 10 11 4.80567 $w=5.58e-07 $l=2.25e-07 $layer=LI1_cond $X=3.315 $Y=1.59
+ $X2=3.315 $Y2=1.815
r31 10 47 1.98274 $w=5.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.315 $Y=1.59
+ $X2=3.315 $Y2=1.565
r32 10 29 0.789345 $w=3.63e-07 $l=2.5e-08 $layer=LI1_cond $X=3.412 $Y=1.505
+ $X2=3.412 $Y2=1.53
r33 9 10 9.94574 $w=3.63e-07 $l=3.15e-07 $layer=LI1_cond $X=3.412 $Y=1.19
+ $X2=3.412 $Y2=1.505
r34 8 9 10.7351 $w=3.63e-07 $l=3.4e-07 $layer=LI1_cond $X=3.412 $Y=0.85
+ $X2=3.412 $Y2=1.19
r35 8 21 6.63049 $w=3.63e-07 $l=2.1e-07 $layer=LI1_cond $X=3.412 $Y=0.85
+ $X2=3.412 $Y2=0.64
r36 7 42 0.987808 $w=3.83e-07 $l=3.3e-08 $layer=LI1_cond $X=3.445 $Y=0.447
+ $X2=3.412 $Y2=0.447
r37 2 35 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=3.05
+ $Y=1.485 $X2=3.19 $Y2=1.96
r38 1 40 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.05
+ $Y=0.235 $X2=3.19 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%VGND 1 2 9 11 13 28 29 32 37 40
r49 39 40 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=0.24
+ $X2=2.845 $Y2=0.24
r50 35 39 2.76018 $w=6.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=0.24
+ $X2=2.68 $Y2=0.24
r51 35 37 12.7821 $w=6.48e-07 $l=2.9e-07 $layer=LI1_cond $X=2.53 $Y=0.24
+ $X2=2.24 $Y2=0.24
r52 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r53 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r54 29 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r55 28 40 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.845
+ $Y2=0
r56 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r57 25 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r58 24 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.24
+ $Y2=0
r59 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r60 22 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r61 22 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r62 21 24 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r63 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r64 19 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.745
+ $Y2=0
r65 19 21 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.15
+ $Y2=0
r66 13 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.745
+ $Y2=0
r67 13 15 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.23
+ $Y2=0
r68 11 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 7 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r71 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.4
r72 2 39 182 $w=1.7e-07 $l=4.65242e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.235 $X2=2.68 $Y2=0.4
r73 1 9 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.745 $Y2=0.4
.ends


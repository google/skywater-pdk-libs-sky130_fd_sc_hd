* File: sky130_fd_sc_hd__mux2_4.pex.spice
* Created: Tue Sep  1 19:14:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX2_4%S 3 6 10 12 15 18 19 20 22 25 27 29 30 33 36
+ 37
r97 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.31
+ $Y=1.16 $X2=3.31 $Y2=1.16
r98 30 37 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.985 $Y=1.16
+ $X2=3.31 $Y2=1.16
r99 29 30 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.85 $Y=1.16
+ $X2=2.985 $Y2=1.16
r100 25 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r101 25 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r102 24 27 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.515 $Y=1.16
+ $X2=0.655 $Y2=1.16
r103 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r104 22 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.765 $Y=0.995
+ $X2=2.85 $Y2=1.16
r105 21 22 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.765 $Y=0.805
+ $X2=2.765 $Y2=0.995
r106 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.68 $Y=0.72
+ $X2=2.765 $Y2=0.805
r107 19 20 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=2.68 $Y=0.72
+ $X2=0.74 $Y2=0.72
r108 18 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.655 $Y=0.995
+ $X2=0.655 $Y2=1.16
r109 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.655 $Y=0.805
+ $X2=0.74 $Y2=0.72
r110 17 18 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.655 $Y=0.805
+ $X2=0.655 $Y2=0.995
r111 13 36 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.37 $Y=1.325
+ $X2=3.37 $Y2=1.16
r112 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.37 $Y=1.325
+ $X2=3.37 $Y2=1.985
r113 10 36 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=1.16
r114 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=0.56
r115 6 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r116 3 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%A_27_47# 1 2 9 13 15 18 20 24 25 28 31 33
c54 24 0 1.44392e-19 $X=0.995 $Y=1.16
r55 28 30 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.217 $Y=0.46
+ $X2=0.217 $Y2=0.625
r56 25 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=1.325
r57 25 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=0.995
r58 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.16 $X2=0.995 $Y2=1.16
r59 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.995 $Y=1.495
+ $X2=0.995 $Y2=1.16
r60 21 31 2.15711 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.58
+ $X2=0.217 $Y2=1.58
r61 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.91 $Y=1.58
+ $X2=0.995 $Y2=1.495
r62 20 21 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.91 $Y=1.58
+ $X2=0.345 $Y2=1.58
r63 16 31 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.217 $Y2=1.58
r64 16 18 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.217 $Y2=1.96
r65 15 31 4.27425 $w=2.12e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.175 $Y=1.495
+ $X2=0.217 $Y2=1.58
r66 15 30 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=0.175 $Y=1.495
+ $X2=0.175 $Y2=0.625
r67 13 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.56
+ $X2=0.955 $Y2=0.995
r68 9 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.945 $Y=1.985
+ $X2=0.945 $Y2=1.325
r69 2 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r70 1 28 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%A0 1 3 6 8 9 16
r34 13 16 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.665 $Y=1.16
+ $X2=1.905 $Y2=1.16
r35 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=1.615 $Y2=1.53
r36 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.16 $X2=1.665 $Y2=1.16
r37 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.325
+ $X2=1.905 $Y2=1.16
r38 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.905 $Y=1.325
+ $X2=1.905 $Y2=1.985
r39 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=0.995
+ $X2=1.905 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.905 $Y=0.995
+ $X2=1.905 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%A1 3 6 8 11 12 13
r34 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.16
+ $X2=2.35 $Y2=1.325
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.16
+ $X2=2.35 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.35
+ $Y=1.16 $X2=2.35 $Y2=1.16
r37 8 12 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.065 $Y=1.16
+ $X2=2.35 $Y2=1.16
r38 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.375 $Y=1.985
+ $X2=2.375 $Y2=1.325
r39 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.375 $Y=0.56
+ $X2=2.375 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%A_396_47# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 35 39 44 45 46 48 50 56 59 65
c127 45 0 1.83477e-19 $X=3.565 $Y=0.74
r128 62 63 61.7195 $w=3.28e-07 $l=4.2e-07 $layer=POLY_cond $X=4.21 $Y=1.16
+ $X2=4.63 $Y2=1.16
r129 57 65 27.186 $w=3.28e-07 $l=1.85e-07 $layer=POLY_cond $X=4.865 $Y=1.16
+ $X2=5.05 $Y2=1.16
r130 57 63 34.5335 $w=3.28e-07 $l=2.35e-07 $layer=POLY_cond $X=4.865 $Y=1.16
+ $X2=4.63 $Y2=1.16
r131 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.865
+ $Y=1.16 $X2=4.865 $Y2=1.16
r132 54 62 53.6372 $w=3.28e-07 $l=3.65e-07 $layer=POLY_cond $X=3.845 $Y=1.16
+ $X2=4.21 $Y2=1.16
r133 54 60 8.08232 $w=3.28e-07 $l=5.5e-08 $layer=POLY_cond $X=3.845 $Y=1.16
+ $X2=3.79 $Y2=1.16
r134 53 56 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.845 $Y=1.16
+ $X2=4.865 $Y2=1.16
r135 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.845
+ $Y=1.16 $X2=3.845 $Y2=1.16
r136 51 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=1.16
+ $X2=3.65 $Y2=1.16
r137 51 53 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.735 $Y=1.16
+ $X2=3.845 $Y2=1.16
r138 49 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=1.245
+ $X2=3.65 $Y2=1.16
r139 49 50 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.65 $Y=1.245
+ $X2=3.65 $Y2=1.595
r140 48 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=1.075
+ $X2=3.65 $Y2=1.16
r141 47 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.65 $Y=0.825
+ $X2=3.65 $Y2=1.075
r142 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.565 $Y=0.74
+ $X2=3.65 $Y2=0.825
r143 45 46 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.565 $Y=0.74
+ $X2=3.23 $Y2=0.74
r144 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.145 $Y=0.655
+ $X2=3.23 $Y2=0.74
r145 43 44 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.145 $Y=0.465
+ $X2=3.145 $Y2=0.655
r146 39 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.565 $Y=1.68
+ $X2=3.65 $Y2=1.595
r147 39 41 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=3.565 $Y=1.68
+ $X2=2.145 $Y2=1.68
r148 35 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=0.38
+ $X2=3.145 $Y2=0.465
r149 35 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.06 $Y=0.38
+ $X2=2.14 $Y2=0.38
r150 31 65 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.16
r151 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.985
r152 28 65 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=1.16
r153 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=0.56
r154 24 63 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=1.325
+ $X2=4.63 $Y2=1.16
r155 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.63 $Y=1.325
+ $X2=4.63 $Y2=1.985
r156 21 63 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=0.995
+ $X2=4.63 $Y2=1.16
r157 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.63 $Y=0.995
+ $X2=4.63 $Y2=0.56
r158 17 62 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.325
+ $X2=4.21 $Y2=1.16
r159 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.21 $Y=1.325
+ $X2=4.21 $Y2=1.985
r160 14 62 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=0.995
+ $X2=4.21 $Y2=1.16
r161 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.21 $Y=0.995
+ $X2=4.21 $Y2=0.56
r162 10 60 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=1.325
+ $X2=3.79 $Y2=1.16
r163 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.79 $Y=1.325
+ $X2=3.79 $Y2=1.985
r164 7 60 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=0.995
+ $X2=3.79 $Y2=1.16
r165 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.79 $Y=0.995
+ $X2=3.79 $Y2=0.56
r166 2 41 600 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.485 $X2=2.145 $Y2=1.68
r167 1 37 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.235 $X2=2.14 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%VPWR 1 2 3 4 15 19 23 25 27 29 31 36 41 46 52
+ 55 58 62
r77 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r78 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r79 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r80 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 50 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r82 50 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r83 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 47 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=2.72
+ $X2=4.42 $Y2=2.72
r85 47 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.585 $Y=2.72
+ $X2=4.83 $Y2=2.72
r86 46 61 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=5.307 $Y2=2.72
r87 46 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=4.83 $Y2=2.72
r88 45 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r89 45 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r90 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r91 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.72
+ $X2=3.58 $Y2=2.72
r92 42 44 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.72
+ $X2=3.91 $Y2=2.72
r93 41 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=4.42 $Y2=2.72
r94 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=3.91 $Y2=2.72
r95 40 56 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r96 40 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r97 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 37 52 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=0.667 $Y2=2.72
r99 37 39 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=1.15 $Y2=2.72
r100 36 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=3.58 $Y2=2.72
r101 36 39 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=1.15 $Y2=2.72
r102 31 52 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.667 $Y2=2.72
r103 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r104 29 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r106 25 61 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=5.26 $Y=2.635
+ $X2=5.307 $Y2=2.72
r107 25 27 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.26 $Y=2.635
+ $X2=5.26 $Y2=2
r108 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=2.635
+ $X2=4.42 $Y2=2.72
r109 21 23 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.42 $Y=2.635
+ $X2=4.42 $Y2=2
r110 17 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=2.635
+ $X2=3.58 $Y2=2.72
r111 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.58 $Y=2.635
+ $X2=3.58 $Y2=2.34
r112 13 52 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.667 $Y=2.635
+ $X2=0.667 $Y2=2.72
r113 13 15 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=0.667 $Y=2.635
+ $X2=0.667 $Y2=2
r114 4 27 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.485 $X2=5.26 $Y2=2
r115 3 23 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.285
+ $Y=1.485 $X2=4.42 $Y2=2
r116 2 19 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.485 $X2=3.58 $Y2=2.34
r117 1 15 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%A_204_297# 1 2 9 12
c23 1 0 1.44392e-19 $X=1.02 $Y=1.485
r24 12 14 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=2.02
+ $X2=1.165 $Y2=2.36
r25 7 14 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.34 $Y=2.36 $X2=1.165
+ $Y2=2.36
r26 7 9 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=1.34 $Y=2.36
+ $X2=2.605 $Y2=2.36
r27 2 9 600 $w=1.7e-07 $l=9.49342e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.485 $X2=2.605 $Y2=2.36
r28 1 12 300 $w=1.7e-07 $l=6.07577e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.485 $X2=1.175 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%A_314_297# 1 2 7 13
r22 11 13 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.16 $Y=2.105
+ $X2=3.16 $Y2=2.3
r23 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=3.16 $Y2=2.105
r24 7 9 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=1.695 $Y2=2.02
r25 2 13 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=1.485 $X2=3.16 $Y2=2.3
r26 1 9 600 $w=1.7e-07 $l=5.94222e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.485 $X2=1.695 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%X 1 2 3 4 15 19 21 22 23 24 27 31 34 36 37 38
+ 39 47 48 50 56
c58 47 0 1.01803e-19 $X=5.315 $Y=0.805
r59 48 56 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.315 $Y=1.575
+ $X2=5.315 $Y2=1.53
r60 47 50 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.315 $Y=0.805
+ $X2=5.315 $Y2=0.85
r61 39 48 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=1.66
+ $X2=5.315 $Y2=1.575
r62 39 56 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=5.315 $Y=1.51
+ $X2=5.315 $Y2=1.53
r63 38 39 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.315 $Y=1.19
+ $X2=5.315 $Y2=1.51
r64 37 47 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=0.72
+ $X2=5.315 $Y2=0.805
r65 37 38 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.315 $Y=0.87
+ $X2=5.315 $Y2=1.19
r66 37 50 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=5.315 $Y=0.87
+ $X2=5.315 $Y2=0.85
r67 35 39 14.9587 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=4.925 $Y=1.66
+ $X2=5.2 $Y2=1.66
r68 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=1.66
+ $X2=4.84 $Y2=1.66
r69 33 37 14.9587 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=4.925 $Y=0.72
+ $X2=5.2 $Y2=0.72
r70 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=0.72
+ $X2=4.84 $Y2=0.72
r71 29 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=1.745
+ $X2=4.84 $Y2=1.66
r72 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.84 $Y=1.745
+ $X2=4.84 $Y2=1.96
r73 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=0.635
+ $X2=4.84 $Y2=0.72
r74 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.84 $Y=0.635
+ $X2=4.84 $Y2=0.42
r75 23 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=1.66
+ $X2=4.84 $Y2=1.66
r76 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.755 $Y=1.66
+ $X2=4.085 $Y2=1.66
r77 21 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=0.72
+ $X2=4.84 $Y2=0.72
r78 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.755 $Y=0.72
+ $X2=4.085 $Y2=0.72
r79 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4 $Y=1.745
+ $X2=4.085 $Y2=1.66
r80 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4 $Y=1.745 $X2=4
+ $Y2=1.96
r81 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4 $Y=0.635
+ $X2=4.085 $Y2=0.72
r82 13 15 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4 $Y=0.635 $X2=4
+ $Y2=0.42
r83 4 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.705
+ $Y=1.485 $X2=4.84 $Y2=1.96
r84 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.865
+ $Y=1.485 $X2=4 $Y2=1.96
r85 2 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.705
+ $Y=0.235 $X2=4.84 $Y2=0.42
r86 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.865
+ $Y=0.235 $X2=4 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_4%VGND 1 2 3 4 15 19 23 25 27 29 31 36 41 46 52
+ 55 58 62
c86 25 0 1.01803e-19 $X=5.26 $Y=0.085
r87 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r88 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r89 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r90 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r91 50 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r92 50 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r93 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r94 47 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.42
+ $Y2=0
r95 47 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.83
+ $Y2=0
r96 46 61 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=5.307
+ $Y2=0
r97 46 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=4.83
+ $Y2=0
r98 45 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r99 45 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r100 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r101 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.58
+ $Y2=0
r102 42 44 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=0
+ $X2=3.91 $Y2=0
r103 41 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.42
+ $Y2=0
r104 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=3.91
+ $Y2=0
r105 40 56 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r106 40 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r107 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r108 37 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r109 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r110 36 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.58
+ $Y2=0
r111 36 39 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=1.15 $Y2=0
r112 31 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r113 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r114 29 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r115 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r116 25 61 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=5.26 $Y=0.085
+ $X2=5.307 $Y2=0
r117 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.26 $Y=0.085
+ $X2=5.26 $Y2=0.38
r118 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=0.085
+ $X2=4.42 $Y2=0
r119 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.42 $Y=0.085
+ $X2=4.42 $Y2=0.38
r120 17 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0
r121 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0.38
r122 13 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r123 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r124 4 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=5.26 $Y2=0.38
r125 3 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.285
+ $Y=0.235 $X2=4.42 $Y2=0.38
r126 2 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.235 $X2=3.58 $Y2=0.38
r127 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


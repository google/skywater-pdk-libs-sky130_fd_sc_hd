* File: sky130_fd_sc_hd__dlrtp_1.spice.SKY130_FD_SC_HD__DLRTP_1.pxi
* Created: Thu Aug 27 14:17:28 2020
* 
x_PM_SKY130_FD_SC_HD__DLRTP_1%GATE N_GATE_c_140_n N_GATE_c_135_n N_GATE_M1019_g
+ N_GATE_c_141_n N_GATE_M1009_g N_GATE_c_136_n N_GATE_c_142_n GATE GATE
+ N_GATE_c_138_n N_GATE_c_139_n PM_SKY130_FD_SC_HD__DLRTP_1%GATE
x_PM_SKY130_FD_SC_HD__DLRTP_1%A_27_47# N_A_27_47#_M1019_s N_A_27_47#_M1009_s
+ N_A_27_47#_M1010_g N_A_27_47#_M1000_g N_A_27_47#_c_179_n N_A_27_47#_M1004_g
+ N_A_27_47#_c_180_n N_A_27_47#_M1015_g N_A_27_47#_c_316_p N_A_27_47#_c_182_n
+ N_A_27_47#_c_183_n N_A_27_47#_c_191_n N_A_27_47#_c_192_n N_A_27_47#_c_184_n
+ N_A_27_47#_c_185_n N_A_27_47#_c_194_n N_A_27_47#_c_195_n N_A_27_47#_c_196_n
+ N_A_27_47#_c_197_n N_A_27_47#_c_198_n N_A_27_47#_c_186_n
+ PM_SKY130_FD_SC_HD__DLRTP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRTP_1%D N_D_c_325_n N_D_M1003_g N_D_M1014_g N_D_c_331_n
+ D N_D_c_327_n N_D_c_328_n PM_SKY130_FD_SC_HD__DLRTP_1%D
x_PM_SKY130_FD_SC_HD__DLRTP_1%A_299_47# N_A_299_47#_M1003_s N_A_299_47#_M1014_s
+ N_A_299_47#_c_374_n N_A_299_47#_M1006_g N_A_299_47#_M1012_g
+ N_A_299_47#_c_382_n N_A_299_47#_c_376_n N_A_299_47#_c_377_n
+ N_A_299_47#_c_378_n N_A_299_47#_c_384_n N_A_299_47#_c_379_n
+ N_A_299_47#_c_380_n PM_SKY130_FD_SC_HD__DLRTP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__DLRTP_1%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1007_g N_A_193_47#_M1001_g N_A_193_47#_c_459_n
+ N_A_193_47#_c_460_n N_A_193_47#_c_467_n N_A_193_47#_c_461_n
+ N_A_193_47#_c_462_n N_A_193_47#_c_468_n N_A_193_47#_c_469_n
+ N_A_193_47#_c_470_n N_A_193_47#_c_471_n N_A_193_47#_c_463_n
+ N_A_193_47#_c_472_n N_A_193_47#_c_473_n PM_SKY130_FD_SC_HD__DLRTP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRTP_1%A_711_21# N_A_711_21#_M1005_s N_A_711_21#_M1002_d
+ N_A_711_21#_M1016_g N_A_711_21#_c_579_n N_A_711_21#_M1018_g
+ N_A_711_21#_M1017_g N_A_711_21#_M1011_g N_A_711_21#_c_580_n
+ N_A_711_21#_c_581_n N_A_711_21#_c_590_n N_A_711_21#_c_582_n
+ N_A_711_21#_c_634_p N_A_711_21#_c_592_n N_A_711_21#_c_583_n
+ N_A_711_21#_c_593_n N_A_711_21#_c_607_p N_A_711_21#_c_608_p
+ N_A_711_21#_c_584_n N_A_711_21#_c_585_n N_A_711_21#_c_586_n
+ PM_SKY130_FD_SC_HD__DLRTP_1%A_711_21#
x_PM_SKY130_FD_SC_HD__DLRTP_1%A_560_425# N_A_560_425#_M1007_d
+ N_A_560_425#_M1004_d N_A_560_425#_c_688_n N_A_560_425#_M1005_g
+ N_A_560_425#_M1002_g N_A_560_425#_c_689_n N_A_560_425#_c_690_n
+ N_A_560_425#_c_704_n N_A_560_425#_c_699_n N_A_560_425#_c_691_n
+ N_A_560_425#_c_697_n N_A_560_425#_c_692_n N_A_560_425#_c_693_n
+ PM_SKY130_FD_SC_HD__DLRTP_1%A_560_425#
x_PM_SKY130_FD_SC_HD__DLRTP_1%RESET_B N_RESET_B_M1008_g N_RESET_B_M1013_g
+ RESET_B RESET_B RESET_B N_RESET_B_c_775_n N_RESET_B_c_776_n N_RESET_B_c_777_n
+ PM_SKY130_FD_SC_HD__DLRTP_1%RESET_B
x_PM_SKY130_FD_SC_HD__DLRTP_1%VPWR N_VPWR_M1009_d N_VPWR_M1014_d N_VPWR_M1018_d
+ N_VPWR_M1013_d N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_814_n
+ N_VPWR_c_815_n VPWR N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n
+ N_VPWR_c_819_n N_VPWR_c_810_n N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n
+ PM_SKY130_FD_SC_HD__DLRTP_1%VPWR
x_PM_SKY130_FD_SC_HD__DLRTP_1%Q N_Q_M1017_d N_Q_M1011_d Q Q Q Q N_Q_c_906_n
+ PM_SKY130_FD_SC_HD__DLRTP_1%Q
x_PM_SKY130_FD_SC_HD__DLRTP_1%VGND N_VGND_M1019_d N_VGND_M1003_d N_VGND_M1016_d
+ N_VGND_M1008_d N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n N_VGND_c_925_n
+ VGND N_VGND_c_926_n N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n
+ N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n N_VGND_c_933_n N_VGND_c_934_n
+ N_VGND_c_935_n PM_SKY130_FD_SC_HD__DLRTP_1%VGND
cc_1 VNB N_GATE_c_135_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_c_136_n 0.0234948f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE 0.0153903f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_GATE_c_138_n 0.0210092f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_GATE_c_139_n 0.0148328f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1010_g 0.0396883f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_179_n 0.00823882f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_8 VNB N_A_27_47#_c_180_n 0.0071182f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_9 VNB N_A_27_47#_M1015_g 0.0454977f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_10 VNB N_A_27_47#_c_182_n 0.0020589f $X=-0.19 $Y=-0.24 $X2=0.205 $Y2=1.53
cc_11 VNB N_A_27_47#_c_183_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_184_n 8.66974e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_185_n 0.00418748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_186_n 0.0238009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_D_c_325_n 0.00566647f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.07
cc_16 VNB N_D_M1003_g 0.025882f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_17 VNB N_D_c_327_n 0.00464339f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_D_c_328_n 0.0428882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_299_47#_c_374_n 0.0170226f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_20 VNB N_A_299_47#_M1012_g 0.0143435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_299_47#_c_376_n 0.00199643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_377_n 0.00552014f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_23 VNB N_A_299_47#_c_378_n 0.00335034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_299_47#_c_379_n 0.00286279f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_25 VNB N_A_299_47#_c_380_n 0.0264162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_c_459_n 0.0139271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_460_n 0.00359704f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_28 VNB N_A_193_47#_c_461_n 0.026888f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_29 VNB N_A_193_47#_c_462_n 0.00327791f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_30 VNB N_A_193_47#_c_463_n 0.0174156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_711_21#_c_579_n 0.0186695f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_32 VNB N_A_711_21#_c_580_n 0.0190662f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_33 VNB N_A_711_21#_c_581_n 0.0120904f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_34 VNB N_A_711_21#_c_582_n 0.00159796f $X=-0.19 $Y=-0.24 $X2=0.205 $Y2=1.53
cc_35 VNB N_A_711_21#_c_583_n 0.00603427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_711_21#_c_584_n 0.00398889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_711_21#_c_585_n 0.0230746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_711_21#_c_586_n 0.0196016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_560_425#_c_688_n 0.0206723f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_40 VNB N_A_560_425#_c_689_n 0.0394607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_560_425#_c_690_n 0.01017f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_42 VNB N_A_560_425#_c_691_n 0.00319466f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_43 VNB N_A_560_425#_c_692_n 0.00298369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_560_425#_c_693_n 0.00368968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB RESET_B 0.00165174f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_46 VNB N_RESET_B_c_775_n 0.0205324f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_47 VNB N_RESET_B_c_776_n 0.00182864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_777_n 0.0173277f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_49 VNB N_VPWR_c_810_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB Q 0.0157845f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_51 VNB N_Q_c_906_n 0.0248025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_922_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_53 VNB N_VGND_c_923_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_54 VNB N_VGND_c_924_n 0.00967467f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_55 VNB N_VGND_c_925_n 0.00269179f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_56 VNB N_VGND_c_926_n 0.0153564f $X=-0.19 $Y=-0.24 $X2=0.205 $Y2=1.53
cc_57 VNB N_VGND_c_927_n 0.0269775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_928_n 0.0423817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_929_n 0.0307951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_930_n 0.0160478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_931_n 0.314468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_932_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_933_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_934_n 0.00516809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_935_n 0.0043871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VPB N_GATE_c_140_n 0.0129143f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_67 VPB N_GATE_c_141_n 0.0186097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_68 VPB N_GATE_c_142_n 0.0239197f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_69 VPB GATE 0.0127706f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_70 VPB N_GATE_c_138_n 0.0106807f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_71 VPB N_A_27_47#_M1000_g 0.0394598f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_72 VPB N_A_27_47#_c_179_n 0.0332204f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_73 VPB N_A_27_47#_M1004_g 0.0340937f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_74 VPB N_A_27_47#_c_180_n 0.0263663f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_75 VPB N_A_27_47#_c_191_n 0.00108837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_192_n 0.0300397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_184_n 6.56074e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_194_n 0.0208829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_195_n 0.00327791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_196_n 0.00545214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_197_n 0.00344459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_198_n 0.00977979f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_186_n 0.0121227f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_D_c_325_n 0.0164643f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.07
cc_85 VPB N_D_M1014_g 0.0212086f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_86 VPB N_D_c_331_n 0.0183374f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_87 VPB N_D_c_327_n 0.00155563f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_88 VPB N_A_299_47#_M1012_g 0.0380048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_299_47#_c_382_n 0.00699762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_299_47#_c_378_n 0.00388743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_299_47#_c_384_n 0.00728202f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_92 VPB N_A_193_47#_M1001_g 0.0231112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_193_47#_c_459_n 0.00769231f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_193_47#_c_460_n 0.00223761f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_95 VPB N_A_193_47#_c_467_n 0.00278943f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_96 VPB N_A_193_47#_c_468_n 0.00795485f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.19
cc_97 VPB N_A_193_47#_c_469_n 0.0024125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_193_47#_c_470_n 0.00681938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_193_47#_c_471_n 0.00364199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_193_47#_c_472_n 0.0292161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_193_47#_c_473_n 0.00802597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_711_21#_c_579_n 0.0146305f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_103 VPB N_A_711_21#_M1018_g 0.0262376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_711_21#_M1011_g 0.0215601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_711_21#_c_590_n 0.044704f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.19
cc_106 VPB N_A_711_21#_c_582_n 0.00232431f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.53
cc_107 VPB N_A_711_21#_c_592_n 0.00139379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_711_21#_c_593_n 0.00423442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_711_21#_c_585_n 0.005118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_560_425#_M1002_g 0.0226618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_560_425#_c_689_n 0.0145732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_560_425#_c_690_n 6.56128e-19 $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_113 VPB N_A_560_425#_c_697_n 0.007565f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_114 VPB N_A_560_425#_c_692_n 0.00167692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_RESET_B_M1013_g 0.0201873f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_116 VPB N_RESET_B_c_775_n 0.00452632f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_117 VPB N_RESET_B_c_776_n 0.00230524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_811_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_119 VPB N_VPWR_c_812_n 0.0036773f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_120 VPB N_VPWR_c_813_n 0.00280379f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_121 VPB N_VPWR_c_814_n 0.0165876f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_122 VPB N_VPWR_c_815_n 0.0454618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_816_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_817_n 0.029347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_818_n 0.0189266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_819_n 0.0151046f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_810_n 0.0523567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_821_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_822_n 0.00407272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_823_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB Q 0.00494099f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_132 VPB Q 0.0252202f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_133 VPB N_Q_c_906_n 0.0151107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 N_GATE_c_135_n N_A_27_47#_M1010_g 0.0187884f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_135 N_GATE_c_139_n N_A_27_47#_M1010_g 0.00412351f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_136 N_GATE_c_142_n N_A_27_47#_M1000_g 0.026381f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_137 N_GATE_c_138_n N_A_27_47#_M1000_g 0.0051869f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_138 N_GATE_c_135_n N_A_27_47#_c_182_n 0.00663338f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_139 N_GATE_c_136_n N_A_27_47#_c_182_n 0.0104883f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_140 N_GATE_c_136_n N_A_27_47#_c_183_n 0.00696191f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_141 GATE N_A_27_47#_c_183_n 0.0125186f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_142 N_GATE_c_138_n N_A_27_47#_c_183_n 3.35813e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_143 N_GATE_c_141_n N_A_27_47#_c_191_n 0.01356f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_144 N_GATE_c_142_n N_A_27_47#_c_191_n 0.00216816f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_145 N_GATE_c_141_n N_A_27_47#_c_192_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_146 N_GATE_c_142_n N_A_27_47#_c_192_n 0.00423203f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_147 GATE N_A_27_47#_c_192_n 0.0217264f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_148 N_GATE_c_138_n N_A_27_47#_c_192_n 5.66731e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_149 N_GATE_c_138_n N_A_27_47#_c_184_n 0.00320294f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_150 N_GATE_c_136_n N_A_27_47#_c_185_n 0.00180622f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_151 GATE N_A_27_47#_c_185_n 0.0288278f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_152 N_GATE_c_139_n N_A_27_47#_c_185_n 0.00152291f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_153 N_GATE_c_140_n N_A_27_47#_c_195_n 0.00339489f $X=0.3 $Y=1.59 $X2=0 $Y2=0
cc_154 N_GATE_c_142_n N_A_27_47#_c_195_n 0.00103052f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_155 GATE N_A_27_47#_c_195_n 0.00639826f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_156 N_GATE_c_140_n N_A_27_47#_c_196_n 7.64926e-19 $X=0.3 $Y=1.59 $X2=0 $Y2=0
cc_157 N_GATE_c_142_n N_A_27_47#_c_196_n 0.00425368f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_158 GATE N_A_27_47#_c_186_n 9.09032e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_159 N_GATE_c_138_n N_A_27_47#_c_186_n 0.0165939f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_160 N_GATE_c_141_n N_VPWR_c_811_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_161 N_GATE_c_141_n N_VPWR_c_816_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_162 N_GATE_c_141_n N_VPWR_c_810_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_163 N_GATE_c_135_n N_VGND_c_922_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_164 N_GATE_c_135_n N_VGND_c_926_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_165 N_GATE_c_136_n N_VGND_c_926_n 4.87495e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_166 N_GATE_c_135_n N_VGND_c_931_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_194_n N_D_c_325_n 0.00200477f $X=2.385 $Y=1.53 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_186_n N_D_c_325_n 0.00328108f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_169 N_A_27_47#_M1000_g N_D_c_331_n 0.00328108f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_194_n N_D_c_327_n 0.00814614f $X=2.385 $Y=1.53 $X2=0 $Y2=0
cc_171 N_A_27_47#_M1010_g N_D_c_328_n 0.00565959f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_194_n N_D_c_328_n 0.00194191f $X=2.385 $Y=1.53 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_179_n N_A_299_47#_M1012_g 0.060232f $X=2.725 $Y=1.69 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_194_n N_A_299_47#_M1012_g 0.00546549f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_197_n N_A_299_47#_M1012_g 0.0014344f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_198_n N_A_299_47#_M1012_g 0.00240655f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_194_n N_A_299_47#_c_382_n 5.24155e-19 $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_198_n N_A_299_47#_c_382_n 5.60149e-19 $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_194_n N_A_299_47#_c_377_n 0.00748499f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_194_n N_A_299_47#_c_378_n 0.0114159f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_197_n N_A_299_47#_c_378_n 0.00124596f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_198_n N_A_299_47#_c_378_n 0.00586183f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_194_n N_A_299_47#_c_384_n 0.0208797f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_197_n N_A_299_47#_c_384_n 0.00130924f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_198_n N_A_299_47#_c_384_n 0.00669529f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_194_n N_A_299_47#_c_380_n 0.0010667f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_M1004_g N_A_193_47#_M1001_g 0.0117482f $X=2.725 $Y=2.305 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1010_g N_A_193_47#_c_459_n 0.00584642f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_182_n N_A_193_47#_c_459_n 0.00977084f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_184_n N_A_193_47#_c_459_n 0.0230475f $X=0.75 $Y=1.235 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_185_n N_A_193_47#_c_459_n 0.0156045f $X=0.72 $Y=1.07 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_194_n N_A_193_47#_c_459_n 0.0183956f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_195_n N_A_193_47#_c_459_n 0.00229404f $X=0.835 $Y=1.53 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_196_n N_A_193_47#_c_459_n 0.0204242f $X=0.69 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_179_n N_A_193_47#_c_460_n 0.00134843f $X=2.725 $Y=1.69 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_180_n N_A_193_47#_c_460_n 0.0110393f $X=3.12 $Y=1.38 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_M1015_g N_A_193_47#_c_460_n 0.00749827f $X=3.195 $Y=0.445
+ $X2=0 $Y2=0
cc_198 N_A_27_47#_c_197_n N_A_193_47#_c_460_n 0.00112777f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_198_n N_A_193_47#_c_460_n 0.0210008f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_194_n N_A_193_47#_c_467_n 0.00177113f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_186_n N_A_193_47#_c_467_n 0.00584642f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_179_n N_A_193_47#_c_461_n 0.0181914f $X=2.725 $Y=1.69 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1015_g N_A_193_47#_c_461_n 0.0213129f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_198_n N_A_193_47#_c_461_n 8.59209e-19 $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_179_n N_A_193_47#_c_462_n 0.00106939f $X=2.725 $Y=1.69 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_180_n N_A_193_47#_c_462_n 0.00390689f $X=3.12 $Y=1.38 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1015_g N_A_193_47#_c_462_n 0.0109049f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_198_n N_A_193_47#_c_462_n 0.00769017f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_M1004_g N_A_193_47#_c_468_n 0.00623292f $X=2.725 $Y=2.305
+ $X2=0 $Y2=0
cc_210 N_A_27_47#_c_180_n N_A_193_47#_c_468_n 5.63902e-19 $X=3.12 $Y=1.38 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_194_n N_A_193_47#_c_468_n 0.0853921f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_197_n N_A_193_47#_c_468_n 0.0266229f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_198_n N_A_193_47#_c_468_n 0.0130908f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1000_g N_A_193_47#_c_469_n 0.00459685f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_191_n N_A_193_47#_c_469_n 0.00552994f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_194_n N_A_193_47#_c_469_n 0.02594f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_196_n N_A_193_47#_c_469_n 0.00110781f $X=0.69 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_M1000_g N_A_193_47#_c_470_n 0.00584642f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_191_n N_A_193_47#_c_470_n 0.00288446f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1004_g N_A_193_47#_c_471_n 0.001487f $X=2.725 $Y=2.305 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_180_n N_A_193_47#_c_471_n 0.00298233f $X=3.12 $Y=1.38 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_M1015_g N_A_193_47#_c_463_n 0.013188f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_179_n N_A_193_47#_c_472_n 0.00153544f $X=2.725 $Y=1.69 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_M1004_g N_A_193_47#_c_472_n 0.015111f $X=2.725 $Y=2.305 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_180_n N_A_193_47#_c_472_n 0.016666f $X=3.12 $Y=1.38 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_179_n N_A_193_47#_c_473_n 8.81078e-19 $X=2.725 $Y=1.69 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_M1004_g N_A_193_47#_c_473_n 0.00454743f $X=2.725 $Y=2.305
+ $X2=0 $Y2=0
cc_228 N_A_27_47#_c_180_n N_A_193_47#_c_473_n 0.00309135f $X=3.12 $Y=1.38 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_198_n N_A_193_47#_c_473_n 0.00289412f $X=2.53 $Y=1.53 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_M1015_g N_A_711_21#_c_579_n 0.0183643f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1015_g N_A_711_21#_c_580_n 0.0344194f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1015_g N_A_560_425#_c_699_n 0.00942169f $X=3.195 $Y=0.445
+ $X2=0 $Y2=0
cc_233 N_A_27_47#_M1015_g N_A_560_425#_c_691_n 0.00629933f $X=3.195 $Y=0.445
+ $X2=0 $Y2=0
cc_234 N_A_27_47#_c_180_n N_A_560_425#_c_697_n 0.00102188f $X=3.12 $Y=1.38 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_M1015_g N_A_560_425#_c_693_n 0.00244306f $X=3.195 $Y=0.445
+ $X2=0 $Y2=0
cc_236 N_A_27_47#_c_191_n N_VPWR_M1009_d 0.00191359f $X=0.605 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_237 N_A_27_47#_M1000_g N_VPWR_c_811_n 0.009762f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_191_n N_VPWR_c_811_n 0.0150624f $X=0.605 $Y=1.88 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_192_n N_VPWR_c_811_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_194_n N_VPWR_c_811_n 2.56192e-19 $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_195_n N_VPWR_c_811_n 0.00313651f $X=0.835 $Y=1.53 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1004_g N_VPWR_c_812_n 0.00384689f $X=2.725 $Y=2.305 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_194_n N_VPWR_c_812_n 0.00166786f $X=2.385 $Y=1.53 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1004_g N_VPWR_c_815_n 0.00585385f $X=2.725 $Y=2.305 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_191_n N_VPWR_c_816_n 0.0018545f $X=0.605 $Y=1.88 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_192_n N_VPWR_c_816_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_247 N_A_27_47#_M1000_g N_VPWR_c_817_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1000_g N_VPWR_c_810_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1004_g N_VPWR_c_810_n 0.00680708f $X=2.725 $Y=2.305 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_191_n N_VPWR_c_810_n 0.00481546f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_192_n N_VPWR_c_810_n 0.00993215f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_182_n N_VGND_M1019_d 0.00164702f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_27_47#_M1010_g N_VGND_c_922_n 0.0118858f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_182_n N_VGND_c_922_n 0.0150545f $X=0.605 $Y=0.72 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_184_n N_VGND_c_922_n 0.00119775f $X=0.75 $Y=1.235 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_186_n N_VGND_c_922_n 5.88506e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_316_p N_VGND_c_926_n 0.00735289f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_182_n N_VGND_c_926_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1010_g N_VGND_c_927_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_260 N_A_27_47#_M1015_g N_VGND_c_928_n 0.0037981f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_M1019_s N_VGND_c_931_n 0.00358206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_M1010_g N_VGND_c_931_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1015_g N_VGND_c_931_n 0.00546293f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_316_p N_VGND_c_931_n 0.00626856f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_182_n N_VGND_c_931_n 0.005471f $X=0.605 $Y=0.72 $X2=0 $Y2=0
cc_266 N_D_M1003_g N_A_299_47#_c_374_n 0.0152919f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_267 N_D_c_325_n N_A_299_47#_M1012_g 0.00785152f $X=1.66 $Y=1.565 $X2=0 $Y2=0
cc_268 N_D_c_331_n N_A_299_47#_M1012_g 0.0197289f $X=1.83 $Y=1.64 $X2=0 $Y2=0
cc_269 N_D_c_328_n N_A_299_47#_M1012_g 0.00438557f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_270 N_D_M1014_g N_A_299_47#_c_382_n 0.0109755f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_271 N_D_c_331_n N_A_299_47#_c_382_n 0.00707117f $X=1.83 $Y=1.64 $X2=0 $Y2=0
cc_272 N_D_M1003_g N_A_299_47#_c_376_n 0.0147009f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_273 N_D_c_327_n N_A_299_47#_c_376_n 0.00446116f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_274 N_D_c_328_n N_A_299_47#_c_376_n 0.00136061f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_275 N_D_M1003_g N_A_299_47#_c_377_n 0.00587811f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_276 N_D_c_327_n N_A_299_47#_c_377_n 0.0108045f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_277 N_D_c_325_n N_A_299_47#_c_378_n 0.00383431f $X=1.66 $Y=1.565 $X2=0 $Y2=0
cc_278 N_D_c_327_n N_A_299_47#_c_378_n 0.0170179f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_279 N_D_c_328_n N_A_299_47#_c_378_n 9.20678e-19 $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_280 N_D_c_325_n N_A_299_47#_c_384_n 0.00399209f $X=1.66 $Y=1.565 $X2=0 $Y2=0
cc_281 N_D_c_331_n N_A_299_47#_c_384_n 0.00876191f $X=1.83 $Y=1.64 $X2=0 $Y2=0
cc_282 N_D_c_327_n N_A_299_47#_c_384_n 0.0218846f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_283 N_D_c_328_n N_A_299_47#_c_384_n 0.00285404f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_284 N_D_M1003_g N_A_299_47#_c_379_n 0.00120862f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_285 N_D_c_327_n N_A_299_47#_c_379_n 0.01591f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_286 N_D_c_328_n N_A_299_47#_c_379_n 0.00539057f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_287 N_D_M1003_g N_A_299_47#_c_380_n 0.0203576f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_288 N_D_c_325_n N_A_193_47#_c_459_n 0.00362589f $X=1.66 $Y=1.565 $X2=0 $Y2=0
cc_289 N_D_M1003_g N_A_193_47#_c_459_n 0.00203361f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_290 N_D_c_327_n N_A_193_47#_c_459_n 0.0224186f $X=1.6 $Y=1.04 $X2=0 $Y2=0
cc_291 N_D_c_328_n N_A_193_47#_c_459_n 0.00258753f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_292 N_D_M1014_g N_A_193_47#_c_467_n 0.00113329f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_293 N_D_M1014_g N_A_193_47#_c_468_n 0.00297192f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_294 N_D_M1014_g N_VPWR_c_812_n 0.00302106f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_295 N_D_M1014_g N_VPWR_c_817_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_296 N_D_M1014_g N_VPWR_c_810_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_297 N_D_M1003_g N_VGND_c_923_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_298 N_D_M1003_g N_VGND_c_927_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_299 N_D_M1003_g N_VGND_c_931_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_300 N_D_c_328_n N_VGND_c_931_n 0.00104112f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_301 N_A_299_47#_c_382_n N_A_193_47#_c_459_n 0.00120694f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_302 N_A_299_47#_c_384_n N_A_193_47#_c_459_n 0.00925144f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_303 N_A_299_47#_c_379_n N_A_193_47#_c_459_n 0.020446f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_304 N_A_299_47#_M1012_g N_A_193_47#_c_460_n 0.00457405f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_305 N_A_299_47#_c_382_n N_A_193_47#_c_467_n 0.051003f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_306 N_A_299_47#_c_377_n N_A_193_47#_c_461_n 0.00114463f $X=2.03 $Y=1.095
+ $X2=0 $Y2=0
cc_307 N_A_299_47#_c_380_n N_A_193_47#_c_461_n 0.0157423f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_308 N_A_299_47#_c_377_n N_A_193_47#_c_462_n 0.0144797f $X=2.03 $Y=1.095 $X2=0
+ $Y2=0
cc_309 N_A_299_47#_c_380_n N_A_193_47#_c_462_n 0.00113059f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_310 N_A_299_47#_M1012_g N_A_193_47#_c_468_n 0.00405325f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_311 N_A_299_47#_c_382_n N_A_193_47#_c_468_n 0.0220246f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_312 N_A_299_47#_c_384_n N_A_193_47#_c_468_n 0.00554627f $X=2.03 $Y=1.58 $X2=0
+ $Y2=0
cc_313 N_A_299_47#_c_382_n N_A_193_47#_c_469_n 0.00276522f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_314 N_A_299_47#_c_374_n N_A_193_47#_c_463_n 0.0233562f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_315 N_A_299_47#_c_374_n N_A_560_425#_c_699_n 6.57184e-19 $X=2.25 $Y=0.765
+ $X2=0 $Y2=0
cc_316 N_A_299_47#_M1012_g N_VPWR_c_812_n 0.021162f $X=2.25 $Y=2.165 $X2=0 $Y2=0
cc_317 N_A_299_47#_c_382_n N_VPWR_c_812_n 0.0234958f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_318 N_A_299_47#_c_384_n N_VPWR_c_812_n 0.0106739f $X=2.03 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A_299_47#_M1012_g N_VPWR_c_815_n 0.00310428f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_320 N_A_299_47#_c_382_n N_VPWR_c_817_n 0.0173028f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_321 N_A_299_47#_M1014_s N_VPWR_c_810_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_322 N_A_299_47#_M1012_g N_VPWR_c_810_n 0.00335906f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_323 N_A_299_47#_c_382_n N_VPWR_c_810_n 0.00621325f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_324 N_A_299_47#_c_377_n N_VGND_M1003_d 0.00209965f $X=2.03 $Y=1.095 $X2=0
+ $Y2=0
cc_325 N_A_299_47#_c_374_n N_VGND_c_923_n 0.00955928f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_326 N_A_299_47#_c_376_n N_VGND_c_923_n 0.0020169f $X=1.945 $Y=0.7 $X2=0 $Y2=0
cc_327 N_A_299_47#_c_377_n N_VGND_c_923_n 0.0151358f $X=2.03 $Y=1.095 $X2=0
+ $Y2=0
cc_328 N_A_299_47#_c_380_n N_VGND_c_923_n 2.06305e-19 $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_329 N_A_299_47#_c_376_n N_VGND_c_927_n 0.00255672f $X=1.945 $Y=0.7 $X2=0
+ $Y2=0
cc_330 N_A_299_47#_c_379_n N_VGND_c_927_n 0.00819232f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_331 N_A_299_47#_c_374_n N_VGND_c_928_n 0.0046653f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_332 N_A_299_47#_c_380_n N_VGND_c_928_n 9.48611e-19 $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_333 N_A_299_47#_M1003_s N_VGND_c_931_n 0.00252595f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_334 N_A_299_47#_c_374_n N_VGND_c_931_n 0.0044965f $X=2.25 $Y=0.765 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_376_n N_VGND_c_931_n 0.00461622f $X=1.945 $Y=0.7 $X2=0
+ $Y2=0
cc_336 N_A_299_47#_c_377_n N_VGND_c_931_n 0.0054616f $X=2.03 $Y=1.095 $X2=0
+ $Y2=0
cc_337 N_A_299_47#_c_379_n N_VGND_c_931_n 0.00698341f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_380_n N_VGND_c_931_n 0.00117722f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_339 N_A_193_47#_c_460_n N_A_711_21#_c_579_n 0.00127278f $X=3.125 $Y=1.635
+ $X2=0 $Y2=0
cc_340 N_A_193_47#_M1001_g N_A_711_21#_M1018_g 0.0162325f $X=3.245 $Y=2.305
+ $X2=0 $Y2=0
cc_341 N_A_193_47#_c_472_n N_A_711_21#_M1018_g 0.00160095f $X=3.245 $Y=1.8 $X2=0
+ $Y2=0
cc_342 N_A_193_47#_c_472_n N_A_711_21#_c_590_n 0.00991944f $X=3.245 $Y=1.8 $X2=0
+ $Y2=0
cc_343 N_A_193_47#_c_473_n N_A_711_21#_c_590_n 3.30195e-19 $X=3.125 $Y=1.815
+ $X2=0 $Y2=0
cc_344 N_A_193_47#_M1001_g N_A_560_425#_c_704_n 0.0100776f $X=3.245 $Y=2.305
+ $X2=0 $Y2=0
cc_345 N_A_193_47#_c_468_n N_A_560_425#_c_704_n 0.00110181f $X=2.865 $Y=1.87
+ $X2=0 $Y2=0
cc_346 N_A_193_47#_c_471_n N_A_560_425#_c_704_n 0.00213959f $X=3.01 $Y=1.87
+ $X2=0 $Y2=0
cc_347 N_A_193_47#_c_472_n N_A_560_425#_c_704_n 7.42338e-19 $X=3.245 $Y=1.8
+ $X2=0 $Y2=0
cc_348 N_A_193_47#_c_473_n N_A_560_425#_c_704_n 0.0157906f $X=3.125 $Y=1.815
+ $X2=0 $Y2=0
cc_349 N_A_193_47#_c_461_n N_A_560_425#_c_699_n 0.00136088f $X=2.775 $Y=0.93
+ $X2=0 $Y2=0
cc_350 N_A_193_47#_c_462_n N_A_560_425#_c_699_n 0.0205447f $X=3.125 $Y=0.93
+ $X2=0 $Y2=0
cc_351 N_A_193_47#_c_463_n N_A_560_425#_c_699_n 0.00410631f $X=2.775 $Y=0.765
+ $X2=0 $Y2=0
cc_352 N_A_193_47#_c_462_n N_A_560_425#_c_691_n 0.0179688f $X=3.125 $Y=0.93
+ $X2=0 $Y2=0
cc_353 N_A_193_47#_M1001_g N_A_560_425#_c_697_n 0.00642569f $X=3.245 $Y=2.305
+ $X2=0 $Y2=0
cc_354 N_A_193_47#_c_460_n N_A_560_425#_c_697_n 0.0200766f $X=3.125 $Y=1.635
+ $X2=0 $Y2=0
cc_355 N_A_193_47#_c_471_n N_A_560_425#_c_697_n 0.00128736f $X=3.01 $Y=1.87
+ $X2=0 $Y2=0
cc_356 N_A_193_47#_c_472_n N_A_560_425#_c_697_n 0.00197109f $X=3.245 $Y=1.8
+ $X2=0 $Y2=0
cc_357 N_A_193_47#_c_473_n N_A_560_425#_c_697_n 0.0236633f $X=3.125 $Y=1.815
+ $X2=0 $Y2=0
cc_358 N_A_193_47#_c_460_n N_A_560_425#_c_693_n 0.0170765f $X=3.125 $Y=1.635
+ $X2=0 $Y2=0
cc_359 N_A_193_47#_c_462_n N_A_560_425#_c_693_n 0.00869845f $X=3.125 $Y=0.93
+ $X2=0 $Y2=0
cc_360 N_A_193_47#_c_468_n N_VPWR_M1014_d 6.81311e-19 $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_361 N_A_193_47#_c_470_n N_VPWR_c_811_n 0.0127345f $X=1.15 $Y=1.87 $X2=0 $Y2=0
cc_362 N_A_193_47#_c_468_n N_VPWR_c_812_n 0.0175545f $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_363 N_A_193_47#_c_473_n N_VPWR_c_812_n 0.00243347f $X=3.125 $Y=1.815 $X2=0
+ $Y2=0
cc_364 N_A_193_47#_M1001_g N_VPWR_c_815_n 0.00366111f $X=3.245 $Y=2.305 $X2=0
+ $Y2=0
cc_365 N_A_193_47#_c_470_n N_VPWR_c_817_n 0.0156296f $X=1.15 $Y=1.87 $X2=0 $Y2=0
cc_366 N_A_193_47#_M1001_g N_VPWR_c_810_n 0.00584911f $X=3.245 $Y=2.305 $X2=0
+ $Y2=0
cc_367 N_A_193_47#_c_468_n N_VPWR_c_810_n 0.075155f $X=2.865 $Y=1.87 $X2=0 $Y2=0
cc_368 N_A_193_47#_c_469_n N_VPWR_c_810_n 0.0151864f $X=1.295 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_193_47#_c_470_n N_VPWR_c_810_n 0.00381175f $X=1.15 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_471_n N_VPWR_c_810_n 0.0147664f $X=3.01 $Y=1.87 $X2=0 $Y2=0
cc_371 N_A_193_47#_c_468_n A_465_369# 0.00395093f $X=2.865 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_372 N_A_193_47#_c_463_n N_VGND_c_923_n 0.00177965f $X=2.775 $Y=0.765 $X2=0
+ $Y2=0
cc_373 N_A_193_47#_c_459_n N_VGND_c_927_n 0.00732874f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_374 N_A_193_47#_c_461_n N_VGND_c_928_n 8.76041e-19 $X=2.775 $Y=0.93 $X2=0
+ $Y2=0
cc_375 N_A_193_47#_c_463_n N_VGND_c_928_n 0.00551122f $X=2.775 $Y=0.765 $X2=0
+ $Y2=0
cc_376 N_A_193_47#_M1010_d N_VGND_c_931_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_c_459_n N_VGND_c_931_n 0.00616598f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_378 N_A_193_47#_c_461_n N_VGND_c_931_n 0.00117722f $X=2.775 $Y=0.93 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_462_n N_VGND_c_931_n 0.00485016f $X=3.125 $Y=0.93 $X2=0
+ $Y2=0
cc_380 N_A_193_47#_c_463_n N_VGND_c_931_n 0.00636171f $X=2.775 $Y=0.765 $X2=0
+ $Y2=0
cc_381 N_A_711_21#_c_582_n N_A_560_425#_c_688_n 0.00449097f $X=4.46 $Y=1.505
+ $X2=0 $Y2=0
cc_382 N_A_711_21#_c_583_n N_A_560_425#_c_688_n 0.00829764f $X=4.36 $Y=0.38
+ $X2=0 $Y2=0
cc_383 N_A_711_21#_M1018_g N_A_560_425#_M1002_g 0.00838165f $X=3.81 $Y=2.275
+ $X2=0 $Y2=0
cc_384 N_A_711_21#_c_590_n N_A_560_425#_M1002_g 0.00737954f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_385 N_A_711_21#_c_582_n N_A_560_425#_M1002_g 0.00757787f $X=4.46 $Y=1.505
+ $X2=0 $Y2=0
cc_386 N_A_711_21#_c_607_p N_A_560_425#_M1002_g 0.0165258f $X=4.795 $Y=1.685
+ $X2=0 $Y2=0
cc_387 N_A_711_21#_c_608_p N_A_560_425#_M1002_g 0.0189805f $X=4.965 $Y=1.685
+ $X2=0 $Y2=0
cc_388 N_A_711_21#_c_579_n N_A_560_425#_c_689_n 0.0214268f $X=3.67 $Y=1.535
+ $X2=0 $Y2=0
cc_389 N_A_711_21#_c_590_n N_A_560_425#_c_689_n 0.00487525f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_390 N_A_711_21#_c_582_n N_A_560_425#_c_689_n 0.015171f $X=4.46 $Y=1.505 $X2=0
+ $Y2=0
cc_391 N_A_711_21#_c_583_n N_A_560_425#_c_689_n 0.00621352f $X=4.36 $Y=0.38
+ $X2=0 $Y2=0
cc_392 N_A_711_21#_c_593_n N_A_560_425#_c_689_n 0.00995575f $X=4.345 $Y=1.685
+ $X2=0 $Y2=0
cc_393 N_A_711_21#_c_608_p N_A_560_425#_c_689_n 6.98066e-19 $X=4.965 $Y=1.685
+ $X2=0 $Y2=0
cc_394 N_A_711_21#_c_582_n N_A_560_425#_c_690_n 0.00454653f $X=4.46 $Y=1.505
+ $X2=0 $Y2=0
cc_395 N_A_711_21#_M1018_g N_A_560_425#_c_704_n 0.00189122f $X=3.81 $Y=2.275
+ $X2=0 $Y2=0
cc_396 N_A_711_21#_c_580_n N_A_560_425#_c_699_n 0.00430566f $X=3.65 $Y=0.755
+ $X2=0 $Y2=0
cc_397 N_A_711_21#_c_579_n N_A_560_425#_c_691_n 0.00230689f $X=3.67 $Y=1.535
+ $X2=0 $Y2=0
cc_398 N_A_711_21#_c_580_n N_A_560_425#_c_691_n 0.0055153f $X=3.65 $Y=0.755
+ $X2=0 $Y2=0
cc_399 N_A_711_21#_c_581_n N_A_560_425#_c_691_n 0.00706322f $X=3.65 $Y=0.905
+ $X2=0 $Y2=0
cc_400 N_A_711_21#_c_583_n N_A_560_425#_c_691_n 0.00568369f $X=4.36 $Y=0.38
+ $X2=0 $Y2=0
cc_401 N_A_711_21#_c_579_n N_A_560_425#_c_697_n 0.0108849f $X=3.67 $Y=1.535
+ $X2=0 $Y2=0
cc_402 N_A_711_21#_M1018_g N_A_560_425#_c_697_n 0.00753204f $X=3.81 $Y=2.275
+ $X2=0 $Y2=0
cc_403 N_A_711_21#_c_590_n N_A_560_425#_c_697_n 0.00982227f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_404 N_A_711_21#_c_593_n N_A_560_425#_c_697_n 0.0228437f $X=4.345 $Y=1.685
+ $X2=0 $Y2=0
cc_405 N_A_711_21#_c_579_n N_A_560_425#_c_692_n 0.0175017f $X=3.67 $Y=1.535
+ $X2=0 $Y2=0
cc_406 N_A_711_21#_c_590_n N_A_560_425#_c_692_n 0.00663133f $X=3.9 $Y=1.7 $X2=0
+ $Y2=0
cc_407 N_A_711_21#_c_582_n N_A_560_425#_c_692_n 0.0255753f $X=4.46 $Y=1.505
+ $X2=0 $Y2=0
cc_408 N_A_711_21#_c_593_n N_A_560_425#_c_692_n 0.02399f $X=4.345 $Y=1.685 $X2=0
+ $Y2=0
cc_409 N_A_711_21#_c_579_n N_A_560_425#_c_693_n 0.00534127f $X=3.67 $Y=1.535
+ $X2=0 $Y2=0
cc_410 N_A_711_21#_c_581_n N_A_560_425#_c_693_n 5.27848e-19 $X=3.65 $Y=0.905
+ $X2=0 $Y2=0
cc_411 N_A_711_21#_M1011_g N_RESET_B_M1013_g 0.0234306f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_412 N_A_711_21#_c_582_n N_RESET_B_M1013_g 6.26375e-19 $X=4.46 $Y=1.505 $X2=0
+ $Y2=0
cc_413 N_A_711_21#_c_634_p N_RESET_B_M1013_g 0.0173865f $X=5.245 $Y=1.62 $X2=0
+ $Y2=0
cc_414 N_A_711_21#_c_592_n N_RESET_B_M1013_g 0.00209445f $X=5.355 $Y=1.505 $X2=0
+ $Y2=0
cc_415 N_A_711_21#_c_583_n RESET_B 0.0372853f $X=4.36 $Y=0.38 $X2=0 $Y2=0
cc_416 N_A_711_21#_c_582_n N_RESET_B_c_775_n 2.99764e-19 $X=4.46 $Y=1.505 $X2=0
+ $Y2=0
cc_417 N_A_711_21#_c_608_p N_RESET_B_c_775_n 7.33678e-19 $X=4.965 $Y=1.685 $X2=0
+ $Y2=0
cc_418 N_A_711_21#_c_584_n N_RESET_B_c_775_n 0.00209445f $X=5.47 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A_711_21#_c_585_n N_RESET_B_c_775_n 0.0201765f $X=5.47 $Y=1.16 $X2=0
+ $Y2=0
cc_420 N_A_711_21#_c_582_n N_RESET_B_c_776_n 0.0372853f $X=4.46 $Y=1.505 $X2=0
+ $Y2=0
cc_421 N_A_711_21#_c_608_p N_RESET_B_c_776_n 0.0233751f $X=4.965 $Y=1.685 $X2=0
+ $Y2=0
cc_422 N_A_711_21#_c_584_n N_RESET_B_c_776_n 0.0259849f $X=5.47 $Y=1.16 $X2=0
+ $Y2=0
cc_423 N_A_711_21#_c_585_n N_RESET_B_c_776_n 3.1902e-19 $X=5.47 $Y=1.16 $X2=0
+ $Y2=0
cc_424 N_A_711_21#_c_583_n N_RESET_B_c_777_n 3.54928e-19 $X=4.36 $Y=0.38 $X2=0
+ $Y2=0
cc_425 N_A_711_21#_c_586_n N_RESET_B_c_777_n 0.0190282f $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_426 N_A_711_21#_c_582_n N_VPWR_M1018_d 6.19838e-19 $X=4.46 $Y=1.505 $X2=0
+ $Y2=0
cc_427 N_A_711_21#_c_593_n N_VPWR_M1018_d 0.00385407f $X=4.345 $Y=1.685 $X2=0
+ $Y2=0
cc_428 N_A_711_21#_c_608_p N_VPWR_M1018_d 0.00201186f $X=4.965 $Y=1.685 $X2=0
+ $Y2=0
cc_429 N_A_711_21#_c_634_p N_VPWR_M1013_d 0.00463173f $X=5.245 $Y=1.62 $X2=0
+ $Y2=0
cc_430 N_A_711_21#_c_592_n N_VPWR_M1013_d 2.61593e-19 $X=5.355 $Y=1.505 $X2=0
+ $Y2=0
cc_431 N_A_711_21#_M1011_g N_VPWR_c_813_n 0.0123636f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_432 N_A_711_21#_c_634_p N_VPWR_c_813_n 0.0187231f $X=5.245 $Y=1.62 $X2=0
+ $Y2=0
cc_433 N_A_711_21#_c_585_n N_VPWR_c_813_n 2.60485e-19 $X=5.47 $Y=1.16 $X2=0
+ $Y2=0
cc_434 N_A_711_21#_M1018_g N_VPWR_c_814_n 0.00349295f $X=3.81 $Y=2.275 $X2=0
+ $Y2=0
cc_435 N_A_711_21#_c_590_n N_VPWR_c_814_n 0.00224307f $X=3.9 $Y=1.7 $X2=0 $Y2=0
cc_436 N_A_711_21#_c_593_n N_VPWR_c_814_n 0.0282685f $X=4.345 $Y=1.685 $X2=0
+ $Y2=0
cc_437 N_A_711_21#_M1018_g N_VPWR_c_815_n 0.00585385f $X=3.81 $Y=2.275 $X2=0
+ $Y2=0
cc_438 N_A_711_21#_c_607_p N_VPWR_c_818_n 0.0167204f $X=4.795 $Y=1.685 $X2=0
+ $Y2=0
cc_439 N_A_711_21#_M1011_g N_VPWR_c_819_n 0.0046653f $X=5.51 $Y=1.985 $X2=0
+ $Y2=0
cc_440 N_A_711_21#_M1002_d N_VPWR_c_810_n 0.00300681f $X=4.645 $Y=1.485 $X2=0
+ $Y2=0
cc_441 N_A_711_21#_M1018_g N_VPWR_c_810_n 0.00959149f $X=3.81 $Y=2.275 $X2=0
+ $Y2=0
cc_442 N_A_711_21#_M1011_g N_VPWR_c_810_n 0.008846f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_443 N_A_711_21#_c_590_n N_VPWR_c_810_n 0.00377972f $X=3.9 $Y=1.7 $X2=0 $Y2=0
cc_444 N_A_711_21#_c_593_n N_VPWR_c_810_n 0.00549701f $X=4.345 $Y=1.685 $X2=0
+ $Y2=0
cc_445 N_A_711_21#_c_607_p N_VPWR_c_810_n 0.0126629f $X=4.795 $Y=1.685 $X2=0
+ $Y2=0
cc_446 N_A_711_21#_c_608_p N_VPWR_c_810_n 0.00560351f $X=4.965 $Y=1.685 $X2=0
+ $Y2=0
cc_447 N_A_711_21#_M1011_g N_Q_c_906_n 0.00665753f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_448 N_A_711_21#_c_634_p N_Q_c_906_n 0.00930834f $X=5.245 $Y=1.62 $X2=0 $Y2=0
cc_449 N_A_711_21#_c_592_n N_Q_c_906_n 0.00947655f $X=5.355 $Y=1.505 $X2=0 $Y2=0
cc_450 N_A_711_21#_c_584_n N_Q_c_906_n 0.0246821f $X=5.47 $Y=1.16 $X2=0 $Y2=0
cc_451 N_A_711_21#_c_585_n N_Q_c_906_n 0.00753248f $X=5.47 $Y=1.16 $X2=0 $Y2=0
cc_452 N_A_711_21#_c_586_n N_Q_c_906_n 0.00828285f $X=5.47 $Y=0.995 $X2=0 $Y2=0
cc_453 N_A_711_21#_c_580_n N_VGND_c_924_n 0.00479349f $X=3.65 $Y=0.755 $X2=0
+ $Y2=0
cc_454 N_A_711_21#_c_583_n N_VGND_c_924_n 0.0261199f $X=4.36 $Y=0.38 $X2=0 $Y2=0
cc_455 N_A_711_21#_c_584_n N_VGND_c_925_n 0.0100737f $X=5.47 $Y=1.16 $X2=0 $Y2=0
cc_456 N_A_711_21#_c_585_n N_VGND_c_925_n 5.23568e-19 $X=5.47 $Y=1.16 $X2=0
+ $Y2=0
cc_457 N_A_711_21#_c_586_n N_VGND_c_925_n 0.013132f $X=5.47 $Y=0.995 $X2=0 $Y2=0
cc_458 N_A_711_21#_c_580_n N_VGND_c_928_n 0.00544232f $X=3.65 $Y=0.755 $X2=0
+ $Y2=0
cc_459 N_A_711_21#_c_581_n N_VGND_c_928_n 8.03613e-19 $X=3.65 $Y=0.905 $X2=0
+ $Y2=0
cc_460 N_A_711_21#_c_583_n N_VGND_c_929_n 0.0192809f $X=4.36 $Y=0.38 $X2=0 $Y2=0
cc_461 N_A_711_21#_c_586_n N_VGND_c_930_n 0.00564095f $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_462 N_A_711_21#_M1005_s N_VGND_c_931_n 0.00211564f $X=4.235 $Y=0.235 $X2=0
+ $Y2=0
cc_463 N_A_711_21#_c_580_n N_VGND_c_931_n 0.011038f $X=3.65 $Y=0.755 $X2=0 $Y2=0
cc_464 N_A_711_21#_c_581_n N_VGND_c_931_n 0.00106884f $X=3.65 $Y=0.905 $X2=0
+ $Y2=0
cc_465 N_A_711_21#_c_583_n N_VGND_c_931_n 0.0137814f $X=4.36 $Y=0.38 $X2=0 $Y2=0
cc_466 N_A_711_21#_c_586_n N_VGND_c_931_n 0.0104943f $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_467 N_A_560_425#_M1002_g N_RESET_B_M1013_g 0.0182457f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_468 N_A_560_425#_c_688_n RESET_B 0.00349673f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_469 N_A_560_425#_c_690_n N_RESET_B_c_775_n 0.0215735f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_470 N_A_560_425#_c_690_n N_RESET_B_c_776_n 0.00349673f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_471 N_A_560_425#_c_688_n N_RESET_B_c_777_n 0.0273635f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_560_425#_M1002_g N_VPWR_c_814_n 0.00345853f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_A_560_425#_c_704_n N_VPWR_c_815_n 0.0382318f $X=3.455 $Y=2.34 $X2=0
+ $Y2=0
cc_474 N_A_560_425#_M1002_g N_VPWR_c_818_n 0.00557327f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_475 N_A_560_425#_M1004_d N_VPWR_c_810_n 0.00247452f $X=2.8 $Y=2.125 $X2=0
+ $Y2=0
cc_476 N_A_560_425#_M1002_g N_VPWR_c_810_n 0.00693619f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_477 N_A_560_425#_c_704_n N_VPWR_c_810_n 0.0220242f $X=3.455 $Y=2.34 $X2=0
+ $Y2=0
cc_478 N_A_560_425#_c_704_n A_664_425# 0.00854179f $X=3.455 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_479 N_A_560_425#_c_697_n A_664_425# 0.00479513f $X=3.54 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_480 N_A_560_425#_c_699_n N_VGND_c_923_n 0.00218059f $X=3.415 $Y=0.45 $X2=0
+ $Y2=0
cc_481 N_A_560_425#_c_688_n N_VGND_c_924_n 0.00295484f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_482 N_A_560_425#_c_689_n N_VGND_c_924_n 0.00140505f $X=4.495 $Y=1.16 $X2=0
+ $Y2=0
cc_483 N_A_560_425#_c_692_n N_VGND_c_924_n 0.0126251f $X=4.09 $Y=1.16 $X2=0
+ $Y2=0
cc_484 N_A_560_425#_c_699_n N_VGND_c_928_n 0.0251685f $X=3.415 $Y=0.45 $X2=0
+ $Y2=0
cc_485 N_A_560_425#_c_688_n N_VGND_c_929_n 0.00469794f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_486 N_A_560_425#_M1007_d N_VGND_c_931_n 0.00237979f $X=2.84 $Y=0.235 $X2=0
+ $Y2=0
cc_487 N_A_560_425#_c_688_n N_VGND_c_931_n 0.00935885f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_A_560_425#_c_699_n N_VGND_c_931_n 0.025963f $X=3.415 $Y=0.45 $X2=0
+ $Y2=0
cc_489 N_A_560_425#_c_699_n A_654_47# 0.00535195f $X=3.415 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_490 N_A_560_425#_c_691_n A_654_47# 0.00135873f $X=3.5 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_491 N_RESET_B_M1013_g N_VPWR_c_813_n 0.00317431f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_492 N_RESET_B_M1013_g N_VPWR_c_818_n 0.00585385f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_493 N_RESET_B_M1013_g N_VPWR_c_810_n 0.0108095f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_494 N_RESET_B_c_777_n N_VGND_c_925_n 0.00358678f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_495 RESET_B N_VGND_c_929_n 0.00894018f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_496 N_RESET_B_c_777_n N_VGND_c_929_n 0.00585385f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_497 RESET_B N_VGND_c_931_n 0.00836812f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_498 N_RESET_B_c_777_n N_VGND_c_931_n 0.01094f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_499 RESET_B A_929_47# 0.0107617f $X=4.745 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_500 N_VPWR_c_810_n A_465_369# 0.00469617f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_501 N_VPWR_c_810_n A_664_425# 0.00473588f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_502 N_VPWR_c_810_n N_Q_M1011_d 0.00383158f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_503 N_VPWR_c_819_n Q 0.0169196f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_504 N_VPWR_c_810_n Q 0.00988906f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_505 Q N_VGND_c_930_n 0.0118336f $X=5.665 $Y=0.425 $X2=0 $Y2=0
cc_506 N_Q_M1017_d N_VGND_c_931_n 0.00308051f $X=5.585 $Y=0.235 $X2=0 $Y2=0
cc_507 Q N_VGND_c_931_n 0.0103153f $X=5.665 $Y=0.425 $X2=0 $Y2=0
cc_508 N_VGND_c_931_n A_465_47# 0.0130138f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_509 N_VGND_c_931_n A_654_47# 0.00242128f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_510 N_VGND_c_931_n A_929_47# 0.00622284f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24

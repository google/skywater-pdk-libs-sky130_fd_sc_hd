* File: sky130_fd_sc_hd__or4bb_1.pex.spice
* Created: Tue Sep  1 19:28:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4BB_1%C_N 3 7 8 9 13 14 15
c32 14 0 3.16902e-20 $X=0.51 $Y=1.16
c33 3 0 1.33412e-19 $X=0.47 $Y=2.26
r34 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r35 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r37 8 9 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.6 $Y=1.19 $X2=0.6
+ $Y2=1.53
r38 8 14 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.6 $Y=1.19 $X2=0.6
+ $Y2=1.16
r39 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=0.675
+ $X2=0.505 $Y2=0.995
r40 3 16 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.47 $Y=2.26
+ $X2=0.47 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%D_N 3 6 8 11 13
r37 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.16
+ $X2=1.03 $Y2=1.325
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.16
+ $X2=1.03 $Y2=0.995
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.16 $X2=1.03 $Y2=1.16
r40 8 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.03
+ $Y2=1.16
r41 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.955 $Y=1.695
+ $X2=0.955 $Y2=1.325
r42 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.95 $Y=0.675
+ $X2=0.95 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%A_205_93# 1 2 9 13 15 20 22 24 29 34
c71 22 0 1.56139e-19 $X=1.49 $Y=1.525
c72 20 0 1.87829e-19 $X=1.49 $Y=1.075
c73 15 0 1.33412e-19 $X=1.405 $Y=1.61
r74 30 34 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.645 $Y=1.16
+ $X2=1.89 $Y2=1.16
r75 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.16 $X2=1.645 $Y2=1.16
r76 26 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.49 $Y=1.16
+ $X2=1.645 $Y2=1.16
r77 24 25 16.8452 $w=2.39e-07 $l=3.3e-07 $layer=LI1_cond $X=1.16 $Y=0.655
+ $X2=1.49 $Y2=0.655
r78 21 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=1.245
+ $X2=1.49 $Y2=1.16
r79 21 22 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.49 $Y=1.245
+ $X2=1.49 $Y2=1.525
r80 20 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=1.075
+ $X2=1.49 $Y2=1.16
r81 19 25 2.73298 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.49 $Y=0.825
+ $X2=1.49 $Y2=0.655
r82 19 20 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.49 $Y=0.825
+ $X2=1.49 $Y2=1.075
r83 15 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.61
+ $X2=1.49 $Y2=1.525
r84 15 17 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.405 $Y=1.61
+ $X2=1.165 $Y2=1.61
r85 11 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.325
+ $X2=1.89 $Y2=1.16
r86 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.89 $Y=1.325
+ $X2=1.89 $Y2=2.275
r87 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=0.995
+ $X2=1.89 $Y2=1.16
r88 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.89 $Y=0.995 $X2=1.89
+ $Y2=0.445
r89 2 17 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.61
r90 1 24 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.465 $X2=1.16 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%A_27_410# 1 2 9 13 16 19 21 24 25 26 29 30
+ 35 37
c89 30 0 3.12278e-19 $X=2.31 $Y=1.16
r90 32 35 3.84148 $w=3.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.17 $Y=0.637
+ $X2=0.295 $Y2=0.637
r91 30 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.16
+ $X2=2.31 $Y2=1.325
r92 30 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.16
+ $X2=2.31 $Y2=0.995
r93 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.16 $X2=2.31 $Y2=1.16
r94 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.31 $Y=1.415
+ $X2=2.31 $Y2=1.16
r95 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.225 $Y=1.5
+ $X2=2.31 $Y2=1.415
r96 25 26 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.225 $Y=1.5
+ $X2=1.915 $Y2=1.5
r97 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.83 $Y=1.585
+ $X2=1.915 $Y2=1.5
r98 23 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.83 $Y=1.585
+ $X2=1.83 $Y2=1.865
r99 22 37 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.95
+ $X2=0.215 $Y2=1.95
r100 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.745 $Y=1.95
+ $X2=1.83 $Y2=1.865
r101 21 22 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.745 $Y=1.95
+ $X2=0.345 $Y2=1.95
r102 17 37 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=1.95
r103 17 19 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=2.29
r104 16 37 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.17 $Y=1.865
+ $X2=0.215 $Y2=1.95
r105 15 32 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.637
r106 15 16 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.865
r107 13 40 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.37 $Y=1.695
+ $X2=2.37 $Y2=1.325
r108 9 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.325 $Y=0.445
+ $X2=2.325 $Y2=0.995
r109 2 19 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r110 1 35 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.465 $X2=0.295 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%B 4 7 8 9 10 13
c43 13 0 1.28784e-20 $X=2.79 $Y=2.335
r44 13 15 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.79 $Y=2.335
+ $X2=2.79 $Y2=2.2
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=2.335 $X2=2.79 $Y2=2.335
r46 10 14 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.99 $Y=2.29 $X2=2.79
+ $Y2=2.29
r47 8 9 65.3429 $w=1.65e-07 $l=1.5e-07 $layer=POLY_cond $X=2.737 $Y=0.76
+ $X2=2.737 $Y2=0.91
r48 7 8 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.745 $Y=0.445
+ $X2=2.745 $Y2=0.76
r49 4 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.73 $Y=1.695
+ $X2=2.73 $Y2=2.2
r50 4 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.73 $Y=1.695
+ $X2=2.73 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%A 3 7 9 12 13
c42 7 0 1.96413e-19 $X=3.165 $Y=1.695
r43 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.16
+ $X2=3.15 $Y2=1.325
r44 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.16
+ $X2=3.15 $Y2=0.995
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.16 $X2=3.15 $Y2=1.16
r46 9 13 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.99 $Y=1.16 $X2=3.15
+ $Y2=1.16
r47 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.165 $Y=1.695
+ $X2=3.165 $Y2=1.325
r48 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.165 $Y=0.445
+ $X2=3.165 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%A_311_413# 1 2 3 12 15 17 23 26 27 28 29 30
+ 33 35 37 42 43 44 49 50 51 54
c114 49 0 1.14153e-19 $X=3.63 $Y=1.16
c115 42 0 1.06604e-19 $X=3.525 $Y=1.495
c116 29 0 1.96413e-19 $X=2.95 $Y=1.87
c117 26 0 1.28784e-20 $X=2.17 $Y=2.205
r118 50 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=1.16
+ $X2=3.63 $Y2=1.325
r119 50 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=1.16
+ $X2=3.63 $Y2=0.995
r120 49 52 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.577 $Y=1.16
+ $X2=3.577 $Y2=1.325
r121 49 51 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.577 $Y=1.16
+ $X2=3.577 $Y2=0.995
r122 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.63
+ $Y=1.16 $X2=3.63 $Y2=1.16
r123 44 46 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.035 $Y=1.58
+ $X2=3.035 $Y2=1.87
r124 42 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.525 $Y=1.495
+ $X2=3.525 $Y2=1.325
r125 39 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.525 $Y=0.825
+ $X2=3.525 $Y2=0.995
r126 38 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=1.58
+ $X2=3.035 $Y2=1.58
r127 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.44 $Y=1.58
+ $X2=3.525 $Y2=1.495
r128 37 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.44 $Y=1.58
+ $X2=3.12 $Y2=1.58
r129 36 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.74
+ $X2=2.955 $Y2=0.74
r130 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.44 $Y=0.74
+ $X2=3.525 $Y2=0.825
r131 35 36 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.44 $Y=0.74 $X2=3.04
+ $Y2=0.74
r132 31 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0.655
+ $X2=2.955 $Y2=0.74
r133 31 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.955 $Y=0.655
+ $X2=2.955 $Y2=0.47
r134 29 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=1.87
+ $X2=3.035 $Y2=1.87
r135 29 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.95 $Y=1.87
+ $X2=2.255 $Y2=1.87
r136 27 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=0.74
+ $X2=2.955 $Y2=0.74
r137 27 28 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.87 $Y=0.74
+ $X2=2.185 $Y2=0.74
r138 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.17 $Y=1.955
+ $X2=2.255 $Y2=1.87
r139 25 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.17 $Y=1.955
+ $X2=2.17 $Y2=2.205
r140 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.1 $Y=0.655
+ $X2=2.185 $Y2=0.74
r141 21 23 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.1 $Y=0.655
+ $X2=2.1 $Y2=0.47
r142 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=2.29
+ $X2=2.17 $Y2=2.205
r143 17 19 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.085 $Y=2.29
+ $X2=1.68 $Y2=2.29
r144 15 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.655 $Y=1.985
+ $X2=3.655 $Y2=1.325
r145 12 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.655 $Y=0.56
+ $X2=3.655 $Y2=0.995
r146 3 19 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=2.065 $X2=1.68 $Y2=2.29
r147 2 33 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.235 $X2=2.955 $Y2=0.47
r148 1 23 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.235 $X2=2.1 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%VPWR 1 2 9 13 15 17 22 32 33 36 39
c52 2 0 1.06604e-19 $X=3.24 $Y=1.485
r53 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r57 30 39 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.57 $Y=2.72 $X2=3.43
+ $Y2=2.72
r58 30 32 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.57 $Y=2.72
+ $X2=3.91 $Y2=2.72
r59 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r61 26 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 25 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r66 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 22 39 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.29 $Y=2.72 $X2=3.43
+ $Y2=2.72
r68 22 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.29 $Y=2.72 $X2=2.99
+ $Y2=2.72
r69 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r70 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 11 39 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.43 $Y2=2.72
r74 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.43 $Y2=2
r75 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.72
r76 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.29
r77 2 13 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=3.24
+ $Y=1.485 $X2=3.44 $Y2=2
r78 1 9 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=0.545 $Y=2.05
+ $X2=0.68 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%X 1 2 12 14 15 16
r18 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=3.917 $Y=1.632
+ $X2=3.917 $Y2=1.845
r19 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=3.917 $Y=1.632
+ $X2=3.917 $Y2=1.495
r20 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=3.865 $Y=0.587
+ $X2=3.97 $Y2=0.587
r21 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.97 $Y=0.76 $X2=3.97
+ $Y2=0.587
r22 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.97 $Y=0.76
+ $X2=3.97 $Y2=1.495
r23 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=3.73
+ $Y=1.485 $X2=3.865 $Y2=1.845
r24 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.865 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_1%VGND 1 2 3 4 17 21 25 29 31 33 38 43 50 51
+ 54 57 60 63
r71 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r72 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r73 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r75 51 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r76 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r77 48 63 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.4
+ $Y2=0
r78 48 50 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.91
+ $Y2=0
r79 47 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r80 47 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r81 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r82 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.535
+ $Y2=0
r83 44 46 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.99
+ $Y2=0
r84 43 63 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.4
+ $Y2=0
r85 43 46 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=2.99
+ $Y2=0
r86 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r87 42 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r88 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r89 39 57 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.657
+ $Y2=0
r90 39 41 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=2.07
+ $Y2=0
r91 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.535
+ $Y2=0
r92 38 41 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.07
+ $Y2=0
r93 37 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r94 37 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r95 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r96 34 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.74
+ $Y2=0
r97 34 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=1.15
+ $Y2=0
r98 33 57 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=1.47 $Y=0 $X2=1.657
+ $Y2=0
r99 33 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.47 $Y=0 $X2=1.15
+ $Y2=0
r100 31 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r101 27 63 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=0.085 $X2=3.4
+ $Y2=0
r102 27 29 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.4 $Y=0.085
+ $X2=3.4 $Y2=0.4
r103 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0
r104 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0.4
r105 19 57 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.657 $Y=0.085
+ $X2=1.657 $Y2=0
r106 19 21 9.68052 $w=3.73e-07 $l=3.15e-07 $layer=LI1_cond $X=1.657 $Y=0.085
+ $X2=1.657 $Y2=0.4
r107 15 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r108 15 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.66
r109 4 29 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.235 $X2=3.425 $Y2=0.4
r110 3 25 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.235 $X2=2.535 $Y2=0.4
r111 2 21 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.68 $Y2=0.4
r112 1 17 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.465 $X2=0.74 $Y2=0.66
.ends


* File: sky130_fd_sc_hd__mux2_8.spice.pex
* Created: Thu Aug 27 14:27:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX2_8%A_79_21# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 41 43 46 48 50 53 55 57 60 62 64 67 69 78 80 81 82 85 89 91 95 96 97
+ 103 116 118 122
c270 122 0 1.38777e-19 $X=7.585 $Y=0.72
c271 103 0 1.98871e-19 $X=7.585 $Y=0.85
c272 91 0 1.56763e-19 $X=7.5 $Y=0.72
r273 113 114 69.2451 $w=3.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.17
+ $X2=2.99 $Y2=1.17
r274 112 113 69.2451 $w=3.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.17
+ $X2=2.57 $Y2=1.17
r275 111 112 69.2451 $w=3.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.73 $Y=1.17
+ $X2=2.15 $Y2=1.17
r276 110 111 69.2451 $w=3.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.17
+ $X2=1.73 $Y2=1.17
r277 106 108 69.2451 $w=3.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.17
+ $X2=0.89 $Y2=1.17
r278 104 122 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.585 $Y=0.85
+ $X2=7.585 $Y2=0.72
r279 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.585 $Y=0.85
+ $X2=7.585 $Y2=0.85
r280 100 118 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.835 $Y=0.85
+ $X2=4.835 $Y2=0.72
r281 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.835 $Y=0.85
+ $X2=4.835 $Y2=0.85
r282 97 99 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.98 $Y=0.85
+ $X2=4.835 $Y2=0.85
r283 96 103 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.44 $Y=0.85
+ $X2=7.585 $Y2=0.85
r284 96 97 3.04455 $w=1.4e-07 $l=2.46e-06 $layer=MET1_cond $X=7.44 $Y=0.85
+ $X2=4.98 $Y2=0.85
r285 91 122 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.72
+ $X2=7.585 $Y2=0.72
r286 91 93 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.5 $Y=0.72
+ $X2=7.28 $Y2=0.72
r287 87 89 178.759 $w=1.68e-07 $l=2.74e-06 $layer=LI1_cond $X=5.32 $Y=1.92
+ $X2=8.06 $Y2=1.92
r288 85 87 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=3.625 $Y=1.92
+ $X2=5.32 $Y2=1.92
r289 82 84 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.625 $Y=0.72
+ $X2=4.54 $Y2=0.72
r290 81 118 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0.72
+ $X2=4.835 $Y2=0.72
r291 81 84 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.75 $Y=0.72
+ $X2=4.54 $Y2=0.72
r292 80 85 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.54 $Y=1.835
+ $X2=3.625 $Y2=1.92
r293 79 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=1.245
+ $X2=3.54 $Y2=1.16
r294 79 80 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.54 $Y=1.245
+ $X2=3.54 $Y2=1.835
r295 78 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=1.075
+ $X2=3.54 $Y2=1.16
r296 77 82 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.54 $Y=0.805
+ $X2=3.625 $Y2=0.72
r297 77 78 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.54 $Y=0.805
+ $X2=3.54 $Y2=1.075
r298 76 116 36.2712 $w=3.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.19 $Y=1.17
+ $X2=3.41 $Y2=1.17
r299 76 114 32.9738 $w=3.5e-07 $l=2e-07 $layer=POLY_cond $X=3.19 $Y=1.17
+ $X2=2.99 $Y2=1.17
r300 75 76 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.19
+ $Y=1.16 $X2=3.19 $Y2=1.16
r301 72 110 26.3791 $w=3.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.15 $Y=1.17
+ $X2=1.31 $Y2=1.17
r302 72 108 42.866 $w=3.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.15 $Y=1.17
+ $X2=0.89 $Y2=1.17
r303 71 75 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=3.19 $Y2=1.16
r304 71 72 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=1.15
+ $Y=1.16 $X2=1.15 $Y2=1.16
r305 69 95 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=1.16
+ $X2=3.54 $Y2=1.16
r306 69 75 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.455 $Y=1.16
+ $X2=3.19 $Y2=1.16
r307 65 116 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.41 $Y=1.345
+ $X2=3.41 $Y2=1.17
r308 65 67 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.41 $Y=1.345
+ $X2=3.41 $Y2=1.985
r309 62 116 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.17
r310 62 64 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r311 58 114 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.99 $Y=1.345
+ $X2=2.99 $Y2=1.17
r312 58 60 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.99 $Y=1.345
+ $X2=2.99 $Y2=1.985
r313 55 114 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.17
r314 55 57 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r315 51 113 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.57 $Y=1.345
+ $X2=2.57 $Y2=1.17
r316 51 53 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.57 $Y=1.345
+ $X2=2.57 $Y2=1.985
r317 48 113 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.17
r318 48 50 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r319 44 112 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.15 $Y=1.345
+ $X2=2.15 $Y2=1.17
r320 44 46 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.15 $Y=1.345
+ $X2=2.15 $Y2=1.985
r321 41 112 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.17
r322 41 43 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
r323 37 111 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.73 $Y=1.345
+ $X2=1.73 $Y2=1.17
r324 37 39 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.73 $Y=1.345
+ $X2=1.73 $Y2=1.985
r325 34 111 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.17
r326 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r327 30 110 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.31 $Y=1.345
+ $X2=1.31 $Y2=1.17
r328 30 32 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.31 $Y=1.345
+ $X2=1.31 $Y2=1.985
r329 27 110 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.17
r330 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r331 23 108 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.89 $Y=1.345
+ $X2=0.89 $Y2=1.17
r332 23 25 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.89 $Y=1.345
+ $X2=0.89 $Y2=1.985
r333 20 108 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.17
r334 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r335 16 106 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.47 $Y=1.345
+ $X2=0.47 $Y2=1.17
r336 16 18 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.47 $Y=1.345
+ $X2=0.47 $Y2=1.985
r337 13 106 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.17
r338 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r339 4 89 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=7.925
+ $Y=1.485 $X2=8.06 $Y2=1.92
r340 3 87 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.485 $X2=5.32 $Y2=1.92
r341 2 93 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.235 $X2=7.28 $Y2=0.72
r342 1 84 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.235 $X2=4.54 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%S 3 6 8 10 13 17 20 24 25 27 28 29 31 32 34
+ 35 40 43 47 48 49
c160 35 0 1.61023e-19 $X=5.9 $Y=1.53
c161 31 0 1.53743e-19 $X=5.95 $Y=1.16
c162 27 0 1.93859e-19 $X=5.67 $Y=1.58
c163 24 0 1.36597e-19 $X=3.88 $Y=1.16
r164 48 54 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=9.362 $Y=1.16
+ $X2=9.362 $Y2=1.53
r165 47 50 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=9.275 $Y=1.16
+ $X2=9.275 $Y2=1.325
r166 47 49 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=9.275 $Y=1.16
+ $X2=9.275 $Y2=0.995
r167 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.3
+ $Y=1.16 $X2=9.3 $Y2=1.16
r168 40 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.425 $Y=1.53
+ $X2=9.425 $Y2=1.53
r169 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.755 $Y=1.53
+ $X2=5.755 $Y2=1.53
r170 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.9 $Y=1.53
+ $X2=5.755 $Y2=1.53
r171 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.28 $Y=1.53
+ $X2=9.425 $Y2=1.53
r172 34 35 4.18316 $w=1.4e-07 $l=3.38e-06 $layer=MET1_cond $X=9.28 $Y=1.53
+ $X2=5.9 $Y2=1.53
r173 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.16 $X2=5.95 $Y2=1.16
r174 29 38 2.56795 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.852 $Y=1.495
+ $X2=5.852 $Y2=1.58
r175 29 31 10.5772 $w=3.63e-07 $l=3.35e-07 $layer=LI1_cond $X=5.852 $Y=1.495
+ $X2=5.852 $Y2=1.16
r176 27 38 5.49844 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=5.67 $Y=1.58
+ $X2=5.852 $Y2=1.58
r177 27 28 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=5.67 $Y=1.58
+ $X2=3.965 $Y2=1.58
r178 25 44 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.882 $Y=1.16
+ $X2=3.882 $Y2=1.325
r179 25 43 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.882 $Y=1.16
+ $X2=3.882 $Y2=0.995
r180 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r181 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.88 $Y=1.495
+ $X2=3.965 $Y2=1.58
r182 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.88 $Y=1.495
+ $X2=3.88 $Y2=1.16
r183 20 50 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.19 $Y=1.985
+ $X2=9.19 $Y2=1.325
r184 17 49 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.19 $Y=0.56
+ $X2=9.19 $Y2=0.995
r185 11 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.325
+ $X2=5.95 $Y2=1.16
r186 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.95 $Y=1.325
+ $X2=5.95 $Y2=1.985
r187 8 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=0.995
+ $X2=5.95 $Y2=1.16
r188 8 10 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=5.95 $Y=0.995
+ $X2=5.95 $Y2=0.555
r189 6 44 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.885 $Y=1.985
+ $X2=3.885 $Y2=1.325
r190 3 43 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.885 $Y=0.555
+ $X2=3.885 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%A1 1 3 4 6 7 9 10 12 13 14 19 25 33 36
c92 14 0 1.83894e-19 $X=4.52 $Y=1.19
r93 31 33 14.7414 $w=4.15e-07 $l=1.1e-07 $layer=POLY_cond $X=8.16 $Y=1.202
+ $X2=8.27 $Y2=1.202
r94 31 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.16
+ $Y=1.16 $X2=8.16 $Y2=1.16
r95 28 31 41.544 $w=4.15e-07 $l=3.1e-07 $layer=POLY_cond $X=7.85 $Y=1.202
+ $X2=8.16 $Y2=1.202
r96 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.39
+ $Y=1.16 $X2=4.39 $Y2=1.16
r97 19 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.045 $Y=1.19
+ $X2=8.045 $Y2=1.19
r98 16 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.375 $Y=1.19
+ $X2=4.375 $Y2=1.19
r99 14 16 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.52 $Y=1.19
+ $X2=4.375 $Y2=1.19
r100 13 19 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.9 $Y=1.19
+ $X2=8.045 $Y2=1.19
r101 13 14 4.18316 $w=1.4e-07 $l=3.38e-06 $layer=MET1_cond $X=7.9 $Y=1.19
+ $X2=4.52 $Y2=1.19
r102 10 33 26.7644 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.27 $Y=1.41
+ $X2=8.27 $Y2=1.202
r103 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.27 $Y=1.41
+ $X2=8.27 $Y2=1.985
r104 7 28 26.7644 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.85 $Y=1.41
+ $X2=7.85 $Y2=1.202
r105 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.85 $Y=1.41
+ $X2=7.85 $Y2=1.985
r106 4 24 56.9138 $w=3.65e-07 $l=3.6e-07 $layer=POLY_cond $X=4.75 $Y=1.142
+ $X2=4.39 $Y2=1.142
r107 4 6 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.75 $Y=0.96 $X2=4.75
+ $Y2=0.555
r108 1 24 9.48563 $w=3.65e-07 $l=6e-08 $layer=POLY_cond $X=4.33 $Y=1.142
+ $X2=4.39 $Y2=1.142
r109 1 3 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.33 $Y=0.96 $X2=4.33
+ $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%A0 1 3 4 6 7 9 10 12 15 18 21 22 23 26 27 33
+ 38 41 43
c118 18 0 1.38777e-19 $X=6.725 $Y=0.73
c119 7 0 1.98871e-19 $X=7.07 $Y=0.96
r120 38 41 1.77299 $w=3.88e-07 $l=6e-08 $layer=LI1_cond $X=5.695 $Y=0.62
+ $X2=5.755 $Y2=0.62
r121 27 43 7.36653 $w=3.88e-07 $l=1.23e-07 $layer=LI1_cond $X=5.767 $Y=0.62
+ $X2=5.89 $Y2=0.62
r122 27 41 0.354598 $w=3.88e-07 $l=1.2e-08 $layer=LI1_cond $X=5.767 $Y=0.62
+ $X2=5.755 $Y2=0.62
r123 27 38 0.384148 $w=3.88e-07 $l=1.3e-08 $layer=LI1_cond $X=5.682 $Y=0.62
+ $X2=5.695 $Y2=0.62
r124 26 37 50.4573 $w=3.63e-07 $l=3.8e-07 $layer=POLY_cond $X=7.11 $Y=1.142
+ $X2=7.49 $Y2=1.142
r125 26 35 5.31129 $w=3.63e-07 $l=4e-08 $layer=POLY_cond $X=7.11 $Y=1.142
+ $X2=7.07 $Y2=1.142
r126 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.11
+ $Y=1.16 $X2=7.11 $Y2=1.16
r127 23 25 16.1233 $w=2.27e-07 $l=3e-07 $layer=LI1_cond $X=6.81 $Y=1.16 $X2=7.11
+ $Y2=1.16
r128 22 27 9.81054 $w=3.88e-07 $l=3.32e-07 $layer=LI1_cond $X=5.35 $Y=0.62
+ $X2=5.682 $Y2=0.62
r129 21 23 2.43258 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.81 $Y=0.995
+ $X2=6.81 $Y2=1.16
r130 20 21 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.81 $Y=0.815
+ $X2=6.81 $Y2=0.995
r131 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.725 $Y=0.73
+ $X2=6.81 $Y2=0.815
r132 18 43 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=6.725 $Y=0.73
+ $X2=5.89 $Y2=0.73
r133 16 33 35.5134 $w=4.15e-07 $l=2.65e-07 $layer=POLY_cond $X=5.265 $Y=1.202
+ $X2=5.53 $Y2=1.202
r134 16 30 20.772 $w=4.15e-07 $l=1.55e-07 $layer=POLY_cond $X=5.265 $Y=1.202
+ $X2=5.11 $Y2=1.202
r135 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.265
+ $Y=1.16 $X2=5.265 $Y2=1.16
r136 13 22 6.17013 $w=3.75e-07 $l=2.33666e-07 $layer=LI1_cond $X=5.265 $Y=0.815
+ $X2=5.35 $Y2=0.62
r137 13 15 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.265 $Y=0.815
+ $X2=5.265 $Y2=1.16
r138 10 37 23.5056 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=7.49 $Y=0.96
+ $X2=7.49 $Y2=1.142
r139 10 12 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=7.49 $Y=0.96
+ $X2=7.49 $Y2=0.555
r140 7 35 23.5056 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=7.07 $Y=0.96
+ $X2=7.07 $Y2=1.142
r141 7 9 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=7.07 $Y=0.96 $X2=7.07
+ $Y2=0.555
r142 4 33 26.7644 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.53 $Y=1.41
+ $X2=5.53 $Y2=1.202
r143 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.53 $Y=1.41
+ $X2=5.53 $Y2=1.985
r144 1 30 26.7644 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.11 $Y=1.41
+ $X2=5.11 $Y2=1.202
r145 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.11 $Y=1.41
+ $X2=5.11 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%A_1259_199# 1 2 9 12 16 19 23 24 26 27 31 32
+ 34 35 36 37 38 41 43 45 47 51 54
c143 51 0 1.56763e-19 $X=6.462 $Y=0.995
c144 31 0 8.18594e-20 $X=8.77 $Y=1.16
c145 23 0 1.04687e-19 $X=6.43 $Y=1.16
r146 43 49 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.4 $Y=2.085
+ $X2=9.4 $Y2=1.94
r147 43 45 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.4 $Y=2.085
+ $X2=9.4 $Y2=2.3
r148 39 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.4 $Y=0.645
+ $X2=9.4 $Y2=0.46
r149 37 49 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.315 $Y=2
+ $X2=9.4 $Y2=1.94
r150 37 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.315 $Y=2
+ $X2=8.855 $Y2=2
r151 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.315 $Y=0.73
+ $X2=9.4 $Y2=0.645
r152 35 36 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.315 $Y=0.73
+ $X2=8.855 $Y2=0.73
r153 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.77 $Y=1.915
+ $X2=8.855 $Y2=2
r154 33 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.77 $Y=1.665
+ $X2=8.77 $Y2=1.58
r155 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.77 $Y=1.665
+ $X2=8.77 $Y2=1.915
r156 32 55 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=1.16
+ $X2=8.76 $Y2=1.325
r157 32 54 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=8.76 $Y=1.16
+ $X2=8.76 $Y2=0.995
r158 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.77
+ $Y=1.16 $X2=8.77 $Y2=1.16
r159 29 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.77 $Y=1.495
+ $X2=8.77 $Y2=1.58
r160 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.77 $Y=1.495
+ $X2=8.77 $Y2=1.16
r161 28 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.77 $Y=0.815
+ $X2=8.855 $Y2=0.73
r162 28 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.77 $Y=0.815
+ $X2=8.77 $Y2=1.16
r163 26 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.685 $Y=1.58
+ $X2=8.77 $Y2=1.58
r164 26 27 141.572 $w=1.68e-07 $l=2.17e-06 $layer=LI1_cond $X=8.685 $Y=1.58
+ $X2=6.515 $Y2=1.58
r165 24 52 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.462 $Y=1.16
+ $X2=6.462 $Y2=1.325
r166 24 51 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.462 $Y=1.16
+ $X2=6.462 $Y2=0.995
r167 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.43
+ $Y=1.16 $X2=6.43 $Y2=1.16
r168 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.43 $Y=1.495
+ $X2=6.515 $Y2=1.58
r169 21 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.43 $Y=1.495
+ $X2=6.43 $Y2=1.16
r170 19 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.69 $Y=1.985
+ $X2=8.69 $Y2=1.325
r171 16 54 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.69 $Y=0.555
+ $X2=8.69 $Y2=0.995
r172 12 52 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.435 $Y=1.985
+ $X2=6.435 $Y2=1.325
r173 9 51 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.435 $Y=0.555
+ $X2=6.435 $Y2=0.995
r174 2 49 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.485 $X2=9.4 $Y2=1.96
r175 2 45 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.485 $X2=9.4 $Y2=2.3
r176 1 41 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=9.265
+ $Y=0.235 $X2=9.4 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48 51
+ 52 54 55 57 58 59 61 76 83 90 91 97 100 103
c133 7 0 8.18594e-20 $X=8.765 $Y=1.485
r134 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r135 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r136 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r137 91 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r138 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r139 88 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=8.98 $Y2=2.72
r140 88 90 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=9.43 $Y2=2.72
r141 87 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r142 87 101 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=6.21 $Y2=2.72
r143 86 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r144 84 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=2.72
+ $X2=6.16 $Y2=2.72
r145 84 86 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=6.245 $Y=2.72
+ $X2=8.51 $Y2=2.72
r146 83 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.815 $Y=2.72
+ $X2=8.98 $Y2=2.72
r147 83 86 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.815 $Y=2.72
+ $X2=8.51 $Y2=2.72
r148 82 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r149 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r150 79 82 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.75 $Y2=2.72
r151 78 81 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.75 $Y2=2.72
r152 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r153 76 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=6.16 $Y2=2.72
r154 76 81 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=5.75 $Y2=2.72
r155 75 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r156 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r157 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r158 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r159 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r160 69 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r161 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r162 66 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.1 $Y2=2.72
r163 66 68 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.61 $Y2=2.72
r164 65 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r165 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r166 62 94 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r167 62 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r168 61 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.1 $Y2=2.72
r169 61 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r170 59 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r171 59 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r172 57 74 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.45 $Y2=2.72
r173 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.62 $Y2=2.72
r174 56 78 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.91 $Y2=2.72
r175 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.62 $Y2=2.72
r176 54 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.53 $Y2=2.72
r177 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.78 $Y2=2.72
r178 53 74 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.45 $Y2=2.72
r179 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.78 $Y2=2.72
r180 51 68 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.61 $Y2=2.72
r181 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.94 $Y2=2.72
r182 50 71 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.53 $Y2=2.72
r183 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=1.94 $Y2=2.72
r184 46 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=2.635
+ $X2=8.98 $Y2=2.72
r185 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.98 $Y=2.635
+ $X2=8.98 $Y2=2.34
r186 42 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.16 $Y=2.635
+ $X2=6.16 $Y2=2.72
r187 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.16 $Y=2.635
+ $X2=6.16 $Y2=2.34
r188 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r189 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.34
r190 34 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r191 34 36 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r192 30 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r193 30 32 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r194 26 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r195 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r196 22 94 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r197 22 24 21.8448 $w=3.33e-07 $l=6.35e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2
r198 7 48 600 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=8.765
+ $Y=1.485 $X2=8.98 $Y2=2.34
r199 6 44 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.025
+ $Y=1.485 $X2=6.16 $Y2=2.34
r200 5 40 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2.34
r201 4 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r202 3 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r203 2 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r204 1 24 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%X 1 2 3 4 5 6 7 8 27 31 33 35 39 43 45 47 51
+ 55 57 59 63 67 70 72 73 74 75 76 77
r88 71 77 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=0.705 $Y=1.575
+ $X2=0.705 $Y2=1.19
r89 71 72 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.575
+ $X2=0.705 $Y2=1.66
r90 69 77 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=0.705 $Y=0.805
+ $X2=0.705 $Y2=1.19
r91 69 70 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.805
+ $X2=0.705 $Y2=0.72
r92 65 67 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.2 $Y=1.745
+ $X2=3.2 $Y2=1.96
r93 61 63 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.2 $Y=0.635
+ $X2=3.2 $Y2=0.46
r94 60 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.66
+ $X2=2.36 $Y2=1.66
r95 59 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.115 $Y=1.66
+ $X2=3.2 $Y2=1.745
r96 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.115 $Y=1.66
+ $X2=2.445 $Y2=1.66
r97 58 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0.72
+ $X2=2.36 $Y2=0.72
r98 57 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.115 $Y=0.72
+ $X2=3.2 $Y2=0.635
r99 57 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.115 $Y=0.72
+ $X2=2.445 $Y2=0.72
r100 53 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=1.745
+ $X2=2.36 $Y2=1.66
r101 53 55 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.36 $Y=1.745
+ $X2=2.36 $Y2=1.96
r102 49 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.635
+ $X2=2.36 $Y2=0.72
r103 49 51 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.36 $Y=0.635
+ $X2=2.36 $Y2=0.42
r104 48 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.66
+ $X2=1.52 $Y2=1.66
r105 47 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=1.66
+ $X2=2.36 $Y2=1.66
r106 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.275 $Y=1.66
+ $X2=1.605 $Y2=1.66
r107 46 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.72
+ $X2=1.52 $Y2=0.72
r108 45 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0.72
+ $X2=2.36 $Y2=0.72
r109 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.275 $Y=0.72
+ $X2=1.605 $Y2=0.72
r110 41 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.745
+ $X2=1.52 $Y2=1.66
r111 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.52 $Y=1.745
+ $X2=1.52 $Y2=1.96
r112 37 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.635
+ $X2=1.52 $Y2=0.72
r113 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.52 $Y=0.635
+ $X2=1.52 $Y2=0.46
r114 36 72 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.815 $Y=1.66
+ $X2=0.705 $Y2=1.66
r115 35 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=1.52 $Y2=1.66
r116 35 36 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=0.815 $Y2=1.66
r117 34 70 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.815 $Y=0.72
+ $X2=0.705 $Y2=0.72
r118 33 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=1.52 $Y2=0.72
r119 33 34 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=0.815 $Y2=0.72
r120 29 72 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=0.68 $Y=1.745
+ $X2=0.705 $Y2=1.66
r121 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=1.745
+ $X2=0.68 $Y2=1.96
r122 25 70 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.705 $Y2=0.72
r123 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.68 $Y2=0.42
r124 8 67 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.96
r125 7 55 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.96
r126 6 43 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r127 5 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
r128 4 63 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.46
r129 3 51 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.42
r130 2 39 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.46
r131 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%A_792_297# 1 2 11
c14 2 0 5.08625e-19 $X=5.605 $Y=1.485
r15 8 11 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=4.12 $Y=2.34 $X2=5.74
+ $Y2=2.34
r16 2 11 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.605
+ $Y=1.485 $X2=5.74 $Y2=2.34
r17 1 8 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.485 $X2=4.12 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%A_1302_297# 1 2 11
r15 8 11 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=6.645 $Y=2.34
+ $X2=8.48 $Y2=2.34
r16 2 11 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.345
+ $Y=1.485 $X2=8.48 $Y2=2.34
r17 1 8 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.51
+ $Y=1.485 $X2=6.645 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48 51
+ 52 54 55 57 58 59 61 76 83 93 94 100 103 106
r151 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r152 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r153 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r154 94 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.97 $Y2=0
r155 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r156 91 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=0
+ $X2=8.98 $Y2=0
r157 91 93 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.145 $Y=0
+ $X2=9.43 $Y2=0
r158 90 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r159 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r160 87 90 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.51 $Y2=0
r161 87 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r162 86 89 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.67 $Y=0 $X2=8.51
+ $Y2=0
r163 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r164 84 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.39 $Y=0
+ $X2=6.225 $Y2=0
r165 84 86 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.39 $Y=0 $X2=6.67
+ $Y2=0
r166 83 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.815 $Y=0
+ $X2=8.98 $Y2=0
r167 83 89 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.815 $Y=0
+ $X2=8.51 $Y2=0
r168 82 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r169 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r170 79 82 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r171 78 81 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.75
+ $Y2=0
r172 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r173 76 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.06 $Y=0
+ $X2=6.225 $Y2=0
r174 76 81 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=5.75
+ $Y2=0
r175 75 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r176 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r177 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r178 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r179 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r180 69 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r181 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r182 66 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r183 66 68 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r184 65 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r185 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r186 62 97 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r187 62 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r188 61 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r189 61 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r190 59 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r191 59 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r192 57 74 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.45
+ $Y2=0
r193 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.62
+ $Y2=0
r194 56 78 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=0
+ $X2=3.91 $Y2=0
r195 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.62
+ $Y2=0
r196 54 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.53
+ $Y2=0
r197 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.78
+ $Y2=0
r198 53 74 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.945 $Y=0
+ $X2=3.45 $Y2=0
r199 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.78
+ $Y2=0
r200 51 68 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.61 $Y2=0
r201 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.94
+ $Y2=0
r202 50 71 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.105 $Y=0
+ $X2=2.53 $Y2=0
r203 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=1.94
+ $Y2=0
r204 46 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=8.98 $Y2=0
r205 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=8.98 $Y2=0.38
r206 42 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.225 $Y2=0
r207 42 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.225 $Y2=0.38
r208 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0
r209 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0.38
r210 34 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r211 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.38
r212 30 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r213 30 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.38
r214 26 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r215 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r216 22 97 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r217 22 24 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r218 7 48 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=8.765
+ $Y=0.235 $X2=8.98 $Y2=0.38
r219 6 44 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=6.025
+ $Y=0.235 $X2=6.225 $Y2=0.38
r220 5 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.38
r221 4 36 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.38
r222 3 32 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r223 2 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r224 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%A_792_47# 1 2 11
r22 8 11 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.12 $Y=0.38 $X2=4.96
+ $Y2=0.38
r23 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.38
r24 1 8 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.96
+ $Y=0.235 $X2=4.12 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_8%A_1302_47# 1 2 11
r21 8 11 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.74 $Y=0.38 $X2=7.7
+ $Y2=0.38
r22 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.565
+ $Y=0.235 $X2=7.7 $Y2=0.38
r23 1 8 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=6.51
+ $Y=0.235 $X2=6.74 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__dfxtp_4.pex.spice
* Created: Tue Sep  1 19:04:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFXTP_4%CLK 1 2 3 5 6 8 11 13 14
c40 1 0 2.71124e-20 $X=0.305 $Y=1.325
r41 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=1.16
+ $X2=0.265 $Y2=1.53
r42 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r43 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r44 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r45 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r46 3 18 88.7086 $w=2.58e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r47 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r48 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r49 1 18 39.2009 $w=2.58e-07 $l=1.75656e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.327 $Y2=1.16
r50 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%A_27_47# 1 2 9 13 17 19 20 25 29 31 35 39 43
+ 44 45 48 50 53 54 55 56 57 64 66 71 74 76 78 82
c214 82 0 1.77381e-19 $X=4.375 $Y=1.41
c215 57 0 1.99186e-19 $X=3.16 $Y=1.87
c216 48 0 1.81794e-19 $X=0.725 $Y=1.795
c217 45 0 3.29888e-20 $X=0.61 $Y=1.88
c218 29 0 4.21632e-20 $X=4.38 $Y=2.275
c219 19 0 1.57835e-19 $X=2.69 $Y=1.32
r220 81 83 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.41
+ $X2=4.375 $Y2=1.575
r221 81 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.375
+ $Y=1.41 $X2=4.375 $Y2=1.41
r222 78 81 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=4.375 $Y=1.32
+ $X2=4.375 $Y2=1.41
r223 74 77 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.74
+ $X2=2.825 $Y2=1.905
r224 74 76 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.74
+ $X2=2.825 $Y2=1.575
r225 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.74 $X2=2.825 $Y2=1.74
r226 67 82 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=4.385 $Y=1.87
+ $X2=4.385 $Y2=1.41
r227 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.395 $Y=1.87
+ $X2=4.395 $Y2=1.87
r228 64 75 6.168 $w=3.53e-07 $l=1.9e-07 $layer=LI1_cond $X=3.015 $Y=1.832
+ $X2=2.825 $Y2=1.832
r229 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.87
+ $X2=3.015 $Y2=1.87
r230 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.87
+ $X2=0.695 $Y2=1.87
r231 57 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.16 $Y=1.87
+ $X2=3.015 $Y2=1.87
r232 56 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.25 $Y=1.87
+ $X2=4.395 $Y2=1.87
r233 56 57 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=4.25 $Y=1.87
+ $X2=3.16 $Y2=1.87
r234 55 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.87
+ $X2=0.695 $Y2=1.87
r235 54 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.87
+ $X2=3.015 $Y2=1.87
r236 54 55 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=2.87 $Y=1.87
+ $X2=0.84 $Y2=1.87
r237 51 71 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r238 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r239 48 60 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r240 48 50 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r241 47 50 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r242 46 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r243 45 60 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r244 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r245 43 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r246 43 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r247 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r248 37 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r249 33 35 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=5.025 $Y=1.245
+ $X2=5.025 $Y2=0.415
r250 32 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.51 $Y=1.32
+ $X2=4.375 $Y2=1.32
r251 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.95 $Y=1.32
+ $X2=5.025 $Y2=1.245
r252 31 32 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.95 $Y=1.32
+ $X2=4.51 $Y2=1.32
r253 29 83 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.38 $Y=2.275
+ $X2=4.38 $Y2=1.575
r254 25 77 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.765 $Y=2.275
+ $X2=2.765 $Y2=1.905
r255 21 76 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.765 $Y=1.395
+ $X2=2.765 $Y2=1.575
r256 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.69 $Y=1.32
+ $X2=2.765 $Y2=1.395
r257 19 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.69 $Y=1.32
+ $X2=2.38 $Y2=1.32
r258 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.305 $Y=1.245
+ $X2=2.38 $Y2=1.32
r259 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.305 $Y=1.245
+ $X2=2.305 $Y2=0.415
r260 11 71 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r261 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r262 7 71 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r263 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r264 2 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r265 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%D 3 7 9 10 17
r40 14 17 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.635 $Y=1.5
+ $X2=1.83 $Y2=1.5
r41 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.5 $X2=1.635 $Y2=1.5
r42 9 10 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.58 $Y=1.19 $X2=1.58
+ $Y2=1.5
r43 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.665
+ $X2=1.83 $Y2=1.5
r44 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.83 $Y=1.665 $X2=1.83
+ $Y2=2.275
r45 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.335
+ $X2=1.83 $Y2=1.5
r46 1 3 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.83 $Y=1.335 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%A_193_47# 1 2 9 13 14 16 19 23 24 27 28 32
+ 33 35 36 37 38 45 47 54 56 61 69
c185 61 0 1.77381e-19 $X=4.605 $Y=0.87
c186 37 0 1.57835e-19 $X=4.25 $Y=0.85
c187 35 0 3.67213e-20 $X=2.41 $Y=0.85
c188 23 0 1.99186e-19 $X=2.315 $Y=1.74
r189 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.605
+ $Y=0.87 $X2=4.605 $Y2=0.87
r190 58 61 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=4.51 $Y=0.87
+ $X2=4.605 $Y2=0.87
r191 54 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=0.87
+ $X2=2.725 $Y2=0.705
r192 48 62 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.395 $Y=0.87
+ $X2=4.605 $Y2=0.87
r193 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.395 $Y=0.85
+ $X2=4.395 $Y2=0.85
r194 45 78 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.555 $Y=0.87
+ $X2=2.35 $Y2=0.87
r195 45 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.725
+ $Y=0.87 $X2=2.725 $Y2=0.87
r196 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=0.85
+ $X2=2.555 $Y2=0.85
r197 41 73 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.96
r198 41 69 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.51
r199 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=0.85
+ $X2=1.155 $Y2=0.85
r200 38 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.7 $Y=0.85
+ $X2=2.555 $Y2=0.85
r201 37 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.25 $Y=0.85
+ $X2=4.395 $Y2=0.85
r202 37 38 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=4.25 $Y=0.85
+ $X2=2.7 $Y2=0.85
r203 36 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=0.85
+ $X2=1.155 $Y2=0.85
r204 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=0.85
+ $X2=2.555 $Y2=0.85
r205 35 36 1.37376 $w=1.4e-07 $l=1.11e-06 $layer=MET1_cond $X=2.41 $Y=0.85
+ $X2=1.3 $Y2=0.85
r206 33 64 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=4.885 $Y=1.74
+ $X2=4.8 $Y2=1.74
r207 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.74 $X2=4.885 $Y2=1.74
r208 29 32 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.745 $Y=1.74
+ $X2=4.885 $Y2=1.74
r209 28 62 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.65 $Y=0.87
+ $X2=4.605 $Y2=0.87
r210 27 29 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=1.575
+ $X2=4.745 $Y2=1.74
r211 26 28 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=4.745 $Y=1.035
+ $X2=4.65 $Y2=0.87
r212 26 27 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=4.745 $Y=1.035
+ $X2=4.745 $Y2=1.575
r213 24 52 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.315 $Y=1.74
+ $X2=2.315 $Y2=1.875
r214 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.315
+ $Y=1.74 $X2=2.315 $Y2=1.74
r215 21 78 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=1.035
+ $X2=2.35 $Y2=0.87
r216 21 23 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=2.35 $Y=1.035
+ $X2=2.35 $Y2=1.74
r217 17 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.8 $Y=1.875
+ $X2=4.8 $Y2=1.74
r218 17 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.8 $Y=1.875 $X2=4.8
+ $Y2=2.275
r219 14 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.51 $Y=0.705
+ $X2=4.51 $Y2=0.87
r220 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.51 $Y=0.705
+ $X2=4.51 $Y2=0.415
r221 13 56 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.785 $Y=0.415
+ $X2=2.785 $Y2=0.705
r222 9 52 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.3 $Y=2.275 $X2=2.3
+ $Y2=1.875
r223 2 73 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r224 1 69 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%A_634_183# 1 2 9 13 15 18 21 23 29 30 32 33
+ 36
r95 35 36 5.54023 $w=2.61e-07 $l=3e-08 $layer=POLY_cond $X=3.245 $Y=0.93
+ $X2=3.275 $Y2=0.93
r96 32 33 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.3
+ $X2=4.075 $Y2=2.135
r97 27 36 24.0077 $w=2.61e-07 $l=1.3e-07 $layer=POLY_cond $X=3.405 $Y=0.93
+ $X2=3.275 $Y2=0.93
r98 26 29 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=0.93
+ $X2=3.49 $Y2=0.93
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.405
+ $Y=0.93 $X2=3.405 $Y2=0.93
r100 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.12 $Y=0.45
+ $X2=4.245 $Y2=0.45
r101 19 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.035 $Y=1.065
+ $X2=4.035 $Y2=0.915
r102 19 33 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.035 $Y=1.065
+ $X2=4.035 $Y2=2.135
r103 18 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.035 $Y=0.765
+ $X2=4.035 $Y2=0.915
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.035 $Y=0.535
+ $X2=4.12 $Y2=0.45
r105 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.035 $Y=0.535
+ $X2=4.035 $Y2=0.765
r106 15 30 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=0.915
+ $X2=4.035 $Y2=0.915
r107 15 29 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.95 $Y=0.915
+ $X2=3.49 $Y2=0.915
r108 11 36 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.275 $Y=0.795
+ $X2=3.275 $Y2=0.93
r109 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.275 $Y=0.795
+ $X2=3.275 $Y2=0.445
r110 7 35 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.245 $Y=1.065
+ $X2=3.245 $Y2=0.93
r111 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=3.245 $Y=1.065
+ $X2=3.245 $Y2=2.275
r112 2 32 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.735 $X2=4.115 $Y2=2.3
r113 1 23 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=4.08
+ $Y=0.235 $X2=4.245 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%A_475_413# 1 2 8 11 13 15 18 20 21 22 26 31
+ 33 35
c109 31 0 1.42307e-19 $X=3.065 $Y=1.315
c110 26 0 3.67213e-20 $X=2.98 $Y=0.45
r111 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.41 $X2=3.695 $Y2=1.41
r112 35 37 17.1405 $w=2.42e-07 $l=3.4e-07 $layer=LI1_cond $X=3.355 $Y=1.41
+ $X2=3.695 $Y2=1.41
r113 32 35 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=1.575
+ $X2=3.355 $Y2=1.41
r114 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.355 $Y=1.575
+ $X2=3.355 $Y2=2.19
r115 31 35 14.6198 $w=2.42e-07 $l=2.9e-07 $layer=LI1_cond $X=3.065 $Y=1.41
+ $X2=3.355 $Y2=1.41
r116 30 31 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.065 $Y=0.535
+ $X2=3.065 $Y2=1.315
r117 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.98 $Y=0.45
+ $X2=3.065 $Y2=0.535
r118 26 28 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.98 $Y=0.45
+ $X2=2.565 $Y2=0.45
r119 22 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=2.275
+ $X2=3.355 $Y2=2.19
r120 22 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.27 $Y=2.275
+ $X2=2.535 $Y2=2.275
r121 20 38 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.41
+ $X2=3.695 $Y2=1.41
r122 20 21 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.83 $Y=1.41
+ $X2=3.905 $Y2=1.41
r123 16 18 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.905 $Y=1.025
+ $X2=4.005 $Y2=1.025
r124 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.005 $Y=0.95
+ $X2=4.005 $Y2=1.025
r125 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.005 $Y=0.95
+ $X2=4.005 $Y2=0.555
r126 9 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.905 $Y=1.545
+ $X2=3.905 $Y2=1.41
r127 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.905 $Y=1.545
+ $X2=3.905 $Y2=2.11
r128 8 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.905 $Y=1.275
+ $X2=3.905 $Y2=1.41
r129 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.905 $Y=1.1
+ $X2=3.905 $Y2=1.025
r130 7 8 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.905 $Y=1.1
+ $X2=3.905 $Y2=1.275
r131 2 24 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=2.065 $X2=2.535 $Y2=2.275
r132 1 28 182 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.565 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%A_1062_300# 1 2 9 13 15 17 20 22 24 27 29 31
+ 34 36 38 41 43 46 50 52 53 55 61 67 69 81
c137 81 0 7.79397e-20 $X=8.215 $Y=1.16
r138 78 79 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=7.36 $Y=1.16
+ $X2=7.795 $Y2=1.16
r139 70 72 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.385 $Y=1.665
+ $X2=5.5 $Y2=1.665
r140 67 68 13.0342 $w=2.34e-07 $l=2.5e-07 $layer=LI1_cond $X=6.255 $Y=1.665
+ $X2=6.505 $Y2=1.665
r141 62 81 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=8.075 $Y=1.16
+ $X2=8.215 $Y2=1.16
r142 62 79 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=8.075 $Y=1.16
+ $X2=7.795 $Y2=1.16
r143 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.075
+ $Y=1.16 $X2=8.075 $Y2=1.16
r144 59 78 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=7.055 $Y=1.16
+ $X2=7.36 $Y2=1.16
r145 59 75 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.055 $Y=1.16
+ $X2=6.94 $Y2=1.16
r146 58 61 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.055 $Y=1.16
+ $X2=8.075 $Y2=1.16
r147 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.055
+ $Y=1.16 $X2=7.055 $Y2=1.16
r148 56 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=1.16
+ $X2=6.505 $Y2=1.16
r149 56 58 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.59 $Y=1.16
+ $X2=7.055 $Y2=1.16
r150 55 68 2.60974 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=1.5
+ $X2=6.505 $Y2=1.665
r151 54 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=1.245
+ $X2=6.505 $Y2=1.16
r152 54 55 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.505 $Y=1.245
+ $X2=6.505 $Y2=1.5
r153 53 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=1.075
+ $X2=6.505 $Y2=1.16
r154 52 65 19.699 $w=3.99e-07 $l=5.86728e-07 $layer=LI1_cond $X=6.505 $Y=0.905
+ $X2=6.34 $Y2=0.395
r155 52 53 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.505 $Y=0.905
+ $X2=6.505 $Y2=1.075
r156 48 67 2.60974 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=1.83
+ $X2=6.255 $Y2=1.665
r157 48 50 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.255 $Y=1.83
+ $X2=6.255 $Y2=1.95
r158 46 72 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=5.565 $Y=1.665
+ $X2=5.5 $Y2=1.665
r159 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.565
+ $Y=1.665 $X2=5.565 $Y2=1.665
r160 43 67 4.19144 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=1.665
+ $X2=6.255 $Y2=1.665
r161 43 45 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=6.17 $Y=1.665
+ $X2=5.565 $Y2=1.665
r162 39 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.215 $Y=1.325
+ $X2=8.215 $Y2=1.16
r163 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.215 $Y=1.325
+ $X2=8.215 $Y2=1.985
r164 36 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.215 $Y=0.995
+ $X2=8.215 $Y2=1.16
r165 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.215 $Y=0.995
+ $X2=8.215 $Y2=0.56
r166 32 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.795 $Y=1.325
+ $X2=7.795 $Y2=1.16
r167 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.795 $Y=1.325
+ $X2=7.795 $Y2=1.985
r168 29 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.795 $Y=0.995
+ $X2=7.795 $Y2=1.16
r169 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.795 $Y=0.995
+ $X2=7.795 $Y2=0.56
r170 25 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.36 $Y=1.325
+ $X2=7.36 $Y2=1.16
r171 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.36 $Y=1.325
+ $X2=7.36 $Y2=1.985
r172 22 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.36 $Y=0.995
+ $X2=7.36 $Y2=1.16
r173 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.36 $Y=0.995
+ $X2=7.36 $Y2=0.56
r174 18 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.325
+ $X2=6.94 $Y2=1.16
r175 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.94 $Y=1.325
+ $X2=6.94 $Y2=1.985
r176 15 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=0.995
+ $X2=6.94 $Y2=1.16
r177 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.94 $Y=0.995
+ $X2=6.94 $Y2=0.56
r178 11 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.5 $X2=5.5
+ $Y2=1.665
r179 11 13 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=5.5 $Y=1.5
+ $X2=5.5 $Y2=0.445
r180 7 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.83
+ $X2=5.385 $Y2=1.665
r181 7 9 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.385 $Y=1.83
+ $X2=5.385 $Y2=2.275
r182 2 67 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.11
+ $Y=1.485 $X2=6.255 $Y2=1.61
r183 2 50 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=6.11
+ $Y=1.485 $X2=6.255 $Y2=1.95
r184 1 65 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=6.13
+ $Y=0.235 $X2=6.255 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%A_891_413# 1 2 7 9 12 14 15 16 20 25 27 30
+ 33
c81 30 0 7.79397e-20 $X=6.065 $Y=1.16
c82 27 0 4.21632e-20 $X=5.225 $Y=2.165
c83 12 0 1.7303e-19 $X=6.465 $Y=1.985
c84 7 0 1.8116e-19 $X=6.465 $Y=0.995
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.16 $X2=6.065 $Y2=1.16
r86 28 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=1.16
+ $X2=5.225 $Y2=1.16
r87 28 30 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.31 $Y=1.16
+ $X2=6.065 $Y2=1.16
r88 26 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=1.245
+ $X2=5.225 $Y2=1.16
r89 26 27 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.225 $Y=1.245
+ $X2=5.225 $Y2=2.165
r90 25 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=1.075
+ $X2=5.225 $Y2=1.16
r91 24 25 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.225 $Y=0.535
+ $X2=5.225 $Y2=1.075
r92 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=0.45
+ $X2=5.225 $Y2=0.535
r93 20 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.14 $Y=0.45
+ $X2=4.805 $Y2=0.45
r94 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=2.25
+ $X2=5.225 $Y2=2.165
r95 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.14 $Y=2.25
+ $X2=4.59 $Y2=2.25
r96 14 31 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=6.39 $Y=1.16
+ $X2=6.065 $Y2=1.16
r97 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.39 $Y=1.16
+ $X2=6.465 $Y2=1.16
r98 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=1.325
+ $X2=6.465 $Y2=1.16
r99 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.465 $Y=1.325
+ $X2=6.465 $Y2=1.985
r100 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=0.995
+ $X2=6.465 $Y2=1.16
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.465 $Y=0.995
+ $X2=6.465 $Y2=0.56
r102 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=2.065 $X2=4.59 $Y2=2.25
r103 1 22 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.235 $X2=4.805 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 51 52 54 55 57 58 59 61 66 84 92 97 100 103 107
c134 107 0 1.81794e-19 $X=8.51 $Y=2.72
c135 1 0 3.29888e-20 $X=0.545 $Y=1.815
r136 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r137 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r138 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r139 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r140 95 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r141 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r142 92 106 3.40825 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=8.34 $Y=2.72 $X2=8.54
+ $Y2=2.72
r143 92 94 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.34 $Y=2.72
+ $X2=8.05 $Y2=2.72
r144 91 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r145 91 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r146 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r147 88 103 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=6.715 $Y2=2.72
r148 88 90 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=7.13 $Y2=2.72
r149 87 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r150 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r151 84 103 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.625 $Y=2.72
+ $X2=6.715 $Y2=2.72
r152 84 86 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=6.625 $Y=2.72
+ $X2=5.75 $Y2=2.72
r153 83 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r155 80 83 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r156 79 82 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r157 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r158 77 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r159 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r160 74 77 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r161 74 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r162 73 76 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r163 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r164 71 100 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.572 $Y2=2.72
r165 71 73 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=2.07 $Y2=2.72
r166 70 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r167 70 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r168 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r169 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r170 67 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r171 66 100 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.572 $Y2=2.72
r172 66 69 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.15 $Y2=2.72
r173 61 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r174 61 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r175 59 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r176 59 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r177 57 90 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.5 $Y=2.72 $X2=7.13
+ $Y2=2.72
r178 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=2.72
+ $X2=7.585 $Y2=2.72
r179 56 94 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.67 $Y=2.72
+ $X2=8.05 $Y2=2.72
r180 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=2.72
+ $X2=7.585 $Y2=2.72
r181 54 82 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.49 $Y=2.72 $X2=5.29
+ $Y2=2.72
r182 54 55 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.49 $Y=2.72
+ $X2=5.597 $Y2=2.72
r183 53 86 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=5.75 $Y2=2.72
r184 53 55 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=5.597 $Y2=2.72
r185 51 76 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r186 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.695 $Y2=2.72
r187 50 79 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.91 $Y2=2.72
r188 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.695 $Y2=2.72
r189 46 106 3.40825 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=8.425 $Y=2.635
+ $X2=8.54 $Y2=2.72
r190 46 48 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.425 $Y=2.635
+ $X2=8.425 $Y2=1.97
r191 42 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=2.635
+ $X2=7.585 $Y2=2.72
r192 42 44 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.585 $Y=2.635
+ $X2=7.585 $Y2=1.97
r193 38 103 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=2.635
+ $X2=6.715 $Y2=2.72
r194 38 40 37.8939 $w=1.78e-07 $l=6.15e-07 $layer=LI1_cond $X=6.715 $Y=2.635
+ $X2=6.715 $Y2=2.02
r195 34 55 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.597 $Y=2.635
+ $X2=5.597 $Y2=2.72
r196 34 36 17.9567 $w=2.13e-07 $l=3.35e-07 $layer=LI1_cond $X=5.597 $Y=2.635
+ $X2=5.597 $Y2=2.3
r197 30 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2.72
r198 30 32 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2
r199 26 100 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.572 $Y=2.635
+ $X2=1.572 $Y2=2.72
r200 26 28 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.572 $Y=2.635
+ $X2=1.572 $Y2=2.34
r201 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r202 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r203 7 48 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=8.29
+ $Y=1.485 $X2=8.425 $Y2=1.97
r204 6 44 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=7.435
+ $Y=1.485 $X2=7.585 $Y2=1.97
r205 5 40 300 $w=1.7e-07 $l=6.14146e-07 $layer=licon1_PDIFF $count=2 $X=6.54
+ $Y=1.485 $X2=6.71 $Y2=2.02
r206 4 36 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=2.065 $X2=5.595 $Y2=2.3
r207 3 32 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=3.32
+ $Y=2.065 $X2=3.695 $Y2=2
r208 2 28 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.065 $X2=1.62 $Y2=2.34
r209 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%A_381_47# 1 2 11 14 15
r30 14 15 11.1996 $w=2.33e-07 $l=2.1e-07 $layer=LI1_cond $X=2.007 $Y=2.275
+ $X2=2.007 $Y2=2.065
r31 7 11 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.535
+ $X2=1.975 $Y2=0.45
r32 7 15 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=1.975 $Y=0.535
+ $X2=1.975 $Y2=2.065
r33 2 14 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.065 $X2=2.04 $Y2=2.275
r34 1 11 182 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.055 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%Q 1 2 3 4 13 14 15 19 23 25 27 30 32 35 37
+ 38 39 40 45
c87 32 0 1.7303e-19 $X=7.152 $Y=1.635
c88 14 0 1.8116e-19 $X=7.32 $Y=0.815
r89 40 54 3.44013 $w=3.33e-07 $l=1e-07 $layer=LI1_cond $X=7.152 $Y=2.21
+ $X2=7.152 $Y2=2.31
r90 39 40 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=7.152 $Y=1.87
+ $X2=7.152 $Y2=2.21
r91 38 45 3.95615 $w=3.33e-07 $l=1.15e-07 $layer=LI1_cond $X=7.152 $Y=0.51
+ $X2=7.152 $Y2=0.395
r92 32 39 8.0843 $w=3.33e-07 $l=2.35e-07 $layer=LI1_cond $X=7.152 $Y=1.635
+ $X2=7.152 $Y2=1.87
r93 32 34 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.152 $Y=1.635
+ $X2=7.152 $Y2=1.55
r94 31 38 7.56828 $w=3.33e-07 $l=2.2e-07 $layer=LI1_cond $X=7.152 $Y=0.73
+ $X2=7.152 $Y2=0.51
r95 29 30 26.5767 $w=2.43e-07 $l=5.65e-07 $layer=LI1_cond $X=8.532 $Y=0.9
+ $X2=8.532 $Y2=1.465
r96 28 35 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.175 $Y=0.815
+ $X2=8.007 $Y2=0.815
r97 27 29 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=8.41 $Y=0.815
+ $X2=8.532 $Y2=0.9
r98 27 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.41 $Y=0.815
+ $X2=8.175 $Y2=0.815
r99 26 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.17 $Y=1.55
+ $X2=8.005 $Y2=1.55
r100 25 30 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=8.41 $Y=1.55
+ $X2=8.532 $Y2=1.465
r101 25 26 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.41 $Y=1.55
+ $X2=8.17 $Y2=1.55
r102 21 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=1.635
+ $X2=8.005 $Y2=1.55
r103 21 23 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.005 $Y=1.635
+ $X2=8.005 $Y2=2.31
r104 17 35 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.007 $Y=0.73
+ $X2=8.007 $Y2=0.815
r105 17 19 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=8.007 $Y=0.73
+ $X2=8.007 $Y2=0.395
r106 16 34 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.32 $Y=1.55
+ $X2=7.152 $Y2=1.55
r107 15 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=1.55
+ $X2=8.005 $Y2=1.55
r108 15 16 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.84 $Y=1.55
+ $X2=7.32 $Y2=1.55
r109 14 31 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=7.32 $Y=0.815
+ $X2=7.152 $Y2=0.73
r110 13 35 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.84 $Y=0.815
+ $X2=8.007 $Y2=0.815
r111 13 14 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.84 $Y=0.815
+ $X2=7.32 $Y2=0.815
r112 4 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.87
+ $Y=1.485 $X2=8.005 $Y2=1.63
r113 4 23 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=7.87
+ $Y=1.485 $X2=8.005 $Y2=2.31
r114 3 54 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=7.015
+ $Y=1.485 $X2=7.15 $Y2=2.31
r115 3 34 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.015
+ $Y=1.485 $X2=7.15 $Y2=1.63
r116 2 19 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=7.87
+ $Y=0.235 $X2=8.005 $Y2=0.395
r117 1 45 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=7.015
+ $Y=0.235 $X2=7.15 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_4%VGND 1 2 3 4 5 6 7 24 28 32 36 38 42 46 48
+ 50 53 54 55 57 62 67 72 84 89 92 95 98 101 105
c140 105 0 2.71124e-20 $X=8.51 $Y=0
r141 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r142 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r143 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r144 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r145 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r146 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r147 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r148 87 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r149 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r150 84 104 3.40825 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=8.345 $Y=0
+ $X2=8.542 $Y2=0
r151 84 86 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.345 $Y=0 $X2=8.05
+ $Y2=0
r152 83 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r153 83 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.67 $Y2=0
r154 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r155 80 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=0 $X2=6.71
+ $Y2=0
r156 80 82 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.795 $Y=0
+ $X2=7.13 $Y2=0
r157 79 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r158 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r159 76 79 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r160 76 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r161 75 78 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r162 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r163 73 95 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.77 $Y=0 $X2=3.585
+ $Y2=0
r164 73 75 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.77 $Y=0 $X2=3.91
+ $Y2=0
r165 72 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=0 $X2=5.71
+ $Y2=0
r166 72 78 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.625 $Y=0
+ $X2=5.29 $Y2=0
r167 71 96 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r168 71 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r169 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r170 68 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.58
+ $Y2=0
r171 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r172 67 95 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.585
+ $Y2=0
r173 67 70 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.4 $Y=0 $X2=2.07
+ $Y2=0
r174 66 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r175 66 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r176 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r177 63 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r178 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r179 62 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.58
+ $Y2=0
r180 62 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r181 57 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r182 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r183 55 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r184 55 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r185 53 82 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.495 $Y=0
+ $X2=7.13 $Y2=0
r186 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=0 $X2=7.58
+ $Y2=0
r187 52 86 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=8.05 $Y2=0
r188 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.58
+ $Y2=0
r189 48 104 3.40825 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.542 $Y2=0
r190 48 50 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0.395
r191 44 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.58 $Y=0.085
+ $X2=7.58 $Y2=0
r192 44 46 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.58 $Y=0.085
+ $X2=7.58 $Y2=0.395
r193 40 101 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.71 $Y=0.085
+ $X2=6.71 $Y2=0
r194 40 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.71 $Y=0.085
+ $X2=6.71 $Y2=0.4
r195 39 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.71
+ $Y2=0
r196 38 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.625 $Y=0 $X2=6.71
+ $Y2=0
r197 38 39 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.625 $Y=0
+ $X2=5.795 $Y2=0
r198 34 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=0.085
+ $X2=5.71 $Y2=0
r199 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.71 $Y=0.085
+ $X2=5.71 $Y2=0.45
r200 30 95 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0
r201 30 32 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0.42
r202 26 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r203 26 28 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.38
r204 22 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r205 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r206 7 50 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=8.29
+ $Y=0.235 $X2=8.43 $Y2=0.395
r207 6 46 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=7.435
+ $Y=0.235 $X2=7.58 $Y2=0.395
r208 5 42 182 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_NDIFF $count=1 $X=6.54
+ $Y=0.235 $X2=6.71 $Y2=0.4
r209 4 36 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.45
r210 3 32 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.235 $X2=3.655 $Y2=0.42
r211 2 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r212 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__clkdlybuf4s25_2.spice.SKY130_FD_SC_HD__CLKDLYBUF4S25_2.pxi
* Created: Thu Aug 27 14:11:53 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A N_A_M1003_g N_A_M1004_g A A N_A_c_67_n
+ N_A_c_68_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_27_47# N_A_27_47#_M1003_s
+ N_A_27_47#_M1004_s N_A_27_47#_M1007_g N_A_27_47#_M1006_g N_A_27_47#_c_99_n
+ N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_118_n N_A_27_47#_c_107_n
+ N_A_27_47#_c_108_n N_A_27_47#_c_102_n N_A_27_47#_c_103_n N_A_27_47#_c_104_n
+ N_A_27_47#_c_105_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_225_47# N_A_225_47#_M1007_d
+ N_A_225_47#_M1006_d N_A_225_47#_c_168_n N_A_225_47#_M1008_g
+ N_A_225_47#_M1001_g N_A_225_47#_c_169_n N_A_225_47#_c_170_n
+ N_A_225_47#_c_177_n N_A_225_47#_c_171_n N_A_225_47#_c_172_n
+ N_A_225_47#_c_173_n N_A_225_47#_c_174_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_225_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_331_47# N_A_331_47#_M1008_s
+ N_A_331_47#_M1001_s N_A_331_47#_M1000_g N_A_331_47#_M1002_g
+ N_A_331_47#_M1009_g N_A_331_47#_M1005_g N_A_331_47#_c_231_n
+ N_A_331_47#_c_246_n N_A_331_47#_c_248_n N_A_331_47#_c_232_n
+ N_A_331_47#_c_237_n N_A_331_47#_c_238_n N_A_331_47#_c_233_n
+ N_A_331_47#_c_234_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%A_331_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%VPWR N_VPWR_M1004_d N_VPWR_M1001_d
+ N_VPWR_M1005_s N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n
+ N_VPWR_c_323_n N_VPWR_c_324_n VPWR N_VPWR_c_325_n N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_318_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%X N_X_M1000_d N_X_M1002_d X X X X X
+ N_X_c_383_n X N_X_c_384_n N_X_c_370_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%VGND N_VGND_M1003_d N_VGND_M1008_d
+ N_VGND_M1009_s N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n N_VGND_c_406_n
+ N_VGND_c_407_n N_VGND_c_408_n VGND N_VGND_c_409_n N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_2%VGND
cc_1 VNB N_A_M1003_g 0.036043f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_c_67_n 0.0325554f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_3 VNB N_A_c_68_n 0.013431f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_4 VNB N_A_27_47#_c_99_n 0.0128214f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=0.97
cc_5 VNB N_A_27_47#_c_100_n 0.0029073f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.19
cc_6 VNB N_A_27_47#_c_101_n 0.0096254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_102_n 0.00238172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_103_n 0.0214347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_104_n 0.00182687f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_105_n 0.0257105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_225_47#_c_168_n 0.0264834f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_12 VNB N_A_225_47#_c_169_n 0.00348322f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.16
cc_13 VNB N_A_225_47#_c_170_n 0.00245472f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.19
cc_14 VNB N_A_225_47#_c_171_n 0.00353577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_225_47#_c_172_n 0.00193376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_225_47#_c_173_n 0.0509187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_225_47#_c_174_n 0.00146857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_331_47#_M1000_g 0.0279888f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_A_331_47#_M1009_g 0.0355782f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.325
cc_20 VNB N_A_331_47#_c_231_n 0.00366043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_331_47#_c_232_n 0.00178379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_331_47#_c_233_n 0.00298931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_331_47#_c_234_n 0.0481066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_318_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 0.00111827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0423317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_403_n 0.00280434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_404_n 0.00280434f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=0.97
cc_29 VNB N_VGND_c_405_n 0.0112316f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.16
cc_30 VNB N_VGND_c_406_n 0.0198232f $X=-0.19 $Y=-0.24 $X2=0.29 $Y2=1.19
cc_31 VNB N_VGND_c_407_n 0.0298131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_408_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_409_n 0.0173049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_410_n 0.021954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_411_n 0.00507198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_412_n 0.207965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_A_M1004_g 0.0238795f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_38 VPB N_A_c_67_n 0.00679192f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_39 VPB N_A_c_68_n 0.0128004f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_40 VPB N_A_27_47#_M1006_g 0.039776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_107_n 9.45936e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_108_n 0.0268938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_103_n 0.00298939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_225_47#_M1001_g 0.0429225f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_45 VPB N_A_225_47#_c_170_n 0.00519831f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.19
cc_46 VPB N_A_225_47#_c_177_n 0.0110201f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.53
cc_47 VPB N_A_225_47#_c_173_n 0.0222854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_331_47#_M1002_g 0.0186006f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_49 VPB N_A_331_47#_M1005_g 0.0250069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_331_47#_c_237_n 0.00269492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_331_47#_c_238_n 0.00303714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_331_47#_c_233_n 0.00174287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_331_47#_c_234_n 0.0138402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_319_n 0.00280434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_320_n 0.00280434f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=0.97
cc_56 VPB N_VPWR_c_321_n 0.0112323f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.16
cc_57 VPB N_VPWR_c_322_n 0.04241f $X=-0.19 $Y=1.305 $X2=0.29 $Y2=1.19
cc_58 VPB N_VPWR_c_323_n 0.0321033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_324_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_325_n 0.0181078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_326_n 0.0223178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_327_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_318_n 0.052879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_370_n 0.00104789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 N_A_c_68_n N_A_27_47#_M1004_s 0.00281283f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_A_27_47#_M1006_g 0.0329299f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_c_68_n N_A_27_47#_M1006_g 2.48091e-19 $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_M1003_g N_A_27_47#_c_100_n 0.0146023f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_69 N_A_c_67_n N_A_27_47#_c_100_n 0.00127344f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_c_68_n N_A_27_47#_c_100_n 0.0106928f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_67_n N_A_27_47#_c_101_n 0.00298745f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_68_n N_A_27_47#_c_101_n 0.0208544f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_A_27_47#_c_118_n 0.0112456f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_c_68_n N_A_27_47#_c_118_n 0.00707115f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_A_27_47#_c_107_n 0.00732996f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_c_68_n N_A_27_47#_c_107_n 0.00278139f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_67_n N_A_27_47#_c_108_n 5.20243e-19 $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_c_68_n N_A_27_47#_c_108_n 0.0223481f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_c_67_n N_A_27_47#_c_102_n 0.00278914f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_68_n N_A_27_47#_c_102_n 0.0470569f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_c_67_n N_A_27_47#_c_103_n 0.0151418f $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_c_68_n N_A_27_47#_c_103_n 2.96489e-19 $X=0.355 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1003_g N_A_27_47#_c_104_n 0.00278914f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_M1003_g N_A_27_47#_c_105_n 0.0185918f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_A_225_47#_c_169_n 5.23262e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_VPWR_c_319_n 0.00320833f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_VPWR_c_325_n 0.00585385f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_VPWR_c_318_n 0.00703811f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VGND_c_403_n 0.00310635f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_M1003_g N_VGND_c_409_n 0.00425831f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_M1003_g N_VGND_c_412_n 0.00681303f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_105_n N_A_225_47#_c_169_n 0.00827634f $X=0.97 $Y=0.995 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_M1006_g N_A_225_47#_c_170_n 0.00326975f $X=1 $Y=2.075 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_107_n N_A_225_47#_c_170_n 0.0171718f $X=0.835 $Y=1.58 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_102_n N_A_225_47#_c_170_n 0.0280463f $X=0.95 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_c_103_n N_A_225_47#_c_170_n 0.00502327f $X=0.95 $Y=1.16 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_M1006_g N_A_225_47#_c_177_n 0.00482969f $X=1 $Y=2.075 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_c_107_n N_A_225_47#_c_177_n 0.0115538f $X=0.835 $Y=1.58 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_104_n N_A_225_47#_c_171_n 0.00651507f $X=0.85 $Y=0.995 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_105_n N_A_225_47#_c_171_n 0.0056534f $X=0.97 $Y=0.995 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_102_n N_A_225_47#_c_173_n 2.66978e-19 $X=0.95 $Y=1.16 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_103_n N_A_225_47#_c_173_n 0.0162828f $X=0.95 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_c_105_n N_A_225_47#_c_174_n 0.00547644f $X=0.97 $Y=0.995 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_105_n N_A_331_47#_c_231_n 7.4634e-19 $X=0.97 $Y=0.995 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_105_n N_A_331_47#_c_232_n 4.35046e-19 $X=0.97 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_118_n N_VPWR_M1004_d 0.00276884f $X=0.665 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_27_47#_c_107_n N_VPWR_M1004_d 0.00496541f $X=0.835 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_27_47#_M1006_g N_VPWR_c_319_n 0.0121164f $X=1 $Y=2.075 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_118_n N_VPWR_c_319_n 0.00455011f $X=0.665 $Y=1.87 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_c_107_n N_VPWR_c_319_n 0.0146125f $X=0.835 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A_27_47#_M1006_g N_VPWR_c_323_n 0.00856787f $X=1 $Y=2.075 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_108_n N_VPWR_c_325_n 0.0174583f $X=0.26 $Y=1.95 $X2=0 $Y2=0
cc_113 N_A_27_47#_M1004_s N_VPWR_c_318_n 0.00242687f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_M1006_g N_VPWR_c_318_n 0.0153846f $X=1 $Y=2.075 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_118_n N_VPWR_c_318_n 0.00753875f $X=0.665 $Y=1.87 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_107_n N_VPWR_c_318_n 6.86822e-19 $X=0.835 $Y=1.58 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_108_n N_VPWR_c_318_n 0.00954569f $X=0.26 $Y=1.95 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_100_n N_VGND_M1003_d 0.00448114f $X=0.665 $Y=0.725 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_27_47#_c_104_n N_VGND_M1003_d 8.53742e-19 $X=0.85 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_27_47#_c_100_n N_VGND_c_403_n 0.0173136f $X=0.665 $Y=0.725 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_102_n N_VGND_c_403_n 0.00152417f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_105_n N_VGND_c_403_n 0.0103613f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_105_n N_VGND_c_407_n 0.00812762f $X=0.97 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_c_99_n N_VGND_c_409_n 0.01293f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_100_n N_VGND_c_409_n 0.00318265f $X=0.665 $Y=0.725 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_M1003_s N_VGND_c_412_n 0.0023646f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_99_n N_VGND_c_412_n 0.00922327f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_100_n N_VGND_c_412_n 0.00694484f $X=0.665 $Y=0.725 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_105_n N_VGND_c_412_n 0.0144398f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_225_47#_c_168_n N_A_331_47#_M1000_g 0.0203508f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_A_225_47#_c_168_n N_A_331_47#_c_231_n 0.00798921f $X=2.04 $Y=0.995
+ $X2=0 $Y2=0
cc_132 N_A_225_47#_c_169_n N_A_331_47#_c_231_n 0.0291839f $X=1.26 $Y=0.515 $X2=0
+ $Y2=0
cc_133 N_A_225_47#_M1001_g N_A_331_47#_c_246_n 0.0148514f $X=2.04 $Y=2.075 $X2=0
+ $Y2=0
cc_134 N_A_225_47#_c_177_n N_A_331_47#_c_246_n 0.0423844f $X=1.26 $Y=1.81 $X2=0
+ $Y2=0
cc_135 N_A_225_47#_c_168_n N_A_331_47#_c_248_n 0.0135859f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_136 N_A_225_47#_c_172_n N_A_331_47#_c_248_n 0.0143404f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_225_47#_c_168_n N_A_331_47#_c_232_n 0.00434319f $X=2.04 $Y=0.995
+ $X2=0 $Y2=0
cc_138 N_A_225_47#_c_172_n N_A_331_47#_c_232_n 0.0222562f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_225_47#_c_173_n N_A_331_47#_c_232_n 0.00666716f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_225_47#_c_174_n N_A_331_47#_c_232_n 0.0138061f $X=1.26 $Y=0.78 $X2=0
+ $Y2=0
cc_141 N_A_225_47#_M1001_g N_A_331_47#_c_237_n 0.0204964f $X=2.04 $Y=2.075 $X2=0
+ $Y2=0
cc_142 N_A_225_47#_c_172_n N_A_331_47#_c_237_n 0.0157354f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_225_47#_M1001_g N_A_331_47#_c_238_n 0.00420324f $X=2.04 $Y=2.075
+ $X2=0 $Y2=0
cc_144 N_A_225_47#_c_170_n N_A_331_47#_c_238_n 0.00374992f $X=1.307 $Y=1.557
+ $X2=0 $Y2=0
cc_145 N_A_225_47#_c_177_n N_A_331_47#_c_238_n 0.0121469f $X=1.26 $Y=1.81 $X2=0
+ $Y2=0
cc_146 N_A_225_47#_c_172_n N_A_331_47#_c_238_n 0.0204549f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A_225_47#_c_173_n N_A_331_47#_c_238_n 0.00509237f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_148 N_A_225_47#_c_168_n N_A_331_47#_c_233_n 0.00444625f $X=2.04 $Y=0.995
+ $X2=0 $Y2=0
cc_149 N_A_225_47#_c_172_n N_A_331_47#_c_233_n 0.0270383f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_225_47#_c_173_n N_A_331_47#_c_233_n 0.0051228f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_225_47#_M1001_g N_A_331_47#_c_234_n 0.0225406f $X=2.04 $Y=2.075 $X2=0
+ $Y2=0
cc_152 N_A_225_47#_c_172_n N_A_331_47#_c_234_n 3.71531e-19 $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_153 N_A_225_47#_c_173_n N_A_331_47#_c_234_n 0.0215873f $X=2.03 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A_225_47#_M1001_g N_VPWR_c_320_n 0.0159008f $X=2.04 $Y=2.075 $X2=0
+ $Y2=0
cc_155 N_A_225_47#_M1001_g N_VPWR_c_323_n 0.00812762f $X=2.04 $Y=2.075 $X2=0
+ $Y2=0
cc_156 N_A_225_47#_c_177_n N_VPWR_c_323_n 0.0183595f $X=1.26 $Y=1.81 $X2=0 $Y2=0
cc_157 N_A_225_47#_M1006_d N_VPWR_c_318_n 0.00382897f $X=1.125 $Y=1.665 $X2=0
+ $Y2=0
cc_158 N_A_225_47#_M1001_g N_VPWR_c_318_n 0.014349f $X=2.04 $Y=2.075 $X2=0 $Y2=0
cc_159 N_A_225_47#_c_177_n N_VPWR_c_318_n 0.0101286f $X=1.26 $Y=1.81 $X2=0 $Y2=0
cc_160 N_A_225_47#_c_169_n N_VGND_c_403_n 0.0147592f $X=1.26 $Y=0.515 $X2=0
+ $Y2=0
cc_161 N_A_225_47#_c_168_n N_VGND_c_404_n 0.00992549f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_225_47#_c_168_n N_VGND_c_407_n 0.00610796f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_225_47#_c_169_n N_VGND_c_407_n 0.0210041f $X=1.26 $Y=0.515 $X2=0
+ $Y2=0
cc_164 N_A_225_47#_M1007_d N_VGND_c_412_n 0.00210122f $X=1.125 $Y=0.235 $X2=0
+ $Y2=0
cc_165 N_A_225_47#_c_168_n N_VGND_c_412_n 0.0080195f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_225_47#_c_169_n N_VGND_c_412_n 0.0124714f $X=1.26 $Y=0.515 $X2=0
+ $Y2=0
cc_167 N_A_331_47#_c_237_n N_VPWR_M1001_d 0.00602621f $X=2.335 $Y=1.622 $X2=0
+ $Y2=0
cc_168 N_A_331_47#_M1002_g N_VPWR_c_320_n 0.00310635f $X=2.565 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_331_47#_c_246_n N_VPWR_c_320_n 0.0369697f $X=1.78 $Y=1.81 $X2=0 $Y2=0
cc_170 N_A_331_47#_c_237_n N_VPWR_c_320_n 0.0204017f $X=2.335 $Y=1.622 $X2=0
+ $Y2=0
cc_171 N_A_331_47#_c_234_n N_VPWR_c_320_n 2.56721e-19 $X=3.065 $Y=1.162 $X2=0
+ $Y2=0
cc_172 N_A_331_47#_M1005_g N_VPWR_c_322_n 0.0218563f $X=3.065 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_331_47#_c_246_n N_VPWR_c_323_n 0.0153589f $X=1.78 $Y=1.81 $X2=0 $Y2=0
cc_174 N_A_331_47#_M1002_g N_VPWR_c_326_n 0.00585385f $X=2.565 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_331_47#_M1005_g N_VPWR_c_326_n 0.00428227f $X=3.065 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_331_47#_M1001_s N_VPWR_c_318_n 0.00351653f $X=1.655 $Y=1.665 $X2=0
+ $Y2=0
cc_177 N_A_331_47#_M1002_g N_VPWR_c_318_n 0.010912f $X=2.565 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_331_47#_M1005_g N_VPWR_c_318_n 0.00823263f $X=3.065 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_331_47#_c_246_n N_VPWR_c_318_n 0.00934584f $X=1.78 $Y=1.81 $X2=0
+ $Y2=0
cc_180 N_A_331_47#_M1000_g X 0.00129929f $X=2.565 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A_331_47#_M1009_g X 0.00850082f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_182 N_A_331_47#_c_248_n X 0.00746791f $X=2.335 $Y=0.72 $X2=0 $Y2=0
cc_183 N_A_331_47#_M1002_g X 0.0101063f $X=2.565 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_331_47#_M1005_g X 0.00291891f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_331_47#_c_237_n X 0.00965697f $X=2.335 $Y=1.622 $X2=0 $Y2=0
cc_186 N_A_331_47#_c_234_n X 0.00372206f $X=3.065 $Y=1.162 $X2=0 $Y2=0
cc_187 N_A_331_47#_M1000_g X 0.0017144f $X=2.565 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_331_47#_M1009_g X 0.0114785f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_331_47#_c_248_n X 0.00245561f $X=2.335 $Y=0.72 $X2=0 $Y2=0
cc_190 N_A_331_47#_c_233_n X 0.026178f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_331_47#_c_234_n X 0.02276f $X=3.065 $Y=1.162 $X2=0 $Y2=0
cc_192 N_A_331_47#_M1005_g N_X_c_383_n 0.0128294f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_331_47#_M1000_g N_X_c_384_n 0.00544414f $X=2.565 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A_331_47#_M1009_g N_X_c_384_n 0.00847502f $X=3.065 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A_331_47#_c_234_n N_X_c_384_n 0.00310423f $X=3.065 $Y=1.162 $X2=0 $Y2=0
cc_196 N_A_331_47#_M1002_g N_X_c_370_n 0.00195285f $X=2.565 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_331_47#_M1005_g N_X_c_370_n 0.0157415f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_331_47#_c_237_n N_X_c_370_n 0.00699251f $X=2.335 $Y=1.622 $X2=0 $Y2=0
cc_199 N_A_331_47#_c_233_n N_X_c_370_n 0.0117143f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_331_47#_c_234_n N_X_c_370_n 0.00660546f $X=3.065 $Y=1.162 $X2=0 $Y2=0
cc_201 N_A_331_47#_c_248_n N_VGND_M1008_d 0.00646208f $X=2.335 $Y=0.72 $X2=0
+ $Y2=0
cc_202 N_A_331_47#_c_233_n N_VGND_M1008_d 9.64575e-19 $X=2.51 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_A_331_47#_M1000_g N_VGND_c_404_n 0.00310635f $X=2.565 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_331_47#_c_231_n N_VGND_c_404_n 0.0144159f $X=1.78 $Y=0.41 $X2=0 $Y2=0
cc_205 N_A_331_47#_c_248_n N_VGND_c_404_n 0.0188777f $X=2.335 $Y=0.72 $X2=0
+ $Y2=0
cc_206 N_A_331_47#_c_234_n N_VGND_c_404_n 2.78268e-19 $X=3.065 $Y=1.162 $X2=0
+ $Y2=0
cc_207 N_A_331_47#_M1009_g N_VGND_c_406_n 0.0113274f $X=3.065 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_331_47#_c_231_n N_VGND_c_407_n 0.0207456f $X=1.78 $Y=0.41 $X2=0 $Y2=0
cc_209 N_A_331_47#_c_248_n N_VGND_c_407_n 0.00309271f $X=2.335 $Y=0.72 $X2=0
+ $Y2=0
cc_210 N_A_331_47#_M1000_g N_VGND_c_410_n 0.00473078f $X=2.565 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_331_47#_M1009_g N_VGND_c_410_n 0.00431806f $X=3.065 $Y=0.445 $X2=0
+ $Y2=0
cc_212 N_A_331_47#_c_248_n N_VGND_c_410_n 0.00212171f $X=2.335 $Y=0.72 $X2=0
+ $Y2=0
cc_213 N_A_331_47#_M1008_s N_VGND_c_412_n 0.00209319f $X=1.655 $Y=0.235 $X2=0
+ $Y2=0
cc_214 N_A_331_47#_M1000_g N_VGND_c_412_n 0.00748898f $X=2.565 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_331_47#_M1009_g N_VGND_c_412_n 0.00687022f $X=3.065 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_A_331_47#_c_231_n N_VGND_c_412_n 0.012358f $X=1.78 $Y=0.41 $X2=0 $Y2=0
cc_217 N_A_331_47#_c_248_n N_VGND_c_412_n 0.00931771f $X=2.335 $Y=0.72 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_318_n N_X_M1002_d 0.00735138f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_c_322_n X 0.0639311f $X=3.35 $Y=1.855 $X2=0 $Y2=0
cc_220 N_VPWR_c_322_n X 0.0173876f $X=3.35 $Y=1.855 $X2=0 $Y2=0
cc_221 N_VPWR_c_326_n N_X_c_383_n 0.019836f $X=3.265 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_318_n N_X_c_383_n 0.0118607f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_223 X N_VGND_c_406_n 0.0234673f $X=3.385 $Y=0.765 $X2=0 $Y2=0
cc_224 N_X_c_384_n N_VGND_c_406_n 0.0205475f $X=2.855 $Y=0.45 $X2=0 $Y2=0
cc_225 N_X_c_384_n N_VGND_c_410_n 0.0166458f $X=2.855 $Y=0.45 $X2=0 $Y2=0
cc_226 N_X_M1000_d N_VGND_c_412_n 0.00737045f $X=2.64 $Y=0.235 $X2=0 $Y2=0
cc_227 X N_VGND_c_412_n 0.00811046f $X=3.385 $Y=0.765 $X2=0 $Y2=0
cc_228 N_X_c_384_n N_VGND_c_412_n 0.0116082f $X=2.855 $Y=0.45 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_4.spice
* Created: Thu Aug 27 14:23:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_4.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_4  VNB VPB A KAPWR X VGND VPWR
* 
* VGND	VGND
* X	X
* KAPWR	KAPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.1113 PD=0.755 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_27_47#_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.07035 PD=0.7 PS=0.755 NRD=0 NRS=15.708 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1000_d N_A_27_47#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_27_47#_M1004_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1004_d N_A_27_47#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1218 PD=0.7 PS=1.42 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_KAPWR_M1006_d N_A_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.265 PD=1.33 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1002_d N_A_27_47#_M1002_g N_KAPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.165 PD=1.28 PS=1.33 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75000.7
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1002_d N_A_27_47#_M1007_g N_KAPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1008 N_X_M1008_d N_A_27_47#_M1008_g N_KAPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1008_d N_A_27_47#_M1009_g N_KAPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.3 PD=1.28 PS=2.6 NRD=0 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.0397 P=9.49
c_31 VNB 0 9.76919e-20 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__lpflow_clkbufkapwr_4.pxi.spice"
*
.ends
*
*

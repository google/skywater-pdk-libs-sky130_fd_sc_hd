* File: sky130_fd_sc_hd__o221a_2.pex.spice
* Created: Tue Sep  1 19:22:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O221A_2%C1 1 3 6 8 9 10 19
c32 9 0 3.65277e-21 $X=0.63 $Y=1.15
r33 13 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r34 10 19 0.823174 $w=3.48e-07 $l=2.5e-08 $layer=LI1_cond $X=0.205 $Y=1.15
+ $X2=0.23 $Y2=1.15
r35 8 13 48.6364 $w=3.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.555 $Y=1.15
+ $X2=0.26 $Y2=1.15
r36 8 9 5.70552 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.555 $Y=1.15 $X2=0.63
+ $Y2=1.15
r37 4 9 38.5496 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.63 $Y=1.325
+ $X2=0.63 $Y2=1.15
r38 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.63 $Y=1.325 $X2=0.63
+ $Y2=1.985
r39 1 9 38.5496 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.63 $Y=0.975
+ $X2=0.63 $Y2=1.15
r40 1 3 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.63 $Y=0.975
+ $X2=0.63 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%B1 1 3 6 8 11
r39 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.16
+ $X2=1.05 $Y2=1.325
r40 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r41 6 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.11 $Y=1.985
+ $X2=1.11 $Y2=1.325
r42 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=0.995
+ $X2=1.05 $Y2=1.16
r43 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.05 $Y=0.995 $X2=1.05
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%B2 3 6 8 9 14 16
c41 14 0 1.39659e-19 $X=1.625 $Y=1.16
c42 9 0 2.99892e-19 $X=1.585 $Y=1.53
c43 8 0 3.65277e-21 $X=1.585 $Y=1.19
r44 14 17 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.577 $Y=1.16
+ $X2=1.577 $Y2=1.325
r45 14 16 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.577 $Y=1.16
+ $X2=1.577 $Y2=0.995
r46 8 9 8.2563 $w=4.58e-07 $l=2.55e-07 $layer=LI1_cond $X=1.645 $Y=1.275
+ $X2=1.645 $Y2=1.53
r47 8 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.16 $X2=1.625 $Y2=1.16
r48 6 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.485 $Y=1.985
+ $X2=1.485 $Y2=1.325
r49 3 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.47 $Y=0.56 $X2=1.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%A2 3 6 8 9 13 14 15
c38 13 0 1.09246e-19 $X=2.25 $Y=1.16
c39 9 0 3.22531e-19 $X=2.065 $Y=1.53
r40 14 17 6.23203 $w=2.08e-07 $l=1.18e-07 $layer=LI1_cond $X=2.25 $Y=1.18
+ $X2=2.132 $Y2=1.18
r41 13 16 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.16 $X2=2.3
+ $Y2=1.325
r42 13 15 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.16 $X2=2.3
+ $Y2=0.995
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r44 9 17 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=2.132 $Y=1.53
+ $X2=2.132 $Y2=1.285
r45 8 17 3.53853 $w=2.08e-07 $l=6.7e-08 $layer=LI1_cond $X=2.065 $Y=1.18
+ $X2=2.132 $Y2=1.18
r46 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.41 $Y=1.985
+ $X2=2.41 $Y2=1.325
r47 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.41 $Y=0.56 $X2=2.41
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%A1 3 5 7 8 11
c35 11 0 3.70702e-19 $X=2.83 $Y=1.16
r36 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.16
+ $X2=2.83 $Y2=1.325
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.16 $X2=2.83 $Y2=1.16
r38 8 12 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=2.985 $Y=1.18
+ $X2=2.83 $Y2=1.18
r39 5 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=0.995
+ $X2=2.83 $Y2=1.16
r40 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.83 $Y=0.995 $X2=2.83
+ $Y2=0.56
r41 3 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.77 $Y=1.985
+ $X2=2.77 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%A_38_47# 1 2 3 10 12 15 17 19 22 26 30 33 34
+ 37 38 39 41 42 43 45 48 51 53 58 64
c136 58 0 1.87831e-19 $X=3.41 $Y=1.16
r137 59 64 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=3.41 $Y=1.16
+ $X2=3.67 $Y2=1.16
r138 59 61 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.41 $Y=1.16
+ $X2=3.25 $Y2=1.16
r139 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.16 $X2=3.41 $Y2=1.16
r140 55 58 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=3.33 $Y=1.18 $X2=3.41
+ $Y2=1.18
r141 44 55 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.33 $Y=1.285
+ $X2=3.33 $Y2=1.18
r142 44 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.33 $Y=1.285
+ $X2=3.33 $Y2=1.455
r143 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=1.54
+ $X2=3.33 $Y2=1.455
r144 42 43 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.245 $Y=1.54
+ $X2=2.625 $Y2=1.54
r145 41 53 8.93966 $w=4.64e-07 $l=4.6465e-07 $layer=LI1_cond $X=2.54 $Y=1.875
+ $X2=2.2 $Y2=2.17
r146 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.54 $Y=1.625
+ $X2=2.625 $Y2=1.54
r147 40 41 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.54 $Y=1.625
+ $X2=2.54 $Y2=1.875
r148 38 53 22.2411 $w=4.64e-07 $l=7.47663e-07 $layer=LI1_cond $X=1.55 $Y=1.96
+ $X2=2.2 $Y2=2.17
r149 38 39 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.55 $Y=1.96
+ $X2=1.33 $Y2=1.96
r150 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.245 $Y=1.875
+ $X2=1.33 $Y2=1.96
r151 36 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.245 $Y=1.67
+ $X2=1.245 $Y2=1.875
r152 35 51 1.72457 $w=2.25e-07 $l=4.9503e-07 $layer=LI1_cond $X=0.715 $Y=1.557
+ $X2=0.25 $Y2=1.495
r153 34 36 6.9898 $w=2.25e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.16 $Y=1.557
+ $X2=1.245 $Y2=1.67
r154 34 35 22.7928 $w=2.23e-07 $l=4.45e-07 $layer=LI1_cond $X=1.16 $Y=1.557
+ $X2=0.715 $Y2=1.557
r155 33 51 4.72821 $w=2.5e-07 $l=4.04228e-07 $layer=LI1_cond $X=0.63 $Y=1.445
+ $X2=0.25 $Y2=1.495
r156 32 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.805
+ $X2=0.63 $Y2=0.72
r157 32 33 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.63 $Y=0.805
+ $X2=0.63 $Y2=1.445
r158 28 51 4.72821 $w=2.5e-07 $l=2.43926e-07 $layer=LI1_cond $X=0.415 $Y=1.67
+ $X2=0.25 $Y2=1.495
r159 28 30 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=0.415 $Y=1.67
+ $X2=0.415 $Y2=2.3
r160 24 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.72
+ $X2=0.63 $Y2=0.72
r161 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.335 $Y=0.635
+ $X2=0.335 $Y2=0.36
r162 20 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r163 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.985
r164 17 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=1.16
r165 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=0.56
r166 13 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.325
+ $X2=3.25 $Y2=1.16
r167 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.25 $Y=1.325
+ $X2=3.25 $Y2=1.985
r168 10 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=1.16
r169 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=0.56
r170 3 53 150 $w=1.7e-07 $l=8.44748e-07 $layer=licon1_PDIFF $count=4 $X=1.56
+ $Y=1.485 $X2=2.2 $Y2=1.96
r171 2 51 400 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.485 $X2=0.415 $Y2=1.62
r172 2 30 400 $w=1.7e-07 $l=9.02773e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.485 $X2=0.415 $Y2=2.3
r173 1 26 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.19
+ $Y=0.235 $X2=0.335 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%VPWR 1 2 3 12 16 18 20 23 24 25 31 38 44 48
+ 52
r60 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 42 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r65 39 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=2.72
+ $X2=2.96 $Y2=2.72
r66 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.125 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 38 47 4.90987 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.927 $Y2=2.72
r68 38 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.45 $Y2=2.72
r69 37 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 34 37 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 33 36 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r73 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.96 $Y2=2.72
r75 31 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r76 29 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r77 29 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 25 52 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 23 28 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.75 $Y=2.72 $X2=0.69
+ $Y2=2.72
r81 23 24 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.75 $Y=2.72 $X2=0.87
+ $Y2=2.72
r82 22 33 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.99 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 22 24 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=0.87
+ $Y2=2.72
r84 18 47 2.94129 $w=3.4e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.885 $Y=2.635
+ $X2=3.927 $Y2=2.72
r85 18 20 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=3.885 $Y=2.635
+ $X2=3.885 $Y2=2.3
r86 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=2.96 $Y2=2.72
r87 14 16 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=2.96 $Y2=1.96
r88 10 24 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=2.635
+ $X2=0.87 $Y2=2.72
r89 10 12 29.7714 $w=2.38e-07 $l=6.2e-07 $layer=LI1_cond $X=0.87 $Y=2.635
+ $X2=0.87 $Y2=2.015
r90 3 20 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=2.3
r91 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.845
+ $Y=1.485 $X2=2.98 $Y2=1.96
r92 1 12 300 $w=1.7e-07 $l=6.09098e-07 $layer=licon1_PDIFF $count=2 $X=0.705
+ $Y=1.485 $X2=0.875 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%X 1 2 9 11 13 15 20 24 27 30
r41 27 30 0.185878 $w=3.08e-07 $l=5e-09 $layer=LI1_cond $X=3.9 $Y=1.875 $X2=3.9
+ $Y2=1.87
r42 24 27 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=1.96 $X2=3.9
+ $Y2=1.875
r43 24 30 1.48702 $w=3.08e-07 $l=4e-08 $layer=LI1_cond $X=3.9 $Y=1.83 $X2=3.9
+ $Y2=1.87
r44 20 24 34.3874 $w=3.08e-07 $l=9.25e-07 $layer=LI1_cond $X=3.9 $Y=0.905
+ $X2=3.9 $Y2=1.83
r45 16 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.545 $Y=1.96
+ $X2=3.42 $Y2=1.96
r46 15 24 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.745 $Y=1.96
+ $X2=3.9 $Y2=1.96
r47 15 16 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.745 $Y=1.96
+ $X2=3.545 $Y2=1.96
r48 11 23 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.045
+ $X2=3.42 $Y2=1.96
r49 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.42 $Y=2.045
+ $X2=3.42 $Y2=2.3
r50 7 20 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.46 $Y=0.82 $X2=3.9
+ $Y2=0.82
r51 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.46 $Y=0.735
+ $X2=3.46 $Y2=0.39
r52 2 23 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=1.485 $X2=3.46 $Y2=1.96
r53 2 13 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=1.485 $X2=3.46 $Y2=2.3
r54 1 9 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.325
+ $Y=0.235 $X2=3.46 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%A_141_47# 1 2 11
r16 8 11 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.84 $Y=0.38 $X2=1.68
+ $Y2=0.38
r17 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.235 $X2=1.68 $Y2=0.38
r18 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.705
+ $Y=0.235 $X2=0.84 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%A_225_47# 1 2 7 11 16
r36 14 16 10.6882 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.26 $Y=0.775
+ $X2=1.47 $Y2=0.775
r37 9 11 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.62 $Y=0.735
+ $X2=2.62 $Y2=0.39
r38 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.455 $Y=0.82
+ $X2=2.62 $Y2=0.735
r39 7 16 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=2.455 $Y=0.82
+ $X2=1.47 $Y2=0.82
r40 2 11 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.235 $X2=2.62 $Y2=0.39
r41 1 14 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.26 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221A_2%VGND 1 2 3 12 14 18 20 22 24 25 26 35 41 45
+ 49
r61 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r62 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r63 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r64 39 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r65 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r66 36 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.04
+ $Y2=0
r67 36 38 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.45
+ $Y2=0
r68 35 44 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.967
+ $Y2=0
r69 35 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.45
+ $Y2=0
r70 34 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r71 34 49 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=0.23
+ $Y2=0
r72 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 29 33 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r74 29 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r75 26 49 0.00711354 $w=4.8e-07 $l=2.5e-08 $layer=MET1_cond $X=0.205 $Y=0
+ $X2=0.23 $Y2=0
r76 24 33 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.07
+ $Y2=0
r77 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.2
+ $Y2=0
r78 20 44 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.967 $Y2=0
r79 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0.39
r80 16 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0
r81 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0.39
r82 15 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.2
+ $Y2=0
r83 14 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0 $X2=3.04
+ $Y2=0
r84 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=2.285
+ $Y2=0
r85 10 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r86 10 12 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.2 $Y=0.085
+ $X2=2.2 $Y2=0.39
r87 3 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.39
r88 2 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.905
+ $Y=0.235 $X2=3.04 $Y2=0.39
r89 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.235 $X2=2.2 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__or4b_2.pxi.spice
* Created: Thu Aug 27 14:44:28 2020
* 
x_PM_SKY130_FD_SC_HD__OR4B_2%D_N N_D_N_M1001_g N_D_N_M1007_g D_N N_D_N_c_72_n
+ PM_SKY130_FD_SC_HD__OR4B_2%D_N
x_PM_SKY130_FD_SC_HD__OR4B_2%A_176_21# N_A_176_21#_M1006_d N_A_176_21#_M1000_d
+ N_A_176_21#_M1005_d N_A_176_21#_c_98_n N_A_176_21#_M1003_g N_A_176_21#_M1008_g
+ N_A_176_21#_c_99_n N_A_176_21#_M1004_g N_A_176_21#_M1011_g N_A_176_21#_c_100_n
+ N_A_176_21#_c_109_n N_A_176_21#_c_101_n N_A_176_21#_c_102_n
+ N_A_176_21#_c_103_n N_A_176_21#_c_104_n N_A_176_21#_c_105_n
+ N_A_176_21#_c_106_n PM_SKY130_FD_SC_HD__OR4B_2%A_176_21#
x_PM_SKY130_FD_SC_HD__OR4B_2%A N_A_M1006_g N_A_M1002_g A N_A_c_210_n
+ PM_SKY130_FD_SC_HD__OR4B_2%A
x_PM_SKY130_FD_SC_HD__OR4B_2%B N_B_M1009_g N_B_M1010_g B N_B_c_248_n
+ PM_SKY130_FD_SC_HD__OR4B_2%B
x_PM_SKY130_FD_SC_HD__OR4B_2%C N_C_M1013_g N_C_M1000_g C C N_C_c_286_n
+ PM_SKY130_FD_SC_HD__OR4B_2%C
x_PM_SKY130_FD_SC_HD__OR4B_2%A_27_53# N_A_27_53#_M1001_s N_A_27_53#_M1007_s
+ N_A_27_53#_M1012_g N_A_27_53#_M1005_g N_A_27_53#_c_315_n N_A_27_53#_c_320_n
+ N_A_27_53#_c_316_n N_A_27_53#_c_317_n N_A_27_53#_c_345_n N_A_27_53#_c_321_n
+ N_A_27_53#_c_322_n N_A_27_53#_c_323_n N_A_27_53#_c_324_n N_A_27_53#_c_318_n
+ N_A_27_53#_c_326_n N_A_27_53#_c_327_n PM_SKY130_FD_SC_HD__OR4B_2%A_27_53#
x_PM_SKY130_FD_SC_HD__OR4B_2%VPWR N_VPWR_M1007_d N_VPWR_M1011_d VPWR
+ N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_417_n N_VPWR_c_422_n
+ N_VPWR_c_423_n PM_SKY130_FD_SC_HD__OR4B_2%VPWR
x_PM_SKY130_FD_SC_HD__OR4B_2%X N_X_M1003_s N_X_M1008_s N_X_c_467_n N_X_c_470_n
+ N_X_c_480_n X PM_SKY130_FD_SC_HD__OR4B_2%X
x_PM_SKY130_FD_SC_HD__OR4B_2%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_M1009_d
+ N_VGND_M1012_d N_VGND_c_503_n N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n
+ N_VGND_c_507_n VGND N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n
+ N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n VGND
+ PM_SKY130_FD_SC_HD__OR4B_2%VGND
cc_1 VNB N_D_N_M1001_g 0.0346312f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB D_N 0.00896472f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_D_N_c_72_n 0.0374744f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_176_21#_c_98_n 0.0168438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_176_21#_c_99_n 0.0163785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_176_21#_c_100_n 0.00416821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_176_21#_c_101_n 8.89549e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_176_21#_c_102_n 0.0126212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_176_21#_c_103_n 9.26975e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_176_21#_c_104_n 0.00327171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_176_21#_c_105_n 0.0354325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_176_21#_c_106_n 0.00133824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_M1006_g 0.027023f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_14 VNB A 0.00567591f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_c_210_n 0.0202916f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_16 VNB N_B_M1009_g 0.03989f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_17 VNB N_C_M1000_g 0.0250329f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.695
cc_18 VNB C 0.0237205f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_C_c_286_n 0.019552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_53#_M1012_g 0.0575627f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_21 VNB N_A_27_53#_c_315_n 0.0165637f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_22 VNB N_A_27_53#_c_316_n 0.00379912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_53#_c_317_n 0.00938726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_53#_c_318_n 0.00665284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_417_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_467_n 8.17626e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_503_n 0.00413572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_504_n 5.88141e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_505_n 8.05577e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_506_n 0.0114996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_507_n 0.0169953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_508_n 0.0162201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_509_n 0.0134689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_510_n 0.0124058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_511_n 0.0222466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_512_n 0.00523295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_513_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_514_n 0.210204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VPB N_D_N_M1007_g 0.0265617f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_40 VPB D_N 0.00773293f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_41 VPB N_D_N_c_72_n 0.00960864f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_42 VPB N_A_176_21#_M1008_g 0.0211083f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_43 VPB N_A_176_21#_M1011_g 0.0209053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_176_21#_c_109_n 0.0284833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_176_21#_c_104_n 0.00237478f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_176_21#_c_105_n 0.0059224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_M1002_g 0.0206731f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_48 VPB N_A_c_210_n 0.00411461f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_B_M1009_g 0.0247431f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.475
cc_50 VPB B 0.0137595f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_51 VPB N_B_c_248_n 0.0349376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_C_M1013_g 0.0190729f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.475
cc_53 VPB N_C_c_286_n 0.00418337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_53#_M1012_g 0.0367708f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_55 VPB N_A_27_53#_c_320_n 0.0183349f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_53#_c_321_n 0.00745379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_53#_c_322_n 0.0044514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_53#_c_323_n 0.00187838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_53#_c_324_n 0.00815442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_53#_c_318_n 0.00299162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_53#_c_326_n 0.00250791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_53#_c_327_n 0.0388337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_418_n 0.0185074f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_64 VPB N_VPWR_c_419_n 0.0168925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_420_n 0.0517936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_417_n 0.0735043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_422_n 0.0163131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_423_n 0.0135969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_X_c_467_n 0.0011611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 N_D_N_M1001_g N_A_176_21#_c_98_n 0.0163129f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_71 N_D_N_M1007_g N_A_176_21#_M1008_g 0.0163129f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_72 N_D_N_c_72_n N_A_176_21#_c_105_n 0.0163129f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_73 N_D_N_M1001_g N_A_27_53#_c_315_n 0.00139995f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_74 N_D_N_M1007_g N_A_27_53#_c_320_n 0.025591f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_75 D_N N_A_27_53#_c_320_n 0.0252458f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_76 N_D_N_c_72_n N_A_27_53#_c_320_n 0.00138357f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_77 N_D_N_M1001_g N_A_27_53#_c_316_n 0.0170526f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_78 D_N N_A_27_53#_c_316_n 0.00547962f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_79 N_D_N_c_72_n N_A_27_53#_c_316_n 0.00110593f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_80 D_N N_A_27_53#_c_317_n 0.0223758f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_81 N_D_N_c_72_n N_A_27_53#_c_317_n 0.00573424f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_82 N_D_N_M1001_g N_A_27_53#_c_318_n 0.00922323f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_83 D_N N_A_27_53#_c_318_n 0.0270768f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_84 N_D_N_M1007_g N_VPWR_c_418_n 0.00253597f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_85 N_D_N_M1007_g N_VPWR_c_417_n 0.00322858f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_86 N_D_N_M1001_g N_X_c_467_n 2.76214e-19 $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_87 N_D_N_M1001_g N_X_c_470_n 2.58841e-19 $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_88 N_D_N_M1001_g X 3.71159e-19 $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_89 N_D_N_M1001_g N_VGND_c_503_n 0.00478714f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_90 N_D_N_M1001_g N_VGND_c_511_n 0.00413798f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_91 N_D_N_M1001_g N_VGND_c_514_n 0.0066853f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_92 N_A_176_21#_c_99_n N_A_M1006_g 0.0177514f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_176_21#_c_100_n N_A_M1006_g 0.0124599f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_94 N_A_176_21#_c_101_n N_A_M1006_g 0.00129218f $X=2.07 $Y=0.47 $X2=0 $Y2=0
cc_95 N_A_176_21#_c_104_n N_A_M1006_g 0.00368162f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_176_21#_M1011_g N_A_M1002_g 0.0249411f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_176_21#_c_109_n N_A_M1002_g 0.0109674f $X=3.225 $Y=1.53 $X2=0 $Y2=0
cc_98 N_A_176_21#_c_104_n N_A_M1002_g 0.00205188f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_176_21#_c_100_n A 0.0161642f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_100 N_A_176_21#_c_109_n A 0.0410544f $X=3.225 $Y=1.53 $X2=0 $Y2=0
cc_101 N_A_176_21#_c_102_n A 0.0121242f $X=2.885 $Y=0.82 $X2=0 $Y2=0
cc_102 N_A_176_21#_c_104_n A 0.0171977f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_176_21#_c_105_n A 6.28947e-19 $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_176_21#_c_106_n A 0.0141021f $X=2.07 $Y=0.82 $X2=0 $Y2=0
cc_105 N_A_176_21#_c_100_n N_A_c_210_n 0.00122978f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_106 N_A_176_21#_c_109_n N_A_c_210_n 0.00285374f $X=3.225 $Y=1.53 $X2=0 $Y2=0
cc_107 N_A_176_21#_c_104_n N_A_c_210_n 0.00239718f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_176_21#_c_105_n N_A_c_210_n 0.0150056f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_176_21#_c_106_n N_A_c_210_n 0.00178723f $X=2.07 $Y=0.82 $X2=0 $Y2=0
cc_110 N_A_176_21#_c_109_n N_B_M1009_g 0.0113059f $X=3.225 $Y=1.53 $X2=0 $Y2=0
cc_111 N_A_176_21#_c_101_n N_B_M1009_g 0.00549939f $X=2.07 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A_176_21#_c_102_n N_B_M1009_g 0.0131801f $X=2.885 $Y=0.82 $X2=0 $Y2=0
cc_113 N_A_176_21#_M1011_g B 0.00370524f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_176_21#_M1011_g N_B_c_248_n 0.00297018f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_176_21#_c_109_n N_C_M1013_g 0.0111483f $X=3.225 $Y=1.53 $X2=0 $Y2=0
cc_116 N_A_176_21#_c_102_n N_C_M1000_g 0.0113262f $X=2.885 $Y=0.82 $X2=0 $Y2=0
cc_117 N_A_176_21#_c_103_n N_C_M1000_g 0.001237f $X=2.97 $Y=0.47 $X2=0 $Y2=0
cc_118 N_A_176_21#_c_109_n C 0.0750642f $X=3.225 $Y=1.53 $X2=0 $Y2=0
cc_119 N_A_176_21#_c_102_n C 0.0382718f $X=2.885 $Y=0.82 $X2=0 $Y2=0
cc_120 N_A_176_21#_c_109_n N_C_c_286_n 0.00310331f $X=3.225 $Y=1.53 $X2=0 $Y2=0
cc_121 N_A_176_21#_c_102_n N_C_c_286_n 0.00322194f $X=2.885 $Y=0.82 $X2=0 $Y2=0
cc_122 N_A_176_21#_c_109_n N_A_27_53#_M1012_g 0.0160163f $X=3.225 $Y=1.53 $X2=0
+ $Y2=0
cc_123 N_A_176_21#_c_102_n N_A_27_53#_M1012_g 0.00538974f $X=2.885 $Y=0.82 $X2=0
+ $Y2=0
cc_124 N_A_176_21#_c_103_n N_A_27_53#_M1012_g 0.001237f $X=2.97 $Y=0.47 $X2=0
+ $Y2=0
cc_125 N_A_176_21#_M1008_g N_A_27_53#_c_320_n 8.57431e-19 $X=0.955 $Y=1.985
+ $X2=0 $Y2=0
cc_126 N_A_176_21#_c_105_n N_A_27_53#_c_320_n 0.00455081f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_127 N_A_176_21#_c_98_n N_A_27_53#_c_316_n 0.001313f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_A_176_21#_M1008_g N_A_27_53#_c_345_n 0.0135374f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_A_176_21#_M1011_g N_A_27_53#_c_345_n 0.0113663f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_176_21#_c_104_n N_A_27_53#_c_345_n 0.00367656f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_131 N_A_176_21#_c_109_n N_A_27_53#_c_321_n 0.0720254f $X=3.225 $Y=1.53 $X2=0
+ $Y2=0
cc_132 N_A_176_21#_c_109_n N_A_27_53#_c_324_n 0.00757798f $X=3.225 $Y=1.53 $X2=0
+ $Y2=0
cc_133 N_A_176_21#_c_98_n N_A_27_53#_c_318_n 0.00455081f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_A_176_21#_M1008_g N_A_27_53#_c_326_n 5.27992e-19 $X=0.955 $Y=1.985
+ $X2=0 $Y2=0
cc_135 N_A_176_21#_M1011_g N_A_27_53#_c_326_n 0.00982358f $X=1.375 $Y=1.985
+ $X2=0 $Y2=0
cc_136 N_A_176_21#_c_109_n N_A_27_53#_c_326_n 0.00376824f $X=3.225 $Y=1.53 $X2=0
+ $Y2=0
cc_137 N_A_176_21#_c_104_n N_A_27_53#_c_326_n 0.0138337f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_176_21#_c_109_n N_A_27_53#_c_327_n 0.00133432f $X=3.225 $Y=1.53 $X2=0
+ $Y2=0
cc_139 N_A_176_21#_c_109_n N_VPWR_M1011_d 6.48779e-19 $X=3.225 $Y=1.53 $X2=0
+ $Y2=0
cc_140 N_A_176_21#_c_104_n N_VPWR_M1011_d 0.00171868f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_176_21#_M1008_g N_VPWR_c_419_n 0.0041283f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_176_21#_M1011_g N_VPWR_c_419_n 0.00413971f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_176_21#_M1008_g N_VPWR_c_417_n 0.00690618f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_176_21#_M1011_g N_VPWR_c_417_n 0.00688158f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_176_21#_M1008_g N_VPWR_c_422_n 0.00623145f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_176_21#_M1011_g N_VPWR_c_423_n 0.00520955f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_176_21#_c_98_n N_X_c_467_n 0.00406091f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_176_21#_M1008_g N_X_c_467_n 0.00362416f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_176_21#_c_99_n N_X_c_467_n 0.00135948f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_176_21#_M1011_g N_X_c_467_n 0.00110132f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_176_21#_c_104_n N_X_c_467_n 0.0397823f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_176_21#_c_105_n N_X_c_467_n 0.0118208f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_176_21#_c_98_n N_X_c_470_n 0.00374785f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_176_21#_c_105_n N_X_c_470_n 0.00371015f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_176_21#_M1008_g N_X_c_480_n 0.00648335f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_176_21#_c_105_n N_X_c_480_n 0.00363828f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_176_21#_c_98_n X 0.00722131f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_176_21#_c_109_n A_387_297# 0.00220477f $X=3.225 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_176_21#_c_109_n A_483_297# 0.00102299f $X=3.225 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_176_21#_c_109_n A_555_297# 0.00230585f $X=3.225 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_176_21#_c_100_n N_VGND_M1004_d 0.0015209f $X=1.985 $Y=0.82 $X2=0
+ $Y2=0
cc_162 N_A_176_21#_c_104_n N_VGND_M1004_d 9.97566e-19 $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_176_21#_c_98_n N_VGND_c_503_n 0.00274665f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_176_21#_c_98_n N_VGND_c_504_n 6.31514e-19 $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A_176_21#_c_99_n N_VGND_c_504_n 0.00688434f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_176_21#_c_100_n N_VGND_c_504_n 0.010792f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_167 N_A_176_21#_c_104_n N_VGND_c_504_n 0.00553109f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_176_21#_c_101_n N_VGND_c_505_n 0.0105328f $X=2.07 $Y=0.47 $X2=0 $Y2=0
cc_169 N_A_176_21#_c_102_n N_VGND_c_505_n 0.0145277f $X=2.885 $Y=0.82 $X2=0
+ $Y2=0
cc_170 N_A_176_21#_c_98_n N_VGND_c_508_n 0.00460147f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_176_21#_c_99_n N_VGND_c_508_n 0.00506536f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_176_21#_c_104_n N_VGND_c_508_n 2.81698e-19 $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_173 N_A_176_21#_c_100_n N_VGND_c_509_n 0.00230538f $X=1.985 $Y=0.82 $X2=0
+ $Y2=0
cc_174 N_A_176_21#_c_101_n N_VGND_c_509_n 0.00869924f $X=2.07 $Y=0.47 $X2=0
+ $Y2=0
cc_175 N_A_176_21#_c_102_n N_VGND_c_509_n 0.00320252f $X=2.885 $Y=0.82 $X2=0
+ $Y2=0
cc_176 N_A_176_21#_c_102_n N_VGND_c_510_n 0.00230538f $X=2.885 $Y=0.82 $X2=0
+ $Y2=0
cc_177 N_A_176_21#_c_103_n N_VGND_c_510_n 0.00854817f $X=2.97 $Y=0.47 $X2=0
+ $Y2=0
cc_178 N_A_176_21#_c_98_n N_VGND_c_514_n 0.0077748f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_179 N_A_176_21#_c_99_n N_VGND_c_514_n 0.00823236f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_176_21#_c_100_n N_VGND_c_514_n 0.00488905f $X=1.985 $Y=0.82 $X2=0
+ $Y2=0
cc_181 N_A_176_21#_c_101_n N_VGND_c_514_n 0.00628404f $X=2.07 $Y=0.47 $X2=0
+ $Y2=0
cc_182 N_A_176_21#_c_102_n N_VGND_c_514_n 0.0107769f $X=2.885 $Y=0.82 $X2=0
+ $Y2=0
cc_183 N_A_176_21#_c_103_n N_VGND_c_514_n 0.00628404f $X=2.97 $Y=0.47 $X2=0
+ $Y2=0
cc_184 N_A_176_21#_c_104_n N_VGND_c_514_n 0.00125691f $X=1.375 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A_M1006_g N_B_M1009_g 0.0172988f $X=1.86 $Y=0.475 $X2=0 $Y2=0
cc_186 N_A_M1002_g N_B_M1009_g 0.0277591f $X=1.86 $Y=1.695 $X2=0 $Y2=0
cc_187 A N_B_M1009_g 0.00595691f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_188 N_A_c_210_n N_B_M1009_g 0.0216491f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_189 A C 0.0138677f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_190 N_A_M1002_g N_A_27_53#_c_321_n 0.0104288f $X=1.86 $Y=1.695 $X2=0 $Y2=0
cc_191 N_A_M1002_g N_A_27_53#_c_326_n 0.0024776f $X=1.86 $Y=1.695 $X2=0 $Y2=0
cc_192 N_A_M1002_g N_VPWR_c_420_n 0.00262341f $X=1.86 $Y=1.695 $X2=0 $Y2=0
cc_193 N_A_M1002_g N_VPWR_c_417_n 0.00336774f $X=1.86 $Y=1.695 $X2=0 $Y2=0
cc_194 N_A_M1002_g N_VPWR_c_423_n 7.40024e-19 $X=1.86 $Y=1.695 $X2=0 $Y2=0
cc_195 N_A_M1006_g N_VGND_c_504_n 0.0073121f $X=1.86 $Y=0.475 $X2=0 $Y2=0
cc_196 N_A_M1006_g N_VGND_c_505_n 5.28608e-19 $X=1.86 $Y=0.475 $X2=0 $Y2=0
cc_197 N_A_M1006_g N_VGND_c_509_n 0.00330296f $X=1.86 $Y=0.475 $X2=0 $Y2=0
cc_198 N_A_M1006_g N_VGND_c_514_n 0.0041734f $X=1.86 $Y=0.475 $X2=0 $Y2=0
cc_199 B N_C_M1013_g 0.00131774f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_200 N_B_M1009_g N_C_M1000_g 0.0250288f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_201 N_B_M1009_g C 0.0013979f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_202 N_B_M1009_g N_C_c_286_n 0.066724f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_203 N_B_M1009_g N_A_27_53#_M1012_g 0.00121851f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_204 N_B_M1009_g N_A_27_53#_c_321_n 0.0102124f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_205 B N_A_27_53#_c_321_n 0.0507965f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_206 N_B_c_248_n N_A_27_53#_c_321_n 0.0011406f $X=2.28 $Y=2.3 $X2=0 $Y2=0
cc_207 N_B_M1009_g N_A_27_53#_c_322_n 0.00179517f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_208 B N_A_27_53#_c_322_n 0.00691653f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_209 B N_A_27_53#_c_323_n 0.0143615f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_210 N_B_c_248_n N_A_27_53#_c_323_n 4.52412e-19 $X=2.28 $Y=2.3 $X2=0 $Y2=0
cc_211 N_B_M1009_g N_A_27_53#_c_326_n 0.00253311f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_212 B N_A_27_53#_c_326_n 0.00246643f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_213 B N_A_27_53#_c_327_n 0.00162833f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_214 N_B_c_248_n N_A_27_53#_c_327_n 0.00560469f $X=2.28 $Y=2.3 $X2=0 $Y2=0
cc_215 B N_VPWR_c_420_n 0.0339392f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_216 N_B_c_248_n N_VPWR_c_420_n 0.00754324f $X=2.28 $Y=2.3 $X2=0 $Y2=0
cc_217 B N_VPWR_c_417_n 0.0248489f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_218 N_B_c_248_n N_VPWR_c_417_n 0.0107433f $X=2.28 $Y=2.3 $X2=0 $Y2=0
cc_219 B N_VPWR_c_423_n 0.00699952f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_220 N_B_c_248_n N_VPWR_c_423_n 7.6396e-19 $X=2.28 $Y=2.3 $X2=0 $Y2=0
cc_221 N_B_M1009_g N_VGND_c_504_n 5.15945e-19 $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_222 N_B_M1009_g N_VGND_c_505_n 0.00733885f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_223 N_B_M1009_g N_VGND_c_509_n 0.00330296f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_224 N_B_M1009_g N_VGND_c_514_n 0.0041734f $X=2.34 $Y=0.475 $X2=0 $Y2=0
cc_225 N_C_M1013_g N_A_27_53#_M1012_g 0.0256158f $X=2.7 $Y=1.695 $X2=0 $Y2=0
cc_226 N_C_M1000_g N_A_27_53#_M1012_g 0.0213843f $X=2.76 $Y=0.475 $X2=0 $Y2=0
cc_227 C N_A_27_53#_M1012_g 0.016761f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_228 N_C_c_286_n N_A_27_53#_M1012_g 0.021893f $X=2.76 $Y=1.16 $X2=0 $Y2=0
cc_229 N_C_M1013_g N_A_27_53#_c_321_n 0.0100804f $X=2.7 $Y=1.695 $X2=0 $Y2=0
cc_230 N_C_M1013_g N_A_27_53#_c_322_n 0.00186808f $X=2.7 $Y=1.695 $X2=0 $Y2=0
cc_231 N_C_M1013_g N_VPWR_c_420_n 0.00232878f $X=2.7 $Y=1.695 $X2=0 $Y2=0
cc_232 N_C_M1013_g N_VPWR_c_417_n 0.00292242f $X=2.7 $Y=1.695 $X2=0 $Y2=0
cc_233 N_C_M1000_g N_VGND_c_505_n 0.00688697f $X=2.76 $Y=0.475 $X2=0 $Y2=0
cc_234 N_C_M1000_g N_VGND_c_507_n 5.53013e-19 $X=2.76 $Y=0.475 $X2=0 $Y2=0
cc_235 C N_VGND_c_507_n 0.0113271f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_236 N_C_M1000_g N_VGND_c_510_n 0.00330296f $X=2.76 $Y=0.475 $X2=0 $Y2=0
cc_237 N_C_M1000_g N_VGND_c_514_n 0.00405984f $X=2.76 $Y=0.475 $X2=0 $Y2=0
cc_238 N_A_27_53#_c_320_n N_VPWR_M1007_d 0.00645115f $X=0.51 $Y=1.747 $X2=-0.19
+ $Y2=-0.24
cc_239 N_A_27_53#_c_345_n N_VPWR_M1007_d 0.0032732f $X=1.44 $Y=2.08 $X2=-0.19
+ $Y2=-0.24
cc_240 N_A_27_53#_c_318_n N_VPWR_M1007_d 0.00116715f $X=0.637 $Y=1.605 $X2=-0.19
+ $Y2=-0.24
cc_241 N_A_27_53#_c_321_n N_VPWR_M1011_d 4.3544e-19 $X=2.86 $Y=1.87 $X2=0 $Y2=0
cc_242 N_A_27_53#_c_326_n N_VPWR_M1011_d 0.00472376f $X=1.577 $Y=1.87 $X2=0
+ $Y2=0
cc_243 N_A_27_53#_c_345_n N_VPWR_c_419_n 0.0108606f $X=1.44 $Y=2.08 $X2=0 $Y2=0
cc_244 N_A_27_53#_c_326_n N_VPWR_c_419_n 5.53374e-19 $X=1.577 $Y=1.87 $X2=0
+ $Y2=0
cc_245 N_A_27_53#_c_323_n N_VPWR_c_420_n 0.00771367f $X=3.03 $Y=2.3 $X2=0 $Y2=0
cc_246 N_A_27_53#_c_324_n N_VPWR_c_420_n 0.0129016f $X=3.105 $Y=2.3 $X2=0 $Y2=0
cc_247 N_A_27_53#_c_327_n N_VPWR_c_420_n 0.00762419f $X=3.18 $Y=2.3 $X2=0 $Y2=0
cc_248 N_A_27_53#_c_320_n N_VPWR_c_417_n 0.0166622f $X=0.51 $Y=1.747 $X2=0 $Y2=0
cc_249 N_A_27_53#_c_345_n N_VPWR_c_417_n 0.0168904f $X=1.44 $Y=2.08 $X2=0 $Y2=0
cc_250 N_A_27_53#_c_321_n N_VPWR_c_417_n 0.0139664f $X=2.86 $Y=1.87 $X2=0 $Y2=0
cc_251 N_A_27_53#_c_323_n N_VPWR_c_417_n 0.00617523f $X=3.03 $Y=2.3 $X2=0 $Y2=0
cc_252 N_A_27_53#_c_324_n N_VPWR_c_417_n 0.010971f $X=3.105 $Y=2.3 $X2=0 $Y2=0
cc_253 N_A_27_53#_c_326_n N_VPWR_c_417_n 0.00246311f $X=1.577 $Y=1.87 $X2=0
+ $Y2=0
cc_254 N_A_27_53#_c_327_n N_VPWR_c_417_n 0.0107433f $X=3.18 $Y=2.3 $X2=0 $Y2=0
cc_255 N_A_27_53#_c_320_n N_VPWR_c_422_n 0.0204248f $X=0.51 $Y=1.747 $X2=0 $Y2=0
cc_256 N_A_27_53#_c_345_n N_VPWR_c_422_n 0.00430549f $X=1.44 $Y=2.08 $X2=0 $Y2=0
cc_257 N_A_27_53#_c_321_n N_VPWR_c_423_n 0.00380528f $X=2.86 $Y=1.87 $X2=0 $Y2=0
cc_258 N_A_27_53#_c_326_n N_VPWR_c_423_n 0.016299f $X=1.577 $Y=1.87 $X2=0 $Y2=0
cc_259 N_A_27_53#_c_345_n N_X_M1008_s 0.00405739f $X=1.44 $Y=2.08 $X2=0 $Y2=0
cc_260 N_A_27_53#_c_316_n N_X_c_467_n 0.00907787f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_261 N_A_27_53#_c_318_n N_X_c_467_n 0.0420777f $X=0.637 $Y=1.605 $X2=0 $Y2=0
cc_262 N_A_27_53#_c_315_n N_X_c_470_n 0.00161347f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_263 N_A_27_53#_c_316_n N_X_c_470_n 0.00454492f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_264 N_A_27_53#_c_345_n N_X_c_480_n 0.018631f $X=1.44 $Y=2.08 $X2=0 $Y2=0
cc_265 N_A_27_53#_c_318_n N_X_c_480_n 0.0247171f $X=0.637 $Y=1.605 $X2=0 $Y2=0
cc_266 N_A_27_53#_c_321_n A_387_297# 0.00221923f $X=2.86 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_267 N_A_27_53#_c_321_n A_483_297# 0.00102299f $X=2.86 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_268 N_A_27_53#_c_321_n A_555_297# 0.00398838f $X=2.86 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_269 N_A_27_53#_c_316_n N_VGND_M1001_d 0.00318579f $X=0.595 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_270 N_A_27_53#_c_316_n N_VGND_c_503_n 0.0116177f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_271 N_A_27_53#_M1012_g N_VGND_c_505_n 5.2354e-19 $X=3.18 $Y=0.475 $X2=0 $Y2=0
cc_272 N_A_27_53#_M1012_g N_VGND_c_507_n 0.0101273f $X=3.18 $Y=0.475 $X2=0 $Y2=0
cc_273 N_A_27_53#_M1012_g N_VGND_c_510_n 0.00442511f $X=3.18 $Y=0.475 $X2=0
+ $Y2=0
cc_274 N_A_27_53#_c_315_n N_VGND_c_511_n 0.0123931f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_275 N_A_27_53#_c_316_n N_VGND_c_511_n 0.00393932f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_276 N_A_27_53#_M1012_g N_VGND_c_514_n 0.00784175f $X=3.18 $Y=0.475 $X2=0
+ $Y2=0
cc_277 N_A_27_53#_c_315_n N_VGND_c_514_n 0.00971608f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_278 N_A_27_53#_c_316_n N_VGND_c_514_n 0.00725735f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_417_n N_X_M1008_s 0.00285156f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_280 X N_VGND_c_503_n 0.0222357f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_281 N_X_c_470_n N_VGND_c_508_n 5.74861e-19 $X=1.11 $Y=0.675 $X2=0 $Y2=0
cc_282 X N_VGND_c_508_n 0.0165263f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_283 N_X_M1003_s N_VGND_c_514_n 0.00393977f $X=1.03 $Y=0.235 $X2=0 $Y2=0
cc_284 N_X_c_470_n N_VGND_c_514_n 8.42631e-19 $X=1.11 $Y=0.675 $X2=0 $Y2=0
cc_285 X N_VGND_c_514_n 0.0103753f $X=1.07 $Y=0.425 $X2=0 $Y2=0

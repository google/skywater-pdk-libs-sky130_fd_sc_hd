* File: sky130_fd_sc_hd__ebufn_2.spice.pex
* Created: Thu Aug 27 14:19:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EBUFN_2%A 3 7 9 10 14
c32 7 0 1.76927e-20 $X=0.47 $Y=2.165
c33 3 0 9.724e-20 $X=0.47 $Y=0.445
r34 14 17 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.552 $Y=1.16
+ $X2=0.552 $Y2=1.325
r35 14 16 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.552 $Y=1.16
+ $X2=0.552 $Y2=0.995
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.16 $X2=0.575 $Y2=1.16
r37 10 15 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.635 $Y=1.53
+ $X2=0.635 $Y2=1.16
r38 9 15 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=0.635 $Y=0.85
+ $X2=0.635 $Y2=1.16
r39 7 17 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=2.165
+ $X2=0.47 $Y2=1.325
r40 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%TE_B 3 7 9 11 13 14 16 18 19 20 23
c61 14 0 3.98363e-20 $X=2.28 $Y=1.395
r62 26 27 32.1566 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=1.1 $Y=1.395 $X2=1.1
+ $Y2=1.47
r63 23 26 37.668 $w=3.6e-07 $l=2.35e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.1
+ $Y2=1.395
r64 23 25 41.774 $w=3.6e-07 $l=1.35e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.1
+ $Y2=1.025
r65 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.16 $X2=1.115 $Y2=1.16
r66 20 24 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.115 $Y=0.85
+ $X2=1.115 $Y2=1.16
r67 16 18 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.355 $Y=1.47
+ $X2=2.355 $Y2=2.015
r68 15 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.01 $Y=1.395
+ $X2=1.935 $Y2=1.395
r69 14 16 27.1723 $w=1.48e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.28 $Y=1.395
+ $X2=2.355 $Y2=1.47
r70 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.28 $Y=1.395
+ $X2=2.01 $Y2=1.395
r71 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.47
+ $X2=1.935 $Y2=1.395
r72 11 13 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.935 $Y=1.47
+ $X2=1.935 $Y2=2.015
r73 10 26 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.28 $Y=1.395
+ $X2=1.1 $Y2=1.395
r74 9 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.86 $Y=1.395
+ $X2=1.935 $Y2=1.395
r75 9 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.86 $Y=1.395
+ $X2=1.28 $Y2=1.395
r76 7 27 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.995 $Y=2.165
+ $X2=0.995 $Y2=1.47
r77 3 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.995 $Y=0.445
+ $X2=0.995 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%A_214_47# 1 2 7 9 10 11 14 15 21 24 26 29 34
+ 36 37 38
c78 38 0 8.87727e-20 $X=2.8 $Y=0.96
c79 37 0 9.7054e-20 $X=2.8 $Y=1.035
c80 34 0 1.76927e-20 $X=1.592 $Y=1.605
c81 29 0 3.98363e-20 $X=2.8 $Y=1.16
c82 15 0 9.724e-20 $X=1.45 $Y=0.425
c83 11 0 1.57709e-19 $X=2.37 $Y=1.035
r84 37 38 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.8 $Y=1.035 $X2=2.8
+ $Y2=0.96
r85 32 34 11.7765 $w=3.18e-07 $l=3.27e-07 $layer=LI1_cond $X=1.265 $Y=1.605
+ $X2=1.592 $Y2=1.605
r86 30 37 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.8 $Y=1.16 $X2=2.8
+ $Y2=1.035
r87 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=1.16 $X2=2.8 $Y2=1.16
r88 27 36 1.78614 $w=2.5e-07 $l=1.43e-07 $layer=LI1_cond $X=1.735 $Y=1.15
+ $X2=1.592 $Y2=1.15
r89 27 29 49.0941 $w=2.48e-07 $l=1.065e-06 $layer=LI1_cond $X=1.735 $Y=1.15
+ $X2=2.8 $Y2=1.15
r90 26 34 1.43246 $w=2.85e-07 $l=1.6e-07 $layer=LI1_cond $X=1.592 $Y=1.445
+ $X2=1.592 $Y2=1.605
r91 25 36 4.66096 $w=2.82e-07 $l=1.25e-07 $layer=LI1_cond $X=1.592 $Y=1.275
+ $X2=1.592 $Y2=1.15
r92 25 26 6.87422 $w=2.83e-07 $l=1.7e-07 $layer=LI1_cond $X=1.592 $Y=1.275
+ $X2=1.592 $Y2=1.445
r93 24 36 4.66096 $w=2.82e-07 $l=1.25996e-07 $layer=LI1_cond $X=1.59 $Y=1.025
+ $X2=1.592 $Y2=1.15
r94 23 24 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=1.59 $Y=0.595
+ $X2=1.59 $Y2=1.025
r95 19 32 1.30983 $w=2.9e-07 $l=1.6e-07 $layer=LI1_cond $X=1.265 $Y=1.765
+ $X2=1.265 $Y2=1.605
r96 19 21 18.0814 $w=2.88e-07 $l=4.55e-07 $layer=LI1_cond $X=1.265 $Y=1.765
+ $X2=1.265 $Y2=2.22
r97 15 23 6.89985 $w=3.4e-07 $l=2.29565e-07 $layer=LI1_cond $X=1.45 $Y=0.425
+ $X2=1.59 $Y2=0.595
r98 15 17 8.30437 $w=3.38e-07 $l=2.45e-07 $layer=LI1_cond $X=1.45 $Y=0.425
+ $X2=1.205 $Y2=0.425
r99 14 38 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.715 $Y=0.56
+ $X2=2.715 $Y2=0.96
r100 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.035
+ $X2=2.8 $Y2=1.035
r101 10 11 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.635 $Y=1.035
+ $X2=2.37 $Y2=1.035
r102 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.295 $Y=0.96
+ $X2=2.37 $Y2=1.035
r103 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.295 $Y=0.96 $X2=2.295
+ $Y2=0.56
r104 2 21 600 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.845 $X2=1.205 $Y2=2.22
r105 1 17 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.205 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%A_27_47# 1 2 9 13 17 21 23 25 29 34 35 38 41
+ 48 49
c81 41 0 9.7054e-20 $X=3.465 $Y=1.19
c82 34 0 3.32593e-19 $X=3.32 $Y=1.19
r83 47 49 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=3.46 $Y=1.16
+ $X2=3.67 $Y2=1.16
r84 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.46
+ $Y=1.16 $X2=3.46 $Y2=1.16
r85 44 47 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=3.25 $Y=1.16
+ $X2=3.46 $Y2=1.16
r86 41 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.465 $Y=1.19
+ $X2=3.465 $Y2=1.19
r87 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=1.19
+ $X2=0.235 $Y2=1.19
r88 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.38 $Y=1.19
+ $X2=0.235 $Y2=1.19
r89 34 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.32 $Y=1.19
+ $X2=3.465 $Y2=1.19
r90 34 35 3.63861 $w=1.4e-07 $l=2.94e-06 $layer=MET1_cond $X=3.32 $Y=1.19
+ $X2=0.38 $Y2=1.19
r91 33 38 32.1213 $w=2.33e-07 $l=6.55e-07 $layer=LI1_cond $X=0.202 $Y=1.845
+ $X2=0.202 $Y2=1.19
r92 31 38 28.1981 $w=2.33e-07 $l=5.75e-07 $layer=LI1_cond $X=0.202 $Y=0.615
+ $X2=0.202 $Y2=1.19
r93 29 31 7.66598 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.215 $Y=0.445
+ $X2=0.215 $Y2=0.615
r94 23 33 5.89299 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.975
+ $X2=0.215 $Y2=1.845
r95 23 25 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=0.215 $Y=1.975
+ $X2=0.215 $Y2=2.22
r96 19 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.67 $Y=1.295
+ $X2=3.67 $Y2=1.16
r97 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.67 $Y=1.295
+ $X2=3.67 $Y2=1.985
r98 15 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.67 $Y=1.025
+ $X2=3.67 $Y2=1.16
r99 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.67 $Y=1.025
+ $X2=3.67 $Y2=0.56
r100 11 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.25 $Y=1.295
+ $X2=3.25 $Y2=1.16
r101 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.25 $Y=1.295
+ $X2=3.25 $Y2=1.985
r102 7 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.25 $Y=1.025
+ $X2=3.25 $Y2=1.16
r103 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.25 $Y=1.025
+ $X2=3.25 $Y2=0.56
r104 2 25 600 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.22
r105 1 29 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%VPWR 1 2 9 13 15 17 22 32 33 36 39
r50 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r53 30 33 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 29 32 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.145 $Y2=2.72
r58 27 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 26 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 23 36 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.95 $Y=2.72
+ $X2=0.732 $Y2=2.72
r63 23 25 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=0.95 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=2.145 $Y2=2.72
r65 22 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=2.72 $X2=1.61
+ $Y2=2.72
r66 17 36 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.732 $Y2=2.72
r67 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.635
+ $X2=2.145 $Y2=2.72
r71 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.145 $Y=2.635
+ $X2=2.145 $Y2=2.36
r72 7 36 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.732 $Y=2.635
+ $X2=0.732 $Y2=2.72
r73 7 9 16.2932 $w=4.33e-07 $l=6.15e-07 $layer=LI1_cond $X=0.732 $Y=2.635
+ $X2=0.732 $Y2=2.02
r74 2 13 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.545 $X2=2.145 $Y2=2.36
r75 1 9 300 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.845 $X2=0.735 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%A_320_309# 1 2 3 12 15 16 20 24 25
r39 23 25 9.59153 $w=5.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.965 $Y=2.2
+ $X2=3.125 $Y2=2.2
r40 23 24 16.926 $w=5.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.965 $Y=2.2
+ $X2=2.48 $Y2=2.2
r41 18 20 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=3.925 $Y=2.295
+ $X2=3.925 $Y2=1.96
r42 16 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.795 $Y=2.38
+ $X2=3.925 $Y2=2.295
r43 16 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.795 $Y=2.38
+ $X2=3.125 $Y2=2.38
r44 15 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.81 $Y=2.02
+ $X2=2.48 $Y2=2.02
r45 10 15 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.705 $Y=2.105
+ $X2=1.81 $Y2=2.02
r46 10 12 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=1.705 $Y=2.105
+ $X2=1.705 $Y2=2.3
r47 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=1.96
r48 2 23 300 $w=1.7e-07 $l=9.86889e-07 $layer=licon1_PDIFF $count=2 $X=2.43
+ $Y=1.545 $X2=2.965 $Y2=2.3
r49 1 12 600 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.545 $X2=1.725 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%Z 1 2 7 11 14 16 17 18 19 20 21 22 23 37 44
c56 44 0 1.01522e-19 $X=3.94 $Y=0.855
c57 16 0 1.91887e-19 $X=3.46 $Y=1.655
c58 14 0 1.57709e-19 $X=3.295 $Y=1.605
c59 7 0 2.29478e-19 $X=3.825 $Y=0.745
r60 22 23 9.41096 $w=3.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.94 $Y=1.19
+ $X2=3.94 $Y2=1.445
r61 21 44 3.33465 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.94 $Y=0.745
+ $X2=3.94 $Y2=0.855
r62 21 22 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.94 $Y=0.895
+ $X2=3.94 $Y2=1.19
r63 21 44 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=3.94 $Y=0.895 $X2=3.94
+ $Y2=0.855
r64 18 19 16.4943 $w=3.18e-07 $l=4.58e-07 $layer=LI1_cond $X=2.547 $Y=1.605
+ $X2=3.005 $Y2=1.605
r65 18 37 0.0720277 $w=3.18e-07 $l=2e-09 $layer=LI1_cond $X=2.547 $Y=1.605
+ $X2=2.545 $Y2=1.605
r66 17 37 16.2062 $w=3.18e-07 $l=4.5e-07 $layer=LI1_cond $X=2.095 $Y=1.605
+ $X2=2.545 $Y2=1.605
r67 14 19 10.444 $w=3.18e-07 $l=2.9e-07 $layer=LI1_cond $X=3.295 $Y=1.605
+ $X2=3.005 $Y2=1.605
r68 14 16 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=1.605
+ $X2=3.46 $Y2=1.605
r69 13 20 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.46 $Y=1.765
+ $X2=3.46 $Y2=1.87
r70 13 16 0.364692 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=3.46 $Y=1.765
+ $X2=3.46 $Y2=1.605
r71 12 16 6.46576 $w=2.5e-07 $l=1.96914e-07 $layer=LI1_cond $X=3.625 $Y=1.535
+ $X2=3.46 $Y2=1.605
r72 11 23 3.89832 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=3.825 $Y=1.535
+ $X2=3.94 $Y2=1.535
r73 11 12 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=3.825 $Y=1.535
+ $X2=3.625 $Y2=1.535
r74 7 21 3.48622 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=3.825 $Y=0.745
+ $X2=3.94 $Y2=0.745
r75 7 9 19.1201 $w=2.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.825 $Y=0.745
+ $X2=3.46 $Y2=0.745
r76 2 16 300 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=1.485 $X2=3.46 $Y2=1.655
r77 1 9 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.46 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%VGND 1 2 9 13 15 17 22 35 36 39 42
c53 35 0 1.01522e-19 $X=3.91 $Y=0
r54 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r55 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r56 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r57 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r58 33 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r59 32 35 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r60 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r61 30 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.505
+ $Y2=0
r62 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.99
+ $Y2=0
r63 29 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r64 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r65 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r66 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r67 25 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r68 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 23 39 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=0.682
+ $Y2=0
r70 23 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=1.15
+ $Y2=0
r71 22 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.505
+ $Y2=0
r72 22 28 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.07
+ $Y2=0
r73 17 39 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.682
+ $Y2=0
r74 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r75 15 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r76 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r77 11 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0
r78 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0.36
r79 7 39 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.682 $Y=0.085
+ $X2=0.682 $Y2=0
r80 7 9 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=0.682 $Y=0.085
+ $X2=0.682 $Y2=0.36
r81 2 13 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.37
+ $Y=0.235 $X2=2.505 $Y2=0.36
r82 1 9 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_2%A_392_47# 1 2 3 10 13 14 19 21
r38 19 21 44.0718 $w=1.88e-07 $l=7.55e-07 $layer=LI1_cond $X=3.125 $Y=0.37
+ $X2=3.88 $Y2=0.37
r39 16 18 3.84148 $w=2.83e-07 $l=9.5e-08 $layer=LI1_cond $X=2.982 $Y=0.655
+ $X2=2.982 $Y2=0.56
r40 15 19 7.17723 $w=1.9e-07 $l=1.84483e-07 $layer=LI1_cond $X=2.982 $Y=0.465
+ $X2=3.125 $Y2=0.37
r41 15 18 3.84148 $w=2.83e-07 $l=9.5e-08 $layer=LI1_cond $X=2.982 $Y=0.465
+ $X2=2.982 $Y2=0.56
r42 13 16 7.09239 $w=2e-07 $l=1.85375e-07 $layer=LI1_cond $X=2.84 $Y=0.755
+ $X2=2.982 $Y2=0.655
r43 13 14 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=2.84 $Y=0.755
+ $X2=2.17 $Y2=0.755
r44 10 14 7.01501 $w=2e-07 $l=1.78115e-07 $layer=LI1_cond $X=2.035 $Y=0.655
+ $X2=2.17 $Y2=0.755
r45 10 12 4.29259 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.035 $Y=0.655
+ $X2=2.035 $Y2=0.56
r46 3 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.38
r47 2 18 182 $w=1.7e-07 $l=4.09115e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.235 $X2=2.98 $Y2=0.56
r48 1 12 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.235 $X2=2.085 $Y2=0.56
.ends


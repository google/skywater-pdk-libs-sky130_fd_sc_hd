* File: sky130_fd_sc_hd__a211o_4.pex.spice
* Created: Thu Aug 27 13:59:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A211O_4%A_79_204# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 56 58 59 60 61 63 67 69 71 75 77 78 79 80 82 95
c163 95 0 2.25268e-20 $X=2.17 $Y=1.185
c164 78 0 3.76681e-19 $X=2.32 $Y=1.505
c165 77 0 1.19052e-19 $X=2.277 $Y=1.185
c166 56 0 1.54492e-19 $X=2.282 $Y=1.045
r167 92 93 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=1.33 $Y=1.185
+ $X2=1.725 $Y2=1.185
r168 91 92 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.295 $Y=1.185
+ $X2=1.33 $Y2=1.185
r169 90 91 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=0.9 $Y=1.185
+ $X2=1.295 $Y2=1.185
r170 89 90 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.865 $Y=1.185
+ $X2=0.9 $Y2=1.185
r171 82 84 10.0081 $w=3.78e-07 $l=3.3e-07 $layer=LI1_cond $X=3.83 $Y=0.38
+ $X2=3.83 $Y2=0.71
r172 78 79 10.2362 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=2.32 $Y=1.505
+ $X2=2.32 $Y2=1.675
r173 73 75 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.325 $Y=0.615
+ $X2=5.325 $Y2=0.36
r174 72 84 4.80115 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.02 $Y=0.71
+ $X2=3.83 $Y2=0.71
r175 71 73 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=5.16 $Y=0.71
+ $X2=5.325 $Y2=0.615
r176 71 72 66.5455 $w=1.88e-07 $l=1.14e-06 $layer=LI1_cond $X=5.16 $Y=0.71
+ $X2=4.02 $Y2=0.71
r177 70 80 6.34807 $w=1.9e-07 $l=1.23e-07 $layer=LI1_cond $X=2.97 $Y=0.71
+ $X2=2.847 $Y2=0.71
r178 69 84 4.80115 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.64 $Y=0.71
+ $X2=3.83 $Y2=0.71
r179 69 70 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=3.64 $Y=0.71 $X2=2.97
+ $Y2=0.71
r180 65 80 0.445202 $w=2.45e-07 $l=9.5e-08 $layer=LI1_cond $X=2.847 $Y=0.615
+ $X2=2.847 $Y2=0.71
r181 65 67 6.115 $w=2.43e-07 $l=1.3e-07 $layer=LI1_cond $X=2.847 $Y=0.615
+ $X2=2.847 $Y2=0.485
r182 61 63 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.455 $Y=1.955
+ $X2=3.345 $Y2=1.955
r183 59 80 6.34807 $w=1.9e-07 $l=1.22e-07 $layer=LI1_cond $X=2.725 $Y=0.71
+ $X2=2.847 $Y2=0.71
r184 59 60 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=2.725 $Y=0.71
+ $X2=2.37 $Y2=0.71
r185 58 61 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=2.367 $Y=1.87
+ $X2=2.455 $Y2=1.955
r186 58 79 12.3584 $w=1.73e-07 $l=1.95e-07 $layer=LI1_cond $X=2.367 $Y=1.87
+ $X2=2.367 $Y2=1.675
r187 56 77 7.33282 $w=1.8e-07 $l=1.42478e-07 $layer=LI1_cond $X=2.282 $Y=1.045
+ $X2=2.277 $Y2=1.185
r188 55 60 6.83148 $w=1.9e-07 $l=1.31852e-07 $layer=LI1_cond $X=2.282 $Y=0.805
+ $X2=2.37 $Y2=0.71
r189 55 56 15.2104 $w=1.73e-07 $l=2.4e-07 $layer=LI1_cond $X=2.282 $Y=0.805
+ $X2=2.282 $Y2=1.045
r190 53 77 7.33282 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=2.277 $Y=1.325
+ $X2=2.277 $Y2=1.185
r191 53 78 10.7912 $w=1.83e-07 $l=1.8e-07 $layer=LI1_cond $X=2.277 $Y=1.325
+ $X2=2.277 $Y2=1.505
r192 52 95 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.76 $Y=1.185
+ $X2=2.17 $Y2=1.185
r193 52 93 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.76 $Y=1.185
+ $X2=1.725 $Y2=1.185
r194 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.76
+ $Y=1.16 $X2=1.76 $Y2=1.16
r195 48 89 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.74 $Y=1.185
+ $X2=0.865 $Y2=1.185
r196 48 86 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.74 $Y=1.185
+ $X2=0.47 $Y2=1.185
r197 47 51 41.9819 $w=2.78e-07 $l=1.02e-06 $layer=LI1_cond $X=0.74 $Y=1.185
+ $X2=1.76 $Y2=1.185
r198 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.74
+ $Y=1.16 $X2=0.74 $Y2=1.16
r199 45 77 0.18844 $w=2.8e-07 $l=9.2e-08 $layer=LI1_cond $X=2.185 $Y=1.185
+ $X2=2.277 $Y2=1.185
r200 45 51 17.4924 $w=2.78e-07 $l=4.25e-07 $layer=LI1_cond $X=2.185 $Y=1.185
+ $X2=1.76 $Y2=1.185
r201 41 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.02
+ $X2=2.17 $Y2=1.185
r202 41 43 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.17 $Y=1.02
+ $X2=2.17 $Y2=0.56
r203 37 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.35
+ $X2=1.76 $Y2=1.185
r204 37 39 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.76 $Y=1.35
+ $X2=1.76 $Y2=1.985
r205 33 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.02
+ $X2=1.725 $Y2=1.185
r206 33 35 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.725 $Y=1.02
+ $X2=1.725 $Y2=0.56
r207 29 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.35
+ $X2=1.33 $Y2=1.185
r208 29 31 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.33 $Y=1.35
+ $X2=1.33 $Y2=1.985
r209 25 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.295 $Y=1.02
+ $X2=1.295 $Y2=1.185
r210 25 27 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.295 $Y=1.02
+ $X2=1.295 $Y2=0.56
r211 21 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=1.35
+ $X2=0.9 $Y2=1.185
r212 21 23 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.9 $Y=1.35
+ $X2=0.9 $Y2=1.985
r213 17 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.865 $Y=1.02
+ $X2=0.865 $Y2=1.185
r214 17 19 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.865 $Y=1.02
+ $X2=0.865 $Y2=0.56
r215 13 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.35
+ $X2=0.47 $Y2=1.185
r216 13 15 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.47 $Y=1.35
+ $X2=0.47 $Y2=1.985
r217 4 63 600 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.485 $X2=3.345 $Y2=1.955
r218 3 75 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.185
+ $Y=0.235 $X2=5.325 $Y2=0.36
r219 2 82 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=3.635
+ $Y=0.235 $X2=3.835 $Y2=0.38
r220 1 67 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.68
+ $Y=0.235 $X2=2.82 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%B1 3 7 11 15 17 18 21 29 30 31 33
c94 30 0 1.9379e-19 $X=4.01 $Y=1.16
c95 29 0 1.31572e-19 $X=4.01 $Y=1.16
c96 18 0 3.37771e-19 $X=2.625 $Y=1.16
c97 17 0 2.25268e-20 $X=2.625 $Y=1.16
c98 11 0 1.86603e-19 $X=4.03 $Y=1.985
c99 3 0 1.02869e-19 $X=2.605 $Y=0.56
r100 29 32 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.01 $Y=1.16
+ $X2=4.01 $Y2=1.35
r101 29 31 47.9601 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.01 $Y=1.16
+ $X2=4.01 $Y2=0.985
r102 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.16 $X2=4.01 $Y2=1.16
r103 21 33 3.9347 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=1.572
+ $X2=3.845 $Y2=1.572
r104 21 30 8.25758 $w=4.83e-07 $l=2.85e-07 $layer=LI1_cond $X=4.01 $Y=1.445
+ $X2=4.01 $Y2=1.16
r105 21 33 0.361551 $w=2.53e-07 $l=8e-09 $layer=LI1_cond $X=3.837 $Y=1.572
+ $X2=3.845 $Y2=1.572
r106 20 21 46.64 $w=2.53e-07 $l=1.032e-06 $layer=LI1_cond $X=2.805 $Y=1.572
+ $X2=3.837 $Y2=1.572
r107 18 27 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.625 $Y=1.16
+ $X2=2.625 $Y2=1.35
r108 18 26 41.84 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.625 $Y=1.16
+ $X2=2.625 $Y2=1.02
r109 17 20 22.8473 $w=2.2e-07 $l=4.12e-07 $layer=LI1_cond $X=2.672 $Y=1.16
+ $X2=2.672 $Y2=1.572
r110 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.16 $X2=2.625 $Y2=1.16
r111 15 31 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.1 $Y=0.56
+ $X2=4.1 $Y2=0.985
r112 11 32 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.03 $Y=1.985
+ $X2=4.03 $Y2=1.35
r113 7 27 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.7 $Y=1.985
+ $X2=2.7 $Y2=1.35
r114 3 26 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.605 $Y=0.56
+ $X2=2.605 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%C1 1 3 6 8 10 13 15
c43 15 0 1.02869e-19 $X=3.455 $Y=1.19
r44 19 21 55.3328 $w=3.65e-07 $l=3.5e-07 $layer=POLY_cond $X=3.13 $Y=1.172
+ $X2=3.48 $Y2=1.172
r45 15 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.48
+ $Y=1.16 $X2=3.48 $Y2=1.16
r46 11 13 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.56 $Y=1.355
+ $X2=3.56 $Y2=1.985
r47 8 11 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.56 $Y=1.172
+ $X2=3.56 $Y2=1.355
r48 8 21 12.6475 $w=3.65e-07 $l=8e-08 $layer=POLY_cond $X=3.56 $Y=1.172 $X2=3.48
+ $Y2=1.172
r49 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.56 $Y=0.99 $X2=3.56
+ $Y2=0.56
r50 4 19 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.13 $Y=1.355
+ $X2=3.13 $Y2=1.172
r51 4 6 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.13 $Y=1.355 $X2=3.13
+ $Y2=1.985
r52 1 19 8.69516 $w=3.65e-07 $l=5.5e-08 $layer=POLY_cond $X=3.075 $Y=1.172
+ $X2=3.13 $Y2=1.172
r53 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.075 $Y=0.99
+ $X2=3.075 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%A2 3 6 10 13 17 18 20 21 26 27 29 34 36 38
c81 29 0 2.26936e-20 $X=5.755 $Y=1.53
c82 17 0 1.86603e-19 $X=4.66 $Y=1.16
c83 6 0 1.9379e-19 $X=4.68 $Y=0.56
r84 29 38 3.24837 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=5.74 $Y=1.605
+ $X2=5.74 $Y2=1.51
r85 29 38 1.74286 $w=2.08e-07 $l=3.3e-08 $layer=LI1_cond $X=5.74 $Y=1.477
+ $X2=5.74 $Y2=1.51
r86 27 37 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=6.06 $Y=1.16 $X2=6.06
+ $Y2=1.35
r87 27 36 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.06 $Y=1.16
+ $X2=6.06 $Y2=1.01
r88 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.06
+ $Y=1.16 $X2=6.06 $Y2=1.16
r89 23 29 8.29177 $w=2.08e-07 $l=1.57e-07 $layer=LI1_cond $X=5.74 $Y=1.32
+ $X2=5.74 $Y2=1.477
r90 22 26 12.2927 $w=2.98e-07 $l=3.2e-07 $layer=LI1_cond $X=5.74 $Y=1.17
+ $X2=6.06 $Y2=1.17
r91 22 23 2.82627 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=5.74 $Y=1.17 $X2=5.74
+ $Y2=1.32
r92 20 29 3.59031 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=5.635 $Y=1.605
+ $X2=5.74 $Y2=1.605
r93 20 21 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=5.635 $Y=1.605
+ $X2=4.825 $Y2=1.605
r94 18 34 59.3261 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.66 $Y=1.16
+ $X2=4.66 $Y2=1.4
r95 18 33 41.84 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.66 $Y=1.16 $X2=4.66
+ $Y2=1.02
r96 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.66
+ $Y=1.16 $X2=4.66 $Y2=1.16
r97 15 21 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=4.66 $Y=1.51
+ $X2=4.825 $Y2=1.605
r98 15 17 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.66 $Y=1.51
+ $X2=4.66 $Y2=1.16
r99 13 37 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.97 $Y=1.985
+ $X2=5.97 $Y2=1.35
r100 10 36 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.97 $Y=0.56 $X2=5.97
+ $Y2=1.01
r101 6 33 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.68 $Y=0.56
+ $X2=4.68 $Y2=1.02
r102 3 34 187.98 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=4.57 $Y=1.985
+ $X2=4.57 $Y2=1.4
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%A1 3 7 11 15 17 24
c49 17 0 1.58656e-19 $X=5.295 $Y=1.19
r50 22 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.2 $Y=1.185
+ $X2=5.54 $Y2=1.185
r51 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.2
+ $Y=1.16 $X2=5.2 $Y2=1.16
r52 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.11 $Y=1.185 $X2=5.2
+ $Y2=1.185
r53 17 23 3.53168 $w=3.08e-07 $l=9.5e-08 $layer=LI1_cond $X=5.295 $Y=1.175
+ $X2=5.2 $Y2=1.175
r54 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=1.35
+ $X2=5.54 $Y2=1.185
r55 13 15 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.54 $Y=1.35
+ $X2=5.54 $Y2=1.985
r56 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=1.02
+ $X2=5.54 $Y2=1.185
r57 9 11 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=5.54 $Y=1.02 $X2=5.54
+ $Y2=0.56
r58 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.11 $Y=1.35
+ $X2=5.11 $Y2=1.185
r59 5 7 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.11 $Y=1.35 $X2=5.11
+ $Y2=1.985
r60 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.11 $Y=1.02
+ $X2=5.11 $Y2=1.185
r61 1 3 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=5.11 $Y=1.02 $X2=5.11
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 39 41
+ 50 57 64 65 71 74 77
c106 5 0 2.26936e-20 $X=5.615 $Y=1.485
c107 1 0 3.98522e-20 $X=0.135 $Y=1.485
r108 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r110 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r111 65 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r112 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r113 62 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=5.755 $Y2=2.72
r114 62 64 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=6.21 $Y2=2.72
r115 61 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r116 61 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r117 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=4.785 $Y2=2.72
r119 58 60 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=5.29 $Y2=2.72
r120 57 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=2.72
+ $X2=5.755 $Y2=2.72
r121 57 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.59 $Y=2.72 $X2=5.29
+ $Y2=2.72
r122 56 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r124 53 56 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=4.37 $Y2=2.72
r125 52 55 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=4.37 $Y2=2.72
r126 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r127 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.785 $Y2=2.72
r128 50 55 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.37 $Y2=2.72
r129 49 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r130 49 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r132 46 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.115 $Y2=2.72
r133 46 48 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.61 $Y2=2.72
r134 45 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r135 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 42 68 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r137 42 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 41 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=2.72
+ $X2=1.115 $Y2=2.72
r139 41 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.95 $Y=2.72
+ $X2=0.69 $Y2=2.72
r140 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r141 39 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r142 37 48 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.81 $Y=2.72 $X2=1.61
+ $Y2=2.72
r143 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=1.935 $Y2=2.72
r144 36 52 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.06 $Y=2.72
+ $X2=2.07 $Y2=2.72
r145 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.06 $Y=2.72
+ $X2=1.935 $Y2=2.72
r146 32 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=2.635
+ $X2=5.755 $Y2=2.72
r147 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.755 $Y=2.635
+ $X2=5.755 $Y2=2.36
r148 28 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.635
+ $X2=4.785 $Y2=2.72
r149 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.785 $Y=2.635
+ $X2=4.785 $Y2=2.36
r150 24 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=2.635
+ $X2=1.935 $Y2=2.72
r151 24 26 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.935 $Y=2.635
+ $X2=1.935 $Y2=2
r152 20 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.635
+ $X2=1.115 $Y2=2.72
r153 20 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.115 $Y=2.635
+ $X2=1.115 $Y2=1.96
r154 16 68 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r155 16 18 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=1.96
r156 5 34 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=5.615
+ $Y=1.485 $X2=5.755 $Y2=2.36
r157 4 30 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.485 $X2=4.785 $Y2=2.36
r158 3 26 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.835
+ $Y=1.485 $X2=1.97 $Y2=2
r159 2 22 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.975
+ $Y=1.485 $X2=1.115 $Y2=1.96
r160 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%X 1 2 3 4 13 15 16 19 21 25 27 31 35 38 39
+ 40 43
c58 40 0 3.98522e-20 $X=0.23 $Y=0.85
r59 40 43 3.30224 $w=2.55e-07 $l=1.2e-07 $layer=LI1_cond $X=0.212 $Y=0.755
+ $X2=0.212 $Y2=0.875
r60 40 43 1.35582 $w=2.53e-07 $l=3e-08 $layer=LI1_cond $X=0.212 $Y=0.905
+ $X2=0.212 $Y2=0.875
r61 37 40 26.6644 $w=2.53e-07 $l=5.9e-07 $layer=LI1_cond $X=0.212 $Y=1.495
+ $X2=0.212 $Y2=0.905
r62 33 35 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.935 $Y=0.615
+ $X2=1.935 $Y2=0.42
r63 29 31 8.75598 $w=1.88e-07 $l=1.5e-07 $layer=LI1_cond $X=1.545 $Y=1.705
+ $X2=1.545 $Y2=1.855
r64 28 39 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=1.175 $Y=0.745
+ $X2=1.08 $Y2=0.745
r65 27 33 7.11373 $w=2.6e-07 $l=1.69115e-07 $layer=LI1_cond $X=1.845 $Y=0.745
+ $X2=1.935 $Y2=0.615
r66 27 28 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=1.845 $Y=0.745
+ $X2=1.175 $Y2=0.745
r67 23 39 2.34704 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=1.08 $Y=0.615
+ $X2=1.08 $Y2=0.745
r68 23 25 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.08 $Y=0.615
+ $X2=1.08 $Y2=0.42
r69 22 38 4.64301 $w=2.1e-07 $l=9.3e-08 $layer=LI1_cond $X=0.78 $Y=1.6 $X2=0.687
+ $Y2=1.6
r70 21 29 6.83868 $w=2.1e-07 $l=1.44914e-07 $layer=LI1_cond $X=1.45 $Y=1.6
+ $X2=1.545 $Y2=1.705
r71 21 22 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.45 $Y=1.6 $X2=0.78
+ $Y2=1.6
r72 17 38 1.80272 $w=1.85e-07 $l=1.05e-07 $layer=LI1_cond $X=0.687 $Y=1.705
+ $X2=0.687 $Y2=1.6
r73 17 19 8.99263 $w=1.83e-07 $l=1.5e-07 $layer=LI1_cond $X=0.687 $Y=1.705
+ $X2=0.687 $Y2=1.855
r74 16 37 6.89985 $w=2.1e-07 $l=1.72696e-07 $layer=LI1_cond $X=0.34 $Y=1.6
+ $X2=0.212 $Y2=1.495
r75 15 38 4.64301 $w=2.1e-07 $l=9.2e-08 $layer=LI1_cond $X=0.595 $Y=1.6
+ $X2=0.687 $Y2=1.6
r76 15 16 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=0.595 $Y=1.6
+ $X2=0.34 $Y2=1.6
r77 14 40 3.52239 $w=2.4e-07 $l=1.28e-07 $layer=LI1_cond $X=0.34 $Y=0.755
+ $X2=0.212 $Y2=0.755
r78 13 39 4.08801 $w=2.5e-07 $l=9.98749e-08 $layer=LI1_cond $X=0.985 $Y=0.755
+ $X2=1.08 $Y2=0.745
r79 13 14 30.9719 $w=2.38e-07 $l=6.45e-07 $layer=LI1_cond $X=0.985 $Y=0.755
+ $X2=0.34 $Y2=0.755
r80 4 31 300 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.545 $Y2=1.855
r81 3 19 300 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.685 $Y2=1.855
r82 2 35 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.8
+ $Y=0.235 $X2=1.94 $Y2=0.42
r83 1 25 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.235 $X2=1.08 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%A_473_297# 1 2 3 4 13 17 21 23 27 31 33 39
+ 40
c67 33 0 1.31572e-19 $X=4.285 $Y=1.992
c68 1 0 1.93402e-19 $X=2.365 $Y=1.485
r69 36 37 11.7689 $w=3.28e-07 $l=3.37e-07 $layer=LI1_cond $X=4.285 $Y=2
+ $X2=4.285 $Y2=2.337
r70 33 36 0.27938 $w=3.28e-07 $l=8e-09 $layer=LI1_cond $X=4.285 $Y=1.992
+ $X2=4.285 $Y2=2
r71 29 40 4.13123 $w=2.92e-07 $l=1.30192e-07 $layer=LI1_cond $X=6.217 $Y=2.105
+ $X2=6.18 $Y2=1.992
r72 29 31 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=6.217 $Y=2.105
+ $X2=6.217 $Y2=2.3
r73 25 40 4.13123 $w=2.92e-07 $l=1.12e-07 $layer=LI1_cond $X=6.18 $Y=1.88
+ $X2=6.18 $Y2=1.992
r74 25 27 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.18 $Y=1.88
+ $X2=6.18 $Y2=1.63
r75 24 39 5.81644 $w=2.25e-07 $l=1.3e-07 $layer=LI1_cond $X=5.42 $Y=1.992
+ $X2=5.29 $Y2=1.992
r76 23 40 2.30226 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=1.992
+ $X2=6.18 $Y2=1.992
r77 23 24 30.4757 $w=2.23e-07 $l=5.95e-07 $layer=LI1_cond $X=6.015 $Y=1.992
+ $X2=5.42 $Y2=1.992
r78 19 39 0.827476 $w=2.6e-07 $l=1.13e-07 $layer=LI1_cond $X=5.29 $Y=2.105
+ $X2=5.29 $Y2=1.992
r79 19 21 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=5.29 $Y=2.105
+ $X2=5.29 $Y2=2.3
r80 18 33 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=4.45 $Y=1.992
+ $X2=4.285 $Y2=1.992
r81 17 39 5.81644 $w=2.25e-07 $l=1.3e-07 $layer=LI1_cond $X=5.16 $Y=1.992
+ $X2=5.29 $Y2=1.992
r82 17 18 36.366 $w=2.23e-07 $l=7.1e-07 $layer=LI1_cond $X=5.16 $Y=1.992
+ $X2=4.45 $Y2=1.992
r83 13 37 2.26808 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=2.337
+ $X2=4.285 $Y2=2.337
r84 13 15 73.666 $w=2.53e-07 $l=1.63e-06 $layer=LI1_cond $X=4.12 $Y=2.337
+ $X2=2.49 $Y2=2.337
r85 4 31 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.485 $X2=6.18 $Y2=2.3
r86 4 27 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.485 $X2=6.18 $Y2=1.63
r87 3 21 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.485 $X2=5.325 $Y2=2.3
r88 2 36 300 $w=1.7e-07 $l=5.98268e-07 $layer=licon1_PDIFF $count=2 $X=4.105
+ $Y=1.485 $X2=4.285 $Y2=2
r89 1 15 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=1.485 $X2=2.49 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_4%VGND 1 2 3 4 5 6 21 25 29 33 35 37 40 41 43
+ 44 46 47 48 50 65 69 78 82 89
r112 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r113 82 85 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.375
+ $Y2=0.36
r114 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r115 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 76 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r117 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r118 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r119 73 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r120 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r121 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r122 70 82 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.375
+ $Y2=0
r123 70 72 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.83
+ $Y2=0
r124 69 88 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=6.015 $Y=0
+ $X2=6.227 $Y2=0
r125 69 75 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.015 $Y=0
+ $X2=5.75 $Y2=0
r126 68 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r127 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r128 65 82 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.375
+ $Y2=0
r129 65 67 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=3.91
+ $Y2=0
r130 64 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r131 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r132 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r133 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r134 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r135 58 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r136 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r137 55 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.65
+ $Y2=0
r138 55 57 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0
+ $X2=1.15 $Y2=0
r139 50 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.485 $Y=0 $X2=0.65
+ $Y2=0
r140 50 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.23 $Y2=0
r141 48 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r142 48 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r143 46 63 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=2.99
+ $Y2=0
r144 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.305
+ $Y2=0
r145 45 67 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.91
+ $Y2=0
r146 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.305
+ $Y2=0
r147 43 60 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.07
+ $Y2=0
r148 43 44 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.387
+ $Y2=0
r149 42 63 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.555 $Y=0
+ $X2=2.99 $Y2=0
r150 42 44 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.555 $Y=0
+ $X2=2.387 $Y2=0
r151 40 57 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.345 $Y=0
+ $X2=1.15 $Y2=0
r152 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.51
+ $Y2=0
r153 39 60 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.675 $Y=0
+ $X2=2.07 $Y2=0
r154 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.51
+ $Y2=0
r155 35 88 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.227 $Y2=0
r156 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.18 $Y2=0.38
r157 31 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0
r158 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0.36
r159 27 44 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.387 $Y=0.085
+ $X2=2.387 $Y2=0
r160 27 29 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=2.387 $Y=0.085
+ $X2=2.387 $Y2=0.36
r161 23 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0
r162 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0.36
r163 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.085
+ $X2=0.65 $Y2=0
r164 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.65 $Y=0.085
+ $X2=0.65 $Y2=0.38
r165 6 37 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.38
r166 5 85 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.235 $X2=4.355 $Y2=0.36
r167 4 33 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.235 $X2=3.305 $Y2=0.36
r168 3 29 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.39 $Y2=0.36
r169 2 25 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.37
+ $Y=0.235 $X2=1.51 $Y2=0.36
r170 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.525
+ $Y=0.235 $X2=0.65 $Y2=0.38
.ends


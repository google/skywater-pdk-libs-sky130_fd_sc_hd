* File: sky130_fd_sc_hd__lpflow_inputisolatch_1.spice.pex
* Created: Thu Aug 27 14:25:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%SLEEP_B 4 5 7 8 10 13 17 19
+ 22 24 28
c40 13 0 2.71124e-20 $X=0.47 $Y=0.805
r41 22 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r42 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r43 22 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r44 19 28 2.01678 $w=2.38e-07 $l=4.2e-08 $layer=LI1_cond $X=0.21 $Y=1.277
+ $X2=0.21 $Y2=1.235
r45 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.75
+ $X2=0.47 $Y2=1.75
r46 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r47 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.825
+ $X2=0.47 $Y2=1.75
r48 8 10 114.073 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.47 $Y=1.825
+ $X2=0.47 $Y2=2.18
r49 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r50 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r51 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.675
+ $X2=0.305 $Y2=1.75
r52 4 25 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.305 $Y=1.675
+ $X2=0.305 $Y2=1.4
r53 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r54 1 24 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_27_47# 1 2 9 13 17 19 20 23
+ 27 30 34 36 37 38 39 43 46 47 50 52 54 57 58 59 61
c138 57 0 8.48005e-20 $X=2.25 $Y=1.52
c139 23 0 1.50999e-19 $X=2.8 $Y=0.415
r140 61 66 10.4675 $w=3.78e-07 $l=1.00623e-07 $layer=POLY_cond $X=0.965 $Y=1.415
+ $X2=0.89 $Y2=1.355
r141 57 59 9.65825 $w=3.38e-07 $l=2e-07 $layer=LI1_cond $X=2.25 $Y=1.525
+ $X2=2.05 $Y2=1.525
r142 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.52 $X2=2.25 $Y2=1.52
r143 53 66 21.0397 $w=3.78e-07 $l=1.65e-07 $layer=POLY_cond $X=0.725 $Y=1.355
+ $X2=0.89 $Y2=1.355
r144 52 55 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.46
r145 52 54 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.13
r146 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.295 $X2=0.725 $Y2=1.295
r147 50 59 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.49 $Y=1.61
+ $X2=2.05 $Y2=1.61
r148 47 61 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=1.405 $Y=1.415
+ $X2=0.965 $Y2=1.415
r149 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=1.415 $X2=1.405 $Y2=1.415
r150 44 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.525
+ $X2=1.49 $Y2=1.61
r151 44 46 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.405 $Y=1.525
+ $X2=1.405 $Y2=1.415
r152 43 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.46
r153 40 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.13
r154 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r155 38 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r156 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r157 36 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r158 32 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.965
+ $X2=0.345 $Y2=1.88
r159 32 34 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=1.965
+ $X2=0.26 $Y2=2.175
r160 28 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r161 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r162 26 58 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.25 $Y=1.55 $X2=2.25
+ $Y2=1.52
r163 26 27 40.8463 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.55
+ $X2=2.25 $Y2=1.685
r164 25 58 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.25 $Y=1.395
+ $X2=2.25 $Y2=1.52
r165 21 23 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.8 $Y=1.245
+ $X2=2.8 $Y2=0.415
r166 20 25 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.385 $Y=1.32
+ $X2=2.25 $Y2=1.395
r167 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.725 $Y=1.32
+ $X2=2.8 $Y2=1.245
r168 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.725 $Y=1.32
+ $X2=2.385 $Y2=1.32
r169 17 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.305 $Y=2.275
+ $X2=2.305 $Y2=1.685
r170 11 66 24.4846 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=0.89 $Y=1.58
+ $X2=0.89 $Y2=1.355
r171 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.89 $Y=1.58 $X2=0.89
+ $Y2=2.18
r172 7 66 24.4846 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=0.89 $Y=1.13
+ $X2=0.89 $Y2=1.355
r173 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.89 $Y=1.13
+ $X2=0.89 $Y2=0.445
r174 2 34 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.905 $X2=0.26 $Y2=2.175
r175 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%D 3 6 8 11 13 18
c43 18 0 1.50999e-19 $X=1.92 $Y=0.925
c44 13 0 1.25524e-19 $X=1.835 $Y=0.73
r45 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=0.93
+ $X2=1.835 $Y2=1.095
r46 11 13 56.192 $w=2.7e-07 $l=2e-07 $layer=POLY_cond $X=1.835 $Y=0.93 $X2=1.835
+ $Y2=0.73
r47 8 18 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.93
+ $X2=1.92 $Y2=0.93
r48 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=0.93 $X2=1.835 $Y2=0.93
r49 6 14 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.83 $Y=2.165
+ $X2=1.83 $Y2=1.095
r50 3 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=0.445 $X2=1.83
+ $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_193_47# 1 2 9 12 15 18 20
+ 23 28 32 34 37 38 39 43
c119 38 0 8.48005e-20 $X=2.76 $Y=1.74
c120 34 0 1.25524e-19 $X=2.59 $Y=0.87
c121 32 0 2.94334e-20 $X=2.38 $Y=0.87
r122 38 47 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=1.74
+ $X2=2.76 $Y2=1.875
r123 37 40 8.8128 $w=3.38e-07 $l=2.6e-07 $layer=LI1_cond $X=2.675 $Y=1.74
+ $X2=2.675 $Y2=2
r124 37 39 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=1.74
+ $X2=2.675 $Y2=1.575
r125 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=1.74 $X2=2.76 $Y2=1.74
r126 32 43 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=2.372 $Y=0.87
+ $X2=2.372 $Y2=0.705
r127 31 34 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.38 $Y=0.87
+ $X2=2.59 $Y2=0.87
r128 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=0.87 $X2=2.38 $Y2=0.87
r129 27 28 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=1.082 $Y=0.74
+ $X2=1.082 $Y2=0.91
r130 25 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=1.035
+ $X2=2.59 $Y2=0.87
r131 25 39 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.59 $Y=1.035
+ $X2=2.59 $Y2=1.575
r132 24 29 1.32297 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.185 $Y=2
+ $X2=1.082 $Y2=2
r133 23 40 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.505 $Y=2 $X2=2.675
+ $Y2=2
r134 23 24 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=2.505 $Y=2
+ $X2=1.185 $Y2=2
r135 20 29 5.65333 $w=1.88e-07 $l=9.35682e-08 $layer=LI1_cond $X=1.1 $Y=2.085
+ $X2=1.082 $Y2=2
r136 20 22 6.45882 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.1 $Y=2.085 $X2=1.1
+ $Y2=2.175
r137 18 27 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.1 $Y=0.51 $X2=1.1
+ $Y2=0.74
r138 15 29 11.4938 $w=1.88e-07 $l=1.83303e-07 $layer=LI1_cond $X=1.065 $Y=1.825
+ $X2=1.082 $Y2=2
r139 15 28 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.065 $Y=1.825
+ $X2=1.065 $Y2=0.91
r140 12 47 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.725 $Y=2.275
+ $X2=2.725 $Y2=1.875
r141 9 43 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.415
+ $X2=2.305 $Y2=0.705
r142 2 22 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.905 $X2=1.1 $Y2=2.175
r143 1 18 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_629_21# 1 2 9 13 15 18 23
+ 25 29
c58 29 0 1.92048e-19 $X=3.96 $Y=1.755
r59 25 27 8.35559 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.98 $Y=0.58
+ $X2=3.98 $Y2=0.745
r60 23 29 6.84016 $w=2.32e-07 $l=1.9139e-07 $layer=LI1_cond $X=4.037 $Y=1.535
+ $X2=3.98 $Y2=1.7
r61 23 27 50.0675 $w=1.73e-07 $l=7.9e-07 $layer=LI1_cond $X=4.037 $Y=1.535
+ $X2=4.037 $Y2=0.745
r62 18 30 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.505 $Y=1.7
+ $X2=3.22 $Y2=1.7
r63 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.505
+ $Y=1.7 $X2=3.505 $Y2=1.7
r64 15 29 0.117566 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=3.835 $Y=1.7
+ $X2=3.98 $Y2=1.7
r65 15 17 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.835 $Y=1.7
+ $X2=3.505 $Y2=1.7
r66 11 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.865
+ $X2=3.22 $Y2=1.7
r67 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.22 $Y=1.865
+ $X2=3.22 $Y2=2.275
r68 7 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.535
+ $X2=3.22 $Y2=1.7
r69 7 9 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=3.22 $Y=1.535
+ $X2=3.22 $Y2=0.415
r70 2 29 300 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=2 $X=3.835
+ $Y=1.485 $X2=3.96 $Y2=1.755
r71 1 25 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=3.96 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_476_47# 1 2 7 9 12 14 16 19
+ 21 23 25 29 34 35 36 39
c100 35 0 1.83571e-19 $X=3.1 $Y=1.325
c101 19 0 1.92048e-19 $X=4.59 $Y=1.985
r102 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.16 $X2=3.695 $Y2=1.16
r103 37 39 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.185 $Y=1.16
+ $X2=3.695 $Y2=1.16
r104 35 37 9.3849 $w=2.44e-07 $l=1.98167e-07 $layer=LI1_cond $X=3.1 $Y=1.325
+ $X2=3.027 $Y2=1.16
r105 35 36 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.1 $Y=1.325
+ $X2=3.1 $Y2=2.255
r106 34 37 9.3849 $w=2.44e-07 $l=1.9775e-07 $layer=LI1_cond $X=2.955 $Y=0.995
+ $X2=3.027 $Y2=1.16
r107 33 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.955 $Y=0.535
+ $X2=2.955 $Y2=0.995
r108 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.87 $Y=0.45
+ $X2=2.955 $Y2=0.535
r109 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.87 $Y=0.45
+ $X2=2.585 $Y2=0.45
r110 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=2.34
+ $X2=3.1 $Y2=2.255
r111 25 27 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.015 $Y=2.34
+ $X2=2.515 $Y2=2.34
r112 22 23 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.17 $Y=1.16
+ $X2=4.59 $Y2=1.16
r113 21 40 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=4.095 $Y=1.16
+ $X2=3.695 $Y2=1.16
r114 21 22 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.095 $Y=1.16
+ $X2=4.17 $Y2=1.16
r115 17 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.16
r116 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.985
r117 14 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=1.16
r118 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=0.56
r119 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=1.325
+ $X2=4.17 $Y2=1.16
r120 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.17 $Y=1.325
+ $X2=4.17 $Y2=1.985
r121 7 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=0.995
+ $X2=4.17 $Y2=1.16
r122 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.17 $Y=0.995
+ $X2=4.17 $Y2=0.56
r123 2 27 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=2.065 $X2=2.515 $Y2=2.34
r124 1 31 182 $w=1.7e-07 $l=3.005e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.585 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%VPWR 1 2 3 4 15 19 21 25 27
+ 29 34 39 49 50 53 56 63 66
r76 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r77 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r78 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r79 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r81 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r82 47 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=2.72
+ $X2=4.38 $Y2=2.72
r83 47 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.465 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 46 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r87 43 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r88 42 45 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r89 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r90 40 42 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=2.07 $Y2=2.72
r91 39 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=2.72
+ $X2=3.44 $Y2=2.72
r92 39 45 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.355 $Y=2.72
+ $X2=2.99 $Y2=2.72
r93 38 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 38 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r96 35 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r97 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 34 40 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.652 $Y=2.72
+ $X2=1.85 $Y2=2.72
r99 34 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r100 34 56 11.0868 $w=3.93e-07 $l=3.8e-07 $layer=LI1_cond $X=1.652 $Y=2.72
+ $X2=1.652 $Y2=2.34
r101 34 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r102 29 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r103 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r104 27 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r106 23 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=2.635
+ $X2=4.38 $Y2=2.72
r107 23 25 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=4.38 $Y=2.635
+ $X2=4.38 $Y2=1.735
r108 22 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.72
+ $X2=3.44 $Y2=2.72
r109 21 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=4.38 $Y2=2.72
r110 21 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=3.525 $Y2=2.72
r111 17 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=2.635
+ $X2=3.44 $Y2=2.72
r112 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.44 $Y=2.635
+ $X2=3.44 $Y2=2.3
r113 13 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r114 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r115 4 25 300 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=2 $X=4.245
+ $Y=1.485 $X2=4.38 $Y2=1.735
r116 3 19 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=2.065 $X2=3.44 $Y2=2.3
r117 2 56 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=2.34
r118 1 15 600 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.905 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%Q 1 2 9 10 11 19 30
r12 28 30 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.89 $Y=0.745
+ $X2=4.89 $Y2=1.67
r13 16 19 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=4.832 $Y=1.812
+ $X2=4.832 $Y2=1.835
r14 10 16 0.566112 $w=2.83e-07 $l=1.4e-08 $layer=LI1_cond $X=4.832 $Y=1.798
+ $X2=4.832 $Y2=1.812
r15 10 30 7.03738 $w=2.83e-07 $l=1.28e-07 $layer=LI1_cond $X=4.832 $Y=1.798
+ $X2=4.832 $Y2=1.67
r16 10 11 13.2228 $w=2.83e-07 $l=3.27e-07 $layer=LI1_cond $X=4.832 $Y=1.883
+ $X2=4.832 $Y2=2.21
r17 10 19 1.94096 $w=2.83e-07 $l=4.8e-08 $layer=LI1_cond $X=4.832 $Y=1.883
+ $X2=4.832 $Y2=1.835
r18 9 28 11.3641 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=4.832 $Y=0.51
+ $X2=4.832 $Y2=0.745
r19 2 19 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=4.665
+ $Y=1.485 $X2=4.8 $Y2=1.835
r20 1 9 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=4.665
+ $Y=0.235 $X2=4.8 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%VGND 1 2 3 4 15 19 23 25 29
+ 31 33 38 43 53 54 57 60 63 66
c78 54 0 2.71124e-20 $X=4.83 $Y=0
r79 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r80 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r81 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r82 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r83 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r84 54 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r85 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r86 51 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.38
+ $Y2=0
r87 51 53 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.83
+ $Y2=0
r88 50 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r89 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r90 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r91 47 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r92 46 49 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r93 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r94 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r95 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=2.07
+ $Y2=0
r96 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.43
+ $Y2=0
r97 43 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=2.99
+ $Y2=0
r98 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r99 42 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r100 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r101 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r102 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r103 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r104 38 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r105 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r106 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r107 31 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r108 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r109 27 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=0.085
+ $X2=4.38 $Y2=0
r110 27 29 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.38 $Y=0.085
+ $X2=4.38 $Y2=0.55
r111 26 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0 $X2=3.43
+ $Y2=0
r112 25 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.38
+ $Y2=0
r113 25 26 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.295 $Y=0 $X2=3.595
+ $Y2=0
r114 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=0.085
+ $X2=3.43 $Y2=0
r115 21 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.43 $Y=0.085
+ $X2=3.43 $Y2=0.445
r116 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r117 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.38
r118 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r119 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r120 4 29 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=4.245
+ $Y=0.235 $X2=4.38 $Y2=0.55
r121 3 23 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.295
+ $Y=0.235 $X2=3.43 $Y2=0.445
r122 2 19 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r123 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


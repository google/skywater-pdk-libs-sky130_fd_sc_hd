* File: sky130_fd_sc_hd__and2b_2.pex.spice
* Created: Thu Aug 27 14:07:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND2B_2%A_N 3 7 9 12 17 22
c30 12 0 1.89169e-19 $X=0.365 $Y=1.16
r31 13 22 1.15244 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=0.3 $Y=1.16 $X2=0.3
+ $Y2=1.19
r32 13 17 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.3 $Y=1.16 $X2=0.3
+ $Y2=0.85
r33 12 15 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.372 $Y=1.16
+ $X2=0.372 $Y2=1.325
r34 12 14 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.372 $Y=1.16
+ $X2=0.372 $Y2=0.995
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.365
+ $Y=1.16 $X2=0.365 $Y2=1.16
r36 9 22 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.3 $Y=1.53 $X2=0.3
+ $Y2=1.19
r37 7 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r38 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_2%A_27_413# 1 2 9 13 17 19 20 22 24 26 33 34
c63 33 0 1.2595e-19 $X=1.09 $Y=0.97
c64 19 0 3.48245e-19 $X=0.62 $Y=1.9
c65 9 0 1.69139e-19 $X=0.985 $Y=2.275
r66 34 36 19.6163 $w=2.58e-07 $l=1.05e-07 $layer=POLY_cond $X=1.09 $Y=0.97
+ $X2=0.985 $Y2=0.97
r67 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=0.97 $X2=1.09 $Y2=0.97
r68 31 33 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=0.737 $Y=0.97
+ $X2=1.09 $Y2=0.97
r69 29 31 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.727 $Y=0.97
+ $X2=0.737 $Y2=0.97
r70 26 28 10.235 $w=2.38e-07 $l=2.1e-07 $layer=LI1_cond $X=0.715 $Y=0.445
+ $X2=0.715 $Y2=0.655
r71 23 31 2.74472 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=0.737 $Y=1.135
+ $X2=0.737 $Y2=0.97
r72 23 24 31.8761 $w=2.33e-07 $l=6.5e-07 $layer=LI1_cond $X=0.737 $Y=1.135
+ $X2=0.737 $Y2=1.785
r73 22 29 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=0.727 $Y=0.805
+ $X2=0.727 $Y2=0.97
r74 22 28 8.0403 $w=2.13e-07 $l=1.5e-07 $layer=LI1_cond $X=0.727 $Y=0.805
+ $X2=0.727 $Y2=0.655
r75 19 24 6.81752 $w=2.3e-07 $l=1.64754e-07 $layer=LI1_cond $X=0.62 $Y=1.9
+ $X2=0.737 $Y2=1.785
r76 19 20 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.62 $Y=1.9
+ $X2=0.345 $Y2=1.9
r77 15 20 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.345 $Y2=1.9
r78 15 17 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.26 $Y2=2.225
r79 11 34 59.7829 $w=2.58e-07 $l=3.93954e-07 $layer=POLY_cond $X=1.41 $Y=0.805
+ $X2=1.09 $Y2=0.97
r80 11 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.41 $Y=0.805
+ $X2=1.41 $Y2=0.445
r81 7 36 15.449 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.135
+ $X2=0.985 $Y2=0.97
r82 7 9 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=0.985 $Y=1.135
+ $X2=0.985 $Y2=2.275
r83 2 17 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.225
r84 1 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_2%B 1 3 7 9 19
c32 19 0 1.69139e-19 $X=2.095 $Y=1.87
c33 7 0 2.58024e-19 $X=1.83 $Y=0.445
c34 1 0 1.16262e-19 $X=1.425 $Y=1.895
r35 13 19 15.7996 $w=3.08e-07 $l=4.25e-07 $layer=LI1_cond $X=1.67 $Y=1.8
+ $X2=2.095 $Y2=1.8
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.73 $X2=1.67 $Y2=1.73
r37 9 13 1.30115 $w=3.08e-07 $l=3.5e-08 $layer=LI1_cond $X=1.635 $Y=1.8 $X2=1.67
+ $Y2=1.8
r38 5 12 83.3829 $w=4.52e-07 $l=6.58726e-07 $layer=POLY_cond $X=1.83 $Y=1.165
+ $X2=1.627 $Y2=1.73
r39 5 7 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.83 $Y=1.165 $X2=1.83
+ $Y2=0.445
r40 1 12 40.728 $w=4.52e-07 $l=2.72276e-07 $layer=POLY_cond $X=1.425 $Y=1.895
+ $X2=1.627 $Y2=1.73
r41 1 3 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.425 $Y=1.895
+ $X2=1.425 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_2%A_212_413# 1 2 7 9 12 14 16 19 23 26 27 29
+ 35 40
r77 39 40 71.2817 $w=3.4e-07 $l=4.2e-07 $layer=POLY_cond $X=2.32 $Y=1.155
+ $X2=2.74 $Y2=1.155
r78 35 36 10.9609 $w=2.56e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=0.44 $X2=1.43
+ $Y2=0.44
r79 30 39 11.8803 $w=3.4e-07 $l=7e-08 $layer=POLY_cond $X=2.25 $Y=1.155 $X2=2.32
+ $Y2=1.155
r80 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r81 27 33 14.4021 $w=4.04e-07 $l=5.11126e-07 $layer=LI1_cond $X=1.905 $Y=1.135
+ $X2=1.43 $Y2=1.21
r82 27 29 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=1.905 $Y=1.135
+ $X2=2.25 $Y2=1.135
r83 26 33 5.83894 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.43 $Y=0.945
+ $X2=1.43 $Y2=1.21
r84 25 36 3.13337 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.43 $Y=0.61 $X2=1.43
+ $Y2=0.44
r85 25 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.43 $Y=0.61
+ $X2=1.43 $Y2=0.945
r86 21 33 7.33812 $w=4.04e-07 $l=3.66906e-07 $layer=LI1_cond $X=1.187 $Y=1.475
+ $X2=1.43 $Y2=1.21
r87 21 23 30.3274 $w=2.83e-07 $l=7.5e-07 $layer=LI1_cond $X=1.187 $Y=1.475
+ $X2=1.187 $Y2=2.225
r88 17 40 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.74 $Y=1.325
+ $X2=2.74 $Y2=1.155
r89 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.74 $Y=1.325
+ $X2=2.74 $Y2=1.985
r90 14 40 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.74 $Y=0.985
+ $X2=2.74 $Y2=1.155
r91 14 16 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.74 $Y=0.985
+ $X2=2.74 $Y2=0.56
r92 10 39 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.32 $Y=1.325
+ $X2=2.32 $Y2=1.155
r93 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.32 $Y=1.325
+ $X2=2.32 $Y2=1.985
r94 7 39 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.32 $Y=0.985
+ $X2=2.32 $Y2=1.155
r95 7 9 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.32 $Y=0.985
+ $X2=2.32 $Y2=0.56
r96 2 23 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=2.065 $X2=1.205 $Y2=2.225
r97 1 35 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_2%VPWR 1 2 3 12 14 16 18 20 30 36 40 44 47
c42 47 0 1.16262e-19 $X=2.99 $Y=2.72
c43 40 0 1.59076e-19 $X=1.51 $Y=2.485
r44 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 42 44 9.66931 $w=6.38e-07 $l=1.25e-07 $layer=LI1_cond $X=2.07 $Y=2.485
+ $X2=2.195 $Y2=2.485
r46 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 39 42 0.840993 $w=6.38e-07 $l=4.5e-08 $layer=LI1_cond $X=2.025 $Y=2.485
+ $X2=2.07 $Y2=2.485
r48 39 40 16.9579 $w=6.38e-07 $l=5.15e-07 $layer=LI1_cond $X=2.025 $Y=2.485
+ $X2=1.51 $Y2=2.485
r49 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 34 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 33 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.195 $Y2=2.72
r53 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 30 46 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.042 $Y2=2.72
r55 30 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 29 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 29 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 28 40 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=1.51 $Y2=2.72
r59 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r61 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 20 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r63 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 14 46 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=3 $Y=2.635
+ $X2=3.042 $Y2=2.72
r67 14 16 33.0794 $w=2.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3 $Y=2.635 $X2=3
+ $Y2=1.86
r68 10 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r69 10 12 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.27
r70 3 16 300 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_PDIFF $count=2 $X=2.815
+ $Y=1.485 $X2=2.95 $Y2=1.86
r71 2 39 300 $w=1.7e-07 $l=6.44011e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.065 $X2=2.025 $Y2=2.33
r72 1 12 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_2%X 1 2 7 9 14 15 16 17 21
c24 15 0 1.32074e-19 $X=2.527 $Y=1.58
r25 17 21 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.527 $Y=2.21
+ $X2=2.527 $Y2=1.835
r26 15 16 51.0182 $w=1.73e-07 $l=8.05e-07 $layer=LI1_cond $X=2.592 $Y=1.58
+ $X2=2.592 $Y2=0.775
r27 14 21 3.89186 $w=3.03e-07 $l=1.03e-07 $layer=LI1_cond $X=2.527 $Y=1.732
+ $X2=2.527 $Y2=1.835
r28 14 15 7.81944 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=2.527 $Y=1.732
+ $X2=2.527 $Y2=1.58
r29 7 16 6.51365 $w=2.33e-07 $l=1.17e-07 $layer=LI1_cond $X=2.562 $Y=0.658
+ $X2=2.562 $Y2=0.775
r30 7 9 7.6834 $w=2.35e-07 $l=1.48e-07 $layer=LI1_cond $X=2.562 $Y=0.658
+ $X2=2.562 $Y2=0.51
r31 2 21 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=2.395
+ $Y=1.485 $X2=2.53 $Y2=1.835
r32 1 9 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.53 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_2%VGND 1 2 3 10 12 16 18 20 22 24 32 41 45
r43 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r44 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r45 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r46 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r47 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r48 33 41 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.075
+ $Y2=0
r49 33 35 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.53
+ $Y2=0
r50 32 44 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.042
+ $Y2=0
r51 32 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.53
+ $Y2=0
r52 31 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r53 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r54 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r55 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r56 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 25 38 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r58 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r59 24 41 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.075
+ $Y2=0
r60 24 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.61
+ $Y2=0
r61 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r62 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r63 18 44 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=3 $Y=0.085
+ $X2=3.042 $Y2=0
r64 18 20 19.8476 $w=2.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0.55
r65 14 41 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0
r66 14 16 11.0923 $w=3.98e-07 $l=3.85e-07 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0.47
r67 10 38 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r68 10 12 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.445
r69 3 20 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.235 $X2=2.95 $Y2=0.55
r70 2 16 182 $w=1.7e-07 $l=3.21559e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.11 $Y2=0.47
r71 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends


* File: sky130_fd_sc_hd__einvn_0.pxi.spice
* Created: Thu Aug 27 14:20:01 2020
* 
x_PM_SKY130_FD_SC_HD__EINVN_0%A_30_47# N_A_30_47#_M1003_s N_A_30_47#_M1000_s
+ N_A_30_47#_M1001_g N_A_30_47#_c_42_n N_A_30_47#_c_47_n N_A_30_47#_c_43_n
+ N_A_30_47#_c_44_n N_A_30_47#_c_48_n N_A_30_47#_c_49_n N_A_30_47#_c_45_n
+ N_A_30_47#_c_46_n PM_SKY130_FD_SC_HD__EINVN_0%A_30_47#
x_PM_SKY130_FD_SC_HD__EINVN_0%TE_B N_TE_B_M1003_g N_TE_B_c_105_n N_TE_B_M1000_g
+ N_TE_B_c_107_n N_TE_B_c_108_n N_TE_B_M1004_g N_TE_B_c_109_n TE_B TE_B
+ N_TE_B_c_103_n N_TE_B_c_104_n PM_SKY130_FD_SC_HD__EINVN_0%TE_B
x_PM_SKY130_FD_SC_HD__EINVN_0%A N_A_M1002_g N_A_M1005_g A A A A N_A_c_149_n
+ PM_SKY130_FD_SC_HD__EINVN_0%A
x_PM_SKY130_FD_SC_HD__EINVN_0%VPWR N_VPWR_M1000_d VPWR N_VPWR_c_175_n
+ N_VPWR_c_176_n N_VPWR_c_174_n N_VPWR_c_178_n PM_SKY130_FD_SC_HD__EINVN_0%VPWR
x_PM_SKY130_FD_SC_HD__EINVN_0%Z N_Z_M1002_d N_Z_M1005_d N_Z_c_205_n Z Z
+ PM_SKY130_FD_SC_HD__EINVN_0%Z
x_PM_SKY130_FD_SC_HD__EINVN_0%VGND N_VGND_M1003_d VGND N_VGND_c_238_n
+ N_VGND_c_239_n N_VGND_c_240_n N_VGND_c_241_n PM_SKY130_FD_SC_HD__EINVN_0%VGND
cc_1 VNB N_A_30_47#_M1001_g 0.0267695f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.445
cc_2 VNB N_A_30_47#_c_42_n 0.0159507f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=0.445
cc_3 VNB N_A_30_47#_c_43_n 0.00856323f $X=-0.19 $Y=-0.24 $X2=0.82 $Y2=0.74
cc_4 VNB N_A_30_47#_c_44_n 0.0101187f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=0.74
cc_5 VNB N_A_30_47#_c_45_n 0.00173964f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_6 VNB N_A_30_47#_c_46_n 0.0244492f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.16
cc_7 VNB N_TE_B_M1003_g 0.038184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_TE_B_c_103_n 0.0243362f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.98
cc_9 VNB N_TE_B_c_104_n 0.0183506f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.825
cc_10 VNB N_A_M1002_g 0.0318754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A 0.0234834f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.445
cc_12 VNB N_A_c_149_n 0.0344588f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=0.74
cc_13 VNB N_VPWR_c_174_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Z_c_205_n 0.0037736f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.445
cc_15 VNB Z 0.0152137f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.445
cc_16 VNB N_VGND_c_238_n 0.0146769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_239_n 0.0224494f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=0.445
cc_18 VNB N_VGND_c_240_n 0.123471f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_241_n 0.00669024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VPB N_A_30_47#_c_47_n 0.0161948f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=2.275
cc_21 VPB N_A_30_47#_c_48_n 0.00153627f $X=-0.19 $Y=1.305 $X2=0.82 $Y2=1.98
cc_22 VPB N_A_30_47#_c_49_n 0.0105622f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.98
cc_23 VPB N_A_30_47#_c_45_n 0.00451862f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_24 VPB N_A_30_47#_c_46_n 0.00643061f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.16
cc_25 VPB N_TE_B_c_105_n 0.021447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_TE_B_M1000_g 0.0344174f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.445
cc_27 VPB N_TE_B_c_107_n 0.028068f $X=-0.19 $Y=1.305 $X2=0.222 $Y2=0.655
cc_28 VPB N_TE_B_c_108_n 0.013884f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=0.445
cc_29 VPB N_TE_B_c_109_n 0.00785214f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=2.275
cc_30 VPB N_TE_B_c_103_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.98
cc_31 VPB N_TE_B_c_104_n 0.0235142f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.825
cc_32 VPB N_A_M1005_g 0.0430028f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.995
cc_33 VPB A 0.0303472f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.445
cc_34 VPB N_A_c_149_n 0.0113274f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=0.74
cc_35 VPB N_VPWR_c_175_n 0.0166274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_176_n 0.022446f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=0.445
cc_37 VPB N_VPWR_c_174_n 0.0435071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_178_n 0.00975765f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=2.275
cc_39 VPB N_Z_c_205_n 0.00363985f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.445
cc_40 VPB Z 0.0152667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 N_A_30_47#_M1001_g N_TE_B_M1003_g 0.0174446f $X=1 $Y=0.445 $X2=0 $Y2=0
cc_42 N_A_30_47#_c_43_n N_TE_B_M1003_g 0.0134831f $X=0.82 $Y=0.74 $X2=0 $Y2=0
cc_43 N_A_30_47#_c_45_n N_TE_B_M1003_g 0.00326217f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_44 N_A_30_47#_c_45_n N_TE_B_c_105_n 0.00166067f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_45 N_A_30_47#_c_48_n N_TE_B_M1000_g 0.0138582f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_46 N_A_30_47#_c_45_n N_TE_B_M1000_g 0.00239355f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_47 N_A_30_47#_c_48_n N_TE_B_c_107_n 0.00609313f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_48 N_A_30_47#_c_45_n N_TE_B_c_107_n 0.00901904f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_49 N_A_30_47#_c_46_n N_TE_B_c_107_n 0.0148379f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_50 N_A_30_47#_c_48_n N_TE_B_c_108_n 0.00560034f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_51 N_A_30_47#_c_45_n N_TE_B_c_108_n 0.00256028f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_30_47#_c_43_n N_TE_B_c_103_n 3.50292e-19 $X=0.82 $Y=0.74 $X2=0 $Y2=0
cc_53 N_A_30_47#_c_44_n N_TE_B_c_103_n 5.4318e-19 $X=0.36 $Y=0.74 $X2=0 $Y2=0
cc_54 N_A_30_47#_c_49_n N_TE_B_c_103_n 3.75655e-19 $X=0.4 $Y=1.98 $X2=0 $Y2=0
cc_55 N_A_30_47#_c_45_n N_TE_B_c_103_n 3.21458e-19 $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_30_47#_c_46_n N_TE_B_c_103_n 0.0203531f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_30_47#_c_43_n N_TE_B_c_104_n 0.0229013f $X=0.82 $Y=0.74 $X2=0 $Y2=0
cc_58 N_A_30_47#_c_44_n N_TE_B_c_104_n 0.0250203f $X=0.36 $Y=0.74 $X2=0 $Y2=0
cc_59 N_A_30_47#_c_48_n N_TE_B_c_104_n 0.0192863f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_60 N_A_30_47#_c_49_n N_TE_B_c_104_n 0.0290371f $X=0.4 $Y=1.98 $X2=0 $Y2=0
cc_61 N_A_30_47#_c_45_n N_TE_B_c_104_n 0.0583396f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_30_47#_c_46_n N_TE_B_c_104_n 0.0021586f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_30_47#_M1001_g N_A_M1002_g 0.0368418f $X=1 $Y=0.445 $X2=0 $Y2=0
cc_64 N_A_30_47#_c_45_n N_A_M1002_g 4.32419e-19 $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_30_47#_c_45_n N_A_M1005_g 0.00177767f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_30_47#_c_46_n N_A_c_149_n 0.0368418f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_30_47#_c_48_n N_VPWR_M1000_d 0.00447929f $X=0.82 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_68 N_A_30_47#_c_45_n N_VPWR_M1000_d 6.08718e-19 $X=0.905 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_69 N_A_30_47#_c_47_n N_VPWR_c_175_n 0.0202523f $X=0.275 $Y=2.275 $X2=0 $Y2=0
cc_70 N_A_30_47#_c_48_n N_VPWR_c_175_n 0.00268635f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_71 N_A_30_47#_M1000_s N_VPWR_c_174_n 0.00213257f $X=0.15 $Y=2.065 $X2=0 $Y2=0
cc_72 N_A_30_47#_c_47_n N_VPWR_c_174_n 0.011999f $X=0.275 $Y=2.275 $X2=0 $Y2=0
cc_73 N_A_30_47#_c_48_n N_VPWR_c_174_n 0.00580114f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_74 N_A_30_47#_c_48_n N_VPWR_c_178_n 0.02623f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_75 N_A_30_47#_M1001_g N_Z_c_205_n 0.00529098f $X=1 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_30_47#_c_43_n N_Z_c_205_n 0.0135843f $X=0.82 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_30_47#_c_48_n N_Z_c_205_n 0.0133617f $X=0.82 $Y=1.98 $X2=0 $Y2=0
cc_78 N_A_30_47#_c_45_n N_Z_c_205_n 0.077436f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_30_47#_M1001_g Z 0.00459872f $X=1 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A_30_47#_c_43_n N_VGND_M1003_d 0.00112182f $X=0.82 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_30_47#_c_42_n N_VGND_c_238_n 0.0188331f $X=0.275 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_30_47#_c_43_n N_VGND_c_238_n 0.00274327f $X=0.82 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A_30_47#_M1001_g N_VGND_c_239_n 0.00331718f $X=1 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_30_47#_M1003_s N_VGND_c_240_n 0.00229009f $X=0.15 $Y=0.235 $X2=0 $Y2=0
cc_85 N_A_30_47#_M1001_g N_VGND_c_240_n 0.00571831f $X=1 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_30_47#_c_42_n N_VGND_c_240_n 0.0104656f $X=0.275 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_30_47#_c_43_n N_VGND_c_240_n 0.00619211f $X=0.82 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_30_47#_M1001_g N_VGND_c_241_n 0.0104712f $X=1 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_30_47#_c_43_n N_VGND_c_241_n 0.0312427f $X=0.82 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_30_47#_c_46_n N_VGND_c_241_n 3.98347e-19 $X=1 $Y=1.16 $X2=0 $Y2=0
cc_91 N_TE_B_c_107_n N_A_M1005_g 0.0604941f $X=0.925 $Y=1.695 $X2=0 $Y2=0
cc_92 N_TE_B_M1000_g N_VPWR_c_175_n 0.00428022f $X=0.485 $Y=2.275 $X2=0 $Y2=0
cc_93 N_TE_B_c_108_n N_VPWR_c_176_n 0.00331718f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_94 N_TE_B_M1000_g N_VPWR_c_174_n 0.00689596f $X=0.485 $Y=2.275 $X2=0 $Y2=0
cc_95 N_TE_B_c_108_n N_VPWR_c_174_n 0.00571831f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_96 N_TE_B_M1000_g N_VPWR_c_178_n 0.00333954f $X=0.485 $Y=2.275 $X2=0 $Y2=0
cc_97 N_TE_B_c_107_n N_VPWR_c_178_n 3.55564e-19 $X=0.925 $Y=1.695 $X2=0 $Y2=0
cc_98 N_TE_B_c_108_n N_VPWR_c_178_n 0.0102986f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_99 N_TE_B_c_107_n N_Z_c_205_n 0.00402483f $X=0.925 $Y=1.695 $X2=0 $Y2=0
cc_100 N_TE_B_c_108_n Z 0.00459872f $X=1 $Y=1.77 $X2=0 $Y2=0
cc_101 N_TE_B_M1003_g N_VGND_c_238_n 0.00342417f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_102 N_TE_B_M1003_g N_VGND_c_240_n 0.00503181f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_103 N_TE_B_M1003_g N_VGND_c_241_n 0.00895265f $X=0.485 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_M1005_g N_VPWR_c_176_n 0.00357877f $X=1.36 $Y=2.165 $X2=0 $Y2=0
cc_105 N_A_M1005_g N_VPWR_c_174_n 0.00605429f $X=1.36 $Y=2.165 $X2=0 $Y2=0
cc_106 N_A_M1005_g N_VPWR_c_178_n 0.00154135f $X=1.36 $Y=2.165 $X2=0 $Y2=0
cc_107 A N_Z_M1005_d 0.0040972f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_108 N_A_M1002_g N_Z_c_205_n 0.0121716f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_M1005_g N_Z_c_205_n 0.0224863f $X=1.36 $Y=2.165 $X2=0 $Y2=0
cc_110 A N_Z_c_205_n 0.0864191f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A_c_149_n N_Z_c_205_n 0.00753413f $X=1.585 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_M1002_g Z 0.0128944f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_113 A Z 0.0213772f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_114 N_A_c_149_n Z 0.00215351f $X=1.585 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_M1005_g Z 0.0128944f $X=1.36 $Y=2.165 $X2=0 $Y2=0
cc_116 A Z 0.0210557f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_117 N_A_M1002_g N_VGND_c_239_n 0.00357877f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_118 N_A_M1002_g N_VGND_c_240_n 0.00605429f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A_M1002_g N_VGND_c_241_n 0.00154984f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_120 N_VPWR_c_174_n A_215_369# 0.0046292f $X=1.61 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_121 N_VPWR_c_174_n N_Z_M1005_d 0.00209344f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_122 N_VPWR_c_176_n Z 0.0356686f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_123 N_VPWR_c_174_n Z 0.0217421f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_124 N_VPWR_c_178_n Z 0.0190336f $X=0.745 $Y=2.36 $X2=0 $Y2=0
cc_125 A_215_369# N_Z_c_205_n 0.00263752f $X=1.075 $Y=1.845 $X2=0.23 $Y2=2.72
cc_126 A_215_369# Z 0.00418839f $X=1.075 $Y=1.845 $X2=0 $Y2=0
cc_127 Z N_VGND_c_239_n 0.0357322f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_128 N_Z_M1002_d N_VGND_c_240_n 0.00209344f $X=1.435 $Y=0.235 $X2=0 $Y2=0
cc_129 Z N_VGND_c_240_n 0.0217513f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_130 Z N_VGND_c_241_n 0.0191591f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_131 N_Z_c_205_n A_215_47# 8.57924e-19 $X=1.245 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_132 Z A_215_47# 0.00419798f $X=1.525 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_133 N_VGND_c_240_n A_215_47# 0.0046292f $X=1.61 $Y=0 $X2=-0.19 $Y2=-0.24

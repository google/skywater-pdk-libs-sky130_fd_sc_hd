* File: sky130_fd_sc_hd__nand2_1.spice.SKY130_FD_SC_HD__NAND2_1.pxi
* Created: Thu Aug 27 14:28:37 2020
* 
x_PM_SKY130_FD_SC_HD__NAND2_1%B N_B_c_28_n N_B_M1002_g N_B_M1000_g B N_B_c_30_n
+ PM_SKY130_FD_SC_HD__NAND2_1%B
x_PM_SKY130_FD_SC_HD__NAND2_1%A N_A_c_51_n N_A_M1001_g N_A_M1003_g A N_A_c_53_n
+ PM_SKY130_FD_SC_HD__NAND2_1%A
x_PM_SKY130_FD_SC_HD__NAND2_1%VPWR N_VPWR_M1000_s N_VPWR_M1003_d N_VPWR_c_75_n
+ N_VPWR_c_76_n N_VPWR_c_77_n N_VPWR_c_78_n VPWR N_VPWR_c_79_n N_VPWR_c_74_n
+ PM_SKY130_FD_SC_HD__NAND2_1%VPWR
x_PM_SKY130_FD_SC_HD__NAND2_1%Y N_Y_M1001_d N_Y_M1000_d N_Y_c_99_n N_Y_c_100_n Y
+ Y N_Y_c_97_n PM_SKY130_FD_SC_HD__NAND2_1%Y
x_PM_SKY130_FD_SC_HD__NAND2_1%VGND N_VGND_M1002_s N_VGND_c_119_n N_VGND_c_120_n
+ VGND N_VGND_c_121_n N_VGND_c_122_n VGND PM_SKY130_FD_SC_HD__NAND2_1%VGND
cc_1 VNB N_B_c_28_n 0.0221895f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB B 0.00939618f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_B_c_30_n 0.0392248f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_4 VNB N_A_c_51_n 0.0221092f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_5 VNB A 0.00855647f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_6 VNB N_A_c_53_n 0.0379831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_VPWR_c_74_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB Y 0.00767174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_Y_c_97_n 0.0276701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_119_n 0.0108751f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_11 VNB N_VGND_c_120_n 0.0328324f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_12 VNB N_VGND_c_121_n 0.0268118f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_13 VNB N_VGND_c_122_n 0.10356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VPB N_B_M1000_g 0.0262407f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_15 VPB B 8.02347e-19 $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_16 VPB N_B_c_30_n 0.0107397f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_17 VPB N_A_M1003_g 0.0262424f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_18 VPB A 7.09926e-19 $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_19 VPB N_A_c_53_n 0.010214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_75_n 0.0102689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_76_n 0.0438743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_77_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_78_n 0.0426603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_79_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_VPWR_c_74_n 0.0419516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB Y 0.00312356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 N_B_c_28_n N_A_c_51_n 0.0217282f $X=0.49 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_28 N_B_M1000_g N_A_M1003_g 0.0217282f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_29 N_B_c_30_n N_A_c_53_n 0.0217282f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_30 N_B_M1000_g N_VPWR_c_76_n 0.00322755f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_31 B N_VPWR_c_76_n 0.0217832f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_32 N_B_c_30_n N_VPWR_c_76_n 0.00601529f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_33 N_B_M1000_g N_VPWR_c_79_n 0.00541359f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_34 N_B_M1000_g N_VPWR_c_74_n 0.0105016f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_35 N_B_M1000_g N_Y_c_99_n 0.00359531f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_36 N_B_M1000_g N_Y_c_100_n 0.00918977f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_37 N_B_c_28_n Y 0.0103495f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_38 B Y 0.0202615f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_39 N_B_c_28_n N_VGND_c_120_n 0.00480583f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_40 B N_VGND_c_120_n 0.0228794f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_41 N_B_c_30_n N_VGND_c_120_n 0.0071164f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_42 N_B_c_28_n N_VGND_c_121_n 0.00585385f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_43 N_B_c_28_n N_VGND_c_122_n 0.0115388f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_44 N_A_M1003_g N_VPWR_c_78_n 0.00321781f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_45 A N_VPWR_c_78_n 0.0191448f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_46 N_A_c_53_n N_VPWR_c_78_n 0.00554938f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_47 N_A_M1003_g N_VPWR_c_79_n 0.00541359f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_48 N_A_M1003_g N_VPWR_c_74_n 0.0104829f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_49 N_A_M1003_g N_Y_c_99_n 0.00288872f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A_M1003_g N_Y_c_100_n 0.00918977f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_51 N_A_c_51_n Y 0.010245f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_52 A Y 0.0187498f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_53 N_A_c_51_n N_Y_c_97_n 0.0211238f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_54 A N_Y_c_97_n 0.0222128f $X=1.06 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A_c_53_n N_Y_c_97_n 0.00712397f $X=1.105 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_c_51_n N_VGND_c_121_n 0.00357877f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_57 N_A_c_51_n N_VGND_c_122_n 0.00620762f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_58 N_VPWR_c_74_n N_Y_M1000_d 0.00215201f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_59 N_VPWR_c_79_n N_Y_c_100_n 0.0189039f $X=1.035 $Y=2.72 $X2=0 $Y2=0
cc_60 N_VPWR_c_74_n N_Y_c_100_n 0.0122217f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_61 N_VPWR_c_78_n N_Y_c_97_n 7.22395e-19 $X=1.12 $Y=1.66 $X2=0 $Y2=0
cc_62 N_VPWR_c_76_n N_VGND_c_120_n 3.44647e-19 $X=0.28 $Y=1.66 $X2=0 $Y2=0
cc_63 N_Y_c_97_n N_VGND_c_121_n 0.0433462f $X=1.12 $Y=0.38 $X2=0 $Y2=0
cc_64 N_Y_M1001_d N_VGND_c_122_n 0.00209344f $X=0.985 $Y=0.235 $X2=0 $Y2=0
cc_65 N_Y_c_97_n N_VGND_c_122_n 0.0259387f $X=1.12 $Y=0.38 $X2=0 $Y2=0
cc_66 Y A_113_47# 4.34665e-19 $X=0.6 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_67 N_Y_c_97_n A_113_47# 0.00325659f $X=1.12 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_68 N_VGND_c_122_n A_113_47# 0.00338335f $X=1.15 $Y=0 $X2=-0.19 $Y2=-0.24

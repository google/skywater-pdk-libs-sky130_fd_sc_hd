* File: sky130_fd_sc_hd__dlclkp_1.pex.spice
* Created: Thu Aug 27 14:16:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%CLK 4 5 7 8 10 13 17 21 25 27 29 30 33 36
+ 37 40 42 45
c135 37 0 1.36988e-19 $X=5.295 $Y=1.19
c136 33 0 6.03924e-20 $X=0.23 $Y=1.19
c137 21 0 9.76047e-20 $X=0.47 $Y=0.805
r138 45 48 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.27
+ $X2=5.38 $Y2=1.435
r139 45 47 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.27
+ $X2=5.38 $Y2=1.105
r140 40 43 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r141 40 42 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r142 37 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.325
+ $Y=1.27 $X2=5.325 $Y2=1.27
r143 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.295 $Y=1.19
+ $X2=5.295 $Y2=1.19
r144 33 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r145 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=1.19
+ $X2=0.23 $Y2=1.19
r146 30 32 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=0.38 $Y=1.19
+ $X2=0.23 $Y2=1.19
r147 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.15 $Y=1.19
+ $X2=5.295 $Y2=1.19
r148 29 30 5.90345 $w=1.4e-07 $l=4.77e-06 $layer=MET1_cond $X=5.15 $Y=1.19
+ $X2=0.38 $Y2=1.19
r149 27 33 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.53
+ $X2=0.207 $Y2=1.19
r150 23 25 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r151 19 21 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r152 17 48 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.495 $Y=2.165
+ $X2=5.495 $Y2=1.435
r153 13 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.495 $Y=0.445
+ $X2=5.495 $Y2=1.105
r154 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=1.665
r155 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r156 5 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.47 $Y2=0.805
r157 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r158 4 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r159 4 43 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r160 1 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r161 1 42 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%GATE 1 3 5 7 8 10 11 12
r44 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.52 $X2=1.765 $Y2=1.52
r45 11 12 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.085 $Y=0.51
+ $X2=2.085 $Y2=0.85
r46 10 18 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=1.61 $Y=1.56
+ $X2=1.765 $Y2=1.56
r47 9 12 32.4409 $w=1.98e-07 $l=5.85e-07 $layer=LI1_cond $X=2.085 $Y=1.435
+ $X2=2.085 $Y2=0.85
r48 8 18 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=1.985 $Y=1.56
+ $X2=1.765 $Y2=1.56
r49 8 9 6.92652 $w=2.5e-07 $l=1.67705e-07 $layer=LI1_cond $X=1.985 $Y=1.56
+ $X2=2.085 $Y2=1.435
r50 5 17 93.6423 $w=2.38e-07 $l=4.77389e-07 $layer=POLY_cond $X=1.905 $Y=1.09
+ $X2=1.805 $Y2=1.52
r51 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.905 $Y=1.09 $X2=1.905
+ $Y2=0.805
r52 1 17 39.9742 $w=2.38e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.83 $Y=1.685
+ $X2=1.805 $Y2=1.52
r53 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.83 $Y=1.685 $X2=1.83
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%A_193_47# 1 2 9 13 17 21 26 27 28 30 34 41
c94 30 0 2.04326e-19 $X=3.055 $Y=0.9
c95 21 0 4.39096e-20 $X=2.39 $Y=1.94
c96 17 0 7.04924e-20 $X=1.1 $Y=0.425
r97 31 41 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=3.055 $Y=0.9
+ $X2=3.18 $Y2=0.9
r98 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.055
+ $Y=0.9 $X2=3.055 $Y2=0.9
r99 28 30 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.59 $Y=0.9
+ $X2=3.055 $Y2=0.9
r100 27 35 37.7695 $w=2.7e-07 $l=1.7e-07 $layer=POLY_cond $X=2.475 $Y=1.74
+ $X2=2.305 $Y2=1.74
r101 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.475
+ $Y=1.74 $X2=2.475 $Y2=1.74
r102 24 26 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=2.49 $Y=1.855
+ $X2=2.49 $Y2=1.74
r103 23 28 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.49 $Y=0.985
+ $X2=2.59 $Y2=0.9
r104 23 26 41.8682 $w=1.98e-07 $l=7.55e-07 $layer=LI1_cond $X=2.49 $Y=0.985
+ $X2=2.49 $Y2=1.74
r105 22 34 2.68609 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.28 $Y=1.94
+ $X2=1.147 $Y2=1.94
r106 21 24 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.39 $Y=1.94
+ $X2=2.49 $Y2=1.855
r107 21 22 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.39 $Y=1.94
+ $X2=1.28 $Y2=1.94
r108 15 34 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.147 $Y=1.855
+ $X2=1.147 $Y2=1.94
r109 15 17 62.1884 $w=2.63e-07 $l=1.43e-06 $layer=LI1_cond $X=1.147 $Y=1.855
+ $X2=1.147 $Y2=0.425
r110 11 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=0.765
+ $X2=3.18 $Y2=0.9
r111 11 13 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.18 $Y=0.765
+ $X2=3.18 $Y2=0.43
r112 7 35 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.305 $Y=1.875
+ $X2=2.305 $Y2=1.74
r113 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.305 $Y=1.875
+ $X2=2.305 $Y2=2.275
r114 2 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r115 1 17 182 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%A_27_47# 1 2 7 9 11 14 16 19 20 21 25 26 27
+ 30 32 35 39 40 41 46 48 50 52 56
c134 27 0 4.39096e-20 $X=2.53 $Y=1.32
c135 14 0 2.6965e-20 $X=0.89 $Y=2.135
c136 11 0 3.34275e-20 $X=0.89 $Y=1.09
r137 51 56 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.225
+ $X2=0.89 $Y2=1.225
r138 50 53 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.225
+ $X2=0.725 $Y2=1.39
r139 50 52 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.225
+ $X2=0.725 $Y2=1.06
r140 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.225 $X2=0.755 $Y2=1.225
r141 46 53 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.39
r142 43 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.695 $Y=0.785
+ $X2=0.695 $Y2=1.06
r143 42 48 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r144 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r145 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r146 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.7
+ $X2=0.695 $Y2=0.785
r147 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.7
+ $X2=0.345 $Y2=0.7
r148 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.345 $Y2=0.7
r149 33 35 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.26 $Y2=0.425
r150 28 30 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.925 $Y=1.395
+ $X2=2.925 $Y2=2.275
r151 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.85 $Y=1.32
+ $X2=2.925 $Y2=1.395
r152 26 27 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.85 $Y=1.32
+ $X2=2.53 $Y2=1.32
r153 23 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.455 $Y=1.245
+ $X2=2.53 $Y2=1.32
r154 23 25 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.455 $Y=1.245
+ $X2=2.455 $Y2=0.54
r155 22 25 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.455 $Y=0.255
+ $X2=2.455 $Y2=0.54
r156 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.38 $Y=0.18
+ $X2=2.455 $Y2=0.255
r157 20 21 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.38 $Y=0.18
+ $X2=1.45 $Y2=0.18
r158 18 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.375 $Y=0.255
+ $X2=1.45 $Y2=0.18
r159 18 19 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.375 $Y=0.255
+ $X2=1.375 $Y2=0.73
r160 17 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.965 $Y=0.805
+ $X2=0.89 $Y2=0.805
r161 16 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.3 $Y=0.805
+ $X2=1.375 $Y2=0.73
r162 16 17 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.3 $Y=0.805
+ $X2=0.965 $Y2=0.805
r163 12 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.36
+ $X2=0.89 $Y2=1.225
r164 12 14 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=0.89 $Y=1.36
+ $X2=0.89 $Y2=2.135
r165 11 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.09
+ $X2=0.89 $Y2=1.225
r166 10 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=0.88
+ $X2=0.89 $Y2=0.805
r167 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.89 $Y=0.88
+ $X2=0.89 $Y2=1.09
r168 7 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=0.73
+ $X2=0.89 $Y2=0.805
r169 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.89 $Y=0.73 $X2=0.89
+ $Y2=0.445
r170 2 48 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r171 1 35 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%A_642_307# 1 2 9 13 15 17 19 21 23 24 31 36
+ 39 42 46 48 53
c109 53 0 7.10306e-21 $X=3.655 $Y=1.7
c110 46 0 1.11073e-19 $X=4.655 $Y=1.16
c111 19 0 3.19209e-20 $X=5.06 $Y=0.805
c112 15 0 1.95495e-19 $X=4.71 $Y=1.325
c113 13 0 1.97223e-19 $X=3.655 $Y=0.445
r114 47 55 79.2176 $w=2.16e-07 $l=3.55e-07 $layer=POLY_cond $X=4.655 $Y=1.16
+ $X2=4.655 $Y2=0.805
r115 46 49 4.89946 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=4.542 $Y=1.16
+ $X2=4.542 $Y2=1.325
r116 46 48 6.68973 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=4.542 $Y=1.16
+ $X2=4.542 $Y2=0.995
r117 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.655
+ $Y=1.16 $X2=4.655 $Y2=1.16
r118 44 48 18.6352 $w=2.33e-07 $l=3.8e-07 $layer=LI1_cond $X=4.462 $Y=0.615
+ $X2=4.462 $Y2=0.995
r119 42 44 7.44435 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.45 $Y=0.45
+ $X2=4.45 $Y2=0.615
r120 37 39 0.196141 $w=3.11e-07 $l=5e-09 $layer=LI1_cond $X=4.02 $Y=1.7
+ $X2=4.025 $Y2=1.7
r121 36 39 19.6926 $w=3.11e-07 $l=5.02e-07 $layer=LI1_cond $X=4.527 $Y=1.7
+ $X2=4.025 $Y2=1.7
r122 36 49 6.63049 $w=3.63e-07 $l=2.1e-07 $layer=LI1_cond $X=4.527 $Y=1.535
+ $X2=4.527 $Y2=1.325
r123 29 37 2.76503 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=1.865
+ $X2=4.02 $Y2=1.7
r124 29 31 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.02 $Y=1.865
+ $X2=4.02 $Y2=2.27
r125 27 53 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.515 $Y=1.7
+ $X2=3.655 $Y2=1.7
r126 27 50 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.515 $Y=1.7
+ $X2=3.285 $Y2=1.7
r127 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.515
+ $Y=1.7 $X2=3.515 $Y2=1.7
r128 24 37 4.12156 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.91 $Y=1.7 $X2=4.02
+ $Y2=1.7
r129 24 26 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.91 $Y=1.7
+ $X2=3.515 $Y2=1.7
r130 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.135 $Y=0.73
+ $X2=5.135 $Y2=0.445
r131 20 55 11.3495 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.79 $Y=0.805
+ $X2=4.655 $Y2=0.805
r132 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.06 $Y=0.805
+ $X2=5.135 $Y2=0.73
r133 19 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.06 $Y=0.805
+ $X2=4.79 $Y2=0.805
r134 15 47 41.3672 $w=2.16e-07 $l=1.90526e-07 $layer=POLY_cond $X=4.71 $Y=1.325
+ $X2=4.655 $Y2=1.16
r135 15 17 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.71 $Y=1.325
+ $X2=4.71 $Y2=2.165
r136 11 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.535
+ $X2=3.655 $Y2=1.7
r137 11 13 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.655 $Y=1.535
+ $X2=3.655 $Y2=0.445
r138 7 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.865
+ $X2=3.285 $Y2=1.7
r139 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.285 $Y=1.865
+ $X2=3.285 $Y2=2.275
r140 2 39 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.485 $X2=4.025 $Y2=1.755
r141 2 31 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.485 $X2=4.025 $Y2=2.27
r142 1 42 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.235 $X2=4.405 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%A_476_413# 1 2 9 12 14 18 23 24 25 27 30 31
+ 33 35
c89 33 0 1.67255e-19 $X=3.64 $Y=1.16
r90 31 36 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=4.132 $Y=1.16
+ $X2=4.132 $Y2=1.325
r91 31 35 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=4.132 $Y=1.16
+ $X2=4.132 $Y2=0.995
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.16 $X2=4.09 $Y2=1.16
r93 28 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=1.16
+ $X2=3.64 $Y2=1.16
r94 28 30 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.725 $Y=1.16
+ $X2=4.09 $Y2=1.16
r95 27 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=0.995
+ $X2=3.64 $Y2=1.16
r96 26 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.64 $Y=0.56
+ $X2=3.64 $Y2=0.995
r97 24 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.555 $Y=1.24
+ $X2=3.64 $Y2=1.16
r98 24 25 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.555 $Y=1.24
+ $X2=3.225 $Y2=1.24
r99 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.14 $Y=1.325
+ $X2=3.225 $Y2=1.24
r100 22 23 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.14 $Y=1.325
+ $X2=3.14 $Y2=2.255
r101 18 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.555 $Y=0.475
+ $X2=3.64 $Y2=0.56
r102 18 20 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.555 $Y=0.475
+ $X2=2.955 $Y2=0.475
r103 14 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.055 $Y=2.34
+ $X2=3.14 $Y2=2.255
r104 14 16 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.055 $Y=2.34
+ $X2=2.64 $Y2=2.34
r105 12 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.235 $Y=1.985
+ $X2=4.235 $Y2=1.325
r106 9 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.195 $Y=0.56
+ $X2=4.195 $Y2=0.995
r107 2 16 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=2.065 $X2=2.64 $Y2=2.34
r108 1 20 182 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.33 $X2=2.955 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%A_957_369# 1 2 9 12 15 18 20 21 22 23 27 28
+ 30 32 35 37
c79 35 0 1.35749e-19 $X=5.875 $Y=1.325
c80 12 0 1.05068e-19 $X=5.97 $Y=1.985
r81 32 34 7.09737 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.997 $Y=0.455
+ $X2=4.997 $Y2=0.62
r82 30 35 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.835 $Y=1.725
+ $X2=5.835 $Y2=1.325
r83 28 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.16
+ $X2=5.915 $Y2=1.325
r84 28 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.16
+ $X2=5.915 $Y2=0.995
r85 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.915
+ $Y=1.16 $X2=5.915 $Y2=1.16
r86 25 35 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.875 $Y=1.2
+ $X2=5.875 $Y2=1.325
r87 25 27 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=5.875 $Y=1.2 $X2=5.875
+ $Y2=1.16
r88 24 27 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=5.875 $Y=0.935
+ $X2=5.875 $Y2=1.16
r89 22 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.75 $Y=1.81
+ $X2=5.835 $Y2=1.725
r90 22 23 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.75 $Y=1.81
+ $X2=5.335 $Y2=1.81
r91 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.75 $Y=0.85
+ $X2=5.875 $Y2=0.935
r92 20 21 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.75 $Y=0.85
+ $X2=5.155 $Y2=0.85
r93 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.17 $Y=1.895
+ $X2=5.335 $Y2=1.81
r94 16 18 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.17 $Y=1.895
+ $X2=5.17 $Y2=2
r95 15 21 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.045 $Y=0.765
+ $X2=5.155 $Y2=0.85
r96 15 34 7.59565 $w=2.18e-07 $l=1.45e-07 $layer=LI1_cond $X=5.045 $Y=0.765
+ $X2=5.045 $Y2=0.62
r97 12 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.97 $Y=1.985
+ $X2=5.97 $Y2=1.325
r98 9 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.97 $Y=0.56 $X2=5.97
+ $Y2=0.995
r99 2 18 300 $w=1.7e-07 $l=4.55961e-07 $layer=licon1_PDIFF $count=2 $X=4.785
+ $Y=1.845 $X2=5.17 $Y2=2
r100 1 32 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=4.8
+ $Y=0.235 $X2=4.925 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%VPWR 1 2 3 4 5 18 22 26 28 32 36 38 40 45
+ 50 55 62 63 66 69 72 75 78
c92 32 0 1.95495e-19 $X=4.46 $Y=2.27
r93 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r94 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r95 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r96 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r97 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r98 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r99 63 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r100 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r101 60 78 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=5.745 $Y2=2.72
r102 60 62 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=6.21 $Y2=2.72
r103 59 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r104 59 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r105 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r106 56 75 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=4.452 $Y2=2.72
r107 56 58 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=5.29 $Y2=2.72
r108 55 78 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.57 $Y=2.72
+ $X2=5.745 $Y2=2.72
r109 55 58 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.57 $Y=2.72
+ $X2=5.29 $Y2=2.72
r110 54 73 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r111 54 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r112 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r113 51 69 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.632 $Y2=2.72
r114 51 53 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=2.07 $Y2=2.72
r115 50 72 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.395 $Y=2.72
+ $X2=3.545 $Y2=2.72
r116 50 53 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.395 $Y=2.72
+ $X2=2.07 $Y2=2.72
r117 49 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r118 49 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r121 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r122 45 69 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=1.632 $Y2=2.72
r123 45 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.45 $Y=2.72 $X2=1.15
+ $Y2=2.72
r124 40 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r125 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 38 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r127 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r128 34 78 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=2.635
+ $X2=5.745 $Y2=2.72
r129 34 36 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.745 $Y=2.635
+ $X2=5.745 $Y2=2.295
r130 30 75 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.452 $Y=2.635
+ $X2=4.452 $Y2=2.72
r131 30 32 14.7594 $w=2.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.452 $Y=2.635
+ $X2=4.452 $Y2=2.27
r132 29 72 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.545 $Y2=2.72
r133 28 75 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.31 $Y=2.72
+ $X2=4.452 $Y2=2.72
r134 28 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.31 $Y=2.72
+ $X2=3.695 $Y2=2.72
r135 24 72 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=2.635
+ $X2=3.545 $Y2=2.72
r136 24 26 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.545 $Y=2.635
+ $X2=3.545 $Y2=2.3
r137 20 69 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.632 $Y=2.635
+ $X2=1.632 $Y2=2.72
r138 20 22 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.632 $Y=2.635
+ $X2=1.632 $Y2=2.34
r139 16 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r140 16 18 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r141 5 36 600 $w=1.7e-07 $l=5.36656e-07 $layer=licon1_PDIFF $count=1 $X=5.57
+ $Y=1.845 $X2=5.76 $Y2=2.295
r142 4 32 600 $w=1.7e-07 $l=8.56723e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.485 $X2=4.46 $Y2=2.27
r143 3 26 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=2.065 $X2=3.495 $Y2=2.3
r144 2 22 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=2.34
r145 1 18 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%GCLK 1 2 8 9 10 11 12 18 31
r17 11 12 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=6.222 $Y=1.87
+ $X2=6.222 $Y2=2.21
r18 11 18 9.13257 $w=2.63e-07 $l=2.1e-07 $layer=LI1_cond $X=6.222 $Y=1.87
+ $X2=6.222 $Y2=1.66
r19 10 31 1.76256 $w=3.38e-07 $l=5.2e-08 $layer=LI1_cond $X=6.21 $Y=0.425
+ $X2=6.262 $Y2=0.425
r20 10 31 4.31807 $w=1.85e-07 $l=1.7e-07 $layer=LI1_cond $X=6.262 $Y=0.595
+ $X2=6.262 $Y2=0.425
r21 10 27 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=6.21 $Y=0.425 $X2=6.18
+ $Y2=0.425
r22 9 10 34.6875 $w=3.08e-07 $l=9e-07 $layer=LI1_cond $X=6.262 $Y=1.495
+ $X2=6.262 $Y2=0.595
r23 8 18 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=6.222 $Y=1.627
+ $X2=6.222 $Y2=1.66
r24 8 9 6.80323 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=6.222 $Y=1.627
+ $X2=6.222 $Y2=1.495
r25 2 18 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=6.045
+ $Y=1.485 $X2=6.18 $Y2=1.66
r26 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_1%VGND 1 2 3 4 15 19 23 27 29 31 36 41 46 53
+ 54 57 60 63 66
c97 54 0 2.71124e-20 $X=6.21 $Y=0
r98 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r99 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r100 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r101 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r102 54 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r103 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r104 51 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.84 $Y=0 $X2=5.755
+ $Y2=0
r105 51 53 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.84 $Y=0 $X2=6.21
+ $Y2=0
r106 50 67 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.75 $Y2=0
r107 50 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r108 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r109 47 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.145 $Y=0 $X2=4.02
+ $Y2=0
r110 47 49 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.145 $Y=0
+ $X2=4.37 $Y2=0
r111 46 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=0 $X2=5.755
+ $Y2=0
r112 46 49 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=5.67 $Y=0 $X2=4.37
+ $Y2=0
r113 45 64 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.91 $Y2=0
r114 45 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r115 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r116 42 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.645
+ $Y2=0
r117 42 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=2.07
+ $Y2=0
r118 41 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.02
+ $Y2=0
r119 41 44 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=2.07 $Y2=0
r120 40 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r121 40 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r122 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r123 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r124 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r125 36 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.645
+ $Y2=0
r126 36 39 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.15
+ $Y2=0
r127 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r128 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r129 29 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r130 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r131 25 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0
r132 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0.38
r133 21 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r134 21 23 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.445
r135 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0
r136 17 19 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0.74
r137 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r138 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r139 4 27 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=5.57
+ $Y=0.235 $X2=5.755 $Y2=0.38
r140 3 23 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.985 $Y2=0.445
r141 2 19 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.525
+ $Y=0.595 $X2=1.65 $Y2=0.74
r142 1 15 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


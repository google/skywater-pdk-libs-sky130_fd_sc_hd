* NGSPICE file created from sky130_fd_sc_hd__inv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=7.9e+11p ps=7.58e+06u
M1001 VPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=3.51e+11p ps=3.68e+06u
M1003 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


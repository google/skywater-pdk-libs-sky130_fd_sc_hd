* File: sky130_fd_sc_hd__o21bai_1.pxi.spice
* Created: Thu Aug 27 14:36:23 2020
* 
x_PM_SKY130_FD_SC_HD__O21BAI_1%B1_N N_B1_N_M1007_g N_B1_N_c_58_n N_B1_N_c_59_n
+ N_B1_N_c_60_n N_B1_N_c_61_n N_B1_N_M1005_g N_B1_N_c_55_n N_B1_N_c_56_n B1_N
+ N_B1_N_c_57_n PM_SKY130_FD_SC_HD__O21BAI_1%B1_N
x_PM_SKY130_FD_SC_HD__O21BAI_1%A_105_352# N_A_105_352#_M1007_d
+ N_A_105_352#_M1005_s N_A_105_352#_c_97_n N_A_105_352#_M1002_g
+ N_A_105_352#_M1000_g N_A_105_352#_c_98_n N_A_105_352#_c_99_n
+ N_A_105_352#_c_107_n N_A_105_352#_c_100_n N_A_105_352#_c_108_n
+ N_A_105_352#_c_101_n N_A_105_352#_c_102_n N_A_105_352#_c_103_n
+ PM_SKY130_FD_SC_HD__O21BAI_1%A_105_352#
x_PM_SKY130_FD_SC_HD__O21BAI_1%A2 N_A2_M1001_g N_A2_M1006_g A2 N_A2_c_164_n
+ N_A2_c_165_n N_A2_c_166_n PM_SKY130_FD_SC_HD__O21BAI_1%A2
x_PM_SKY130_FD_SC_HD__O21BAI_1%A1 N_A1_M1003_g N_A1_M1004_g A1 N_A1_c_202_n
+ N_A1_c_203_n PM_SKY130_FD_SC_HD__O21BAI_1%A1
x_PM_SKY130_FD_SC_HD__O21BAI_1%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_227_n
+ N_VPWR_c_228_n N_VPWR_c_229_n VPWR N_VPWR_c_230_n N_VPWR_c_231_n
+ N_VPWR_c_232_n N_VPWR_c_226_n PM_SKY130_FD_SC_HD__O21BAI_1%VPWR
x_PM_SKY130_FD_SC_HD__O21BAI_1%Y N_Y_M1002_s N_Y_M1000_d N_Y_c_266_n N_Y_c_269_n
+ N_Y_c_279_n N_Y_c_268_n Y PM_SKY130_FD_SC_HD__O21BAI_1%Y
x_PM_SKY130_FD_SC_HD__O21BAI_1%VGND N_VGND_M1007_s N_VGND_M1006_d N_VGND_c_314_n
+ N_VGND_c_315_n N_VGND_c_316_n VGND N_VGND_c_317_n N_VGND_c_318_n
+ N_VGND_c_319_n N_VGND_c_320_n PM_SKY130_FD_SC_HD__O21BAI_1%VGND
x_PM_SKY130_FD_SC_HD__O21BAI_1%A_297_47# N_A_297_47#_M1002_d N_A_297_47#_M1004_d
+ N_A_297_47#_c_368_n N_A_297_47#_c_352_n N_A_297_47#_c_353_n
+ N_A_297_47#_c_354_n N_A_297_47#_c_362_n PM_SKY130_FD_SC_HD__O21BAI_1%A_297_47#
cc_1 VNB N_B1_N_c_55_n 0.0146653f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_2 VNB N_B1_N_c_56_n 0.0277812f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_3 VNB N_B1_N_c_57_n 0.0409554f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=0.995
cc_4 VNB N_A_105_352#_c_97_n 0.020544f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.61
cc_5 VNB N_A_105_352#_c_98_n 0.0381959f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.17
cc_6 VNB N_A_105_352#_c_99_n 0.0104469f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_7 VNB N_A_105_352#_c_100_n 0.00580428f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.325
cc_8 VNB N_A_105_352#_c_101_n 9.91781e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_105_352#_c_102_n 0.00296816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_105_352#_c_103_n 0.00246355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_164_n 0.0195954f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.17
cc_12 VNB N_A2_c_165_n 0.00806639f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.345
cc_13 VNB N_A2_c_166_n 0.0165907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB A1 0.0130114f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.685
cc_15 VNB N_A1_c_202_n 0.031218f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.17
cc_16 VNB N_A1_c_203_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_226_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_266_n 0.00101686f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.17
cc_19 VNB N_VGND_c_314_n 0.0102019f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.61
cc_20 VNB N_VGND_c_315_n 0.0323671f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=1.97
cc_21 VNB N_VGND_c_316_n 0.00465632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_317_n 0.044593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_318_n 0.0174529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_319_n 0.174774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_320_n 0.00324149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_297_47#_c_352_n 0.0162553f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.17
cc_27 VNB N_A_297_47#_c_353_n 0.0016561f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.345
cc_28 VNB N_A_297_47#_c_354_n 0.0182532f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_29 VPB N_B1_N_c_58_n 0.0124051f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.535
cc_30 VPB N_B1_N_c_59_n 0.0236736f $X=-0.19 $Y=1.305 $X2=0.785 $Y2=1.61
cc_31 VPB N_B1_N_c_60_n 0.012679f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.61
cc_32 VPB N_B1_N_c_61_n 0.0394899f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.685
cc_33 VPB N_B1_N_c_55_n 0.00538841f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_34 VPB N_B1_N_c_56_n 0.00490307f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_35 VPB B1_N 0.0608071f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_36 VPB N_A_105_352#_M1000_g 0.0214777f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.345
cc_37 VPB N_A_105_352#_c_98_n 0.0147051f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.17
cc_38 VPB N_A_105_352#_c_99_n 6.77422e-19 $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_39 VPB N_A_105_352#_c_107_n 0.004229f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_40 VPB N_A_105_352#_c_108_n 0.00265927f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.53
cc_41 VPB N_A_105_352#_c_101_n 0.00297611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A2_M1001_g 0.0191712f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.675
cc_43 VPB N_A2_c_164_n 0.00534709f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.17
cc_44 VPB N_A1_M1003_g 0.0249935f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.675
cc_45 VPB N_A1_c_202_n 0.00709581f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.17
cc_46 VPB N_VPWR_c_227_n 0.00872967f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.97
cc_47 VPB N_VPWR_c_228_n 0.0115474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_229_n 0.0395329f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_49 VPB N_VPWR_c_230_n 0.0290164f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=0.995
cc_50 VPB N_VPWR_c_231_n 0.0264806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_232_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_226_n 0.0567651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_Y_c_266_n 0.0014004f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.17
cc_54 VPB N_Y_c_268_n 0.00406896f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_B1_N_c_59_n N_A_105_352#_M1000_g 0.0259763f $X=0.785 $Y=1.61 $X2=0 $Y2=0
cc_56 N_B1_N_c_59_n N_A_105_352#_c_98_n 0.00912069f $X=0.785 $Y=1.61 $X2=0 $Y2=0
cc_57 N_B1_N_c_55_n N_A_105_352#_c_98_n 3.27378e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_58 N_B1_N_c_56_n N_A_105_352#_c_98_n 0.0203188f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_59 N_B1_N_c_60_n N_A_105_352#_c_107_n 0.003689f $X=0.585 $Y=1.61 $X2=0 $Y2=0
cc_60 N_B1_N_c_61_n N_A_105_352#_c_107_n 0.00914228f $X=0.86 $Y=1.685 $X2=0
+ $Y2=0
cc_61 B1_N N_A_105_352#_c_107_n 0.0402303f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_62 N_B1_N_c_55_n N_A_105_352#_c_100_n 0.0262483f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_63 N_B1_N_c_56_n N_A_105_352#_c_100_n 0.00336656f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B1_N_c_59_n N_A_105_352#_c_108_n 0.0149797f $X=0.785 $Y=1.61 $X2=0 $Y2=0
cc_65 N_B1_N_c_60_n N_A_105_352#_c_108_n 0.00506859f $X=0.585 $Y=1.61 $X2=0
+ $Y2=0
cc_66 N_B1_N_c_61_n N_A_105_352#_c_108_n 0.00680822f $X=0.86 $Y=1.685 $X2=0
+ $Y2=0
cc_67 N_B1_N_c_55_n N_A_105_352#_c_108_n 6.56352e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_68 B1_N N_A_105_352#_c_108_n 0.0136248f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_69 N_B1_N_c_58_n N_A_105_352#_c_101_n 0.00336656f $X=0.51 $Y=1.535 $X2=0
+ $Y2=0
cc_70 N_B1_N_c_59_n N_A_105_352#_c_101_n 0.00231499f $X=0.785 $Y=1.61 $X2=0
+ $Y2=0
cc_71 B1_N N_A_105_352#_c_101_n 0.00907541f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_72 N_B1_N_c_57_n N_A_105_352#_c_103_n 0.00523341f $X=0.45 $Y=0.995 $X2=0
+ $Y2=0
cc_73 N_B1_N_c_61_n N_VPWR_c_227_n 0.0101118f $X=0.86 $Y=1.685 $X2=0 $Y2=0
cc_74 B1_N N_VPWR_c_227_n 0.00779366f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_75 N_B1_N_c_61_n N_VPWR_c_230_n 0.00568582f $X=0.86 $Y=1.685 $X2=0 $Y2=0
cc_76 B1_N N_VPWR_c_230_n 0.0170586f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_77 N_B1_N_c_61_n N_VPWR_c_226_n 0.0118663f $X=0.86 $Y=1.685 $X2=0 $Y2=0
cc_78 B1_N N_VPWR_c_226_n 0.010222f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_79 N_B1_N_c_57_n N_Y_c_269_n 0.00566071f $X=0.45 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B1_N_c_59_n N_Y_c_268_n 3.04461e-19 $X=0.785 $Y=1.61 $X2=0 $Y2=0
cc_81 N_B1_N_c_61_n Y 6.48481e-19 $X=0.86 $Y=1.685 $X2=0 $Y2=0
cc_82 N_B1_N_c_55_n N_VGND_c_315_n 0.0227306f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B1_N_c_56_n N_VGND_c_315_n 9.6102e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B1_N_c_57_n N_VGND_c_315_n 0.0142191f $X=0.45 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B1_N_c_57_n N_VGND_c_317_n 0.00585385f $X=0.45 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B1_N_c_57_n N_VGND_c_319_n 0.013019f $X=0.45 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_105_352#_M1000_g N_A2_M1001_g 0.0125647f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_105_352#_c_99_n N_A2_c_164_n 0.0200991f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_105_352#_c_99_n N_A2_c_165_n 0.00183882f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_105_352#_c_97_n N_A2_c_166_n 0.0102028f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_105_352#_c_108_n N_VPWR_M1005_d 0.00190565f $X=0.867 $Y=1.535
+ $X2=-0.19 $Y2=-0.24
cc_92 N_A_105_352#_c_101_n N_VPWR_M1005_d 4.49946e-19 $X=0.93 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_105_352#_M1000_g N_VPWR_c_227_n 0.00678258f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_94 N_A_105_352#_c_98_n N_VPWR_c_227_n 0.00511275f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_95 N_A_105_352#_c_107_n N_VPWR_c_227_n 0.0134303f $X=0.65 $Y=1.96 $X2=0 $Y2=0
cc_96 N_A_105_352#_c_108_n N_VPWR_c_227_n 0.00265269f $X=0.867 $Y=1.535 $X2=0
+ $Y2=0
cc_97 N_A_105_352#_c_107_n N_VPWR_c_230_n 0.00718354f $X=0.65 $Y=1.96 $X2=0
+ $Y2=0
cc_98 N_A_105_352#_M1000_g N_VPWR_c_231_n 0.00564131f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_99 N_A_105_352#_M1000_g N_VPWR_c_226_n 0.010531f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_105_352#_c_107_n N_VPWR_c_226_n 0.00880775f $X=0.65 $Y=1.96 $X2=0
+ $Y2=0
cc_101 N_A_105_352#_c_97_n N_Y_c_266_n 0.00529755f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_105_352#_M1000_g N_Y_c_266_n 0.00450555f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_105_352#_c_98_n N_Y_c_266_n 0.0149192f $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_105_352#_c_99_n N_Y_c_266_n 0.0039934f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_105_352#_c_100_n N_Y_c_266_n 0.0335338f $X=0.867 $Y=1.142 $X2=0 $Y2=0
cc_106 N_A_105_352#_c_103_n N_Y_c_266_n 0.00856928f $X=0.867 $Y=0.995 $X2=0
+ $Y2=0
cc_107 N_A_105_352#_c_102_n N_Y_c_269_n 0.00697618f $X=0.68 $Y=0.66 $X2=0 $Y2=0
cc_108 N_A_105_352#_c_97_n N_Y_c_279_n 0.00396136f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_105_352#_c_98_n N_Y_c_279_n 0.00297982f $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_105_352#_c_102_n N_Y_c_279_n 0.0110893f $X=0.68 $Y=0.66 $X2=0 $Y2=0
cc_111 N_A_105_352#_M1000_g N_Y_c_268_n 0.0168639f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_105_352#_c_98_n N_Y_c_268_n 8.40343e-19 $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_105_352#_c_108_n N_Y_c_268_n 0.00768253f $X=0.867 $Y=1.535 $X2=0
+ $Y2=0
cc_114 N_A_105_352#_c_101_n N_Y_c_268_n 0.0067118f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_105_352#_M1000_g Y 0.0104038f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_105_352#_c_107_n Y 0.00399131f $X=0.65 $Y=1.96 $X2=0 $Y2=0
cc_117 N_A_105_352#_c_108_n Y 0.00296084f $X=0.867 $Y=1.535 $X2=0 $Y2=0
cc_118 N_A_105_352#_c_97_n N_VGND_c_317_n 0.00565249f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_119 N_A_105_352#_c_102_n N_VGND_c_317_n 0.00701298f $X=0.68 $Y=0.66 $X2=0
+ $Y2=0
cc_120 N_A_105_352#_c_97_n N_VGND_c_319_n 0.0116132f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_121 N_A_105_352#_c_102_n N_VGND_c_319_n 0.00974798f $X=0.68 $Y=0.66 $X2=0
+ $Y2=0
cc_122 N_A_105_352#_c_97_n N_A_297_47#_c_353_n 8.50418e-19 $X=1.41 $Y=0.995
+ $X2=0 $Y2=0
cc_123 N_A2_M1001_g N_A1_M1003_g 0.0611398f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A2_c_164_n A1 2.3931e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A2_c_165_n A1 0.0176496f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A2_c_164_n N_A1_c_202_n 0.0224569f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A2_c_165_n N_A1_c_202_n 7.34602e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A2_c_166_n N_A1_c_203_n 0.0259398f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_M1001_g N_VPWR_c_229_n 0.00420581f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A2_M1001_g N_VPWR_c_231_n 0.00579312f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A2_M1001_g N_VPWR_c_226_n 0.0106978f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A2_M1001_g N_Y_c_266_n 6.22251e-19 $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A2_c_164_n N_Y_c_266_n 7.96886e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A2_c_165_n N_Y_c_266_n 0.0163414f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A2_c_166_n N_Y_c_266_n 4.30902e-19 $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A2_M1001_g N_Y_c_268_n 0.0031615f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A2_c_164_n N_Y_c_268_n 0.00176257f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A2_c_165_n N_Y_c_268_n 0.0203331f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A2_M1001_g Y 0.0126219f $X=1.865 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A2_c_166_n N_VGND_c_316_n 0.00268723f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A2_c_166_n N_VGND_c_317_n 0.0042616f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A2_c_166_n N_VGND_c_319_n 0.00592935f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A2_c_164_n N_A_297_47#_c_352_n 0.00236039f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A2_c_165_n N_A_297_47#_c_352_n 0.020259f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A2_c_166_n N_A_297_47#_c_352_n 0.0100958f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A2_c_164_n N_A_297_47#_c_353_n 6.3983e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A2_c_165_n N_A_297_47#_c_353_n 0.014417f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_166_n N_A_297_47#_c_354_n 5.66403e-19 $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_165_n N_A_297_47#_c_362_n 0.00115914f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_166_n N_A_297_47#_c_362_n 0.00289352f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_M1003_g N_VPWR_c_229_n 0.027322f $X=2.27 $Y=1.985 $X2=0 $Y2=0
cc_152 A1 N_VPWR_c_229_n 0.0204754f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A1_c_202_n N_VPWR_c_229_n 0.00452834f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A1_M1003_g N_VPWR_c_231_n 0.00290915f $X=2.27 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A1_M1003_g N_VPWR_c_226_n 0.00525288f $X=2.27 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A1_M1003_g N_Y_c_268_n 6.13891e-19 $X=2.27 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A1_M1003_g Y 0.00228854f $X=2.27 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A1_c_203_n N_VGND_c_316_n 0.00268723f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A1_c_203_n N_VGND_c_318_n 0.00425021f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A1_c_203_n N_VGND_c_319_n 0.00671814f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_161 A1 N_A_297_47#_c_352_n 0.0368575f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A1_c_202_n N_A_297_47#_c_352_n 0.00518233f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A1_c_203_n N_A_297_47#_c_352_n 0.00972538f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A1_c_203_n N_A_297_47#_c_354_n 0.00658829f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_165 N_VPWR_c_226_n N_Y_M1000_d 0.00243306f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_166 N_VPWR_M1005_d N_Y_c_268_n 0.00246556f $X=0.935 $Y=1.76 $X2=0 $Y2=0
cc_167 N_VPWR_c_227_n N_Y_c_268_n 0.00568599f $X=1.135 $Y=1.96 $X2=0 $Y2=0
cc_168 N_VPWR_c_229_n N_Y_c_268_n 0.00307433f $X=2.48 $Y=1.62 $X2=0 $Y2=0
cc_169 N_VPWR_c_229_n Y 0.0275777f $X=2.48 $Y=1.62 $X2=0 $Y2=0
cc_170 N_VPWR_c_231_n Y 0.0186379f $X=2.27 $Y=2.72 $X2=0 $Y2=0
cc_171 N_VPWR_c_226_n Y 0.0122121f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_172 N_VPWR_c_226_n A_388_297# 0.0109087f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_173 N_Y_c_269_n N_VGND_c_317_n 0.0115427f $X=1.235 $Y=0.645 $X2=0 $Y2=0
cc_174 N_Y_c_279_n N_VGND_c_317_n 8.03473e-19 $X=1.235 $Y=0.825 $X2=0 $Y2=0
cc_175 N_Y_M1002_s N_VGND_c_319_n 0.00370545f $X=1.075 $Y=0.235 $X2=0 $Y2=0
cc_176 N_Y_c_269_n N_VGND_c_319_n 0.00645781f $X=1.235 $Y=0.645 $X2=0 $Y2=0
cc_177 N_Y_c_279_n N_VGND_c_319_n 0.00194999f $X=1.235 $Y=0.825 $X2=0 $Y2=0
cc_178 N_Y_c_279_n N_A_297_47#_c_368_n 0.00538187f $X=1.235 $Y=0.825 $X2=0 $Y2=0
cc_179 N_Y_c_279_n N_A_297_47#_c_353_n 0.0113451f $X=1.235 $Y=0.825 $X2=0 $Y2=0
cc_180 N_VGND_c_319_n N_A_297_47#_M1002_d 0.00264678f $X=2.53 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_181 N_VGND_c_319_n N_A_297_47#_M1004_d 0.00209863f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_182 N_VGND_M1006_d N_A_297_47#_c_352_n 0.00165819f $X=1.945 $Y=0.235 $X2=0
+ $Y2=0
cc_183 N_VGND_c_316_n N_A_297_47#_c_352_n 0.0116529f $X=2.08 $Y=0.39 $X2=0 $Y2=0
cc_184 N_VGND_c_317_n N_A_297_47#_c_352_n 0.00202181f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_185 N_VGND_c_318_n N_A_297_47#_c_352_n 0.00193763f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_319_n N_A_297_47#_c_352_n 0.00857256f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_187 N_VGND_c_318_n N_A_297_47#_c_354_n 0.0191165f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_188 N_VGND_c_319_n N_A_297_47#_c_354_n 0.0123122f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_c_317_n N_A_297_47#_c_362_n 0.0189202f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_190 N_VGND_c_319_n N_A_297_47#_c_362_n 0.0122874f $X=2.53 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a2bb2o_4.spice.SKY130_FD_SC_HD__A2BB2O_4.pxi
* Created: Thu Aug 27 14:03:24 2020
* 
x_PM_SKY130_FD_SC_HD__A2BB2O_4%B1 N_B1_M1016_g N_B1_M1019_g N_B1_c_131_n
+ N_B1_M1027_g N_B1_M1025_g N_B1_c_140_n N_B1_c_132_n N_B1_c_133_n N_B1_c_134_n
+ B1 N_B1_c_135_n N_B1_c_136_n N_B1_c_137_n PM_SKY130_FD_SC_HD__A2BB2O_4%B1
x_PM_SKY130_FD_SC_HD__A2BB2O_4%B2 N_B2_c_214_n N_B2_M1013_g N_B2_M1001_g
+ N_B2_c_215_n N_B2_M1018_g N_B2_M1003_g B2 N_B2_c_217_n
+ PM_SKY130_FD_SC_HD__A2BB2O_4%B2
x_PM_SKY130_FD_SC_HD__A2BB2O_4%A_415_21# N_A_415_21#_M1008_d N_A_415_21#_M1014_s
+ N_A_415_21#_M1012_s N_A_415_21#_c_259_n N_A_415_21#_M1020_g
+ N_A_415_21#_M1004_g N_A_415_21#_c_260_n N_A_415_21#_M1024_g
+ N_A_415_21#_M1022_g N_A_415_21#_c_261_n N_A_415_21#_c_262_n
+ N_A_415_21#_c_263_n N_A_415_21#_c_264_n N_A_415_21#_c_265_n
+ N_A_415_21#_c_266_n N_A_415_21#_c_280_p N_A_415_21#_c_303_p
+ N_A_415_21#_c_267_n N_A_415_21#_c_282_p N_A_415_21#_c_268_n
+ N_A_415_21#_c_269_n N_A_415_21#_c_287_p PM_SKY130_FD_SC_HD__A2BB2O_4%A_415_21#
x_PM_SKY130_FD_SC_HD__A2BB2O_4%A1_N N_A1_N_M1008_g N_A1_N_M1009_g N_A1_N_c_398_n
+ N_A1_N_M1021_g N_A1_N_M1023_g N_A1_N_c_406_n A1_N A1_N N_A1_N_c_401_n
+ N_A1_N_c_402_n N_A1_N_c_403_n PM_SKY130_FD_SC_HD__A2BB2O_4%A1_N
x_PM_SKY130_FD_SC_HD__A2BB2O_4%A2_N N_A2_N_c_488_n N_A2_N_M1007_g N_A2_N_M1012_g
+ N_A2_N_c_489_n N_A2_N_M1014_g N_A2_N_M1015_g A2_N N_A2_N_c_490_n
+ N_A2_N_c_491_n PM_SKY130_FD_SC_HD__A2BB2O_4%A2_N
x_PM_SKY130_FD_SC_HD__A2BB2O_4%A_193_47# N_A_193_47#_M1013_d N_A_193_47#_M1020_s
+ N_A_193_47#_M1004_s N_A_193_47#_c_536_n N_A_193_47#_M1006_g
+ N_A_193_47#_M1000_g N_A_193_47#_c_537_n N_A_193_47#_M1010_g
+ N_A_193_47#_M1002_g N_A_193_47#_c_538_n N_A_193_47#_M1011_g
+ N_A_193_47#_M1005_g N_A_193_47#_c_539_n N_A_193_47#_M1017_g
+ N_A_193_47#_M1026_g N_A_193_47#_c_540_n N_A_193_47#_c_560_n
+ N_A_193_47#_c_541_n N_A_193_47#_c_607_n N_A_193_47#_c_653_p
+ N_A_193_47#_c_542_n N_A_193_47#_c_543_n N_A_193_47#_c_550_n
+ N_A_193_47#_c_551_n N_A_193_47#_c_552_n N_A_193_47#_c_553_n
+ N_A_193_47#_c_544_n N_A_193_47#_c_555_n PM_SKY130_FD_SC_HD__A2BB2O_4%A_193_47#
x_PM_SKY130_FD_SC_HD__A2BB2O_4%A_27_297# N_A_27_297#_M1019_s N_A_27_297#_M1001_s
+ N_A_27_297#_M1025_s N_A_27_297#_M1022_d N_A_27_297#_c_753_p
+ N_A_27_297#_c_718_n N_A_27_297#_c_714_n N_A_27_297#_c_754_p
+ N_A_27_297#_c_723_n N_A_27_297#_c_715_n N_A_27_297#_c_734_n
+ N_A_27_297#_c_751_p N_A_27_297#_c_730_n N_A_27_297#_c_743_n
+ PM_SKY130_FD_SC_HD__A2BB2O_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A2BB2O_4%VPWR N_VPWR_M1019_d N_VPWR_M1003_d N_VPWR_M1009_d
+ N_VPWR_M1023_d N_VPWR_M1002_s N_VPWR_M1026_s N_VPWR_c_767_n N_VPWR_c_768_n
+ N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n
+ N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n N_VPWR_c_777_n VPWR
+ N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_766_n
+ N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n
+ PM_SKY130_FD_SC_HD__A2BB2O_4%VPWR
x_PM_SKY130_FD_SC_HD__A2BB2O_4%A_717_297# N_A_717_297#_M1009_s
+ N_A_717_297#_M1015_d N_A_717_297#_c_885_n N_A_717_297#_c_891_n
+ N_A_717_297#_c_888_n PM_SKY130_FD_SC_HD__A2BB2O_4%A_717_297#
x_PM_SKY130_FD_SC_HD__A2BB2O_4%X N_X_M1006_d N_X_M1011_d N_X_M1000_d N_X_M1005_d
+ N_X_c_913_n N_X_c_954_n N_X_c_916_n N_X_c_920_n N_X_c_901_n N_X_c_902_n
+ N_X_c_934_n N_X_c_959_n N_X_c_903_n N_X_c_904_n N_X_c_906_n X X N_X_c_909_n
+ PM_SKY130_FD_SC_HD__A2BB2O_4%X
x_PM_SKY130_FD_SC_HD__A2BB2O_4%VGND N_VGND_M1016_d N_VGND_M1027_d N_VGND_M1024_d
+ N_VGND_M1007_d N_VGND_M1021_s N_VGND_M1010_s N_VGND_M1017_s N_VGND_c_982_n
+ N_VGND_c_983_n N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n
+ N_VGND_c_988_n N_VGND_c_989_n N_VGND_c_990_n N_VGND_c_991_n N_VGND_c_992_n
+ N_VGND_c_993_n N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n
+ VGND N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n
+ N_VGND_c_1002_n PM_SKY130_FD_SC_HD__A2BB2O_4%VGND
x_PM_SKY130_FD_SC_HD__A2BB2O_4%A_109_47# N_A_109_47#_M1016_s N_A_109_47#_M1018_s
+ N_A_109_47#_c_1103_n N_A_109_47#_c_1102_n N_A_109_47#_c_1107_n
+ PM_SKY130_FD_SC_HD__A2BB2O_4%A_109_47#
cc_1 VNB N_B1_c_131_n 0.0162054f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_2 VNB N_B1_c_132_n 6.86943e-19 $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.445
cc_3 VNB N_B1_c_133_n 0.00383856f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_4 VNB N_B1_c_134_n 0.0194119f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_5 VNB N_B1_c_135_n 0.0281636f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_6 VNB N_B1_c_136_n 0.0155878f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_7 VNB N_B1_c_137_n 0.021834f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_8 VNB N_B2_c_214_n 0.0161301f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_9 VNB N_B2_c_215_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_10 VNB B2 0.00164887f $X=-0.19 $Y=-0.24 $X2=1.515 $Y2=1.53
cc_11 VNB N_B2_c_217_n 0.0307903f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_12 VNB N_A_415_21#_c_259_n 0.0159859f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_13 VNB N_A_415_21#_c_260_n 0.0193955f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.245
cc_14 VNB N_A_415_21#_c_261_n 2.36777e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_415_21#_c_262_n 0.0523147f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_16 VNB N_A_415_21#_c_263_n 0.00331986f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_17 VNB N_A_415_21#_c_264_n 8.80236e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_18 VNB N_A_415_21#_c_265_n 0.0028719f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_19 VNB N_A_415_21#_c_266_n 2.65295e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_415_21#_c_267_n 0.00512232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_415_21#_c_268_n 0.00108817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_415_21#_c_269_n 0.00307597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A1_N_c_398_n 0.0163564f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_24 VNB A1_N 0.00309127f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.445
cc_25 VNB A1_N 0.00375531f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.16
cc_26 VNB N_A1_N_c_401_n 0.0243367f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_27 VNB N_A1_N_c_402_n 0.0196134f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_28 VNB N_A1_N_c_403_n 0.0204281f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_29 VNB N_A2_N_c_488_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_30 VNB N_A2_N_c_489_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_31 VNB N_A2_N_c_490_n 0.00327879f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_32 VNB N_A2_N_c_491_n 0.0286689f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_33 VNB N_A_193_47#_c_536_n 0.0161454f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_34 VNB N_A_193_47#_c_537_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.6 $Y2=1.245
cc_35 VNB N_A_193_47#_c_538_n 0.0157972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_539_n 0.0191608f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.325
cc_37 VNB N_A_193_47#_c_540_n 0.00660331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_541_n 0.0015888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_193_47#_c_542_n 0.00219064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_543_n 9.74694e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_193_47#_c_544_n 0.0657261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_766_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_X_c_901_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_44 VNB N_X_c_902_n 0.00210954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_903_n 0.0113532f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_46 VNB N_X_c_904_n 0.00221468f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.19
cc_47 VNB X 0.0216602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_982_n 0.0110494f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_49 VNB N_VGND_c_983_n 0.0064991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_984_n 0.00410177f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_51 VNB N_VGND_c_985_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_52 VNB N_VGND_c_986_n 0.00630241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_987_n 0.0176493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_988_n 0.00359433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_989_n 0.00416791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_990_n 0.0359188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_991_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_992_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_993_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_994_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_995_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_996_n 0.017009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_997_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_998_n 0.0210665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_999_n 0.369023f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1000_n 0.0173211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1001_n 0.0197313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1002_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_109_47#_c_1102_n 0.00331844f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_70 VPB N_B1_M1019_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_71 VPB N_B1_M1025_g 0.0181922f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_72 VPB N_B1_c_140_n 0.0085411f $X=-0.19 $Y=1.305 $X2=1.515 $Y2=1.53
cc_73 VPB N_B1_c_132_n 0.00130166f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.445
cc_74 VPB N_B1_c_134_n 0.00452287f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_75 VPB N_B1_c_135_n 0.00483422f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_76 VPB N_B1_c_136_n 0.0160332f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_77 VPB N_B2_M1001_g 0.018362f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_78 VPB N_B2_M1003_g 0.018351f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_79 VPB N_B2_c_217_n 0.00405312f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_80 VPB N_A_415_21#_M1004_g 0.0187684f $X=-0.19 $Y=1.305 $X2=1.515 $Y2=1.53
cc_81 VPB N_A_415_21#_M1022_g 0.0226996f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_82 VPB N_A_415_21#_c_262_n 0.0160069f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_83 VPB N_A_415_21#_c_264_n 0.0178087f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_84 VPB N_A1_N_M1009_g 0.0219574f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_85 VPB N_A1_N_M1023_g 0.0172429f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_86 VPB N_A1_N_c_406_n 0.00788908f $X=-0.19 $Y=1.305 $X2=1.515 $Y2=1.53
cc_87 VPB A1_N 0.00279337f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.445
cc_88 VPB A1_N 0.00228101f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.16
cc_89 VPB N_A1_N_c_401_n 0.00638236f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_90 VPB N_A1_N_c_403_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_91 VPB N_A2_N_M1012_g 0.0183411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_92 VPB N_A2_N_M1015_g 0.0183385f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_93 VPB N_A2_N_c_491_n 0.00400438f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_94 VPB N_A_193_47#_M1000_g 0.017975f $X=-0.19 $Y=1.305 $X2=1.515 $Y2=1.53
cc_95 VPB N_A_193_47#_M1002_g 0.0184401f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_96 VPB N_A_193_47#_M1005_g 0.0184597f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_97 VPB N_A_193_47#_M1026_g 0.022036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_193_47#_c_541_n 0.00154937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_193_47#_c_550_n 0.00938894f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_193_47#_c_551_n 0.00117154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_193_47#_c_552_n 0.0010614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_193_47#_c_553_n 0.00153686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_193_47#_c_544_n 0.0111799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_193_47#_c_555_n 9.22248e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_297#_c_714_n 0.00692367f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.445
cc_106 VPB N_A_27_297#_c_715_n 0.00353338f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.325
cc_107 VPB N_VPWR_c_767_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_108 VPB N_VPWR_c_768_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_109 VPB N_VPWR_c_769_n 0.00517963f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_110 VPB N_VPWR_c_770_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_111 VPB N_VPWR_c_771_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.19
cc_112 VPB N_VPWR_c_772_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_773_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_774_n 0.0379753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_775_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_776_n 0.0343319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_777_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_778_n 0.0174714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_779_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_780_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_781_n 0.0204409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_766_n 0.0753335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_783_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_784_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_785_n 0.00478125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_786_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_X_c_906_n 0.00297629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB X 0.00597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB X 0.00130197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_X_c_909_n 0.0163194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 N_B1_c_137_n N_B2_c_214_n 0.0241442f $X=0.41 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_132 N_B1_M1019_g N_B2_M1001_g 0.0241442f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_133 N_B1_c_140_n N_B2_M1001_g 0.00995634f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_134 N_B1_c_131_n N_B2_c_215_n 0.0269014f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B1_M1025_g N_B2_M1003_g 0.0424827f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B1_c_140_n N_B2_M1003_g 0.0107507f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_137 N_B1_c_140_n B2 0.0381541f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_138 N_B1_c_132_n B2 0.00227533f $X=1.6 $Y=1.445 $X2=0 $Y2=0
cc_139 N_B1_c_133_n B2 0.014073f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B1_c_135_n B2 7.59344e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B1_c_136_n B2 0.0143152f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B1_c_140_n N_B2_c_217_n 0.00214031f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_143 N_B1_c_132_n N_B2_c_217_n 0.00386559f $X=1.6 $Y=1.445 $X2=0 $Y2=0
cc_144 N_B1_c_133_n N_B2_c_217_n 0.0011131f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B1_c_134_n N_B2_c_217_n 0.0222997f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B1_c_135_n N_B2_c_217_n 0.0241442f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B1_c_136_n N_B2_c_217_n 0.00483648f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B1_c_131_n N_A_415_21#_c_259_n 0.0261706f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_149 N_B1_M1025_g N_A_415_21#_M1004_g 0.0133907f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B1_c_132_n N_A_415_21#_c_262_n 6.19192e-19 $X=1.6 $Y=1.445 $X2=0 $Y2=0
cc_151 N_B1_c_133_n N_A_415_21#_c_262_n 0.00141851f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_152 N_B1_c_134_n N_A_415_21#_c_262_n 0.0225703f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_153 N_B1_c_131_n N_A_193_47#_c_540_n 0.0118089f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B1_c_140_n N_A_193_47#_c_540_n 0.0054287f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_155 N_B1_c_133_n N_A_193_47#_c_540_n 0.0270322f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B1_c_134_n N_A_193_47#_c_540_n 0.00295767f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B1_c_131_n N_A_193_47#_c_560_n 9.11043e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B1_c_132_n N_A_193_47#_c_541_n 0.00476267f $X=1.6 $Y=1.445 $X2=0 $Y2=0
cc_159 N_B1_c_133_n N_A_193_47#_c_541_n 0.00780783f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B1_c_134_n N_A_193_47#_c_541_n 8.02928e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B1_c_131_n N_A_193_47#_c_542_n 5.32265e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B1_c_140_n N_A_193_47#_c_555_n 3.47224e-19 $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_163 N_B1_c_132_n N_A_193_47#_c_555_n 9.35155e-19 $X=1.6 $Y=1.445 $X2=0 $Y2=0
cc_164 N_B1_c_136_n N_A_27_297#_M1019_s 0.00271779f $X=0.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_165 N_B1_c_140_n N_A_27_297#_M1001_s 0.00165831f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_166 N_B1_M1019_g N_A_27_297#_c_718_n 0.0095558f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_167 N_B1_c_140_n N_A_27_297#_c_718_n 0.021464f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_168 N_B1_c_136_n N_A_27_297#_c_718_n 0.0111744f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B1_c_135_n N_A_27_297#_c_714_n 3.79492e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_c_136_n N_A_27_297#_c_714_n 0.0179952f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B1_M1025_g N_A_27_297#_c_723_n 0.0109901f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_172 N_B1_c_140_n N_A_27_297#_c_723_n 0.0239693f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_173 N_B1_c_133_n N_A_27_297#_c_723_n 0.00330156f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B1_M1025_g N_A_27_297#_c_715_n 2.0859e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_175 N_B1_c_140_n N_A_27_297#_c_715_n 0.00787128f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_176 N_B1_c_133_n N_A_27_297#_c_715_n 0.00280327f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B1_c_134_n N_A_27_297#_c_715_n 2.26413e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B1_c_140_n N_A_27_297#_c_730_n 0.0126919f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_179 N_B1_c_140_n N_VPWR_M1019_d 0.00166235f $X=1.515 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_180 N_B1_c_140_n N_VPWR_M1003_d 0.00166017f $X=1.515 $Y=1.53 $X2=0 $Y2=0
cc_181 N_B1_M1019_g N_VPWR_c_767_n 0.00302074f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B1_M1025_g N_VPWR_c_768_n 0.00302074f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_M1025_g N_VPWR_c_774_n 0.00585385f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_M1019_g N_VPWR_c_778_n 0.00585385f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_M1019_g N_VPWR_c_766_n 0.00686624f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_M1025_g N_VPWR_c_766_n 0.00593924f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B1_c_135_n N_VGND_c_983_n 0.00176179f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B1_c_136_n N_VGND_c_983_n 0.0145468f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B1_c_137_n N_VGND_c_983_n 0.00460417f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B1_c_131_n N_VGND_c_984_n 0.00268723f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B1_c_131_n N_VGND_c_990_n 0.0042294f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B1_c_137_n N_VGND_c_990_n 0.00539841f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B1_c_131_n N_VGND_c_999_n 0.00579958f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B1_c_137_n N_VGND_c_999_n 0.010446f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B1_c_137_n N_A_109_47#_c_1103_n 0.00266812f $X=0.41 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_B1_c_140_n N_A_109_47#_c_1102_n 0.00711902f $X=1.515 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_B1_c_136_n N_A_109_47#_c_1102_n 0.00506593f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B1_c_137_n N_A_109_47#_c_1102_n 0.00561701f $X=0.41 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_B1_c_131_n N_A_109_47#_c_1107_n 0.00303739f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_B2_c_215_n N_A_193_47#_c_540_n 0.00871206f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_201 B2 N_A_193_47#_c_540_n 0.00514788f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_202 N_B2_c_214_n N_A_193_47#_c_542_n 0.00371029f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B2_c_215_n N_A_193_47#_c_542_n 0.00389925f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_204 B2 N_A_193_47#_c_542_n 0.0248173f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_205 N_B2_c_217_n N_A_193_47#_c_542_n 0.00224391f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B2_M1001_g N_A_27_297#_c_718_n 0.00956194f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B2_M1003_g N_A_27_297#_c_723_n 0.00956194f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B2_M1001_g N_VPWR_c_767_n 0.00157837f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B2_M1003_g N_VPWR_c_768_n 0.00157837f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B2_M1001_g N_VPWR_c_779_n 0.00585385f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B2_M1003_g N_VPWR_c_779_n 0.00585385f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B2_M1001_g N_VPWR_c_766_n 0.00591203f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B2_M1003_g N_VPWR_c_766_n 0.00591203f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B2_c_214_n N_VGND_c_990_n 0.00357877f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B2_c_215_n N_VGND_c_990_n 0.00357877f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B2_c_214_n N_VGND_c_999_n 0.00525237f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B2_c_215_n N_VGND_c_999_n 0.00524329f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B2_c_214_n N_A_109_47#_c_1107_n 0.0105795f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B2_c_215_n N_A_109_47#_c_1107_n 0.00931565f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_220 B2 N_A_109_47#_c_1107_n 0.00315795f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_221 N_A_415_21#_c_264_n N_A1_N_M1009_g 0.0111914f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_222 N_A_415_21#_c_280_p N_A1_N_M1009_g 0.014345f $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_223 N_A_415_21#_c_267_n N_A1_N_c_398_n 0.00258856f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_224 N_A_415_21#_c_282_p N_A1_N_c_398_n 0.00513121f $X=4.56 $Y=0.39 $X2=0
+ $Y2=0
cc_225 N_A_415_21#_M1012_s N_A1_N_c_406_n 0.00165831f $X=4.005 $Y=1.485 $X2=0
+ $Y2=0
cc_226 N_A_415_21#_c_280_p N_A1_N_c_406_n 0.0193381f $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_227 N_A_415_21#_c_267_n N_A1_N_c_406_n 0.00495999f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_228 N_A_415_21#_c_269_n N_A1_N_c_406_n 0.00495999f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_229 N_A_415_21#_c_287_p N_A1_N_c_406_n 0.0108571f $X=4.14 $Y=1.875 $X2=0
+ $Y2=0
cc_230 N_A_415_21#_c_264_n A1_N 0.0216817f $X=3.05 $Y=1.495 $X2=0 $Y2=0
cc_231 N_A_415_21#_c_265_n A1_N 0.0172107f $X=3.555 $Y=0.815 $X2=0 $Y2=0
cc_232 N_A_415_21#_c_280_p A1_N 0.00974891f $X=4.015 $Y=1.875 $X2=0 $Y2=0
cc_233 N_A_415_21#_c_268_n A1_N 0.0141173f $X=3.05 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_415_21#_c_269_n A1_N 0.00750214f $X=3.72 $Y=0.815 $X2=0 $Y2=0
cc_235 N_A_415_21#_c_267_n A1_N 0.0100882f $X=4.395 $Y=0.815 $X2=0 $Y2=0
cc_236 N_A_415_21#_c_262_n N_A1_N_c_401_n 0.010016f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_415_21#_c_263_n N_A1_N_c_401_n 0.00181398f $X=3.05 $Y=1.075 $X2=0
+ $Y2=0
cc_238 N_A_415_21#_c_264_n N_A1_N_c_401_n 2.75171e-19 $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_239 N_A_415_21#_c_265_n N_A1_N_c_401_n 0.00296008f $X=3.555 $Y=0.815 $X2=0
+ $Y2=0
cc_240 N_A_415_21#_c_280_p N_A1_N_c_401_n 6.45198e-19 $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_241 N_A_415_21#_c_268_n N_A1_N_c_401_n 6.90629e-19 $X=3.05 $Y=1.16 $X2=0
+ $Y2=0
cc_242 N_A_415_21#_c_269_n N_A1_N_c_401_n 0.00153445f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_243 N_A_415_21#_c_263_n N_A1_N_c_402_n 0.00271538f $X=3.05 $Y=1.075 $X2=0
+ $Y2=0
cc_244 N_A_415_21#_c_265_n N_A1_N_c_402_n 0.0106092f $X=3.555 $Y=0.815 $X2=0
+ $Y2=0
cc_245 N_A_415_21#_c_303_p N_A1_N_c_402_n 0.0109565f $X=3.72 $Y=0.39 $X2=0 $Y2=0
cc_246 N_A_415_21#_c_269_n N_A1_N_c_402_n 0.00112502f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_247 N_A_415_21#_c_267_n N_A1_N_c_403_n 0.00153445f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_248 N_A_415_21#_c_303_p N_A2_N_c_488_n 0.00630972f $X=3.72 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_249 N_A_415_21#_c_267_n N_A2_N_c_488_n 0.00869748f $X=4.395 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_250 N_A_415_21#_c_282_p N_A2_N_c_488_n 5.22228e-19 $X=4.56 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_251 N_A_415_21#_c_269_n N_A2_N_c_488_n 0.00112628f $X=3.72 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_252 N_A_415_21#_c_280_p N_A2_N_M1012_g 0.00938242f $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_253 N_A_415_21#_c_303_p N_A2_N_c_489_n 5.22228e-19 $X=3.72 $Y=0.39 $X2=0
+ $Y2=0
cc_254 N_A_415_21#_c_267_n N_A2_N_c_489_n 0.00982376f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_255 N_A_415_21#_c_282_p N_A2_N_c_489_n 0.00630972f $X=4.56 $Y=0.39 $X2=0
+ $Y2=0
cc_256 N_A_415_21#_c_267_n N_A2_N_c_490_n 0.0381033f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_257 N_A_415_21#_c_269_n N_A2_N_c_490_n 0.00552894f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_258 N_A_415_21#_c_267_n N_A2_N_c_491_n 0.00222133f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_259 N_A_415_21#_c_259_n N_A_193_47#_c_540_n 0.0120921f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_415_21#_c_259_n N_A_193_47#_c_560_n 0.00667227f $X=2.15 $Y=0.995
+ $X2=0 $Y2=0
cc_261 N_A_415_21#_c_260_n N_A_193_47#_c_560_n 0.0111581f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_415_21#_c_266_n N_A_193_47#_c_560_n 3.85524e-19 $X=3.145 $Y=0.815
+ $X2=0 $Y2=0
cc_263 N_A_415_21#_c_259_n N_A_193_47#_c_541_n 0.00232906f $X=2.15 $Y=0.995
+ $X2=0 $Y2=0
cc_264 N_A_415_21#_M1004_g N_A_193_47#_c_541_n 0.0011752f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_265 N_A_415_21#_c_260_n N_A_193_47#_c_541_n 0.00104304f $X=2.57 $Y=0.995
+ $X2=0 $Y2=0
cc_266 N_A_415_21#_M1022_g N_A_193_47#_c_541_n 0.00104304f $X=2.57 $Y=1.985
+ $X2=0 $Y2=0
cc_267 N_A_415_21#_c_261_n N_A_193_47#_c_541_n 0.0127231f $X=2.955 $Y=1.16 $X2=0
+ $Y2=0
cc_268 N_A_415_21#_c_262_n N_A_193_47#_c_541_n 0.0214396f $X=2.78 $Y=1.16 $X2=0
+ $Y2=0
cc_269 N_A_415_21#_c_263_n N_A_193_47#_c_541_n 0.00572741f $X=3.05 $Y=1.075
+ $X2=0 $Y2=0
cc_270 N_A_415_21#_c_264_n N_A_193_47#_c_541_n 0.00574524f $X=3.05 $Y=1.495
+ $X2=0 $Y2=0
cc_271 N_A_415_21#_c_259_n N_A_193_47#_c_543_n 0.00218377f $X=2.15 $Y=0.995
+ $X2=0 $Y2=0
cc_272 N_A_415_21#_c_260_n N_A_193_47#_c_543_n 0.00389811f $X=2.57 $Y=0.995
+ $X2=0 $Y2=0
cc_273 N_A_415_21#_c_266_n N_A_193_47#_c_543_n 0.0072611f $X=3.145 $Y=0.815
+ $X2=0 $Y2=0
cc_274 N_A_415_21#_c_261_n N_A_193_47#_c_550_n 0.0109126f $X=2.955 $Y=1.16 $X2=0
+ $Y2=0
cc_275 N_A_415_21#_c_262_n N_A_193_47#_c_550_n 0.00651916f $X=2.78 $Y=1.16 $X2=0
+ $Y2=0
cc_276 N_A_415_21#_c_264_n N_A_193_47#_c_550_n 0.0324576f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_277 N_A_415_21#_c_265_n N_A_193_47#_c_550_n 0.00402343f $X=3.555 $Y=0.815
+ $X2=0 $Y2=0
cc_278 N_A_415_21#_c_280_p N_A_193_47#_c_550_n 0.00878769f $X=4.015 $Y=1.875
+ $X2=0 $Y2=0
cc_279 N_A_415_21#_c_267_n N_A_193_47#_c_550_n 0.00185612f $X=4.395 $Y=0.815
+ $X2=0 $Y2=0
cc_280 N_A_415_21#_c_269_n N_A_193_47#_c_550_n 0.0017748f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_281 N_A_415_21#_c_287_p N_A_193_47#_c_550_n 0.00196365f $X=4.14 $Y=1.875
+ $X2=0 $Y2=0
cc_282 N_A_415_21#_M1022_g N_A_193_47#_c_551_n 0.00866873f $X=2.57 $Y=1.985
+ $X2=0 $Y2=0
cc_283 N_A_415_21#_c_261_n N_A_193_47#_c_551_n 0.00257646f $X=2.955 $Y=1.16
+ $X2=0 $Y2=0
cc_284 N_A_415_21#_c_262_n N_A_193_47#_c_551_n 9.49442e-19 $X=2.78 $Y=1.16 $X2=0
+ $Y2=0
cc_285 N_A_415_21#_c_264_n N_A_193_47#_c_551_n 0.00251936f $X=3.05 $Y=1.495
+ $X2=0 $Y2=0
cc_286 N_A_415_21#_M1004_g N_A_193_47#_c_555_n 8.22863e-19 $X=2.15 $Y=1.985
+ $X2=0 $Y2=0
cc_287 N_A_415_21#_M1022_g N_A_193_47#_c_555_n 0.0177845f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_415_21#_c_261_n N_A_193_47#_c_555_n 3.03251e-19 $X=2.955 $Y=1.16
+ $X2=0 $Y2=0
cc_289 N_A_415_21#_c_264_n N_A_193_47#_c_555_n 0.0190269f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_290 N_A_415_21#_M1004_g N_A_27_297#_c_715_n 2.27076e-19 $X=2.15 $Y=1.985
+ $X2=0 $Y2=0
cc_291 N_A_415_21#_M1004_g N_A_27_297#_c_734_n 0.0121306f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_292 N_A_415_21#_M1022_g N_A_27_297#_c_734_n 0.00905298f $X=2.57 $Y=1.985
+ $X2=0 $Y2=0
cc_293 N_A_415_21#_c_264_n N_VPWR_M1009_d 0.00783975f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_294 N_A_415_21#_c_280_p N_VPWR_M1009_d 0.00165272f $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_295 N_A_415_21#_M1022_g N_VPWR_c_769_n 0.00214938f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_415_21#_c_264_n N_VPWR_c_769_n 0.0105983f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_297 N_A_415_21#_c_280_p N_VPWR_c_769_n 0.00554231f $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_298 N_A_415_21#_M1004_g N_VPWR_c_774_n 0.00357877f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A_415_21#_M1022_g N_VPWR_c_774_n 0.00357877f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_A_415_21#_c_264_n N_VPWR_c_774_n 6.22982e-19 $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_301 N_A_415_21#_c_280_p N_VPWR_c_776_n 0.00204269f $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_302 N_A_415_21#_M1012_s N_VPWR_c_766_n 0.0021603f $X=4.005 $Y=1.485 $X2=0
+ $Y2=0
cc_303 N_A_415_21#_M1004_g N_VPWR_c_766_n 0.00525237f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_A_415_21#_M1022_g N_VPWR_c_766_n 0.00655123f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_A_415_21#_c_264_n N_VPWR_c_766_n 0.0016194f $X=3.05 $Y=1.495 $X2=0
+ $Y2=0
cc_306 N_A_415_21#_c_280_p N_VPWR_c_766_n 0.00486744f $X=4.015 $Y=1.875 $X2=0
+ $Y2=0
cc_307 N_A_415_21#_c_280_p N_A_717_297#_M1009_s 0.0031158f $X=4.015 $Y=1.875
+ $X2=-0.19 $Y2=-0.24
cc_308 N_A_415_21#_M1012_s N_A_717_297#_c_885_n 0.00312348f $X=4.005 $Y=1.485
+ $X2=0 $Y2=0
cc_309 N_A_415_21#_c_280_p N_A_717_297#_c_885_n 0.00522481f $X=4.015 $Y=1.875
+ $X2=0 $Y2=0
cc_310 N_A_415_21#_c_287_p N_A_717_297#_c_885_n 0.0112811f $X=4.14 $Y=1.875
+ $X2=0 $Y2=0
cc_311 N_A_415_21#_c_280_p N_A_717_297#_c_888_n 0.0112635f $X=4.015 $Y=1.875
+ $X2=0 $Y2=0
cc_312 N_A_415_21#_c_267_n N_X_c_902_n 3.42999e-19 $X=4.395 $Y=0.815 $X2=0 $Y2=0
cc_313 N_A_415_21#_c_265_n N_VGND_M1024_d 0.00337553f $X=3.555 $Y=0.815 $X2=0
+ $Y2=0
cc_314 N_A_415_21#_c_266_n N_VGND_M1024_d 0.00592929f $X=3.145 $Y=0.815 $X2=0
+ $Y2=0
cc_315 N_A_415_21#_c_267_n N_VGND_M1007_d 0.00162089f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_316 N_A_415_21#_c_259_n N_VGND_c_984_n 0.00146339f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_415_21#_c_267_n N_VGND_c_985_n 0.0122559f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_318 N_A_415_21#_c_267_n N_VGND_c_986_n 0.00750114f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_319 N_A_415_21#_c_265_n N_VGND_c_992_n 0.00198695f $X=3.555 $Y=0.815 $X2=0
+ $Y2=0
cc_320 N_A_415_21#_c_303_p N_VGND_c_992_n 0.0188551f $X=3.72 $Y=0.39 $X2=0 $Y2=0
cc_321 N_A_415_21#_c_267_n N_VGND_c_992_n 0.00198695f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_322 N_A_415_21#_c_267_n N_VGND_c_994_n 0.00198695f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_323 N_A_415_21#_c_282_p N_VGND_c_994_n 0.0188551f $X=4.56 $Y=0.39 $X2=0 $Y2=0
cc_324 N_A_415_21#_M1008_d N_VGND_c_999_n 0.00215201f $X=3.585 $Y=0.235 $X2=0
+ $Y2=0
cc_325 N_A_415_21#_M1014_s N_VGND_c_999_n 0.00215201f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_415_21#_c_259_n N_VGND_c_999_n 0.00576327f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_415_21#_c_260_n N_VGND_c_999_n 0.0108251f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_A_415_21#_c_265_n N_VGND_c_999_n 0.00475876f $X=3.555 $Y=0.815 $X2=0
+ $Y2=0
cc_329 N_A_415_21#_c_266_n N_VGND_c_999_n 8.23161e-19 $X=3.145 $Y=0.815 $X2=0
+ $Y2=0
cc_330 N_A_415_21#_c_303_p N_VGND_c_999_n 0.0122069f $X=3.72 $Y=0.39 $X2=0 $Y2=0
cc_331 N_A_415_21#_c_267_n N_VGND_c_999_n 0.00835832f $X=4.395 $Y=0.815 $X2=0
+ $Y2=0
cc_332 N_A_415_21#_c_282_p N_VGND_c_999_n 0.0122069f $X=4.56 $Y=0.39 $X2=0 $Y2=0
cc_333 N_A_415_21#_c_259_n N_VGND_c_1000_n 0.00424416f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_415_21#_c_260_n N_VGND_c_1000_n 0.00541359f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A_415_21#_c_260_n N_VGND_c_1001_n 0.00335921f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_A_415_21#_c_261_n N_VGND_c_1001_n 0.00843619f $X=2.955 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_A_415_21#_c_262_n N_VGND_c_1001_n 0.0049954f $X=2.78 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_A_415_21#_c_265_n N_VGND_c_1001_n 0.0181768f $X=3.555 $Y=0.815 $X2=0
+ $Y2=0
cc_339 N_A_415_21#_c_266_n N_VGND_c_1001_n 0.0163451f $X=3.145 $Y=0.815 $X2=0
+ $Y2=0
cc_340 N_A1_N_c_402_n N_A2_N_c_488_n 0.0124239f $X=3.48 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_341 N_A1_N_M1009_g N_A2_N_M1012_g 0.0433788f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A1_N_c_406_n N_A2_N_M1012_g 0.0103235f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_343 A1_N N_A2_N_M1012_g 0.00235723f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_344 N_A1_N_c_398_n N_A2_N_c_489_n 0.0124239f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A1_N_M1023_g N_A2_N_M1015_g 0.0277801f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A1_N_c_406_n N_A2_N_M1015_g 0.0149047f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_347 N_A1_N_c_406_n N_A2_N_c_490_n 0.0399588f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_348 A1_N N_A2_N_c_490_n 0.0166516f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_349 A1_N N_A2_N_c_490_n 0.0174911f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_350 N_A1_N_c_401_n N_A2_N_c_490_n 7.27271e-19 $X=3.48 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A1_N_c_403_n N_A2_N_c_490_n 6.80324e-19 $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A1_N_c_406_n N_A2_N_c_491_n 0.00214031f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_353 A1_N N_A2_N_c_491_n 6.10557e-19 $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_354 A1_N N_A2_N_c_491_n 0.00465908f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_355 N_A1_N_c_401_n N_A2_N_c_491_n 0.022499f $X=3.48 $Y=1.16 $X2=0 $Y2=0
cc_356 N_A1_N_c_403_n N_A2_N_c_491_n 0.0223771f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_357 N_A1_N_c_398_n N_A_193_47#_c_536_n 0.01227f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A1_N_M1023_g N_A_193_47#_M1000_g 0.0279096f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_359 N_A1_N_c_406_n N_A_193_47#_M1000_g 8.81365e-19 $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_360 A1_N N_A_193_47#_c_607_n 0.0143593f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_361 N_A1_N_M1009_g N_A_193_47#_c_550_n 0.0029652f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_362 N_A1_N_c_406_n N_A_193_47#_c_550_n 0.0698351f $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_363 A1_N N_A_193_47#_c_550_n 0.0138643f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_364 N_A1_N_c_406_n N_A_193_47#_c_552_n 2.316e-19 $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_365 A1_N N_A_193_47#_c_552_n 2.15773e-19 $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_366 N_A1_N_M1023_g N_A_193_47#_c_553_n 3.60782e-19 $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_367 N_A1_N_c_406_n N_A_193_47#_c_553_n 0.0118726f $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_368 A1_N N_A_193_47#_c_553_n 0.0155882f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_369 A1_N N_A_193_47#_c_544_n 0.00235611f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_370 N_A1_N_c_403_n N_A_193_47#_c_544_n 0.02273f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_371 N_A1_N_c_406_n N_VPWR_M1023_d 0.0013609f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_372 N_A1_N_M1009_g N_VPWR_c_769_n 0.00502497f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_373 N_A1_N_M1023_g N_VPWR_c_770_n 0.00302074f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A1_N_c_406_n N_VPWR_c_770_n 0.0048223f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_375 N_A1_N_M1009_g N_VPWR_c_776_n 0.00441875f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_376 N_A1_N_M1023_g N_VPWR_c_776_n 0.00585385f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_377 N_A1_N_M1009_g N_VPWR_c_766_n 0.00721346f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_378 N_A1_N_M1023_g N_VPWR_c_766_n 0.0104912f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A1_N_c_406_n N_A_717_297#_M1009_s 0.00161973f $X=4.605 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_380 N_A1_N_c_406_n N_A_717_297#_M1015_d 0.00164852f $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_381 N_A1_N_c_406_n N_A_717_297#_c_891_n 0.0116235f $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_382 N_A1_N_c_398_n N_VGND_c_986_n 0.0015308f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_383 A1_N N_VGND_c_986_n 0.0057781f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_384 N_A1_N_c_403_n N_VGND_c_986_n 2.29798e-19 $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A1_N_c_402_n N_VGND_c_992_n 0.00423334f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A1_N_c_398_n N_VGND_c_994_n 0.00541359f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A1_N_c_398_n N_VGND_c_999_n 0.00955595f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_388 N_A1_N_c_402_n N_VGND_c_999_n 0.00706711f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_389 N_A1_N_c_402_n N_VGND_c_1001_n 0.00335921f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_390 N_A2_N_c_490_n N_A_193_47#_c_550_n 0.00443567f $X=4.145 $Y=1.16 $X2=0
+ $Y2=0
cc_391 N_A2_N_M1012_g N_VPWR_c_776_n 0.00357877f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A2_N_M1015_g N_VPWR_c_776_n 0.00357877f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A2_N_M1012_g N_VPWR_c_766_n 0.00525237f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A2_N_M1015_g N_VPWR_c_766_n 0.00525237f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_395 N_A2_N_M1012_g N_A_717_297#_c_885_n 0.00846708f $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_396 N_A2_N_M1015_g N_A_717_297#_c_885_n 0.0121306f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_397 N_A2_N_c_488_n N_VGND_c_985_n 0.00146339f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A2_N_c_489_n N_VGND_c_985_n 0.00146448f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A2_N_c_488_n N_VGND_c_992_n 0.00423334f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_400 N_A2_N_c_489_n N_VGND_c_994_n 0.00423334f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A2_N_c_488_n N_VGND_c_999_n 0.0057435f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A2_N_c_489_n N_VGND_c_999_n 0.0057435f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_403 N_A_193_47#_c_550_n N_A_27_297#_M1022_d 0.00324704f $X=5.17 $Y=1.53 $X2=0
+ $Y2=0
cc_404 N_A_193_47#_c_551_n N_A_27_297#_M1022_d 0.00116111f $X=2.68 $Y=1.53 $X2=0
+ $Y2=0
cc_405 N_A_193_47#_c_540_n N_A_27_297#_c_715_n 0.00630624f $X=2.195 $Y=0.82
+ $X2=0 $Y2=0
cc_406 N_A_193_47#_c_551_n N_A_27_297#_c_715_n 9.77976e-19 $X=2.68 $Y=1.53 $X2=0
+ $Y2=0
cc_407 N_A_193_47#_c_555_n N_A_27_297#_c_715_n 0.00223004f $X=2.36 $Y=1.62 $X2=0
+ $Y2=0
cc_408 N_A_193_47#_M1004_s N_A_27_297#_c_734_n 0.00312348f $X=2.225 $Y=1.485
+ $X2=0 $Y2=0
cc_409 N_A_193_47#_c_555_n N_A_27_297#_c_734_n 0.0166196f $X=2.36 $Y=1.62 $X2=0
+ $Y2=0
cc_410 N_A_193_47#_c_550_n N_A_27_297#_c_743_n 0.00769272f $X=5.17 $Y=1.53 $X2=0
+ $Y2=0
cc_411 N_A_193_47#_c_551_n N_A_27_297#_c_743_n 9.00065e-19 $X=2.68 $Y=1.53 $X2=0
+ $Y2=0
cc_412 N_A_193_47#_c_550_n N_VPWR_M1009_d 0.00104312f $X=5.17 $Y=1.53 $X2=0
+ $Y2=0
cc_413 N_A_193_47#_c_550_n N_VPWR_M1023_d 0.00154493f $X=5.17 $Y=1.53 $X2=0
+ $Y2=0
cc_414 N_A_193_47#_c_550_n N_VPWR_c_769_n 5.37033e-19 $X=5.17 $Y=1.53 $X2=0
+ $Y2=0
cc_415 N_A_193_47#_M1000_g N_VPWR_c_770_n 0.00157837f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_A_193_47#_c_550_n N_VPWR_c_770_n 0.00805046f $X=5.17 $Y=1.53 $X2=0
+ $Y2=0
cc_417 N_A_193_47#_M1000_g N_VPWR_c_771_n 0.00585385f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_A_193_47#_M1002_g N_VPWR_c_771_n 0.00585385f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_419 N_A_193_47#_M1002_g N_VPWR_c_772_n 0.00157837f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A_193_47#_M1005_g N_VPWR_c_772_n 0.00157837f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_421 N_A_193_47#_M1026_g N_VPWR_c_773_n 0.00338128f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_422 N_A_193_47#_M1005_g N_VPWR_c_780_n 0.00585385f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_423 N_A_193_47#_M1026_g N_VPWR_c_780_n 0.00585385f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_424 N_A_193_47#_M1004_s N_VPWR_c_766_n 0.00216833f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_425 N_A_193_47#_M1000_g N_VPWR_c_766_n 0.010464f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_426 N_A_193_47#_M1002_g N_VPWR_c_766_n 0.00588483f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_427 N_A_193_47#_M1005_g N_VPWR_c_766_n 0.00588483f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_428 N_A_193_47#_M1026_g N_VPWR_c_766_n 0.0117628f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_429 N_A_193_47#_c_550_n N_A_717_297#_c_891_n 0.00207359f $X=5.17 $Y=1.53
+ $X2=0 $Y2=0
cc_430 N_A_193_47#_c_552_n N_X_M1000_d 0.00470536f $X=5.315 $Y=1.53 $X2=0 $Y2=0
cc_431 N_A_193_47#_c_553_n N_X_M1000_d 0.00242139f $X=5.315 $Y=1.53 $X2=0 $Y2=0
cc_432 N_A_193_47#_c_536_n N_X_c_913_n 0.00494802f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_433 N_A_193_47#_c_537_n N_X_c_913_n 0.00612654f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A_193_47#_c_538_n N_X_c_913_n 5.16334e-19 $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_435 N_A_193_47#_M1002_g N_X_c_916_n 0.0113688f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_436 N_A_193_47#_M1005_g N_X_c_916_n 0.0113688f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_437 N_A_193_47#_c_653_p N_X_c_916_n 0.0140663f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_438 N_A_193_47#_c_544_n N_X_c_916_n 0.00166652f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_439 N_A_193_47#_c_653_p N_X_c_920_n 0.0011835f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_440 N_A_193_47#_c_552_n N_X_c_920_n 0.00546229f $X=5.315 $Y=1.53 $X2=0 $Y2=0
cc_441 N_A_193_47#_c_553_n N_X_c_920_n 0.0107118f $X=5.315 $Y=1.53 $X2=0 $Y2=0
cc_442 N_A_193_47#_c_544_n N_X_c_920_n 3.77487e-19 $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A_193_47#_c_537_n N_X_c_901_n 0.00870364f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_444 N_A_193_47#_c_538_n N_X_c_901_n 0.00870364f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_445 N_A_193_47#_c_653_p N_X_c_901_n 0.0356734f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_446 N_A_193_47#_c_544_n N_X_c_901_n 0.00222133f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_447 N_A_193_47#_c_536_n N_X_c_902_n 0.00259239f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_448 N_A_193_47#_c_537_n N_X_c_902_n 0.00113229f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_449 N_A_193_47#_c_607_n N_X_c_902_n 0.018801f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_450 N_A_193_47#_c_653_p N_X_c_902_n 0.00824993f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_451 N_A_193_47#_c_552_n N_X_c_902_n 9.35813e-19 $X=5.315 $Y=1.53 $X2=0 $Y2=0
cc_452 N_A_193_47#_c_544_n N_X_c_902_n 0.00229945f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_453 N_A_193_47#_c_537_n N_X_c_934_n 5.16334e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_454 N_A_193_47#_c_538_n N_X_c_934_n 0.00612654f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_455 N_A_193_47#_c_539_n N_X_c_934_n 0.0107369f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_456 N_A_193_47#_c_539_n N_X_c_903_n 0.011353f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_457 N_A_193_47#_c_653_p N_X_c_903_n 0.00234861f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_458 N_A_193_47#_c_538_n N_X_c_904_n 0.00113229f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_459 N_A_193_47#_c_539_n N_X_c_904_n 0.00113229f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_460 N_A_193_47#_c_653_p N_X_c_904_n 0.0261859f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_461 N_A_193_47#_c_544_n N_X_c_904_n 0.00230115f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_193_47#_M1005_g N_X_c_906_n 0.00102706f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_463 N_A_193_47#_M1026_g N_X_c_906_n 2.9179e-19 $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_464 N_A_193_47#_c_653_p N_X_c_906_n 0.0200119f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_465 N_A_193_47#_c_553_n N_X_c_906_n 0.00239492f $X=5.315 $Y=1.53 $X2=0 $Y2=0
cc_466 N_A_193_47#_c_544_n N_X_c_906_n 0.00231083f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_467 N_A_193_47#_c_539_n X 0.019973f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_468 N_A_193_47#_c_653_p X 0.0140302f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_193_47#_M1026_g X 0.0184691f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_470 N_A_193_47#_c_653_p X 0.00526128f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_471 N_A_193_47#_c_540_n N_VGND_M1027_d 0.00165819f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_472 N_A_193_47#_c_540_n N_VGND_c_984_n 0.0116529f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_473 N_A_193_47#_c_536_n N_VGND_c_986_n 0.0015308f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_193_47#_c_550_n N_VGND_c_986_n 0.00388941f $X=5.17 $Y=1.53 $X2=0
+ $Y2=0
cc_475 N_A_193_47#_c_536_n N_VGND_c_987_n 0.00542163f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_A_193_47#_c_537_n N_VGND_c_987_n 0.00424138f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_477 N_A_193_47#_c_537_n N_VGND_c_988_n 0.00146448f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_193_47#_c_538_n N_VGND_c_988_n 0.00146448f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_A_193_47#_c_539_n N_VGND_c_989_n 0.00316354f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_A_193_47#_c_540_n N_VGND_c_990_n 0.00194318f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_481 N_A_193_47#_c_538_n N_VGND_c_996_n 0.00424138f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_482 N_A_193_47#_c_539_n N_VGND_c_996_n 0.00424138f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_193_47#_M1013_d N_VGND_c_999_n 0.00216833f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_484 N_A_193_47#_M1020_s N_VGND_c_999_n 0.00215201f $X=2.225 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_193_47#_c_536_n N_VGND_c_999_n 0.00952972f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_486 N_A_193_47#_c_537_n N_VGND_c_999_n 0.00571728f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_487 N_A_193_47#_c_538_n N_VGND_c_999_n 0.00571728f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_A_193_47#_c_539_n N_VGND_c_999_n 0.00704335f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_489 N_A_193_47#_c_540_n N_VGND_c_999_n 0.00922137f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_490 N_A_193_47#_c_560_n N_VGND_c_999_n 0.0122165f $X=2.36 $Y=0.39 $X2=0 $Y2=0
cc_491 N_A_193_47#_c_540_n N_VGND_c_1000_n 0.00193763f $X=2.195 $Y=0.82 $X2=0
+ $Y2=0
cc_492 N_A_193_47#_c_560_n N_VGND_c_1000_n 0.0188914f $X=2.36 $Y=0.39 $X2=0
+ $Y2=0
cc_493 N_A_193_47#_c_540_n N_A_109_47#_M1018_s 0.00195168f $X=2.195 $Y=0.82
+ $X2=0 $Y2=0
cc_494 N_A_193_47#_c_542_n N_A_109_47#_c_1102_n 0.0105363f $X=1.1 $Y=0.73 $X2=0
+ $Y2=0
cc_495 N_A_193_47#_M1013_d N_A_109_47#_c_1107_n 0.00304656f $X=0.965 $Y=0.235
+ $X2=0 $Y2=0
cc_496 N_A_193_47#_c_540_n N_A_109_47#_c_1107_n 0.0141805f $X=2.195 $Y=0.82
+ $X2=0 $Y2=0
cc_497 N_A_193_47#_c_542_n N_A_109_47#_c_1107_n 0.0156278f $X=1.1 $Y=0.73 $X2=0
+ $Y2=0
cc_498 N_A_27_297#_c_718_n N_VPWR_M1019_d 0.00328796f $X=0.975 $Y=1.87 $X2=-0.19
+ $Y2=1.305
cc_499 N_A_27_297#_c_723_n N_VPWR_M1003_d 0.00325391f $X=1.815 $Y=1.87 $X2=0
+ $Y2=0
cc_500 N_A_27_297#_c_718_n N_VPWR_c_767_n 0.0123301f $X=0.975 $Y=1.87 $X2=0
+ $Y2=0
cc_501 N_A_27_297#_c_723_n N_VPWR_c_768_n 0.0123301f $X=1.815 $Y=1.87 $X2=0
+ $Y2=0
cc_502 N_A_27_297#_c_743_n N_VPWR_c_769_n 0.0180653f $X=2.78 $Y=2.3 $X2=0 $Y2=0
cc_503 N_A_27_297#_c_734_n N_VPWR_c_774_n 0.0330174f $X=2.655 $Y=2.38 $X2=0
+ $Y2=0
cc_504 N_A_27_297#_c_751_p N_VPWR_c_774_n 0.0143053f $X=2.065 $Y=2.38 $X2=0
+ $Y2=0
cc_505 N_A_27_297#_c_743_n N_VPWR_c_774_n 0.0151213f $X=2.78 $Y=2.3 $X2=0 $Y2=0
cc_506 N_A_27_297#_c_753_p N_VPWR_c_778_n 0.0158369f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_507 N_A_27_297#_c_754_p N_VPWR_c_779_n 0.0142343f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_508 N_A_27_297#_M1019_s N_VPWR_c_766_n 0.00212725f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_509 N_A_27_297#_M1001_s N_VPWR_c_766_n 0.00223619f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_510 N_A_27_297#_M1025_s N_VPWR_c_766_n 0.00220214f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_511 N_A_27_297#_M1022_d N_VPWR_c_766_n 0.00207714f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_512 N_A_27_297#_c_753_p N_VPWR_c_766_n 0.00955092f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_513 N_A_27_297#_c_718_n N_VPWR_c_766_n 0.0109281f $X=0.975 $Y=1.87 $X2=0
+ $Y2=0
cc_514 N_A_27_297#_c_754_p N_VPWR_c_766_n 0.00955092f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_515 N_A_27_297#_c_723_n N_VPWR_c_766_n 0.0109281f $X=1.815 $Y=1.87 $X2=0
+ $Y2=0
cc_516 N_A_27_297#_c_734_n N_VPWR_c_766_n 0.0204667f $X=2.655 $Y=2.38 $X2=0
+ $Y2=0
cc_517 N_A_27_297#_c_751_p N_VPWR_c_766_n 0.00962271f $X=2.065 $Y=2.38 $X2=0
+ $Y2=0
cc_518 N_A_27_297#_c_743_n N_VPWR_c_766_n 0.00938089f $X=2.78 $Y=2.3 $X2=0 $Y2=0
cc_519 N_VPWR_c_766_n N_A_717_297#_M1009_s 0.00219818f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_520 N_VPWR_c_766_n N_A_717_297#_M1015_d 0.00246446f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_776_n N_A_717_297#_c_885_n 0.0473226f $X=4.855 $Y=2.72 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_766_n N_A_717_297#_c_885_n 0.0300947f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_776_n N_A_717_297#_c_888_n 0.0136817f $X=4.855 $Y=2.72 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_766_n N_A_717_297#_c_888_n 0.00938089f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_766_n N_X_M1000_d 0.00254126f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_526 N_VPWR_c_766_n N_X_M1005_d 0.00254126f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_527 N_VPWR_c_771_n N_X_c_954_n 0.0142343f $X=5.695 $Y=2.72 $X2=0 $Y2=0
cc_528 N_VPWR_c_766_n N_X_c_954_n 0.00955092f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_529 N_VPWR_M1002_s N_X_c_916_n 0.00441488f $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_530 N_VPWR_c_772_n N_X_c_916_n 0.0102703f $X=5.82 $Y=2.33 $X2=0 $Y2=0
cc_531 N_VPWR_c_766_n N_X_c_916_n 0.0110299f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_532 N_VPWR_c_780_n N_X_c_959_n 0.0142343f $X=6.535 $Y=2.72 $X2=0 $Y2=0
cc_533 N_VPWR_c_766_n N_X_c_959_n 0.00955092f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_534 N_VPWR_M1026_s X 2.90082e-19 $X=6.525 $Y=1.485 $X2=0 $Y2=0
cc_535 N_VPWR_c_773_n X 0.00229378f $X=6.66 $Y=1.99 $X2=0 $Y2=0
cc_536 N_VPWR_M1026_s N_X_c_909_n 0.00267829f $X=6.525 $Y=1.485 $X2=0 $Y2=0
cc_537 N_VPWR_c_773_n N_X_c_909_n 0.0156881f $X=6.66 $Y=1.99 $X2=0 $Y2=0
cc_538 N_X_c_901_n N_VGND_M1010_s 0.00162089f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_539 N_X_c_903_n N_VGND_M1017_s 0.00324195f $X=6.61 $Y=0.815 $X2=0 $Y2=0
cc_540 N_X_c_902_n N_VGND_c_986_n 0.00750114f $X=5.565 $Y=0.815 $X2=0 $Y2=0
cc_541 N_X_c_913_n N_VGND_c_987_n 0.0167046f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_542 N_X_c_901_n N_VGND_c_987_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_543 N_X_c_901_n N_VGND_c_988_n 0.0122559f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_544 N_X_c_903_n N_VGND_c_989_n 0.013754f $X=6.61 $Y=0.815 $X2=0 $Y2=0
cc_545 N_X_c_901_n N_VGND_c_996_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_546 N_X_c_934_n N_VGND_c_996_n 0.0167046f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_547 N_X_c_903_n N_VGND_c_996_n 0.00198695f $X=6.61 $Y=0.815 $X2=0 $Y2=0
cc_548 N_X_c_903_n N_VGND_c_998_n 0.00293286f $X=6.61 $Y=0.815 $X2=0 $Y2=0
cc_549 N_X_M1006_d N_VGND_c_999_n 0.00216035f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_550 N_X_M1011_d N_VGND_c_999_n 0.00216035f $X=6.105 $Y=0.235 $X2=0 $Y2=0
cc_551 N_X_c_913_n N_VGND_c_999_n 0.0120721f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_552 N_X_c_901_n N_VGND_c_999_n 0.00835832f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_553 N_X_c_934_n N_VGND_c_999_n 0.0120721f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_554 N_X_c_903_n N_VGND_c_999_n 0.00953573f $X=6.61 $Y=0.815 $X2=0 $Y2=0
cc_555 N_VGND_c_999_n N_A_109_47#_M1016_s 0.00215206f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_556 N_VGND_c_999_n N_A_109_47#_M1018_s 0.00215227f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_990_n N_A_109_47#_c_1103_n 0.015211f $X=1.855 $Y=0 $X2=0 $Y2=0
cc_558 N_VGND_c_999_n N_A_109_47#_c_1103_n 0.00940707f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_983_n N_A_109_47#_c_1102_n 0.0154056f $X=0.26 $Y=0.39 $X2=0
+ $Y2=0
cc_560 N_VGND_c_990_n N_A_109_47#_c_1107_n 0.0504977f $X=1.855 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_999_n N_A_109_47#_c_1107_n 0.0327385f $X=7.13 $Y=0 $X2=0 $Y2=0

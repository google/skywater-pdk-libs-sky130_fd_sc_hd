* File: sky130_fd_sc_hd__nand4_1.pex.spice
* Created: Thu Aug 27 14:30:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4_1%D 1 3 6 8 14
r25 11 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r26 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r27 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r29 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_1%C 1 3 6 8 9 10 15 16
r39 17 24 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=0.702 $Y=0.995
+ $X2=0.702 $Y2=1.16
r40 16 24 6.56543 $w=3.28e-07 $l=1.88e-07 $layer=LI1_cond $X=0.89 $Y=1.16
+ $X2=0.702 $Y2=1.16
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r42 10 24 0.244458 $w=3.28e-07 $l=7e-09 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.702 $Y2=1.16
r43 9 17 7.77229 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=0.702 $Y=0.85
+ $X2=0.702 $Y2=0.995
r44 8 9 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=0.702 $Y=0.51
+ $X2=0.702 $Y2=0.85
r45 4 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r46 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r47 1 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_1%B 3 6 9 13 14 16 19
r43 16 24 12.3335 $w=3.48e-07 $l=3.15e-07 $layer=LI1_cond $X=1.175 $Y=0.51
+ $X2=1.175 $Y2=0.825
r44 14 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.37 $Y2=1.325
r45 14 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.37 $Y2=0.995
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r47 10 13 4.29547 $w=3.28e-07 $l=1.23e-07 $layer=LI1_cond $X=1.247 $Y=1.16
+ $X2=1.37 $Y2=1.16
r48 9 10 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=1.247 $Y=0.995
+ $X2=1.247 $Y2=1.16
r49 9 24 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=1.247 $Y=0.995
+ $X2=1.247 $Y2=0.825
r50 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.985
+ $X2=1.31 $Y2=1.325
r51 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.56 $X2=1.31
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_1%A 1 3 6 8 9 15
r28 12 15 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.79 $Y=1.16
+ $X2=2.06 $Y2=1.16
r29 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.095 $Y=1.16
+ $X2=2.095 $Y2=1.53
r30 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r31 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.325
+ $X2=1.79 $Y2=1.16
r32 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.79 $Y=1.325 $X2=1.79
+ $Y2=1.985
r33 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=0.995
+ $X2=1.79 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.79 $Y=0.995 $X2=1.79
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_1%VPWR 1 2 3 10 12 18 20 22 25 26 27 33 42
r36 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r39 33 41 4.29523 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.107 $Y2=2.72
r40 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.61 $Y2=2.72
r41 32 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 29 38 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r44 29 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 27 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 27 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r47 25 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72 $X2=1.1
+ $Y2=2.72
r49 24 35 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72 $X2=1.1
+ $Y2=2.72
r51 20 41 3.06482 $w=2.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.107 $Y2=2.72
r52 20 22 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2
r53 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r54 16 18 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r55 12 15 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r56 10 38 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r57 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r58 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.485 $X2=2 $Y2=2
r59 2 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r60 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r61 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_1%Y 1 2 3 10 12 14 18 21 25 26 29
c46 21 0 1.04363e-19 $X=1.71 $Y=1.495
r47 26 33 13.3545 $w=6.93e-07 $l=3.15e-07 $layer=LI1_cond $X=1.867 $Y=0.51
+ $X2=1.867 $Y2=0.825
r48 26 29 2.23727 $w=6.93e-07 $l=1.3e-07 $layer=LI1_cond $X=1.867 $Y=0.51
+ $X2=1.867 $Y2=0.38
r49 21 25 3.70735 $w=2.5e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.71 $Y=1.495
+ $X2=1.59 $Y2=1.58
r50 21 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.71 $Y=1.495
+ $X2=1.71 $Y2=0.825
r51 16 25 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.55 $Y=1.665
+ $X2=1.59 $Y2=1.58
r52 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.55 $Y=1.665
+ $X2=1.55 $Y2=2.34
r53 15 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.58
+ $X2=0.68 $Y2=1.58
r54 14 25 2.76166 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.385 $Y=1.58
+ $X2=1.59 $Y2=1.58
r55 14 15 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.385 $Y=1.58
+ $X2=0.845 $Y2=1.58
r56 10 23 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.665 $X2=0.68
+ $Y2=1.58
r57 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r58 3 25 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.55 $Y2=1.66
r59 3 18 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.55 $Y2=2.34
r60 2 23 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r61 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r62 1 29 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.865
+ $Y=0.235 $X2=2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_1%VGND 1 4 6 8 15 16
r27 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r28 13 16 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r29 12 15 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r30 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r31 10 19 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r32 10 12 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r33 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r34 8 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r35 4 19 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r36 4 6 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r37 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a311o_4.spice.pex
* Created: Thu Aug 27 14:04:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A311O_4%C1 1 3 6 8 10 13 15 16 17 26
r43 25 26 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r44 22 25 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r45 16 17 19.8327 $w=2.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.16
+ $X2=0.242 $Y2=1.53
r46 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r47 15 16 16.6166 $w=2.13e-07 $l=3.1e-07 $layer=LI1_cond $X=0.242 $Y=0.85
+ $X2=0.242 $Y2=1.16
r48 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r50 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r52 4 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r54 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%B1 1 3 6 8 10 13 15 16 23 24
c54 24 0 2.54221e-20 $X=1.73 $Y=1.135
c55 23 0 3.79813e-20 $X=1.34 $Y=1.16
c56 6 0 2.2886e-20 $X=1.31 $Y=1.985
r57 26 32 1.19342 $w=1.95e-07 $l=1.05e-07 $layer=LI1_cond $X=1.157 $Y=1.285
+ $X2=1.157 $Y2=1.18
r58 23 32 9.66494 $w=2.08e-07 $l=1.83e-07 $layer=LI1_cond $X=1.34 $Y=1.18
+ $X2=1.157 $Y2=1.18
r59 22 24 70.327 $w=3.2e-07 $l=3.9e-07 $layer=POLY_cond $X=1.34 $Y=1.135
+ $X2=1.73 $Y2=1.135
r60 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=1.16 $X2=1.34 $Y2=1.16
r61 19 22 5.40977 $w=3.2e-07 $l=3e-08 $layer=POLY_cond $X=1.31 $Y=1.135 $X2=1.34
+ $Y2=1.135
r62 16 26 13.9347 $w=1.93e-07 $l=2.45e-07 $layer=LI1_cond $X=1.157 $Y=1.53
+ $X2=1.157 $Y2=1.285
r63 15 32 0.105628 $w=2.08e-07 $l=2e-09 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=1.157 $Y2=1.18
r64 11 24 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.135
r65 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r66 8 24 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.73 $Y=0.975
+ $X2=1.73 $Y2=1.135
r67 8 10 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.73 $Y=0.975
+ $X2=1.73 $Y2=0.56
r68 4 19 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.135
r69 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295 $X2=1.31
+ $Y2=1.985
r70 1 19 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.31 $Y=0.975
+ $X2=1.31 $Y2=1.135
r71 1 3 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.31 $Y=0.975
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A_109_47# 1 2 3 4 15 17 18 19 21 24 26 28 31
+ 33 35 36 38 39 41 47 48 52 55 56 58 61 64 67 68 69 71 73 76 81 84 87
c201 64 0 2.37016e-19 $X=3.78 $Y=1.16
c202 47 0 2.2886e-20 $X=0.68 $Y=1.7
c203 18 0 2.63538e-20 $X=2.225 $Y=1.16
c204 15 0 9.19584e-20 $X=2.15 $Y=0.56
r205 94 95 11.9012 $w=3.24e-07 $l=8e-08 $layer=POLY_cond $X=3.43 $Y=1.202
+ $X2=3.51 $Y2=1.202
r206 70 87 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.6 $Y=0.825 $X2=6.6
+ $Y2=0.735
r207 70 71 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.6 $Y=0.825
+ $X2=6.6 $Y2=1.455
r208 68 71 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.515 $Y=1.54
+ $X2=6.6 $Y2=1.455
r209 68 69 143.203 $w=1.68e-07 $l=2.195e-06 $layer=LI1_cond $X=6.515 $Y=1.54
+ $X2=4.32 $Y2=1.54
r210 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.235 $Y=1.455
+ $X2=4.32 $Y2=1.54
r211 66 67 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.235 $Y=1.245
+ $X2=4.235 $Y2=1.455
r212 64 97 22.3148 $w=3.24e-07 $l=1.5e-07 $layer=POLY_cond $X=3.78 $Y=1.202
+ $X2=3.93 $Y2=1.202
r213 64 95 40.1667 $w=3.24e-07 $l=2.7e-07 $layer=POLY_cond $X=3.78 $Y=1.202
+ $X2=3.51 $Y2=1.202
r214 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.78
+ $Y=1.16 $X2=3.78 $Y2=1.16
r215 61 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.15 $Y=1.16
+ $X2=4.235 $Y2=1.245
r216 61 63 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.15 $Y=1.16
+ $X2=3.78 $Y2=1.16
r217 59 90 7.43827 $w=3.24e-07 $l=5e-08 $layer=POLY_cond $X=2.54 $Y=1.202
+ $X2=2.59 $Y2=1.202
r218 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.54
+ $Y=1.16 $X2=2.54 $Y2=1.16
r219 56 58 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.025 $Y=1.16
+ $X2=2.54 $Y2=1.16
r220 55 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=1.075
+ $X2=2.025 $Y2=1.16
r221 54 55 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.94 $Y=0.885
+ $X2=1.94 $Y2=1.075
r222 53 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.8
+ $X2=1.52 $Y2=0.8
r223 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.855 $Y=0.8
+ $X2=1.94 $Y2=0.885
r224 52 53 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.855 $Y=0.8
+ $X2=1.605 $Y2=0.8
r225 51 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.715
+ $X2=1.52 $Y2=0.8
r226 50 81 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.465
+ $X2=1.52 $Y2=0.38
r227 50 51 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.52 $Y=0.465
+ $X2=1.52 $Y2=0.715
r228 49 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.8
+ $X2=0.68 $Y2=0.8
r229 48 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0.8
+ $X2=1.52 $Y2=0.8
r230 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=0.8
+ $X2=0.765 $Y2=0.8
r231 45 76 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.955
+ $X2=0.68 $Y2=2.04
r232 45 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.68 $Y=1.955
+ $X2=0.68 $Y2=1.7
r233 44 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.885
+ $X2=0.68 $Y2=0.8
r234 44 47 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=0.68 $Y=0.885
+ $X2=0.68 $Y2=1.7
r235 43 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.715
+ $X2=0.68 $Y2=0.8
r236 42 73 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.465
+ $X2=0.68 $Y2=0.38
r237 42 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.68 $Y=0.465
+ $X2=0.68 $Y2=0.715
r238 39 97 20.7868 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.93 $Y=1.41
+ $X2=3.93 $Y2=1.202
r239 39 41 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.93 $Y=1.41
+ $X2=3.93 $Y2=1.985
r240 36 95 20.7868 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.51 $Y=1.41
+ $X2=3.51 $Y2=1.202
r241 36 38 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.51 $Y=1.41
+ $X2=3.51 $Y2=1.985
r242 33 94 20.7868 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.202
r243 33 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
r244 29 94 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=3.09 $Y=1.202
+ $X2=3.43 $Y2=1.202
r245 29 92 11.9012 $w=3.24e-07 $l=8e-08 $layer=POLY_cond $X=3.09 $Y=1.202
+ $X2=3.01 $Y2=1.202
r246 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.985
r247 26 92 20.7868 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=1.202
r248 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r249 22 92 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=2.67 $Y=1.202
+ $X2=3.01 $Y2=1.202
r250 22 90 11.9012 $w=3.24e-07 $l=8e-08 $layer=POLY_cond $X=2.67 $Y=1.202
+ $X2=2.59 $Y2=1.202
r251 22 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.985
r252 19 90 20.7868 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.202
r253 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r254 17 59 5.20011 $w=3.24e-07 $l=5.30471e-08 $layer=POLY_cond $X=2.515 $Y=1.16
+ $X2=2.54 $Y2=1.202
r255 17 18 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.515 $Y=1.16
+ $X2=2.225 $Y2=1.16
r256 13 18 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.225 $Y2=1.16
r257 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r258 4 76 600 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.04
r259 4 47 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.7
r260 3 87 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=6.545
+ $Y=0.235 $X2=6.68 $Y2=0.74
r261 2 84 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.72
r262 2 81 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r263 1 79 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.72
r264 1 73 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A3 1 3 4 6 7 9 10 12 13 19
c51 13 0 9.4401e-20 $X=4.855 $Y=1.19
r52 19 21 10.927 $w=3.97e-07 $l=9e-08 $layer=POLY_cond $X=4.68 $Y=1.185 $X2=4.77
+ $Y2=1.185
r53 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.68
+ $Y=1.16 $X2=4.68 $Y2=1.16
r54 17 19 3.64232 $w=3.97e-07 $l=3e-08 $layer=POLY_cond $X=4.65 $Y=1.185
+ $X2=4.68 $Y2=1.185
r55 16 17 36.4232 $w=3.97e-07 $l=3e-07 $layer=POLY_cond $X=4.35 $Y=1.185
+ $X2=4.65 $Y2=1.185
r56 13 20 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=4.855 $Y=1.18
+ $X2=4.68 $Y2=1.18
r57 10 21 25.678 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.77 $Y=1.41
+ $X2=4.77 $Y2=1.185
r58 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.77 $Y=1.41
+ $X2=4.77 $Y2=1.985
r59 7 17 25.678 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.65 $Y=0.96 $X2=4.65
+ $Y2=1.185
r60 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.65 $Y=0.96 $X2=4.65
+ $Y2=0.56
r61 4 16 25.678 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.35 $Y=1.41 $X2=4.35
+ $Y2=1.185
r62 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.35 $Y=1.41 $X2=4.35
+ $Y2=1.985
r63 1 16 14.5693 $w=3.97e-07 $l=2.78613e-07 $layer=POLY_cond $X=4.23 $Y=0.96
+ $X2=4.35 $Y2=1.185
r64 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.23 $Y=0.96 $X2=4.23
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A2 3 7 11 15 17 18 28
r46 26 28 38.8804 $w=2.7e-07 $l=1.75e-07 $layer=POLY_cond $X=5.875 $Y=1.16
+ $X2=6.05 $Y2=1.16
r47 24 26 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=5.67 $Y=1.16
+ $X2=5.875 $Y2=1.16
r48 23 24 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=5.63 $Y=1.16 $X2=5.67
+ $Y2=1.16
r49 21 23 84.426 $w=2.7e-07 $l=3.8e-07 $layer=POLY_cond $X=5.25 $Y=1.16 $X2=5.63
+ $Y2=1.16
r50 18 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.875
+ $Y=1.16 $X2=5.875 $Y2=1.16
r51 17 18 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=5.375 $Y=1.18
+ $X2=5.835 $Y2=1.18
r52 13 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.05 $Y=1.025
+ $X2=6.05 $Y2=1.16
r53 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.05 $Y=1.025
+ $X2=6.05 $Y2=0.56
r54 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.67 $Y=1.295
+ $X2=5.67 $Y2=1.16
r55 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.67 $Y=1.295
+ $X2=5.67 $Y2=1.985
r56 5 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.63 $Y=1.025
+ $X2=5.63 $Y2=1.16
r57 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.63 $Y=1.025
+ $X2=5.63 $Y2=0.56
r58 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.25 $Y=1.295
+ $X2=5.25 $Y2=1.16
r59 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.25 $Y=1.295 $X2=5.25
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A1 1 3 6 8 10 13 15 16 23
r49 21 23 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=6.89 $Y=1.16
+ $X2=7.11 $Y2=1.16
r50 19 21 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.47 $Y=1.16
+ $X2=6.89 $Y2=1.16
r51 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.11 $Y=1.16
+ $X2=7.11 $Y2=1.53
r52 15 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.11
+ $Y=1.16 $X2=7.11 $Y2=1.16
r53 11 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.16
r54 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.985
r55 8 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=1.16
r56 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=0.56
r57 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.47 $Y=1.325
+ $X2=6.47 $Y2=1.16
r58 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.47 $Y=1.325 $X2=6.47
+ $Y2=1.985
r59 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.47 $Y=0.995
+ $X2=6.47 $Y2=1.16
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.47 $Y=0.995 $X2=6.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A_27_297# 1 2 3 12 14 15 18 20 24 26
c33 18 0 6.34034e-20 $X=1.1 $Y=1.96
r34 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=1.94 $Y2=1.96
r35 21 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.38 $X2=1.1
+ $Y2=2.38
r36 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.855 $Y=2.38
+ $X2=1.94 $Y2=2.295
r37 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=2.38
+ $X2=1.185 $Y2=2.38
r38 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.295 $X2=1.1
+ $Y2=2.38
r39 16 18 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=2.295
+ $X2=1.1 $Y2=1.96
r40 14 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.38 $X2=1.1
+ $Y2=2.38
r41 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=2.38
+ $X2=0.345 $Y2=2.38
r42 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.345 $Y2=2.38
r43 10 12 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=1.96
r44 3 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r45 2 18 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r46 1 12 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A_277_297# 1 2 3 4 15 17 18 20 21 22 25 27
+ 31 33 35 37 40 42
c90 21 0 1.42615e-19 $X=4.475 $Y=2
r91 35 44 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.68 $Y=2.085
+ $X2=6.68 $Y2=1.94
r92 35 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.68 $Y=2.085
+ $X2=6.68 $Y2=2.3
r93 34 42 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.545 $Y=2
+ $X2=5.46 $Y2=1.94
r94 33 44 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=6.595 $Y=2
+ $X2=6.68 $Y2=1.94
r95 33 34 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=6.595 $Y=2
+ $X2=5.545 $Y2=2
r96 29 42 1.34256 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.46 $Y=2.085
+ $X2=5.46 $Y2=1.94
r97 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.46 $Y=2.085
+ $X2=5.46 $Y2=2.3
r98 28 40 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.645 $Y=2
+ $X2=4.56 $Y2=1.94
r99 27 42 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.375 $Y=2
+ $X2=5.46 $Y2=1.94
r100 27 28 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.375 $Y=2
+ $X2=4.645 $Y2=2
r101 23 40 1.34256 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.56 $Y=2.085
+ $X2=4.56 $Y2=1.94
r102 23 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.56 $Y=2.085
+ $X2=4.56 $Y2=2.3
r103 21 40 5.16603 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.475 $Y=2
+ $X2=4.56 $Y2=1.94
r104 21 22 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=4.475 $Y=2
+ $X2=2.385 $Y2=2
r105 20 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.29 $Y=1.915
+ $X2=2.385 $Y2=2
r106 19 20 16.9282 $w=1.88e-07 $l=2.9e-07 $layer=LI1_cond $X=2.29 $Y=1.625
+ $X2=2.29 $Y2=1.915
r107 17 19 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.195 $Y=1.54
+ $X2=2.29 $Y2=1.625
r108 17 18 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.195 $Y=1.54
+ $X2=1.605 $Y2=1.54
r109 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.52 $Y=1.625
+ $X2=1.605 $Y2=1.54
r110 13 15 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=1.625
+ $X2=1.52 $Y2=1.96
r111 4 44 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=6.545
+ $Y=1.485 $X2=6.68 $Y2=1.96
r112 4 37 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.545
+ $Y=1.485 $X2=6.68 $Y2=2.3
r113 3 42 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.485 $X2=5.46 $Y2=1.96
r114 3 31 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.485 $X2=5.46 $Y2=2.3
r115 2 40 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.96
r116 2 25 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2.3
r117 1 15 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 37 41 43 45
+ 48 49 50 51 52 54 69 75 78 81 85
r126 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r127 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r128 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r129 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r130 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r131 73 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r132 73 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r133 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r134 70 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.045 $Y=2.72
+ $X2=5.88 $Y2=2.72
r135 70 72 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.045 $Y=2.72
+ $X2=6.67 $Y2=2.72
r136 69 84 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=6.935 $Y=2.72
+ $X2=7.147 $Y2=2.72
r137 69 72 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.935 $Y=2.72
+ $X2=6.67 $Y2=2.72
r138 68 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r139 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r140 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r141 65 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r142 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r143 62 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=2.72
+ $X2=2.46 $Y2=2.72
r144 62 64 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=2.72
+ $X2=2.99 $Y2=2.72
r145 61 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r146 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r147 56 60 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r148 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.46 $Y2=2.72
r149 54 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.07 $Y2=2.72
r150 52 61 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r151 52 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r152 50 67 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=3.91 $Y2=2.72
r153 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=4.14 $Y2=2.72
r154 48 64 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=2.99 $Y2=2.72
r155 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.3 $Y2=2.72
r156 47 67 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.91 $Y2=2.72
r157 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.3 $Y2=2.72
r158 43 84 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=7.102 $Y=2.635
+ $X2=7.147 $Y2=2.72
r159 43 45 25.973 $w=3.33e-07 $l=7.55e-07 $layer=LI1_cond $X=7.102 $Y=2.635
+ $X2=7.102 $Y2=1.88
r160 39 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.88 $Y=2.635
+ $X2=5.88 $Y2=2.72
r161 39 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.88 $Y=2.635
+ $X2=5.88 $Y2=2.34
r162 38 78 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.175 $Y=2.72
+ $X2=4.995 $Y2=2.72
r163 37 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=2.72
+ $X2=5.88 $Y2=2.72
r164 37 38 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.715 $Y=2.72
+ $X2=5.175 $Y2=2.72
r165 33 78 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=2.635
+ $X2=4.995 $Y2=2.72
r166 33 35 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=4.995 $Y=2.635
+ $X2=4.995 $Y2=2.34
r167 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.14 $Y2=2.72
r168 31 78 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.815 $Y=2.72
+ $X2=4.995 $Y2=2.72
r169 31 32 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.815 $Y=2.72
+ $X2=4.305 $Y2=2.72
r170 27 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.72
r171 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.34
r172 23 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.635 $X2=3.3
+ $Y2=2.72
r173 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.3 $Y=2.635
+ $X2=3.3 $Y2=2.34
r174 19 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.72
r175 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.34
r176 6 45 300 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_PDIFF $count=2 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=1.88
r177 5 41 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=1.485 $X2=5.88 $Y2=2.34
r178 4 35 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2.34
r179 3 29 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2.34
r180 2 25 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=2.34
r181 1 21 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%X 1 2 3 4 14 15 19 24 30 32 33 39 43 48
c56 32 0 9.19584e-20 $X=3.015 $Y=0.85
r57 39 43 0.853147 $w=1.93e-07 $l=1.5e-08 $layer=LI1_cond $X=3.007 $Y=1.545
+ $X2=3.007 $Y2=1.53
r58 33 39 3.31084 $w=1.95e-07 $l=1.32868e-07 $layer=LI1_cond $X=2.91 $Y=1.63
+ $X2=3.007 $Y2=1.545
r59 33 43 1.99068 $w=1.93e-07 $l=3.5e-08 $layer=LI1_cond $X=3.007 $Y=1.495
+ $X2=3.007 $Y2=1.53
r60 32 48 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.015 $Y=0.8
+ $X2=3.22 $Y2=0.8
r61 32 38 0.521925 $w=1.68e-07 $l=8e-09 $layer=LI1_cond $X=3.015 $Y=0.8
+ $X2=3.007 $Y2=0.8
r62 32 33 33.2727 $w=1.93e-07 $l=5.85e-07 $layer=LI1_cond $X=3.007 $Y=0.91
+ $X2=3.007 $Y2=1.495
r63 32 38 1.42191 $w=1.93e-07 $l=2.5e-08 $layer=LI1_cond $X=3.007 $Y=0.91
+ $X2=3.007 $Y2=0.885
r64 24 26 5.85433 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=0.38
+ $X2=2.37 $Y2=0.465
r65 22 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.715
+ $X2=3.22 $Y2=0.8
r66 21 30 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.465
+ $X2=3.22 $Y2=0.38
r67 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.22 $Y=0.465
+ $X2=3.22 $Y2=0.715
r68 17 33 3.54733 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.105 $Y=1.63
+ $X2=2.91 $Y2=1.63
r69 17 19 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.105 $Y=1.63
+ $X2=3.72 $Y2=1.63
r70 16 28 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.8 $X2=2.38
+ $Y2=0.8
r71 15 38 6.32834 $w=1.68e-07 $l=9.7e-08 $layer=LI1_cond $X=2.91 $Y=0.8
+ $X2=3.007 $Y2=0.8
r72 15 16 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.91 $Y=0.8
+ $X2=2.465 $Y2=0.8
r73 14 28 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=0.715
+ $X2=2.38 $Y2=0.8
r74 14 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.38 $Y=0.715
+ $X2=2.38 $Y2=0.465
r75 4 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=1.63
r76 3 33 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.63
r77 2 48 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.72
r78 2 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.38
r79 1 28 182 $w=1.7e-07 $l=5.57136e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.38 $Y2=0.72
r80 1 24 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.38 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%VGND 1 2 3 4 5 6 19 21 25 29 33 35 39 42 43
+ 45 46 48 49 50 62 71 72 79 85
c110 29 0 2.63538e-20 $X=1.94 $Y=0.38
r111 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r112 80 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r113 79 82 8.91196 $w=5.08e-07 $l=3.8e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.81
+ $Y2=0.38
r114 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r115 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r116 69 72 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=7.13 $Y2=0
r117 69 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r118 68 71 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.29 $Y=0 $X2=7.13
+ $Y2=0
r119 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r120 66 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=0 $X2=4.86
+ $Y2=0
r121 66 68 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.945 $Y=0 $X2=5.29
+ $Y2=0
r122 65 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r123 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r124 62 79 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.81
+ $Y2=0
r125 62 64 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.45 $Y2=0
r126 61 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r127 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r128 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r129 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r130 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r131 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r132 52 75 4.03846 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r133 52 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r134 50 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r135 50 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r136 48 60 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0
+ $X2=2.53 $Y2=0
r137 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.8
+ $Y2=0
r138 47 64 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.45
+ $Y2=0
r139 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.8
+ $Y2=0
r140 45 57 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r141 45 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.94
+ $Y2=0
r142 44 60 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.53 $Y2=0
r143 44 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.94
+ $Y2=0
r144 42 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r145 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r146 41 57 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r147 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r148 37 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.86 $Y=0.085
+ $X2=4.86 $Y2=0
r149 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.86 $Y=0.085
+ $X2=4.86 $Y2=0.38
r150 36 79 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=3.81
+ $Y2=0
r151 35 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.775 $Y=0 $X2=4.86
+ $Y2=0
r152 35 36 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.775 $Y=0
+ $X2=4.065 $Y2=0
r153 31 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r154 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.38
r155 27 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r156 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.38
r157 23 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r158 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r159 19 75 3.10471 $w=2.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.172 $Y2=0
r160 19 21 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.22 $Y2=0.4
r161 6 39 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.725
+ $Y=0.235 $X2=4.86 $Y2=0.38
r162 5 82 91 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.235 $X2=3.98 $Y2=0.38
r163 4 33 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.38
r164 3 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r165 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r166 1 21 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A_861_47# 1 2 8 12 17 18
r32 17 18 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.84 $Y=0.765
+ $X2=5.675 $Y2=0.765
r33 10 15 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=0.8 $X2=4.44
+ $Y2=0.8
r34 10 18 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=4.525 $Y=0.8
+ $X2=5.675 $Y2=0.8
r35 8 15 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0.715 $X2=4.44
+ $Y2=0.8
r36 7 12 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0.465
+ $X2=4.44 $Y2=0.38
r37 7 8 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.44 $Y=0.465 $X2=4.44
+ $Y2=0.715
r38 2 17 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.84 $Y2=0.73
r39 1 15 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.44 $Y2=0.72
r40 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.44 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_4%A_1059_47# 1 2 3 10 16 22 25 28 29
r34 27 29 1.97562 $w=2.43e-07 $l=4.2e-08 $layer=LI1_cond $X=7.1 $Y=0.377
+ $X2=7.142 $Y2=0.377
r35 27 28 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.1 $Y=0.377
+ $X2=6.935 $Y2=0.377
r36 20 29 0.495957 $w=2.55e-07 $l=1.23e-07 $layer=LI1_cond $X=7.142 $Y=0.5
+ $X2=7.142 $Y2=0.377
r37 20 22 10.8465 $w=2.53e-07 $l=2.4e-07 $layer=LI1_cond $X=7.142 $Y=0.5
+ $X2=7.142 $Y2=0.74
r38 19 25 4.70473 $w=1.9e-07 $l=9.44722e-08 $layer=LI1_cond $X=6.345 $Y=0.34
+ $X2=6.26 $Y2=0.36
r39 19 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.345 $Y=0.34
+ $X2=6.935 $Y2=0.34
r40 14 25 1.74598 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.26 $Y=0.465
+ $X2=6.26 $Y2=0.36
r41 14 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.26 $Y=0.465
+ $X2=6.26 $Y2=0.72
r42 10 25 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.36
+ $X2=6.26 $Y2=0.36
r43 10 12 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=6.175 $Y=0.36
+ $X2=5.42 $Y2=0.36
r44 3 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.965
+ $Y=0.235 $X2=7.1 $Y2=0.38
r45 3 22 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=6.965
+ $Y=0.235 $X2=7.1 $Y2=0.74
r46 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.125
+ $Y=0.235 $X2=6.26 $Y2=0.38
r47 2 16 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.125
+ $Y=0.235 $X2=6.26 $Y2=0.72
r48 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.42 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__mux4_2.spice
* Created: Thu Aug 27 14:28:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux4_2.spice.pex"
.subckt sky130_fd_sc_hd__mux4_2  VNB VPB S0 A2 A3 S1 A1 A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* A1	A1
* S1	S1
* A3	A3
* A2	A2
* S0	S0
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_S0_M1025_g N_A_27_47#_M1025_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1013 A_193_47# N_A2_M1013_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.0567 PD=0.802308 PS=0.69 NRD=32.628 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_288_47#_M1004_d N_A_27_47#_M1004_g A_193_47# VNB NSHORT L=0.15 W=0.36
+ AD=0.0711 AS=0.0609231 PD=0.755 PS=0.687692 NRD=18.324 NRS=38.076 M=1 R=2.4
+ SA=75001.1 SB=75001.8 A=0.054 P=1.02 MULT=1
MM1002 A_397_47# N_S0_M1002_g N_A_288_47#_M1004_d VNB NSHORT L=0.15 W=0.36
+ AD=0.0618923 AS=0.0711 PD=0.692308 PS=0.755 NRD=38.964 NRS=19.992 M=1 R=2.4
+ SA=75001.6 SB=75001.2 A=0.054 P=1.02 MULT=1
MM1007 N_VGND_M1007_d N_A3_M1007_g A_397_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0722077 PD=0.81 PS=0.807692 NRD=14.28 NRS=33.396 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1014 N_A_600_345#_M1014_d N_S1_M1014_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0819 PD=1.38 PS=0.81 NRD=1.428 NRS=17.136 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_788_316#_M1019_d N_S1_M1019_g N_A_288_47#_M1019_s VNB NSHORT L=0.15
+ W=0.42 AD=0.05775 AS=0.1092 PD=0.695 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_872_316#_M1012_d N_A_600_345#_M1012_g N_A_788_316#_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.05775 PD=1.36 PS=0.695 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 A_1064_47# N_A1_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0846462 AS=0.1092 PD=0.866923 PS=1.36 NRD=41.868 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1015 N_A_872_316#_M1015_d N_S0_M1015_g A_1064_47# VNB NSHORT L=0.15 W=0.36
+ AD=0.072 AS=0.0725538 PD=0.76 PS=0.743077 NRD=19.992 NRS=48.84 M=1 R=2.4
+ SA=75000.7 SB=75002.2 A=0.054 P=1.02 MULT=1
MM1005 A_1281_47# N_A_27_47#_M1005_g N_A_872_316#_M1015_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.072 PD=0.687692 PS=0.76 NRD=38.076 NRS=19.992 M=1
+ R=2.4 SA=75001.3 SB=75001.7 A=0.054 P=1.02 MULT=1
MM1024 N_VGND_M1024_d N_A0_M1024_g A_1281_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0838037 AS=0.0710769 PD=0.788972 PS=0.802308 NRD=22.848 NRS=32.628 M=1
+ R=2.8 SA=75001.5 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1024_d N_A_788_316#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.129696 AS=0.08775 PD=1.22103 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_788_316#_M1010_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.221 AS=0.08775 PD=1.98 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75001.8
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1016 N_VPWR_M1016_d N_S0_M1016_g N_A_27_47#_M1016_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1000 A_193_369# N_A2_M1000_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.115623 AS=0.0864 PD=1.16528 PS=0.91 NRD=38.6711 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1023 N_A_288_47#_M1023_d N_S0_M1023_g A_193_369# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.0758774 PD=0.69 PS=0.764717 NRD=0 NRS=58.9227 M=1 R=2.8
+ SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1017 A_372_413# N_A_27_47#_M1017_g N_A_288_47#_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.130358 AS=0.0567 PD=1.05396 PS=0.69 NRD=119.776 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A3_M1003_g A_372_413# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.198642 PD=0.91 PS=1.60604 NRD=0 NRS=78.603 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1026 N_A_600_345#_M1026_d N_S1_M1026_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_A_788_316#_M1020_d N_A_600_345#_M1020_g N_A_288_47#_M1020_s VPB PHIGHVT
+ L=0.15 W=0.54 AD=0.0729 AS=0.1404 PD=0.81 PS=1.6 NRD=0 NRS=0 M=1 R=3.6
+ SA=75000.2 SB=75000.6 A=0.081 P=1.38 MULT=1
MM1008 N_A_872_316#_M1008_d N_S1_M1008_g N_A_788_316#_M1020_d VPB PHIGHVT L=0.15
+ W=0.54 AD=0.1404 AS=0.0729 PD=1.6 PS=0.81 NRD=0 NRS=0 M=1 R=3.6 SA=75000.6
+ SB=75000.2 A=0.081 P=1.38 MULT=1
MM1001 A_1060_369# N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.16634 AS=0.1664 PD=1.40679 PS=1.8 NRD=63.0597 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1022 N_A_872_316#_M1022_d N_A_27_47#_M1022_g A_1060_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.10916 PD=0.69 PS=0.923208 NRD=0 NRS=96.0966 M=1 R=2.8
+ SA=75000.9 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1018 A_1279_413# N_S0_M1018_g N_A_872_316#_M1022_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0834849 AS=0.0567 PD=0.788491 PS=0.69 NRD=67.4331 NRS=0 M=1 R=2.8
+ SA=75001.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A0_M1021_g A_1279_413# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.120195 AS=0.127215 PD=1.04195 PS=1.20151 NRD=18.4589 NRS=44.2462 M=1
+ R=4.26667 SA=75001.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1021_d N_A_788_316#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.187805 AS=0.135 PD=1.62805 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_788_316#_M1011_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.34 AS=0.135 PD=2.68 PS=1.27 NRD=14.775 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.8993 P=20.53
*
.include "sky130_fd_sc_hd__mux4_2.spice.SKY130_FD_SC_HD__MUX4_2.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a311o_1.spice
* Created: Tue Sep  1 18:54:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a311o_1.pex.spice"
.subckt sky130_fd_sc_hd__a311o_1  VNB VPB A3 A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_75_199#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.112125 AS=0.169 PD=0.995 PS=1.82 NRD=12.912 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1009 A_208_47# N_A3_M1009_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.125125 AS=0.112125 PD=1.035 PS=0.995 NRD=25.38 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1005 A_315_47# N_A2_M1005_g A_208_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.125125 PD=1.17 PS=1.035 NRD=37.836 NRS=25.38 M=1 R=4.33333 SA=75001.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1008 N_A_75_199#_M1008_d N_A1_M1008_g A_315_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.169 PD=0.975 PS=1.17 NRD=4.608 NRS=37.836 M=1 R=4.33333
+ SA=75001.9 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_B1_M1001_g N_A_75_199#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.134875 AS=0.105625 PD=1.065 PS=0.975 NRD=12.912 NRS=3.684 M=1 R=4.33333
+ SA=75002.4 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_A_75_199#_M1010_d N_C1_M1010_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.134875 PD=1.82 PS=1.065 NRD=0 NRS=11.988 M=1 R=4.33333
+ SA=75002.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_75_199#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1425 AS=0.285 PD=1.285 PS=2.57 NRD=0 NRS=3.9203 M=1 R=6.66667 SA=75000.2
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1006 N_A_201_297#_M1006_d N_A3_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.1425 PD=1.33 PS=1.285 NRD=6.8753 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_201_297#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.305 AS=0.165 PD=1.61 PS=1.33 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75001.1
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1007 N_A_201_297#_M1007_d N_A1_M1007_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1625 AS=0.305 PD=1.325 PS=1.61 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1003 A_544_297# N_B1_M1003_g N_A_201_297#_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.2075 AS=0.1625 PD=1.415 PS=1.325 NRD=30.0228 NRS=3.9203 M=1 R=6.66667
+ SA=75002.4 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1000 N_A_75_199#_M1000_d N_C1_M1000_g A_544_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.2075 PD=2.52 PS=1.415 NRD=0 NRS=30.0228 M=1 R=6.66667 SA=75002.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_58 VPB 0 1.12853e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a311o_1.pxi.spice"
*
.ends
*
*

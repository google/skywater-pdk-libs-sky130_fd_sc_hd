* File: sky130_fd_sc_hd__mux4_4.pxi.spice
* Created: Thu Aug 27 14:28:30 2020
* 
x_PM_SKY130_FD_SC_HD__MUX4_4%S0 N_S0_M1029_g N_S0_M1021_g N_S0_c_190_n
+ N_S0_M1025_g N_S0_c_191_n N_S0_M1026_g N_S0_M1010_g N_S0_c_194_n N_S0_c_195_n
+ N_S0_M1016_g S0 S0 N_S0_c_208_n N_S0_c_209_n N_S0_c_210_n N_S0_c_211_n
+ N_S0_c_197_n N_S0_c_213_n N_S0_c_214_n N_S0_c_198_n N_S0_c_199_n
+ PM_SKY130_FD_SC_HD__MUX4_4%S0
x_PM_SKY130_FD_SC_HD__MUX4_4%A2 N_A2_M1018_g N_A2_M1001_g A2 A2 N_A2_c_393_n
+ N_A2_c_394_n PM_SKY130_FD_SC_HD__MUX4_4%A2
x_PM_SKY130_FD_SC_HD__MUX4_4%A_27_47# N_A_27_47#_M1029_s N_A_27_47#_M1021_s
+ N_A_27_47#_c_447_n N_A_27_47#_M1006_g N_A_27_47#_M1017_g N_A_27_47#_M1023_g
+ N_A_27_47#_c_448_n N_A_27_47#_M1028_g N_A_27_47#_c_671_p N_A_27_47#_c_606_p
+ N_A_27_47#_c_449_n N_A_27_47#_c_460_n N_A_27_47#_c_461_n N_A_27_47#_c_450_n
+ N_A_27_47#_c_451_n N_A_27_47#_c_452_n N_A_27_47#_c_453_n N_A_27_47#_c_462_n
+ N_A_27_47#_c_463_n N_A_27_47#_c_464_n N_A_27_47#_c_465_n N_A_27_47#_c_466_n
+ N_A_27_47#_c_467_n N_A_27_47#_c_454_n N_A_27_47#_c_455_n N_A_27_47#_c_456_n
+ PM_SKY130_FD_SC_HD__MUX4_4%A_27_47#
x_PM_SKY130_FD_SC_HD__MUX4_4%A3 N_A3_M1030_g N_A3_c_688_n N_A3_c_694_n
+ N_A3_M1002_g N_A3_c_695_n A3 A3 N_A3_c_691_n N_A3_c_692_n
+ PM_SKY130_FD_SC_HD__MUX4_4%A3
x_PM_SKY130_FD_SC_HD__MUX4_4%S1 N_S1_c_747_n N_S1_M1027_g N_S1_c_749_n
+ N_S1_M1009_g N_S1_c_754_n N_S1_c_755_n N_S1_c_750_n N_S1_c_751_n N_S1_M1012_g
+ N_S1_M1013_g S1 S1 PM_SKY130_FD_SC_HD__MUX4_4%S1
x_PM_SKY130_FD_SC_HD__MUX4_4%A_601_345# N_A_601_345#_M1009_d
+ N_A_601_345#_M1027_d N_A_601_345#_M1019_g N_A_601_345#_c_833_n
+ N_A_601_345#_M1007_g N_A_601_345#_c_835_n N_A_601_345#_c_836_n
+ N_A_601_345#_c_837_n N_A_601_345#_c_838_n N_A_601_345#_c_839_n
+ PM_SKY130_FD_SC_HD__MUX4_4%A_601_345#
x_PM_SKY130_FD_SC_HD__MUX4_4%A1 N_A1_M1000_g N_A1_M1024_g A1 A1 N_A1_c_904_n
+ PM_SKY130_FD_SC_HD__MUX4_4%A1
x_PM_SKY130_FD_SC_HD__MUX4_4%A0 N_A0_M1020_g N_A0_M1022_g N_A0_c_943_n
+ N_A0_c_944_n A0 A0 PM_SKY130_FD_SC_HD__MUX4_4%A0
x_PM_SKY130_FD_SC_HD__MUX4_4%A_789_316# N_A_789_316#_M1012_d
+ N_A_789_316#_M1019_d N_A_789_316#_c_991_n N_A_789_316#_M1003_g
+ N_A_789_316#_M1004_g N_A_789_316#_c_992_n N_A_789_316#_M1005_g
+ N_A_789_316#_M1008_g N_A_789_316#_c_993_n N_A_789_316#_c_994_n
+ N_A_789_316#_c_995_n N_A_789_316#_M1011_g N_A_789_316#_M1014_g
+ N_A_789_316#_c_996_n N_A_789_316#_M1031_g N_A_789_316#_M1015_g
+ N_A_789_316#_c_997_n N_A_789_316#_c_998_n N_A_789_316#_c_1008_n
+ N_A_789_316#_c_1009_n N_A_789_316#_c_1010_n N_A_789_316#_c_1011_n
+ N_A_789_316#_c_1012_n N_A_789_316#_c_999_n N_A_789_316#_c_1014_n
+ N_A_789_316#_c_1015_n N_A_789_316#_c_1016_n N_A_789_316#_c_1030_n
+ N_A_789_316#_c_1031_n PM_SKY130_FD_SC_HD__MUX4_4%A_789_316#
x_PM_SKY130_FD_SC_HD__MUX4_4%VPWR N_VPWR_M1021_d N_VPWR_M1002_d N_VPWR_M1000_s
+ N_VPWR_M1022_d N_VPWR_M1008_d N_VPWR_M1015_d N_VPWR_c_1178_n N_VPWR_c_1179_n
+ N_VPWR_c_1180_n N_VPWR_c_1181_n N_VPWR_c_1182_n N_VPWR_c_1183_n
+ N_VPWR_c_1184_n N_VPWR_c_1185_n N_VPWR_c_1186_n N_VPWR_c_1187_n
+ N_VPWR_c_1188_n VPWR N_VPWR_c_1189_n N_VPWR_c_1190_n N_VPWR_c_1191_n
+ N_VPWR_c_1192_n N_VPWR_c_1193_n N_VPWR_c_1194_n N_VPWR_c_1195_n
+ N_VPWR_c_1177_n PM_SKY130_FD_SC_HD__MUX4_4%VPWR
x_PM_SKY130_FD_SC_HD__MUX4_4%A_288_47# N_A_288_47#_M1006_d N_A_288_47#_M1012_s
+ N_A_288_47#_M1025_d N_A_288_47#_M1019_s N_A_288_47#_c_1337_n
+ N_A_288_47#_c_1338_n N_A_288_47#_c_1325_n N_A_288_47#_c_1329_n
+ N_A_288_47#_c_1341_n N_A_288_47#_c_1330_n N_A_288_47#_c_1331_n
+ N_A_288_47#_c_1326_n N_A_288_47#_c_1327_n N_A_288_47#_c_1328_n
+ N_A_288_47#_c_1334_n N_A_288_47#_c_1374_n N_A_288_47#_c_1335_n
+ PM_SKY130_FD_SC_HD__MUX4_4%A_288_47#
x_PM_SKY130_FD_SC_HD__MUX4_4%A_873_316# N_A_873_316#_M1007_d
+ N_A_873_316#_M1010_d N_A_873_316#_M1013_d N_A_873_316#_M1023_d
+ N_A_873_316#_c_1463_n N_A_873_316#_c_1466_n N_A_873_316#_c_1464_n
+ N_A_873_316#_c_1468_n N_A_873_316#_c_1540_p N_A_873_316#_c_1475_n
+ N_A_873_316#_c_1513_n N_A_873_316#_c_1476_n N_A_873_316#_c_1514_n
+ N_A_873_316#_c_1469_n PM_SKY130_FD_SC_HD__MUX4_4%A_873_316#
x_PM_SKY130_FD_SC_HD__MUX4_4%X N_X_M1003_s N_X_M1011_s N_X_M1004_s N_X_M1014_s
+ N_X_c_1565_n N_X_c_1561_n N_X_c_1574_n N_X_c_1577_n N_X_c_1580_n N_X_c_1582_n
+ N_X_c_1563_n N_X_c_1590_n X X X X X X PM_SKY130_FD_SC_HD__MUX4_4%X
x_PM_SKY130_FD_SC_HD__MUX4_4%VGND N_VGND_M1029_d N_VGND_M1030_d N_VGND_M1024_s
+ N_VGND_M1020_d N_VGND_M1005_d N_VGND_M1031_d N_VGND_c_1619_n N_VGND_c_1620_n
+ N_VGND_c_1621_n N_VGND_c_1622_n N_VGND_c_1623_n N_VGND_c_1624_n
+ N_VGND_c_1625_n VGND N_VGND_c_1626_n N_VGND_c_1627_n N_VGND_c_1628_n
+ N_VGND_c_1629_n N_VGND_c_1630_n N_VGND_c_1631_n N_VGND_c_1632_n
+ N_VGND_c_1633_n N_VGND_c_1634_n N_VGND_c_1635_n N_VGND_c_1636_n
+ N_VGND_c_1637_n PM_SKY130_FD_SC_HD__MUX4_4%VGND
cc_1 VNB N_S0_M1029_g 0.0352159f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_S0_c_190_n 0.00810316f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.615
cc_3 VNB N_S0_c_191_n 0.0148947f $X=-0.19 $Y=-0.24 $X2=1.84 $Y2=1.32
cc_4 VNB N_S0_M1026_g 0.04359f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.415
cc_5 VNB N_S0_M1010_g 0.0457627f $X=-0.19 $Y=-0.24 $X2=5.785 $Y2=0.415
cc_6 VNB N_S0_c_194_n 0.0107197f $X=-0.19 $Y=-0.24 $X2=6.25 $Y2=1.32
cc_7 VNB N_S0_c_195_n 0.00201541f $X=-0.19 $Y=-0.24 $X2=5.86 $Y2=1.32
cc_8 VNB S0 0.00247953f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_9 VNB N_S0_c_197_n 0.00205509f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.53
cc_10 VNB N_S0_c_198_n 0.0432497f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_11 VNB N_S0_c_199_n 0.0110759f $X=-0.19 $Y=-0.24 $X2=6.385 $Y2=1.32
cc_12 VNB N_A2_M1001_g 0.0128595f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_13 VNB A2 0.00268806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB A2 0.0042355f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.615
cc_15 VNB N_A2_c_393_n 0.0275156f $X=-0.19 $Y=-0.24 $X2=1.445 $Y2=1.32
cc_16 VNB N_A2_c_394_n 0.0166422f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.415
cc_17 VNB N_A_27_47#_c_447_n 0.0180404f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_18 VNB N_A_27_47#_c_448_n 0.0180623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_449_n 0.00401519f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_20 VNB N_A_27_47#_c_450_n 0.0100323f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_21 VNB N_A_27_47#_c_451_n 0.0313728f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.53
cc_22 VNB N_A_27_47#_c_452_n 0.0030285f $X=-0.19 $Y=-0.24 $X2=6.215 $Y2=1.53
cc_23 VNB N_A_27_47#_c_453_n 0.00540154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_454_n 0.00906583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_455_n 0.032928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_456_n 0.00415242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A3_c_688_n 0.0112092f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_28 VNB A3 0.00653171f $X=-0.19 $Y=-0.24 $X2=1.84 $Y2=1.32
cc_29 VNB A3 0.00177632f $X=-0.19 $Y=-0.24 $X2=1.445 $Y2=1.32
cc_30 VNB N_A3_c_691_n 0.0241632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A3_c_692_n 0.0172648f $X=-0.19 $Y=-0.24 $X2=5.785 $Y2=0.415
cc_32 VNB N_S1_c_747_n 0.0288831f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_33 VNB N_S1_M1027_g 0.00924061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_S1_c_749_n 0.0184815f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_35 VNB N_S1_c_750_n 0.0513215f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=2.275
cc_36 VNB N_S1_c_751_n 0.0179541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB S1 0.00677138f $X=-0.19 $Y=-0.24 $X2=5.785 $Y2=1.245
cc_38 VNB N_A_601_345#_c_833_n 0.0321009f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=2.275
cc_39 VNB N_A_601_345#_M1007_g 0.0381718f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=1.245
cc_40 VNB N_A_601_345#_c_835_n 0.0234246f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.415
cc_41 VNB N_A_601_345#_c_836_n 0.00740591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_601_345#_c_837_n 0.00626684f $X=-0.19 $Y=-0.24 $X2=5.785 $Y2=0.415
cc_43 VNB N_A_601_345#_c_838_n 0.00114392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_601_345#_c_839_n 0.00367345f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_45 VNB N_A1_M1024_g 0.0386874f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_46 VNB A1 0.0121957f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.615
cc_47 VNB N_A1_c_904_n 0.0312386f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.415
cc_48 VNB N_A0_M1020_g 0.0291922f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_49 VNB N_A0_c_943_n 0.0139105f $X=-0.19 $Y=-0.24 $X2=1.37 $Y2=1.615
cc_50 VNB N_A0_c_944_n 0.0257079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB A0 0.00260222f $X=-0.19 $Y=-0.24 $X2=1.84 $Y2=1.32
cc_52 VNB N_A_789_316#_c_991_n 0.0166938f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_53 VNB N_A_789_316#_c_992_n 0.016273f $X=-0.19 $Y=-0.24 $X2=1.445 $Y2=1.32
cc_54 VNB N_A_789_316#_c_993_n 0.0165671f $X=-0.19 $Y=-0.24 $X2=5.785 $Y2=0.415
cc_55 VNB N_A_789_316#_c_994_n 0.0259285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_789_316#_c_995_n 0.0164536f $X=-0.19 $Y=-0.24 $X2=6.25 $Y2=1.32
cc_57 VNB N_A_789_316#_c_996_n 0.0215005f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_58 VNB N_A_789_316#_c_997_n 0.0384602f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_59 VNB N_A_789_316#_c_998_n 0.00865735f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.53
cc_60 VNB N_A_789_316#_c_999_n 0.00267682f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.45
cc_61 VNB N_VPWR_c_1177_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_288_47#_c_1325_n 0.0043778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_288_47#_c_1326_n 0.00668781f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.53
cc_64 VNB N_A_288_47#_c_1327_n 0.00364533f $X=-0.19 $Y=-0.24 $X2=6.07 $Y2=1.53
cc_65 VNB N_A_288_47#_c_1328_n 7.8042e-19 $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_66 VNB N_A_873_316#_c_1463_n 0.0132662f $X=-0.19 $Y=-0.24 $X2=1.445 $Y2=1.32
cc_67 VNB N_A_873_316#_c_1464_n 0.0123599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_X_c_1561_n 0.00108687f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB X 8.78104e-19 $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.53
cc_70 VNB N_VGND_c_1619_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=5.785 $Y2=0.415
cc_71 VNB N_VGND_c_1620_n 0.00290102f $X=-0.19 $Y=-0.24 $X2=6.325 $Y2=1.575
cc_72 VNB N_VGND_c_1621_n 0.010332f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_73 VNB N_VGND_c_1622_n 0.00229342f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.53
cc_74 VNB N_VGND_c_1623_n 0.00282952f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_75 VNB N_VGND_c_1624_n 0.01004f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_76 VNB N_VGND_c_1625_n 0.0329454f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.53
cc_77 VNB N_VGND_c_1626_n 0.0150758f $X=-0.19 $Y=-0.24 $X2=6.215 $Y2=1.53
cc_78 VNB N_VGND_c_1627_n 0.0419673f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_79 VNB N_VGND_c_1628_n 0.0541513f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.45
cc_80 VNB N_VGND_c_1629_n 0.0497635f $X=-0.19 $Y=-0.24 $X2=6.385 $Y2=1.41
cc_81 VNB N_VGND_c_1630_n 0.0171682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1631_n 0.0170713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1632_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1633_n 0.00516502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1634_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1635_n 0.00356594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1636_n 0.00356594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1637_n 0.438322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VPB N_S0_M1021_g 0.0433759f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_90 VPB N_S0_c_190_n 0.0227389f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=1.615
cc_91 VPB N_S0_M1025_g 0.0331485f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=2.275
cc_92 VPB N_S0_c_191_n 0.0167376f $X=-0.19 $Y=1.305 $X2=1.84 $Y2=1.32
cc_93 VPB N_S0_c_194_n 0.01241f $X=-0.19 $Y=1.305 $X2=6.25 $Y2=1.32
cc_94 VPB N_S0_c_195_n 0.0045458f $X=-0.19 $Y=1.305 $X2=5.86 $Y2=1.32
cc_95 VPB N_S0_M1016_g 0.0376059f $X=-0.19 $Y=1.305 $X2=6.325 $Y2=2.275
cc_96 VPB S0 0.0145413f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_97 VPB N_S0_c_208_n 0.00666793f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.53
cc_98 VPB N_S0_c_209_n 0.0141389f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.53
cc_99 VPB N_S0_c_210_n 0.0435336f $X=-0.19 $Y=1.305 $X2=6.07 $Y2=1.53
cc_100 VPB N_S0_c_211_n 0.00423102f $X=-0.19 $Y=1.305 $X2=1.3 $Y2=1.53
cc_101 VPB N_S0_c_197_n 0.00302522f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.53
cc_102 VPB N_S0_c_213_n 0.00246888f $X=-0.19 $Y=1.305 $X2=6.215 $Y2=1.53
cc_103 VPB N_S0_c_214_n 0.00362396f $X=-0.19 $Y=1.305 $X2=6.215 $Y2=1.53
cc_104 VPB N_S0_c_198_n 0.0110719f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_105 VPB N_S0_c_199_n 0.0215929f $X=-0.19 $Y=1.305 $X2=6.385 $Y2=1.32
cc_106 VPB N_A2_M1001_g 0.0369519f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_107 VPB N_A_27_47#_M1017_g 0.02251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_47#_M1023_g 0.0226804f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.415
cc_109 VPB N_A_27_47#_c_449_n 0.00368949f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_110 VPB N_A_27_47#_c_460_n 0.00646631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_461_n 0.00677133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_27_47#_c_462_n 0.0085993f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.32
cc_113 VPB N_A_27_47#_c_463_n 0.0027247f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.45
cc_114 VPB N_A_27_47#_c_464_n 0.00188091f $X=-0.19 $Y=1.305 $X2=6.385 $Y2=1.41
cc_115 VPB N_A_27_47#_c_465_n 0.0277359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_466_n 0.00526335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_467_n 0.0275765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_c_454_n 0.00474478f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_456_n 0.00201397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A3_c_688_n 0.0117778f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_121 VPB N_A3_c_694_n 0.0237103f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_122 VPB N_A3_c_695_n 0.0181615f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=2.275
cc_123 VPB A3 9.23002e-19 $X=-0.19 $Y=1.305 $X2=1.445 $Y2=1.32
cc_124 VPB N_S1_M1027_g 0.0332464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_S1_c_754_n 0.096695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_S1_c_755_n 0.00958866f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=1.615
cc_127 VPB N_S1_M1013_g 0.0364991f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.415
cc_128 VPB S1 0.00178367f $X=-0.19 $Y=1.305 $X2=5.785 $Y2=1.245
cc_129 VPB N_A_601_345#_M1019_g 0.0238152f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=1.615
cc_130 VPB N_A_601_345#_c_835_n 0.0207466f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.415
cc_131 VPB N_A_601_345#_c_836_n 0.00224568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_601_345#_c_838_n 0.0132075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A1_M1000_g 0.0458456f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_134 VPB A1 0.0035535f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=1.615
cc_135 VPB N_A1_c_904_n 0.0156887f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.415
cc_136 VPB N_A0_M1022_g 0.0377501f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_137 VPB N_A0_c_943_n 0.00286793f $X=-0.19 $Y=1.305 $X2=1.37 $Y2=1.615
cc_138 VPB N_A0_c_944_n 0.00429793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_789_316#_M1004_g 0.0185811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_789_316#_M1008_g 0.0187212f $X=-0.19 $Y=1.305 $X2=5.785 $Y2=1.245
cc_141 VPB N_A_789_316#_c_993_n 0.00594691f $X=-0.19 $Y=1.305 $X2=5.785
+ $Y2=0.415
cc_142 VPB N_A_789_316#_c_994_n 0.00449786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_789_316#_M1014_g 0.0191153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_789_316#_M1015_g 0.025294f $X=-0.19 $Y=1.305 $X2=6.07 $Y2=1.53
cc_145 VPB N_A_789_316#_c_997_n 0.0048883f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.53
cc_146 VPB N_A_789_316#_c_998_n 0.00438187f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.53
cc_147 VPB N_A_789_316#_c_1008_n 0.00187498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_789_316#_c_1009_n 0.00313433f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.16
cc_149 VPB N_A_789_316#_c_1010_n 0.00173284f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.16
cc_150 VPB N_A_789_316#_c_1011_n 0.00185715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_789_316#_c_1012_n 0.00258066f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_152 VPB N_A_789_316#_c_999_n 3.66738e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.45
cc_153 VPB N_A_789_316#_c_1014_n 0.00232217f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_789_316#_c_1015_n 0.00114749f $X=-0.19 $Y=1.305 $X2=6.385
+ $Y2=1.41
cc_155 VPB N_A_789_316#_c_1016_n 0.00329434f $X=-0.19 $Y=1.305 $X2=6.385
+ $Y2=1.575
cc_156 VPB N_VPWR_c_1178_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=5.785 $Y2=0.415
cc_157 VPB N_VPWR_c_1179_n 0.00835502f $X=-0.19 $Y=1.305 $X2=6.325 $Y2=1.575
cc_158 VPB N_VPWR_c_1180_n 0.013457f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_159 VPB N_VPWR_c_1181_n 0.00468459f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.53
cc_160 VPB N_VPWR_c_1182_n 0.00226048f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.53
cc_161 VPB N_VPWR_c_1183_n 0.0100141f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.53
cc_162 VPB N_VPWR_c_1184_n 0.0422332f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.53
cc_163 VPB N_VPWR_c_1185_n 0.0491497f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_164 VPB N_VPWR_c_1186_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_165 VPB N_VPWR_c_1187_n 0.0519215f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1188_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_167 VPB N_VPWR_c_1189_n 0.0150788f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.45
cc_168 VPB N_VPWR_c_1190_n 0.0543338f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.53
cc_169 VPB N_VPWR_c_1191_n 0.0200388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1192_n 0.0170713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1193_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1194_n 0.0066101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1195_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1177_n 0.0497858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_288_47#_c_1329_n 0.00997171f $X=-0.19 $Y=1.305 $X2=5.86 $Y2=1.32
cc_176 VPB N_A_288_47#_c_1330_n 0.00983477f $X=-0.19 $Y=1.305 $X2=6.325
+ $Y2=2.275
cc_177 VPB N_A_288_47#_c_1331_n 4.38222e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_288_47#_c_1326_n 0.00277353f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.53
cc_179 VPB N_A_288_47#_c_1327_n 0.00136736f $X=-0.19 $Y=1.305 $X2=6.07 $Y2=1.53
cc_180 VPB N_A_288_47#_c_1334_n 3.67896e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_288_47#_c_1335_n 0.00406359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_873_316#_c_1463_n 0.00645389f $X=-0.19 $Y=1.305 $X2=1.445
+ $Y2=1.32
cc_183 VPB N_A_873_316#_c_1466_n 0.0111242f $X=-0.19 $Y=1.305 $X2=1.915
+ $Y2=1.245
cc_184 VPB N_A_873_316#_c_1464_n 0.00454907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_873_316#_c_1468_n 0.00168598f $X=-0.19 $Y=1.305 $X2=5.785
+ $Y2=0.415
cc_186 VPB N_A_873_316#_c_1469_n 0.00105233f $X=-0.19 $Y=1.305 $X2=6.07 $Y2=1.53
cc_187 VPB N_X_c_1563_n 0.0011999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB X 0.0012809f $X=-0.19 $Y=1.305 $X2=1.3 $Y2=1.53
cc_189 N_S0_c_190_n N_A2_M1001_g 0.0230379f $X=1.37 $Y=1.615 $X2=0 $Y2=0
cc_190 N_S0_M1025_g N_A2_M1001_g 0.0383473f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_191 N_S0_c_208_n N_A2_M1001_g 0.00594683f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_192 N_S0_c_211_n N_A2_M1001_g 9.9583e-19 $X=1.3 $Y=1.53 $X2=0 $Y2=0
cc_193 N_S0_c_197_n N_A2_M1001_g 0.00193624f $X=1.155 $Y=1.53 $X2=0 $Y2=0
cc_194 N_S0_c_198_n N_A2_M1001_g 0.0528485f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_195 N_S0_M1029_g A2 3.057e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_196 N_S0_c_190_n A2 0.00133318f $X=1.37 $Y=1.615 $X2=0 $Y2=0
cc_197 N_S0_c_208_n A2 0.00572305f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_198 N_S0_c_211_n A2 0.0054611f $X=1.3 $Y=1.53 $X2=0 $Y2=0
cc_199 N_S0_c_197_n A2 0.00784362f $X=1.155 $Y=1.53 $X2=0 $Y2=0
cc_200 N_S0_M1029_g N_A2_c_393_n 0.0165033f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_201 N_S0_c_208_n N_A2_c_393_n 0.00149712f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_202 N_S0_c_211_n N_A2_c_393_n 0.00118428f $X=1.3 $Y=1.53 $X2=0 $Y2=0
cc_203 N_S0_c_197_n N_A2_c_393_n 9.40361e-19 $X=1.155 $Y=1.53 $X2=0 $Y2=0
cc_204 N_S0_M1029_g N_A2_c_394_n 0.0142481f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_205 N_S0_M1026_g N_A_27_47#_c_447_n 0.0177394f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_206 N_S0_M1025_g N_A_27_47#_M1017_g 0.0201836f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_207 N_S0_M1016_g N_A_27_47#_M1023_g 0.0187022f $X=6.325 $Y=2.275 $X2=0 $Y2=0
cc_208 N_S0_M1010_g N_A_27_47#_c_448_n 0.0184915f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_209 N_S0_M1029_g N_A_27_47#_c_449_n 0.00862509f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_210 N_S0_M1021_g N_A_27_47#_c_449_n 0.00911908f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_211 S0 N_A_27_47#_c_449_n 0.0525762f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_212 N_S0_c_208_n N_A_27_47#_c_449_n 0.0235359f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_213 N_S0_c_209_n N_A_27_47#_c_449_n 0.00268638f $X=0.38 $Y=1.53 $X2=0 $Y2=0
cc_214 N_S0_c_211_n N_A_27_47#_c_449_n 0.00228258f $X=1.3 $Y=1.53 $X2=0 $Y2=0
cc_215 N_S0_c_197_n N_A_27_47#_c_449_n 0.0102687f $X=1.155 $Y=1.53 $X2=0 $Y2=0
cc_216 N_S0_c_198_n N_A_27_47#_c_449_n 0.00796989f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_217 N_S0_c_190_n N_A_27_47#_c_460_n 8.45937e-19 $X=1.37 $Y=1.615 $X2=0 $Y2=0
cc_218 N_S0_M1025_g N_A_27_47#_c_460_n 0.01066f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_219 N_S0_c_191_n N_A_27_47#_c_460_n 0.00281568f $X=1.84 $Y=1.32 $X2=0 $Y2=0
cc_220 N_S0_c_208_n N_A_27_47#_c_460_n 0.014054f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_221 N_S0_c_210_n N_A_27_47#_c_460_n 0.00431952f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_222 N_S0_c_211_n N_A_27_47#_c_460_n 0.00821549f $X=1.3 $Y=1.53 $X2=0 $Y2=0
cc_223 N_S0_c_197_n N_A_27_47#_c_460_n 0.024961f $X=1.155 $Y=1.53 $X2=0 $Y2=0
cc_224 N_S0_M1021_g N_A_27_47#_c_461_n 0.0184821f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_225 S0 N_A_27_47#_c_461_n 0.0148027f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_226 N_S0_c_208_n N_A_27_47#_c_461_n 0.00395767f $X=1.01 $Y=1.53 $X2=0 $Y2=0
cc_227 N_S0_c_209_n N_A_27_47#_c_461_n 0.0041868f $X=0.38 $Y=1.53 $X2=0 $Y2=0
cc_228 N_S0_c_198_n N_A_27_47#_c_461_n 0.00200422f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_229 N_S0_M1029_g N_A_27_47#_c_450_n 0.0142655f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_230 S0 N_A_27_47#_c_450_n 0.0147211f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_231 N_S0_c_209_n N_A_27_47#_c_450_n 0.00268817f $X=0.38 $Y=1.53 $X2=0 $Y2=0
cc_232 N_S0_c_198_n N_A_27_47#_c_450_n 0.0041992f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_233 N_S0_c_190_n N_A_27_47#_c_451_n 0.0234927f $X=1.37 $Y=1.615 $X2=0 $Y2=0
cc_234 N_S0_M1026_g N_A_27_47#_c_451_n 0.019381f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_235 N_S0_c_210_n N_A_27_47#_c_451_n 2.32311e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_236 N_S0_c_197_n N_A_27_47#_c_451_n 7.38135e-19 $X=1.155 $Y=1.53 $X2=0 $Y2=0
cc_237 N_S0_c_190_n N_A_27_47#_c_452_n 0.00107346f $X=1.37 $Y=1.615 $X2=0 $Y2=0
cc_238 N_S0_c_191_n N_A_27_47#_c_452_n 4.97671e-19 $X=1.84 $Y=1.32 $X2=0 $Y2=0
cc_239 N_S0_M1026_g N_A_27_47#_c_452_n 0.00191472f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_240 N_S0_c_210_n N_A_27_47#_c_452_n 0.00565103f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_241 N_S0_M1010_g N_A_27_47#_c_453_n 0.0126611f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_242 N_S0_c_194_n N_A_27_47#_c_453_n 0.00529488f $X=6.25 $Y=1.32 $X2=0 $Y2=0
cc_243 N_S0_c_210_n N_A_27_47#_c_453_n 0.00494576f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_244 N_S0_c_213_n N_A_27_47#_c_453_n 0.00305817f $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_245 N_S0_c_214_n N_A_27_47#_c_453_n 0.00943055f $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_246 N_S0_c_210_n N_A_27_47#_c_462_n 0.301644f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_247 N_S0_M1025_g N_A_27_47#_c_463_n 0.0010293f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_248 N_S0_c_210_n N_A_27_47#_c_463_n 0.0259379f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_249 N_S0_c_210_n N_A_27_47#_c_464_n 0.0255939f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_250 N_S0_c_190_n N_A_27_47#_c_465_n 0.0163856f $X=1.37 $Y=1.615 $X2=0 $Y2=0
cc_251 N_S0_c_191_n N_A_27_47#_c_465_n 0.0206876f $X=1.84 $Y=1.32 $X2=0 $Y2=0
cc_252 N_S0_c_210_n N_A_27_47#_c_465_n 3.65383e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_253 N_S0_M1025_g N_A_27_47#_c_466_n 0.00425396f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_254 N_S0_c_191_n N_A_27_47#_c_466_n 0.00300332f $X=1.84 $Y=1.32 $X2=0 $Y2=0
cc_255 N_S0_c_210_n N_A_27_47#_c_466_n 0.0103825f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_256 N_S0_c_211_n N_A_27_47#_c_466_n 0.00138334f $X=1.3 $Y=1.53 $X2=0 $Y2=0
cc_257 N_S0_c_195_n N_A_27_47#_c_467_n 0.0215228f $X=5.86 $Y=1.32 $X2=0 $Y2=0
cc_258 N_S0_M1016_g N_A_27_47#_c_467_n 0.0168768f $X=6.325 $Y=2.275 $X2=0 $Y2=0
cc_259 N_S0_c_210_n N_A_27_47#_c_467_n 5.96199e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_260 N_S0_c_213_n N_A_27_47#_c_467_n 6.73758e-19 $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_261 N_S0_c_214_n N_A_27_47#_c_467_n 2.32403e-19 $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_262 N_S0_M1010_g N_A_27_47#_c_454_n 0.00816658f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_263 N_S0_c_194_n N_A_27_47#_c_454_n 0.0061637f $X=6.25 $Y=1.32 $X2=0 $Y2=0
cc_264 N_S0_c_195_n N_A_27_47#_c_454_n 0.00451376f $X=5.86 $Y=1.32 $X2=0 $Y2=0
cc_265 N_S0_M1016_g N_A_27_47#_c_454_n 0.00197425f $X=6.325 $Y=2.275 $X2=0 $Y2=0
cc_266 N_S0_c_210_n N_A_27_47#_c_454_n 0.0165427f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_267 N_S0_c_213_n N_A_27_47#_c_454_n 0.00278449f $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_268 N_S0_c_214_n N_A_27_47#_c_454_n 0.028941f $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_269 N_S0_c_199_n N_A_27_47#_c_454_n 0.00105544f $X=6.385 $Y=1.32 $X2=0 $Y2=0
cc_270 N_S0_M1010_g N_A_27_47#_c_455_n 0.0213388f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_271 N_S0_c_194_n N_A_27_47#_c_455_n 0.0224415f $X=6.25 $Y=1.32 $X2=0 $Y2=0
cc_272 N_S0_c_214_n N_A_27_47#_c_455_n 0.0014931f $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_273 N_S0_c_190_n N_A_27_47#_c_456_n 0.00407077f $X=1.37 $Y=1.615 $X2=0 $Y2=0
cc_274 N_S0_c_191_n N_A_27_47#_c_456_n 0.0117963f $X=1.84 $Y=1.32 $X2=0 $Y2=0
cc_275 N_S0_M1026_g N_A_27_47#_c_456_n 0.00433144f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_276 N_S0_c_210_n N_A_27_47#_c_456_n 0.00800201f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_277 N_S0_c_211_n N_A_27_47#_c_456_n 2.65465e-19 $X=1.3 $Y=1.53 $X2=0 $Y2=0
cc_278 N_S0_c_197_n N_A_27_47#_c_456_n 0.0226549f $X=1.155 $Y=1.53 $X2=0 $Y2=0
cc_279 N_S0_M1026_g N_A3_c_688_n 0.00975299f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_280 N_S0_c_210_n N_A3_c_688_n 0.00281616f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_281 N_S0_c_210_n N_A3_c_695_n 0.00588092f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_282 N_S0_M1026_g A3 8.90548e-19 $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_283 N_S0_c_210_n A3 0.00539843f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_284 N_S0_M1026_g A3 2.79419e-19 $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_285 N_S0_c_210_n A3 0.0104635f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_286 N_S0_M1026_g N_A3_c_691_n 0.0143597f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_287 N_S0_c_210_n N_A3_c_691_n 9.68438e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_288 N_S0_M1026_g N_A3_c_692_n 0.0238303f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_289 N_S0_c_210_n N_S1_c_747_n 7.7475e-19 $X=6.07 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_290 N_S0_c_210_n N_S1_M1027_g 0.00682163f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_291 N_S0_c_210_n N_S1_c_750_n 0.00336531f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_292 N_S0_c_210_n N_S1_M1013_g 0.00625641f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_293 N_S0_c_210_n S1 0.0121766f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_294 N_S0_c_210_n N_A_601_345#_M1019_g 0.00412283f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_295 N_S0_c_210_n N_A_601_345#_c_833_n 0.00309622f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_296 N_S0_c_210_n N_A_601_345#_c_835_n 0.00452009f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_297 N_S0_c_210_n N_A_601_345#_c_838_n 0.0266831f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_298 N_S0_c_210_n N_A1_M1000_g 0.00948456f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_299 N_S0_M1010_g N_A1_M1024_g 0.029526f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_300 N_S0_c_210_n A1 0.0107577f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_301 N_S0_M1010_g N_A1_c_904_n 0.00455685f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_302 N_S0_c_210_n N_A1_c_904_n 0.00145767f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_303 N_S0_M1016_g N_A0_M1022_g 0.0345762f $X=6.325 $Y=2.275 $X2=0 $Y2=0
cc_304 N_S0_c_214_n N_A0_M1022_g 9.18038e-19 $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_305 N_S0_c_199_n N_A0_M1022_g 0.0136507f $X=6.385 $Y=1.32 $X2=0 $Y2=0
cc_306 N_S0_M1010_g N_A0_c_943_n 2.01922e-19 $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_307 N_S0_c_214_n N_A0_c_943_n 0.00629593f $X=6.215 $Y=1.53 $X2=0 $Y2=0
cc_308 N_S0_c_199_n N_A0_c_943_n 5.65638e-19 $X=6.385 $Y=1.32 $X2=0 $Y2=0
cc_309 N_S0_c_199_n N_A0_c_944_n 0.00525853f $X=6.385 $Y=1.32 $X2=0 $Y2=0
cc_310 N_S0_c_210_n N_A_789_316#_M1019_d 6.16189e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_311 N_S0_c_210_n N_A_789_316#_c_998_n 0.0139892f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_312 N_S0_M1016_g N_A_789_316#_c_1008_n 0.00848933f $X=6.325 $Y=2.275 $X2=0
+ $Y2=0
cc_313 N_S0_M1016_g N_A_789_316#_c_1010_n 7.58543e-19 $X=6.325 $Y=2.275 $X2=0
+ $Y2=0
cc_314 N_S0_c_213_n N_A_789_316#_c_1010_n 9.4687e-19 $X=6.215 $Y=1.53 $X2=0
+ $Y2=0
cc_315 N_S0_c_214_n N_A_789_316#_c_1010_n 0.00987457f $X=6.215 $Y=1.53 $X2=0
+ $Y2=0
cc_316 N_S0_c_199_n N_A_789_316#_c_1010_n 5.56235e-19 $X=6.385 $Y=1.32 $X2=0
+ $Y2=0
cc_317 N_S0_c_214_n N_A_789_316#_c_1011_n 0.00454895f $X=6.215 $Y=1.53 $X2=0
+ $Y2=0
cc_318 N_S0_M1016_g N_A_789_316#_c_1014_n 0.00380986f $X=6.325 $Y=2.275 $X2=0
+ $Y2=0
cc_319 N_S0_c_210_n N_A_789_316#_c_1014_n 0.00774624f $X=6.07 $Y=1.53 $X2=0
+ $Y2=0
cc_320 N_S0_c_213_n N_A_789_316#_c_1014_n 0.0150323f $X=6.215 $Y=1.53 $X2=0
+ $Y2=0
cc_321 N_S0_c_214_n N_A_789_316#_c_1014_n 0.00544375f $X=6.215 $Y=1.53 $X2=0
+ $Y2=0
cc_322 N_S0_c_199_n N_A_789_316#_c_1014_n 9.57678e-19 $X=6.385 $Y=1.32 $X2=0
+ $Y2=0
cc_323 N_S0_M1016_g N_A_789_316#_c_1030_n 0.00100458f $X=6.325 $Y=2.275 $X2=0
+ $Y2=0
cc_324 N_S0_M1016_g N_A_789_316#_c_1031_n 0.00151791f $X=6.325 $Y=2.275 $X2=0
+ $Y2=0
cc_325 N_S0_M1021_g N_VPWR_c_1178_n 0.01126f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_326 N_S0_M1025_g N_VPWR_c_1178_n 0.00199783f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_327 N_S0_M1025_g N_VPWR_c_1185_n 0.00546481f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_328 N_S0_M1016_g N_VPWR_c_1187_n 0.00545391f $X=6.325 $Y=2.275 $X2=0 $Y2=0
cc_329 N_S0_M1021_g N_VPWR_c_1189_n 0.0033925f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_330 N_S0_M1021_g N_VPWR_c_1177_n 0.004976f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_331 N_S0_M1025_g N_VPWR_c_1177_n 0.00624711f $X=1.37 $Y=2.275 $X2=0 $Y2=0
cc_332 N_S0_M1016_g N_VPWR_c_1177_n 0.00557212f $X=6.325 $Y=2.275 $X2=0 $Y2=0
cc_333 N_S0_c_210_n N_A_288_47#_M1019_s 6.75395e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_334 N_S0_M1025_g N_A_288_47#_c_1337_n 0.00428325f $X=1.37 $Y=2.275 $X2=0
+ $Y2=0
cc_335 N_S0_M1026_g N_A_288_47#_c_1338_n 0.0106725f $X=1.915 $Y=0.415 $X2=0
+ $Y2=0
cc_336 N_S0_M1026_g N_A_288_47#_c_1325_n 0.016315f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_337 N_S0_c_210_n N_A_288_47#_c_1329_n 0.0139277f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_338 N_S0_c_210_n N_A_288_47#_c_1341_n 5.58339e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_339 N_S0_c_191_n N_A_288_47#_c_1326_n 0.00510606f $X=1.84 $Y=1.32 $X2=0 $Y2=0
cc_340 N_S0_M1026_g N_A_288_47#_c_1326_n 4.69181e-19 $X=1.915 $Y=0.415 $X2=0
+ $Y2=0
cc_341 N_S0_c_210_n N_A_288_47#_c_1326_n 0.0104059f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_342 N_S0_c_210_n N_A_288_47#_c_1327_n 0.0127493f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_343 N_S0_c_210_n N_A_873_316#_M1013_d 2.14086e-19 $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_344 N_S0_c_210_n N_A_873_316#_c_1463_n 0.0203392f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_345 N_S0_c_210_n N_A_873_316#_c_1466_n 0.0198601f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_346 N_S0_M1010_g N_A_873_316#_c_1464_n 0.00712483f $X=5.785 $Y=0.415 $X2=0
+ $Y2=0
cc_347 N_S0_c_210_n N_A_873_316#_c_1464_n 0.0155282f $X=6.07 $Y=1.53 $X2=0 $Y2=0
cc_348 N_S0_M1010_g N_A_873_316#_c_1475_n 0.0110411f $X=5.785 $Y=0.415 $X2=0
+ $Y2=0
cc_349 N_S0_M1016_g N_A_873_316#_c_1476_n 0.00246628f $X=6.325 $Y=2.275 $X2=0
+ $Y2=0
cc_350 N_S0_c_210_n N_A_873_316#_c_1476_n 9.00069e-19 $X=6.07 $Y=1.53 $X2=0
+ $Y2=0
cc_351 N_S0_c_213_n N_A_873_316#_c_1476_n 0.00117806f $X=6.215 $Y=1.53 $X2=0
+ $Y2=0
cc_352 N_S0_c_214_n N_A_873_316#_c_1476_n 0.00270797f $X=6.215 $Y=1.53 $X2=0
+ $Y2=0
cc_353 N_S0_c_210_n N_A_873_316#_c_1469_n 0.00369858f $X=6.07 $Y=1.53 $X2=0
+ $Y2=0
cc_354 N_S0_M1029_g N_VGND_c_1619_n 0.0112612f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_355 N_S0_M1026_g N_VGND_c_1620_n 0.00171495f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_356 N_S0_M1029_g N_VGND_c_1626_n 0.00339367f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_357 N_S0_M1026_g N_VGND_c_1627_n 0.00379702f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_358 N_S0_M1010_g N_VGND_c_1629_n 0.00366111f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_359 N_S0_M1029_g N_VGND_c_1637_n 0.00497794f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_360 N_S0_M1026_g N_VGND_c_1637_n 0.00584218f $X=1.915 $Y=0.415 $X2=0 $Y2=0
cc_361 N_S0_M1010_g N_VGND_c_1637_n 0.00589952f $X=5.785 $Y=0.415 $X2=0 $Y2=0
cc_362 A2 N_A_27_47#_c_447_n 0.0030487f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_363 N_A2_c_394_n N_A_27_47#_c_447_n 0.0221703f $X=0.925 $Y=0.765 $X2=0 $Y2=0
cc_364 N_A2_M1001_g N_A_27_47#_c_449_n 0.0102831f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_365 A2 N_A_27_47#_c_449_n 0.0221499f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_366 N_A2_c_393_n N_A_27_47#_c_449_n 0.00180072f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_367 N_A2_M1001_g N_A_27_47#_c_460_n 0.0120729f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_368 N_A2_c_393_n N_A_27_47#_c_460_n 0.00158391f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_369 N_A2_M1001_g N_A_27_47#_c_461_n 0.00346204f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_370 A2 N_A_27_47#_c_450_n 0.00642654f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_371 A2 N_A_27_47#_c_450_n 0.00319986f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_372 N_A2_c_393_n N_A_27_47#_c_450_n 2.8911e-19 $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_373 N_A2_c_394_n N_A_27_47#_c_450_n 0.00118376f $X=0.925 $Y=0.765 $X2=0 $Y2=0
cc_374 A2 N_A_27_47#_c_451_n 0.00207962f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_375 N_A2_c_393_n N_A_27_47#_c_451_n 0.0148435f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_376 A2 N_A_27_47#_c_452_n 0.0045313f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_377 A2 N_A_27_47#_c_452_n 0.0217225f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_378 N_A2_c_393_n N_A_27_47#_c_452_n 2.04707e-19 $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_379 N_A2_M1001_g N_A_27_47#_c_456_n 0.00344585f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_380 A2 N_A_27_47#_c_456_n 0.00304052f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_381 N_A2_c_393_n N_A_27_47#_c_456_n 2.60449e-19 $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_382 N_A2_M1001_g N_VPWR_c_1178_n 0.00982614f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_383 N_A2_M1001_g N_VPWR_c_1185_n 0.0046653f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_384 N_A2_M1001_g N_VPWR_c_1177_n 0.00442041f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_385 N_A2_M1001_g N_A_288_47#_c_1337_n 7.34665e-19 $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_386 A2 N_A_288_47#_c_1325_n 0.00346292f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_387 A2 N_VGND_c_1619_n 0.00503234f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_388 N_A2_c_394_n N_VGND_c_1619_n 0.0101171f $X=0.925 $Y=0.765 $X2=0 $Y2=0
cc_389 A2 N_VGND_c_1627_n 0.00740795f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_390 N_A2_c_393_n N_VGND_c_1627_n 0.00115507f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_391 N_A2_c_394_n N_VGND_c_1627_n 0.0046653f $X=0.925 $Y=0.765 $X2=0 $Y2=0
cc_392 A2 N_VGND_c_1637_n 0.00741879f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_393 A2 N_VGND_c_1637_n 0.00599839f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_394 N_A2_c_393_n N_VGND_c_1637_n 0.00143621f $X=0.925 $Y=0.93 $X2=0 $Y2=0
cc_395 N_A2_c_394_n N_VGND_c_1637_n 0.00440885f $X=0.925 $Y=0.765 $X2=0 $Y2=0
cc_396 A2 A_193_47# 0.00752768f $X=1.07 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_397 N_A_27_47#_c_456_n N_A3_c_688_n 2.69784e-19 $X=1.735 $Y=1.575 $X2=0 $Y2=0
cc_398 N_A_27_47#_M1017_g N_A3_c_694_n 0.0138424f $X=1.79 $Y=2.275 $X2=0 $Y2=0
cc_399 N_A_27_47#_c_462_n N_A3_c_694_n 0.00580906f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_400 N_A_27_47#_c_465_n N_A3_c_694_n 0.00498599f $X=1.82 $Y=1.74 $X2=0 $Y2=0
cc_401 N_A_27_47#_c_462_n N_A3_c_695_n 0.00220307f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_402 N_A_27_47#_c_465_n N_A3_c_695_n 0.00134881f $X=1.82 $Y=1.74 $X2=0 $Y2=0
cc_403 N_A_27_47#_c_462_n N_S1_M1027_g 0.00310138f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_404 N_A_27_47#_c_462_n N_S1_c_754_n 7.54852e-19 $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_405 N_A_27_47#_c_462_n N_S1_M1013_g 0.00272158f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_406 N_A_27_47#_c_462_n N_A_601_345#_M1019_g 0.00263087f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_462_n N_A_601_345#_c_838_n 0.0185991f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_M1023_g N_A1_M1000_g 0.0154632f $X=5.905 $Y=2.275 $X2=0 $Y2=0
cc_409 N_A_27_47#_c_462_n N_A1_M1000_g 0.00637365f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_410 N_A_27_47#_c_467_n N_A1_M1000_g 0.00734459f $X=5.875 $Y=1.74 $X2=0 $Y2=0
cc_411 N_A_27_47#_c_454_n N_A1_M1000_g 0.00131494f $X=5.875 $Y=1.74 $X2=0 $Y2=0
cc_412 N_A_27_47#_c_448_n N_A0_M1020_g 0.0317614f $X=6.335 $Y=0.705 $X2=0 $Y2=0
cc_413 N_A_27_47#_c_453_n N_A0_M1020_g 2.38614e-19 $X=6.205 $Y=0.87 $X2=0 $Y2=0
cc_414 N_A_27_47#_c_453_n N_A0_c_943_n 0.00248128f $X=6.205 $Y=0.87 $X2=0 $Y2=0
cc_415 N_A_27_47#_c_454_n N_A0_c_943_n 0.00143247f $X=5.875 $Y=1.74 $X2=0 $Y2=0
cc_416 N_A_27_47#_c_455_n N_A0_c_943_n 3.79122e-19 $X=6.335 $Y=0.87 $X2=0 $Y2=0
cc_417 N_A_27_47#_c_455_n N_A0_c_944_n 0.00142667f $X=6.335 $Y=0.87 $X2=0 $Y2=0
cc_418 N_A_27_47#_c_448_n A0 0.00936228f $X=6.335 $Y=0.705 $X2=0 $Y2=0
cc_419 N_A_27_47#_c_453_n A0 0.0178996f $X=6.205 $Y=0.87 $X2=0 $Y2=0
cc_420 N_A_27_47#_c_462_n N_A_789_316#_M1019_d 0.00139404f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_462_n N_A_789_316#_c_998_n 0.0146457f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1023_g N_A_789_316#_c_1014_n 0.00125658f $X=5.905 $Y=2.275
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_462_n N_A_789_316#_c_1014_n 0.0865979f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_464_n N_A_789_316#_c_1014_n 0.0265153f $X=5.755 $Y=1.87
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_c_467_n N_A_789_316#_c_1014_n 9.1661e-19 $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_454_n N_A_789_316#_c_1014_n 0.00140404f $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_427 N_A_27_47#_c_462_n N_A_789_316#_c_1015_n 0.0274654f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_462_n N_A_789_316#_c_1016_n 0.00376868f $X=5.61 $Y=1.87
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_460_n N_VPWR_M1021_d 0.00116722f $X=1.565 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_430 N_A_27_47#_c_461_n N_VPWR_M1021_d 0.00242809f $X=0.67 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_431 N_A_27_47#_c_462_n N_VPWR_M1002_d 0.00361504f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_462_n N_VPWR_M1000_s 0.00166679f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_433 N_A_27_47#_c_460_n N_VPWR_c_1178_n 0.00538445f $X=1.565 $Y=1.87 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_461_n N_VPWR_c_1178_n 0.00798323f $X=0.67 $Y=1.87 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_c_462_n N_VPWR_c_1179_n 0.0081452f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_436 N_A_27_47#_c_462_n N_VPWR_c_1180_n 0.00382585f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_M1017_g N_VPWR_c_1185_n 0.00390868f $X=1.79 $Y=2.275 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_M1023_g N_VPWR_c_1187_n 0.00385416f $X=5.905 $Y=2.275 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_c_606_p N_VPWR_c_1189_n 0.00886455f $X=0.26 $Y=2.21 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_c_461_n N_VPWR_c_1189_n 0.00246701f $X=0.67 $Y=1.87 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_M1021_s N_VPWR_c_1177_n 0.00233501f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_M1017_g N_VPWR_c_1177_n 0.0059629f $X=1.79 $Y=2.275 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_M1023_g N_VPWR_c_1177_n 0.00539892f $X=5.905 $Y=2.275 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_606_p N_VPWR_c_1177_n 0.00753677f $X=0.26 $Y=2.21 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_460_n N_VPWR_c_1177_n 0.0200614f $X=1.565 $Y=1.87 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_c_461_n N_VPWR_c_1177_n 0.00504f $X=0.67 $Y=1.87 $X2=0 $Y2=0
cc_447 N_A_27_47#_c_462_n N_VPWR_c_1177_n 0.0370753f $X=5.61 $Y=1.87 $X2=0 $Y2=0
cc_448 N_A_27_47#_c_463_n N_VPWR_c_1177_n 0.0160199f $X=1.76 $Y=1.87 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_460_n A_193_369# 0.00373969f $X=1.565 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_450 N_A_27_47#_c_462_n N_A_288_47#_M1019_s 0.00112767f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_M1017_g N_A_288_47#_c_1337_n 0.00945162f $X=1.79 $Y=2.275
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_c_460_n N_A_288_47#_c_1337_n 0.00793212f $X=1.565 $Y=1.87
+ $X2=0 $Y2=0
cc_453 N_A_27_47#_c_462_n N_A_288_47#_c_1337_n 0.00239538f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_463_n N_A_288_47#_c_1337_n 0.00325767f $X=1.76 $Y=1.87 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_465_n N_A_288_47#_c_1337_n 0.00203367f $X=1.82 $Y=1.74 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_466_n N_A_288_47#_c_1337_n 0.019174f $X=1.82 $Y=1.74 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_451_n N_A_288_47#_c_1338_n 0.00342692f $X=1.495 $Y=0.87
+ $X2=0 $Y2=0
cc_458 N_A_27_47#_c_452_n N_A_288_47#_c_1338_n 0.0180135f $X=1.65 $Y=0.87 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_447_n N_A_288_47#_c_1325_n 5.93063e-19 $X=1.365 $Y=0.705
+ $X2=0 $Y2=0
cc_460 N_A_27_47#_c_451_n N_A_288_47#_c_1325_n 3.02207e-19 $X=1.495 $Y=0.87
+ $X2=0 $Y2=0
cc_461 N_A_27_47#_c_452_n N_A_288_47#_c_1325_n 0.024855f $X=1.65 $Y=0.87 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_456_n N_A_288_47#_c_1325_n 0.0143036f $X=1.735 $Y=1.575
+ $X2=0 $Y2=0
cc_463 N_A_27_47#_M1017_g N_A_288_47#_c_1329_n 0.00391048f $X=1.79 $Y=2.275
+ $X2=0 $Y2=0
cc_464 N_A_27_47#_c_462_n N_A_288_47#_c_1329_n 0.0132084f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_463_n N_A_288_47#_c_1329_n 0.00147315f $X=1.76 $Y=1.87 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_465_n N_A_288_47#_c_1329_n 0.0023745f $X=1.82 $Y=1.74 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_466_n N_A_288_47#_c_1329_n 0.0274922f $X=1.82 $Y=1.74 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_456_n N_A_288_47#_c_1329_n 0.00661642f $X=1.735 $Y=1.575
+ $X2=0 $Y2=0
cc_469 N_A_27_47#_c_462_n N_A_288_47#_c_1341_n 0.00744441f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_462_n N_A_288_47#_c_1330_n 0.00187686f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_462_n N_A_288_47#_c_1331_n 0.00418499f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_465_n N_A_288_47#_c_1326_n 0.00156489f $X=1.82 $Y=1.74 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_456_n N_A_288_47#_c_1326_n 0.0121557f $X=1.735 $Y=1.575
+ $X2=0 $Y2=0
cc_474 N_A_27_47#_c_462_n N_A_288_47#_c_1327_n 0.00302831f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_462_n N_A_288_47#_c_1334_n 0.0865557f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_M1017_g N_A_288_47#_c_1374_n 0.00114372f $X=1.79 $Y=2.275
+ $X2=0 $Y2=0
cc_477 N_A_27_47#_c_462_n N_A_288_47#_c_1374_n 0.0263636f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_465_n N_A_288_47#_c_1374_n 2.73637e-19 $X=1.82 $Y=1.74 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_462_n N_A_288_47#_c_1335_n 0.0276035f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_c_462_n A_373_413# 0.00325861f $X=5.61 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_481 N_A_27_47#_c_462_n N_A_873_316#_M1013_d 0.00209072f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_462_n N_A_873_316#_c_1463_n 0.0108836f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_462_n N_A_873_316#_c_1466_n 0.0143232f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_c_453_n N_A_873_316#_c_1464_n 0.0274865f $X=6.205 $Y=0.87
+ $X2=0 $Y2=0
cc_485 N_A_27_47#_c_454_n N_A_873_316#_c_1464_n 0.0406897f $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_486 N_A_27_47#_M1023_g N_A_873_316#_c_1468_n 0.00337169f $X=5.905 $Y=2.275
+ $X2=0 $Y2=0
cc_487 N_A_27_47#_c_462_n N_A_873_316#_c_1468_n 0.0140427f $X=5.61 $Y=1.87 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_464_n N_A_873_316#_c_1468_n 0.00275409f $X=5.755 $Y=1.87
+ $X2=0 $Y2=0
cc_489 N_A_27_47#_c_467_n N_A_873_316#_c_1468_n 4.04648e-19 $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_490 N_A_27_47#_c_454_n N_A_873_316#_c_1468_n 0.0172732f $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_491 N_A_27_47#_c_453_n N_A_873_316#_c_1475_n 0.0259764f $X=6.205 $Y=0.87
+ $X2=0 $Y2=0
cc_492 N_A_27_47#_c_455_n N_A_873_316#_c_1475_n 0.00325712f $X=6.335 $Y=0.87
+ $X2=0 $Y2=0
cc_493 N_A_27_47#_M1023_g N_A_873_316#_c_1476_n 0.00887377f $X=5.905 $Y=2.275
+ $X2=0 $Y2=0
cc_494 N_A_27_47#_c_462_n N_A_873_316#_c_1476_n 7.78043e-19 $X=5.61 $Y=1.87
+ $X2=0 $Y2=0
cc_495 N_A_27_47#_c_464_n N_A_873_316#_c_1476_n 7.97005e-19 $X=5.755 $Y=1.87
+ $X2=0 $Y2=0
cc_496 N_A_27_47#_c_467_n N_A_873_316#_c_1476_n 0.00193698f $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_497 N_A_27_47#_c_454_n N_A_873_316#_c_1476_n 0.0189711f $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_498 N_A_27_47#_c_467_n N_A_873_316#_c_1469_n 5.13754e-19 $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_499 N_A_27_47#_c_454_n N_A_873_316#_c_1469_n 0.0142775f $X=5.875 $Y=1.74
+ $X2=0 $Y2=0
cc_500 N_A_27_47#_c_462_n A_1061_369# 4.93895e-19 $X=5.61 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_501 N_A_27_47#_c_450_n N_VGND_M1029_d 9.16826e-19 $X=0.585 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_502 N_A_27_47#_c_447_n N_VGND_c_1619_n 0.00170713f $X=1.365 $Y=0.705 $X2=0
+ $Y2=0
cc_503 N_A_27_47#_c_450_n N_VGND_c_1619_n 0.00721829f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_c_671_p N_VGND_c_1626_n 0.00859955f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_c_450_n N_VGND_c_1626_n 0.0024638f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_c_447_n N_VGND_c_1627_n 0.00555329f $X=1.365 $Y=0.705 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_451_n N_VGND_c_1627_n 6.43063e-19 $X=1.495 $Y=0.87 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_452_n N_VGND_c_1627_n 9.49253e-19 $X=1.65 $Y=0.87 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_c_448_n N_VGND_c_1629_n 0.00555329f $X=6.335 $Y=0.705 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_c_453_n N_VGND_c_1629_n 9.49253e-19 $X=6.205 $Y=0.87 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_c_455_n N_VGND_c_1629_n 6.11083e-19 $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_512 N_A_27_47#_M1029_s N_VGND_c_1637_n 0.00234741f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_c_447_n N_VGND_c_1637_n 0.0103474f $X=1.365 $Y=0.705 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_448_n N_VGND_c_1637_n 0.0103474f $X=6.335 $Y=0.705 $X2=0
+ $Y2=0
cc_515 N_A_27_47#_c_671_p N_VGND_c_1637_n 0.00743105f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_c_450_n N_VGND_c_1637_n 0.00497314f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_451_n N_VGND_c_1637_n 8.53329e-19 $X=1.495 $Y=0.87 $X2=0
+ $Y2=0
cc_518 N_A_27_47#_c_452_n N_VGND_c_1637_n 0.00205647f $X=1.65 $Y=0.87 $X2=0
+ $Y2=0
cc_519 N_A_27_47#_c_453_n N_VGND_c_1637_n 0.00295441f $X=6.205 $Y=0.87 $X2=0
+ $Y2=0
cc_520 N_A_27_47#_c_455_n N_VGND_c_1637_n 8.53329e-19 $X=6.335 $Y=0.87 $X2=0
+ $Y2=0
cc_521 A3 N_S1_c_747_n 0.00214806f $X=2.45 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_522 N_A3_c_691_n N_S1_c_747_n 0.0207417f $X=2.41 $Y=0.93 $X2=-0.19 $Y2=-0.24
cc_523 N_A3_c_692_n N_S1_c_747_n 0.00103795f $X=2.41 $Y=0.765 $X2=-0.19
+ $Y2=-0.24
cc_524 N_A3_c_688_n N_S1_M1027_g 0.0126585f $X=2.395 $Y=1.5 $X2=0 $Y2=0
cc_525 N_A3_c_695_n N_S1_M1027_g 0.0187074f $X=2.51 $Y=1.575 $X2=0 $Y2=0
cc_526 A3 N_S1_M1027_g 6.79827e-19 $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_527 N_A3_c_692_n N_S1_c_749_n 0.0137149f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_528 N_A3_c_694_n N_S1_c_755_n 0.0187074f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_529 N_A3_c_688_n S1 5.90277e-19 $X=2.395 $Y=1.5 $X2=0 $Y2=0
cc_530 A3 S1 0.0478665f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_531 N_A3_c_691_n S1 3.38407e-19 $X=2.41 $Y=0.93 $X2=0 $Y2=0
cc_532 N_A3_c_694_n N_A_601_345#_c_838_n 0.00125935f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_533 N_A3_c_694_n N_VPWR_c_1179_n 0.0064285f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_534 N_A3_c_694_n N_VPWR_c_1185_n 0.00585385f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_535 N_A3_c_694_n N_VPWR_c_1177_n 0.00587666f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_536 N_A3_c_692_n N_A_288_47#_c_1338_n 0.00145818f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_537 N_A3_c_688_n N_A_288_47#_c_1325_n 9.61953e-19 $X=2.395 $Y=1.5 $X2=0 $Y2=0
cc_538 A3 N_A_288_47#_c_1325_n 0.0240227f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_539 A3 N_A_288_47#_c_1325_n 0.00948099f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_540 N_A3_c_691_n N_A_288_47#_c_1325_n 0.00133579f $X=2.41 $Y=0.93 $X2=0 $Y2=0
cc_541 N_A3_c_692_n N_A_288_47#_c_1325_n 0.00349406f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_542 N_A3_c_688_n N_A_288_47#_c_1329_n 0.00798315f $X=2.395 $Y=1.5 $X2=0 $Y2=0
cc_543 N_A3_c_694_n N_A_288_47#_c_1329_n 0.0105472f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_544 N_A3_c_688_n N_A_288_47#_c_1326_n 0.00307277f $X=2.395 $Y=1.5 $X2=0 $Y2=0
cc_545 A3 N_A_288_47#_c_1326_n 0.00647251f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_546 N_A3_c_694_n N_A_288_47#_c_1334_n 0.00410206f $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_547 N_A3_c_694_n N_A_288_47#_c_1374_n 4.9262e-19 $X=2.51 $Y=1.65 $X2=0 $Y2=0
cc_548 A3 N_VGND_c_1620_n 0.0115245f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_549 N_A3_c_691_n N_VGND_c_1620_n 3.61231e-19 $X=2.41 $Y=0.93 $X2=0 $Y2=0
cc_550 N_A3_c_692_n N_VGND_c_1620_n 0.00975119f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_551 A3 N_VGND_c_1627_n 0.00314583f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_552 N_A3_c_692_n N_VGND_c_1627_n 0.00391931f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_553 A3 N_VGND_c_1637_n 0.00579556f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_554 N_A3_c_692_n N_VGND_c_1637_n 0.00476517f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_555 N_S1_c_754_n N_A_601_345#_M1019_g 0.00975169f $X=4.215 $Y=2.54 $X2=0
+ $Y2=0
cc_556 N_S1_M1013_g N_A_601_345#_M1019_g 0.0197432f $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_557 N_S1_M1013_g N_A_601_345#_c_833_n 0.0120884f $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_558 N_S1_c_751_n N_A_601_345#_M1007_g 0.0192711f $X=3.885 $Y=0.73 $X2=0 $Y2=0
cc_559 N_S1_c_747_n N_A_601_345#_c_835_n 3.3029e-19 $X=2.93 $Y=1.095 $X2=0 $Y2=0
cc_560 N_S1_M1027_g N_A_601_345#_c_835_n 0.0156633f $X=2.93 $Y=2.045 $X2=0 $Y2=0
cc_561 N_S1_c_750_n N_A_601_345#_c_835_n 0.0490984f $X=3.81 $Y=0.805 $X2=0 $Y2=0
cc_562 S1 N_A_601_345#_c_835_n 0.00152957f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_563 N_S1_c_747_n N_A_601_345#_c_837_n 0.00109538f $X=2.93 $Y=1.095 $X2=0
+ $Y2=0
cc_564 N_S1_c_749_n N_A_601_345#_c_837_n 0.00538776f $X=2.935 $Y=0.73 $X2=0
+ $Y2=0
cc_565 N_S1_c_750_n N_A_601_345#_c_837_n 0.0116555f $X=3.81 $Y=0.805 $X2=0 $Y2=0
cc_566 N_S1_c_751_n N_A_601_345#_c_837_n 6.32935e-19 $X=3.885 $Y=0.73 $X2=0
+ $Y2=0
cc_567 S1 N_A_601_345#_c_837_n 0.0258653f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_568 N_S1_M1027_g N_A_601_345#_c_838_n 0.0179348f $X=2.93 $Y=2.045 $X2=0 $Y2=0
cc_569 N_S1_c_754_n N_A_601_345#_c_838_n 0.00578358f $X=4.215 $Y=2.54 $X2=0
+ $Y2=0
cc_570 N_S1_c_750_n N_A_601_345#_c_838_n 0.00300126f $X=3.81 $Y=0.805 $X2=0
+ $Y2=0
cc_571 S1 N_A_601_345#_c_838_n 0.0214342f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_572 N_S1_c_749_n N_A_601_345#_c_839_n 0.00233282f $X=2.935 $Y=0.73 $X2=0
+ $Y2=0
cc_573 N_S1_c_750_n N_A_601_345#_c_839_n 0.00530393f $X=3.81 $Y=0.805 $X2=0
+ $Y2=0
cc_574 N_S1_c_751_n N_A_601_345#_c_839_n 0.00108928f $X=3.885 $Y=0.73 $X2=0
+ $Y2=0
cc_575 S1 N_A_601_345#_c_839_n 0.00330055f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_576 N_S1_c_751_n N_A_789_316#_c_998_n 0.00191245f $X=3.885 $Y=0.73 $X2=0
+ $Y2=0
cc_577 N_S1_M1013_g N_A_789_316#_c_998_n 0.00238534f $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_578 N_S1_c_754_n N_A_789_316#_c_1012_n 0.00293376f $X=4.215 $Y=2.54 $X2=0
+ $Y2=0
cc_579 N_S1_M1013_g N_A_789_316#_c_1015_n 0.00411296f $X=4.29 $Y=1.85 $X2=0
+ $Y2=0
cc_580 N_S1_M1013_g N_A_789_316#_c_1016_n 0.0125788f $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_581 N_S1_M1027_g N_VPWR_c_1179_n 0.00655497f $X=2.93 $Y=2.045 $X2=0 $Y2=0
cc_582 N_S1_M1013_g N_VPWR_c_1180_n 0.0110777f $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_583 N_S1_c_755_n N_VPWR_c_1190_n 0.0435688f $X=3.005 $Y=2.54 $X2=0 $Y2=0
cc_584 N_S1_c_754_n N_VPWR_c_1177_n 0.0304569f $X=4.215 $Y=2.54 $X2=0 $Y2=0
cc_585 N_S1_c_755_n N_VPWR_c_1177_n 0.00442783f $X=3.005 $Y=2.54 $X2=0 $Y2=0
cc_586 N_S1_M1027_g N_A_288_47#_c_1330_n 0.0024883f $X=2.93 $Y=2.045 $X2=0 $Y2=0
cc_587 N_S1_c_754_n N_A_288_47#_c_1330_n 0.0101272f $X=4.215 $Y=2.54 $X2=0 $Y2=0
cc_588 N_S1_M1013_g N_A_288_47#_c_1330_n 2.99929e-19 $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_589 N_S1_M1027_g N_A_288_47#_c_1331_n 0.00263002f $X=2.93 $Y=2.045 $X2=0
+ $Y2=0
cc_590 N_S1_c_750_n N_A_288_47#_c_1327_n 0.00890714f $X=3.81 $Y=0.805 $X2=0
+ $Y2=0
cc_591 N_S1_c_751_n N_A_288_47#_c_1327_n 0.00142837f $X=3.885 $Y=0.73 $X2=0
+ $Y2=0
cc_592 N_S1_c_750_n N_A_288_47#_c_1328_n 0.00269638f $X=3.81 $Y=0.805 $X2=0
+ $Y2=0
cc_593 N_S1_c_751_n N_A_288_47#_c_1328_n 0.00362535f $X=3.885 $Y=0.73 $X2=0
+ $Y2=0
cc_594 N_S1_M1027_g N_A_288_47#_c_1334_n 0.0049068f $X=2.93 $Y=2.045 $X2=0 $Y2=0
cc_595 N_S1_c_754_n N_A_288_47#_c_1334_n 0.00260084f $X=4.215 $Y=2.54 $X2=0
+ $Y2=0
cc_596 N_S1_M1027_g N_A_288_47#_c_1335_n 0.00136441f $X=2.93 $Y=2.045 $X2=0
+ $Y2=0
cc_597 N_S1_c_754_n N_A_288_47#_c_1335_n 0.00358607f $X=4.215 $Y=2.54 $X2=0
+ $Y2=0
cc_598 N_S1_M1013_g N_A_288_47#_c_1335_n 5.70583e-19 $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_599 N_S1_M1013_g N_A_873_316#_c_1463_n 0.0028409f $X=4.29 $Y=1.85 $X2=0 $Y2=0
cc_600 N_S1_c_747_n N_VGND_c_1620_n 0.00120134f $X=2.93 $Y=1.095 $X2=0 $Y2=0
cc_601 N_S1_c_749_n N_VGND_c_1620_n 0.00710898f $X=2.935 $Y=0.73 $X2=0 $Y2=0
cc_602 N_S1_c_747_n N_VGND_c_1628_n 3.27123e-19 $X=2.93 $Y=1.095 $X2=0 $Y2=0
cc_603 N_S1_c_749_n N_VGND_c_1628_n 0.00426984f $X=2.935 $Y=0.73 $X2=0 $Y2=0
cc_604 N_S1_c_750_n N_VGND_c_1628_n 0.0030174f $X=3.81 $Y=0.805 $X2=0 $Y2=0
cc_605 N_S1_c_751_n N_VGND_c_1628_n 0.00565823f $X=3.885 $Y=0.73 $X2=0 $Y2=0
cc_606 S1 N_VGND_c_1628_n 0.00312826f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_607 N_S1_c_749_n N_VGND_c_1637_n 0.00749741f $X=2.935 $Y=0.73 $X2=0 $Y2=0
cc_608 N_S1_c_750_n N_VGND_c_1637_n 0.00370828f $X=3.81 $Y=0.805 $X2=0 $Y2=0
cc_609 N_S1_c_751_n N_VGND_c_1637_n 0.0117171f $X=3.885 $Y=0.73 $X2=0 $Y2=0
cc_610 S1 N_VGND_c_1637_n 0.00521238f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_611 N_A_601_345#_M1007_g N_A1_c_904_n 0.00306719f $X=4.31 $Y=0.445 $X2=0
+ $Y2=0
cc_612 N_A_601_345#_c_833_n N_A_789_316#_c_998_n 0.015488f $X=4.235 $Y=1.165
+ $X2=0 $Y2=0
cc_613 N_A_601_345#_M1007_g N_A_789_316#_c_998_n 0.00651443f $X=4.31 $Y=0.445
+ $X2=0 $Y2=0
cc_614 N_A_601_345#_c_836_n N_A_789_316#_c_998_n 0.007437f $X=3.87 $Y=1.225
+ $X2=0 $Y2=0
cc_615 N_A_601_345#_M1019_g N_A_789_316#_c_1012_n 9.91098e-19 $X=3.87 $Y=1.85
+ $X2=0 $Y2=0
cc_616 N_A_601_345#_M1019_g N_VPWR_c_1177_n 4.46264e-19 $X=3.87 $Y=1.85 $X2=0
+ $Y2=0
cc_617 N_A_601_345#_M1019_g N_A_288_47#_c_1341_n 8.98734e-19 $X=3.87 $Y=1.85
+ $X2=0 $Y2=0
cc_618 N_A_601_345#_c_835_n N_A_288_47#_c_1341_n 0.00184988f $X=3.795 $Y=1.225
+ $X2=0 $Y2=0
cc_619 N_A_601_345#_c_838_n N_A_288_47#_c_1341_n 0.00702473f $X=3.4 $Y=1.225
+ $X2=0 $Y2=0
cc_620 N_A_601_345#_M1019_g N_A_288_47#_c_1330_n 0.00424598f $X=3.87 $Y=1.85
+ $X2=0 $Y2=0
cc_621 N_A_601_345#_c_838_n N_A_288_47#_c_1330_n 0.00300039f $X=3.4 $Y=1.225
+ $X2=0 $Y2=0
cc_622 N_A_601_345#_M1019_g N_A_288_47#_c_1331_n 0.00202398f $X=3.87 $Y=1.85
+ $X2=0 $Y2=0
cc_623 N_A_601_345#_M1019_g N_A_288_47#_c_1327_n 0.0114548f $X=3.87 $Y=1.85
+ $X2=0 $Y2=0
cc_624 N_A_601_345#_c_835_n N_A_288_47#_c_1327_n 0.0117196f $X=3.795 $Y=1.225
+ $X2=0 $Y2=0
cc_625 N_A_601_345#_c_836_n N_A_288_47#_c_1327_n 0.00405971f $X=3.87 $Y=1.225
+ $X2=0 $Y2=0
cc_626 N_A_601_345#_c_837_n N_A_288_47#_c_1327_n 0.021905f $X=3.335 $Y=1.06
+ $X2=0 $Y2=0
cc_627 N_A_601_345#_c_838_n N_A_288_47#_c_1327_n 0.0454283f $X=3.4 $Y=1.225
+ $X2=0 $Y2=0
cc_628 N_A_601_345#_c_837_n N_A_288_47#_c_1328_n 0.0159402f $X=3.335 $Y=1.06
+ $X2=0 $Y2=0
cc_629 N_A_601_345#_c_839_n N_A_288_47#_c_1328_n 0.00973816f $X=3.335 $Y=0.38
+ $X2=0 $Y2=0
cc_630 N_A_601_345#_M1027_d N_A_288_47#_c_1334_n 0.00287178f $X=3.005 $Y=1.725
+ $X2=0 $Y2=0
cc_631 N_A_601_345#_c_838_n N_A_288_47#_c_1334_n 0.00945466f $X=3.4 $Y=1.225
+ $X2=0 $Y2=0
cc_632 N_A_601_345#_M1007_g N_A_873_316#_c_1463_n 0.0130074f $X=4.31 $Y=0.445
+ $X2=0 $Y2=0
cc_633 N_A_601_345#_c_837_n N_VGND_c_1620_n 0.00289962f $X=3.335 $Y=1.06 $X2=0
+ $Y2=0
cc_634 N_A_601_345#_c_839_n N_VGND_c_1620_n 0.0115629f $X=3.335 $Y=0.38 $X2=0
+ $Y2=0
cc_635 N_A_601_345#_M1007_g N_VGND_c_1621_n 0.00319988f $X=4.31 $Y=0.445 $X2=0
+ $Y2=0
cc_636 N_A_601_345#_M1007_g N_VGND_c_1628_n 0.00585385f $X=4.31 $Y=0.445 $X2=0
+ $Y2=0
cc_637 N_A_601_345#_c_839_n N_VGND_c_1628_n 0.0205768f $X=3.335 $Y=0.38 $X2=0
+ $Y2=0
cc_638 N_A_601_345#_M1009_d N_VGND_c_1637_n 0.0021994f $X=3.01 $Y=0.235 $X2=0
+ $Y2=0
cc_639 N_A_601_345#_M1007_g N_VGND_c_1637_n 0.0121029f $X=4.31 $Y=0.445 $X2=0
+ $Y2=0
cc_640 N_A_601_345#_c_839_n N_VGND_c_1637_n 0.0154649f $X=3.335 $Y=0.38 $X2=0
+ $Y2=0
cc_641 N_A1_M1000_g N_A_789_316#_c_1014_n 0.00368747f $X=5.23 $Y=2.165 $X2=0
+ $Y2=0
cc_642 N_A1_M1000_g N_VPWR_c_1180_n 0.00712348f $X=5.23 $Y=2.165 $X2=0 $Y2=0
cc_643 N_A1_M1000_g N_VPWR_c_1187_n 0.00585385f $X=5.23 $Y=2.165 $X2=0 $Y2=0
cc_644 N_A1_M1000_g N_VPWR_c_1177_n 0.00724353f $X=5.23 $Y=2.165 $X2=0 $Y2=0
cc_645 N_A1_M1000_g N_A_873_316#_c_1463_n 0.00559084f $X=5.23 $Y=2.165 $X2=0
+ $Y2=0
cc_646 N_A1_M1024_g N_A_873_316#_c_1463_n 0.00319248f $X=5.25 $Y=0.445 $X2=0
+ $Y2=0
cc_647 A1 N_A_873_316#_c_1463_n 0.0522563f $X=4.75 $Y=0.765 $X2=0 $Y2=0
cc_648 N_A1_c_904_n N_A_873_316#_c_1463_n 0.00121365f $X=5.23 $Y=1.23 $X2=0
+ $Y2=0
cc_649 N_A1_M1000_g N_A_873_316#_c_1466_n 0.0143119f $X=5.23 $Y=2.165 $X2=0
+ $Y2=0
cc_650 A1 N_A_873_316#_c_1466_n 0.0257056f $X=4.75 $Y=0.765 $X2=0 $Y2=0
cc_651 N_A1_c_904_n N_A_873_316#_c_1466_n 0.00325922f $X=5.23 $Y=1.23 $X2=0
+ $Y2=0
cc_652 N_A1_M1024_g N_A_873_316#_c_1464_n 0.00793917f $X=5.25 $Y=0.445 $X2=0
+ $Y2=0
cc_653 A1 N_A_873_316#_c_1464_n 0.0454654f $X=4.75 $Y=0.765 $X2=0 $Y2=0
cc_654 N_A1_c_904_n N_A_873_316#_c_1464_n 0.0082757f $X=5.23 $Y=1.23 $X2=0 $Y2=0
cc_655 N_A1_M1000_g N_A_873_316#_c_1468_n 0.00579011f $X=5.23 $Y=2.165 $X2=0
+ $Y2=0
cc_656 N_A1_M1000_g N_A_873_316#_c_1513_n 0.00141938f $X=5.23 $Y=2.165 $X2=0
+ $Y2=0
cc_657 N_A1_M1024_g N_A_873_316#_c_1514_n 9.53828e-19 $X=5.25 $Y=0.445 $X2=0
+ $Y2=0
cc_658 N_A1_M1024_g N_VGND_c_1621_n 0.00461751f $X=5.25 $Y=0.445 $X2=0 $Y2=0
cc_659 A1 N_VGND_c_1621_n 0.0281027f $X=4.75 $Y=0.765 $X2=0 $Y2=0
cc_660 N_A1_c_904_n N_VGND_c_1621_n 8.19449e-19 $X=5.23 $Y=1.23 $X2=0 $Y2=0
cc_661 A1 N_VGND_c_1628_n 8.41908e-19 $X=4.75 $Y=0.765 $X2=0 $Y2=0
cc_662 N_A1_M1024_g N_VGND_c_1629_n 0.00585385f $X=5.25 $Y=0.445 $X2=0 $Y2=0
cc_663 N_A1_M1024_g N_VGND_c_1637_n 0.0122213f $X=5.25 $Y=0.445 $X2=0 $Y2=0
cc_664 A1 N_VGND_c_1637_n 0.00283021f $X=4.75 $Y=0.765 $X2=0 $Y2=0
cc_665 N_A0_M1020_g N_A_789_316#_c_991_n 0.021383f $X=6.81 $Y=0.445 $X2=0 $Y2=0
cc_666 A0 N_A_789_316#_c_991_n 0.00118764f $X=6.59 $Y=0.425 $X2=0 $Y2=0
cc_667 N_A0_M1022_g N_A_789_316#_M1004_g 0.030867f $X=6.83 $Y=2.165 $X2=0 $Y2=0
cc_668 N_A0_c_943_n N_A_789_316#_c_994_n 3.12326e-19 $X=6.695 $Y=0.995 $X2=0
+ $Y2=0
cc_669 N_A0_c_944_n N_A_789_316#_c_994_n 0.0203102f $X=6.865 $Y=1.16 $X2=0 $Y2=0
cc_670 N_A0_M1022_g N_A_789_316#_c_1008_n 0.011716f $X=6.83 $Y=2.165 $X2=0 $Y2=0
cc_671 N_A0_M1022_g N_A_789_316#_c_1009_n 0.00624325f $X=6.83 $Y=2.165 $X2=0
+ $Y2=0
cc_672 N_A0_c_943_n N_A_789_316#_c_1009_n 0.00731293f $X=6.695 $Y=0.995 $X2=0
+ $Y2=0
cc_673 N_A0_c_944_n N_A_789_316#_c_1009_n 0.00219554f $X=6.865 $Y=1.16 $X2=0
+ $Y2=0
cc_674 N_A0_M1022_g N_A_789_316#_c_1010_n 0.00383803f $X=6.83 $Y=2.165 $X2=0
+ $Y2=0
cc_675 N_A0_c_943_n N_A_789_316#_c_1010_n 0.01487f $X=6.695 $Y=0.995 $X2=0 $Y2=0
cc_676 N_A0_M1022_g N_A_789_316#_c_1011_n 0.00168903f $X=6.83 $Y=2.165 $X2=0
+ $Y2=0
cc_677 N_A0_c_943_n N_A_789_316#_c_999_n 0.0260946f $X=6.695 $Y=0.995 $X2=0
+ $Y2=0
cc_678 N_A0_c_944_n N_A_789_316#_c_999_n 0.00197607f $X=6.865 $Y=1.16 $X2=0
+ $Y2=0
cc_679 N_A0_M1022_g N_A_789_316#_c_1030_n 7.65852e-19 $X=6.83 $Y=2.165 $X2=0
+ $Y2=0
cc_680 N_A0_M1022_g N_A_789_316#_c_1031_n 0.00569174f $X=6.83 $Y=2.165 $X2=0
+ $Y2=0
cc_681 N_A0_M1022_g N_VPWR_c_1181_n 0.00989024f $X=6.83 $Y=2.165 $X2=0 $Y2=0
cc_682 N_A0_M1022_g N_VPWR_c_1187_n 0.00462191f $X=6.83 $Y=2.165 $X2=0 $Y2=0
cc_683 N_A0_M1022_g N_VPWR_c_1177_n 0.00751757f $X=6.83 $Y=2.165 $X2=0 $Y2=0
cc_684 N_A0_M1022_g N_A_873_316#_c_1476_n 2.89316e-19 $X=6.83 $Y=2.165 $X2=0
+ $Y2=0
cc_685 N_A0_M1020_g N_VGND_c_1622_n 0.00886296f $X=6.81 $Y=0.445 $X2=0 $Y2=0
cc_686 A0 N_VGND_c_1622_n 0.0332811f $X=6.59 $Y=0.425 $X2=0 $Y2=0
cc_687 N_A0_M1020_g N_VGND_c_1629_n 0.00430438f $X=6.81 $Y=0.445 $X2=0 $Y2=0
cc_688 A0 N_VGND_c_1629_n 0.0109051f $X=6.59 $Y=0.425 $X2=0 $Y2=0
cc_689 N_A0_M1020_g N_VGND_c_1637_n 0.00705731f $X=6.81 $Y=0.445 $X2=0 $Y2=0
cc_690 A0 N_VGND_c_1637_n 0.0105489f $X=6.59 $Y=0.425 $X2=0 $Y2=0
cc_691 A0 A_1282_47# 0.0052103f $X=6.59 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_692 N_A_789_316#_c_1014_n N_VPWR_M1000_s 5.58164e-19 $X=6.53 $Y=2.21 $X2=0
+ $Y2=0
cc_693 N_A_789_316#_c_1009_n N_VPWR_M1022_d 0.00805037f $X=7.12 $Y=1.58 $X2=0
+ $Y2=0
cc_694 N_A_789_316#_c_998_n N_VPWR_c_1180_n 0.00185641f $X=4.1 $Y=0.51 $X2=0
+ $Y2=0
cc_695 N_A_789_316#_c_1014_n N_VPWR_c_1180_n 0.0179356f $X=6.53 $Y=2.21 $X2=0
+ $Y2=0
cc_696 N_A_789_316#_c_1015_n N_VPWR_c_1180_n 0.00275185f $X=4.52 $Y=2.21 $X2=0
+ $Y2=0
cc_697 N_A_789_316#_c_1016_n N_VPWR_c_1180_n 0.00868777f $X=4.375 $Y=2.21 $X2=0
+ $Y2=0
cc_698 N_A_789_316#_M1004_g N_VPWR_c_1181_n 0.00278284f $X=7.315 $Y=1.985 $X2=0
+ $Y2=0
cc_699 N_A_789_316#_c_1008_n N_VPWR_c_1181_n 0.0201657f $X=6.765 $Y=2.125 $X2=0
+ $Y2=0
cc_700 N_A_789_316#_c_1009_n N_VPWR_c_1181_n 0.0133801f $X=7.12 $Y=1.58 $X2=0
+ $Y2=0
cc_701 N_A_789_316#_c_1030_n N_VPWR_c_1181_n 0.00268915f $X=6.675 $Y=2.21 $X2=0
+ $Y2=0
cc_702 N_A_789_316#_c_1031_n N_VPWR_c_1181_n 0.0113595f $X=6.765 $Y=2.21 $X2=0
+ $Y2=0
cc_703 N_A_789_316#_M1008_g N_VPWR_c_1182_n 0.00987804f $X=7.735 $Y=1.985 $X2=0
+ $Y2=0
cc_704 N_A_789_316#_c_993_n N_VPWR_c_1182_n 0.00304775f $X=8.16 $Y=1.16 $X2=0
+ $Y2=0
cc_705 N_A_789_316#_M1014_g N_VPWR_c_1182_n 0.0148958f $X=8.235 $Y=1.985 $X2=0
+ $Y2=0
cc_706 N_A_789_316#_M1015_g N_VPWR_c_1182_n 9.06352e-19 $X=8.655 $Y=1.985 $X2=0
+ $Y2=0
cc_707 N_A_789_316#_M1015_g N_VPWR_c_1184_n 0.0230564f $X=8.655 $Y=1.985 $X2=0
+ $Y2=0
cc_708 N_A_789_316#_c_1014_n N_VPWR_c_1187_n 0.00322607f $X=6.53 $Y=2.21 $X2=0
+ $Y2=0
cc_709 N_A_789_316#_c_1030_n N_VPWR_c_1187_n 8.0313e-19 $X=6.675 $Y=2.21 $X2=0
+ $Y2=0
cc_710 N_A_789_316#_c_1031_n N_VPWR_c_1187_n 0.0101875f $X=6.765 $Y=2.21 $X2=0
+ $Y2=0
cc_711 N_A_789_316#_c_1012_n N_VPWR_c_1190_n 0.00647892f $X=4.185 $Y=2.21 $X2=0
+ $Y2=0
cc_712 N_A_789_316#_c_1014_n N_VPWR_c_1190_n 0.00125241f $X=6.53 $Y=2.21 $X2=0
+ $Y2=0
cc_713 N_A_789_316#_c_1015_n N_VPWR_c_1190_n 7.76522e-19 $X=4.52 $Y=2.21 $X2=0
+ $Y2=0
cc_714 N_A_789_316#_c_1016_n N_VPWR_c_1190_n 0.0111567f $X=4.375 $Y=2.21 $X2=0
+ $Y2=0
cc_715 N_A_789_316#_M1004_g N_VPWR_c_1191_n 0.00541763f $X=7.315 $Y=1.985 $X2=0
+ $Y2=0
cc_716 N_A_789_316#_M1008_g N_VPWR_c_1191_n 0.00421428f $X=7.735 $Y=1.985 $X2=0
+ $Y2=0
cc_717 N_A_789_316#_M1014_g N_VPWR_c_1192_n 0.0046653f $X=8.235 $Y=1.985 $X2=0
+ $Y2=0
cc_718 N_A_789_316#_M1015_g N_VPWR_c_1192_n 0.00428949f $X=8.655 $Y=1.985 $X2=0
+ $Y2=0
cc_719 N_A_789_316#_M1004_g N_VPWR_c_1177_n 0.00968077f $X=7.315 $Y=1.985 $X2=0
+ $Y2=0
cc_720 N_A_789_316#_M1008_g N_VPWR_c_1177_n 0.00694799f $X=7.735 $Y=1.985 $X2=0
+ $Y2=0
cc_721 N_A_789_316#_M1014_g N_VPWR_c_1177_n 0.00789179f $X=8.235 $Y=1.985 $X2=0
+ $Y2=0
cc_722 N_A_789_316#_M1015_g N_VPWR_c_1177_n 0.00798572f $X=8.655 $Y=1.985 $X2=0
+ $Y2=0
cc_723 N_A_789_316#_c_1012_n N_VPWR_c_1177_n 0.00286413f $X=4.185 $Y=2.21 $X2=0
+ $Y2=0
cc_724 N_A_789_316#_c_1014_n N_VPWR_c_1177_n 0.17108f $X=6.53 $Y=2.21 $X2=0
+ $Y2=0
cc_725 N_A_789_316#_c_1015_n N_VPWR_c_1177_n 0.0297601f $X=4.52 $Y=2.21 $X2=0
+ $Y2=0
cc_726 N_A_789_316#_c_1016_n N_VPWR_c_1177_n 0.00197276f $X=4.375 $Y=2.21 $X2=0
+ $Y2=0
cc_727 N_A_789_316#_c_1030_n N_VPWR_c_1177_n 0.0297101f $X=6.675 $Y=2.21 $X2=0
+ $Y2=0
cc_728 N_A_789_316#_c_1031_n N_VPWR_c_1177_n 0.00215271f $X=6.765 $Y=2.21 $X2=0
+ $Y2=0
cc_729 N_A_789_316#_c_1012_n N_A_288_47#_c_1330_n 0.0131455f $X=4.185 $Y=2.21
+ $X2=0 $Y2=0
cc_730 N_A_789_316#_c_1015_n N_A_288_47#_c_1330_n 7.53591e-19 $X=4.52 $Y=2.21
+ $X2=0 $Y2=0
cc_731 N_A_789_316#_c_998_n N_A_288_47#_c_1328_n 0.0987706f $X=4.1 $Y=0.51 $X2=0
+ $Y2=0
cc_732 N_A_789_316#_c_1012_n N_A_288_47#_c_1335_n 8.20074e-19 $X=4.185 $Y=2.21
+ $X2=0 $Y2=0
cc_733 N_A_789_316#_c_1015_n N_A_873_316#_M1013_d 0.00107375f $X=4.52 $Y=2.21
+ $X2=0 $Y2=0
cc_734 N_A_789_316#_c_1014_n N_A_873_316#_M1023_d 0.00299297f $X=6.53 $Y=2.21
+ $X2=0 $Y2=0
cc_735 N_A_789_316#_c_998_n N_A_873_316#_c_1463_n 0.0611274f $X=4.1 $Y=0.51
+ $X2=0 $Y2=0
cc_736 N_A_789_316#_c_1014_n N_A_873_316#_c_1463_n 4.40444e-19 $X=6.53 $Y=2.21
+ $X2=0 $Y2=0
cc_737 N_A_789_316#_c_1015_n N_A_873_316#_c_1463_n 3.97141e-19 $X=4.52 $Y=2.21
+ $X2=0 $Y2=0
cc_738 N_A_789_316#_c_1016_n N_A_873_316#_c_1463_n 0.00600827f $X=4.375 $Y=2.21
+ $X2=0 $Y2=0
cc_739 N_A_789_316#_c_1014_n N_A_873_316#_c_1468_n 0.00351097f $X=6.53 $Y=2.21
+ $X2=0 $Y2=0
cc_740 N_A_789_316#_c_1014_n N_A_873_316#_c_1513_n 0.00522075f $X=6.53 $Y=2.21
+ $X2=0 $Y2=0
cc_741 N_A_789_316#_c_1014_n N_A_873_316#_c_1476_n 0.0249706f $X=6.53 $Y=2.21
+ $X2=0 $Y2=0
cc_742 N_A_789_316#_c_1030_n N_A_873_316#_c_1476_n 0.00153799f $X=6.675 $Y=2.21
+ $X2=0 $Y2=0
cc_743 N_A_789_316#_c_1031_n N_A_873_316#_c_1476_n 0.0062331f $X=6.765 $Y=2.21
+ $X2=0 $Y2=0
cc_744 N_A_789_316#_c_1014_n A_1061_369# 0.00249485f $X=6.53 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_745 N_A_789_316#_c_1008_n A_1280_413# 0.00367035f $X=6.765 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_746 N_A_789_316#_c_1014_n A_1280_413# 0.00278888f $X=6.53 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_747 N_A_789_316#_c_1030_n A_1280_413# 0.00833367f $X=6.675 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_748 N_A_789_316#_c_1031_n A_1280_413# 0.00590254f $X=6.765 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_749 N_A_789_316#_M1004_g N_X_c_1565_n 0.00297963f $X=7.315 $Y=1.985 $X2=0
+ $Y2=0
cc_750 N_A_789_316#_M1008_g N_X_c_1565_n 0.00375653f $X=7.735 $Y=1.985 $X2=0
+ $Y2=0
cc_751 N_A_789_316#_c_994_n N_X_c_1565_n 0.00399972f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_752 N_A_789_316#_c_1009_n N_X_c_1565_n 0.0137876f $X=7.12 $Y=1.58 $X2=0 $Y2=0
cc_753 N_A_789_316#_c_991_n N_X_c_1561_n 0.00403664f $X=7.315 $Y=0.995 $X2=0
+ $Y2=0
cc_754 N_A_789_316#_c_992_n N_X_c_1561_n 0.00698416f $X=7.735 $Y=0.995 $X2=0
+ $Y2=0
cc_755 N_A_789_316#_c_994_n N_X_c_1561_n 0.00381421f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_756 N_A_789_316#_c_995_n N_X_c_1561_n 3.91723e-19 $X=8.235 $Y=0.995 $X2=0
+ $Y2=0
cc_757 N_A_789_316#_c_999_n N_X_c_1561_n 0.00489457f $X=7.345 $Y=1.16 $X2=0
+ $Y2=0
cc_758 N_A_789_316#_c_993_n N_X_c_1574_n 0.02343f $X=8.16 $Y=1.16 $X2=0 $Y2=0
cc_759 N_A_789_316#_c_994_n N_X_c_1574_n 0.00446442f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_760 N_A_789_316#_c_997_n N_X_c_1574_n 0.0209498f $X=8.655 $Y=1.16 $X2=0 $Y2=0
cc_761 N_A_789_316#_M1004_g N_X_c_1577_n 0.00750243f $X=7.315 $Y=1.985 $X2=0
+ $Y2=0
cc_762 N_A_789_316#_M1008_g N_X_c_1577_n 0.0107776f $X=7.735 $Y=1.985 $X2=0
+ $Y2=0
cc_763 N_A_789_316#_c_999_n N_X_c_1577_n 0.00153049f $X=7.345 $Y=1.16 $X2=0
+ $Y2=0
cc_764 N_A_789_316#_M1008_g N_X_c_1580_n 0.00351969f $X=7.735 $Y=1.985 $X2=0
+ $Y2=0
cc_765 N_A_789_316#_c_1008_n N_X_c_1580_n 0.00454339f $X=6.765 $Y=2.125 $X2=0
+ $Y2=0
cc_766 N_A_789_316#_c_992_n N_X_c_1582_n 0.00948419f $X=7.735 $Y=0.995 $X2=0
+ $Y2=0
cc_767 N_A_789_316#_c_994_n N_X_c_1582_n 0.00339791f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_768 N_A_789_316#_M1004_g N_X_c_1563_n 0.00109594f $X=7.315 $Y=1.985 $X2=0
+ $Y2=0
cc_769 N_A_789_316#_M1008_g N_X_c_1563_n 0.00488658f $X=7.735 $Y=1.985 $X2=0
+ $Y2=0
cc_770 N_A_789_316#_c_994_n N_X_c_1563_n 0.00104072f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_771 N_A_789_316#_M1014_g N_X_c_1563_n 5.83519e-19 $X=8.235 $Y=1.985 $X2=0
+ $Y2=0
cc_772 N_A_789_316#_c_1011_n N_X_c_1563_n 0.00769733f $X=7.205 $Y=1.495 $X2=0
+ $Y2=0
cc_773 N_A_789_316#_c_999_n N_X_c_1563_n 0.0013231f $X=7.345 $Y=1.16 $X2=0 $Y2=0
cc_774 N_A_789_316#_c_994_n N_X_c_1590_n 0.0071976f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_775 N_A_789_316#_c_999_n N_X_c_1590_n 0.0191717f $X=7.345 $Y=1.16 $X2=0 $Y2=0
cc_776 N_A_789_316#_c_995_n X 0.00242114f $X=8.235 $Y=0.995 $X2=0 $Y2=0
cc_777 N_A_789_316#_c_996_n X 0.019213f $X=8.655 $Y=0.995 $X2=0 $Y2=0
cc_778 N_A_789_316#_c_997_n X 0.00889892f $X=8.655 $Y=1.16 $X2=0 $Y2=0
cc_779 N_A_789_316#_c_997_n X 0.0178209f $X=8.655 $Y=1.16 $X2=0 $Y2=0
cc_780 N_A_789_316#_M1014_g X 0.00313845f $X=8.235 $Y=1.985 $X2=0 $Y2=0
cc_781 N_A_789_316#_M1015_g X 0.0281322f $X=8.655 $Y=1.985 $X2=0 $Y2=0
cc_782 N_A_789_316#_c_997_n X 0.00405549f $X=8.655 $Y=1.16 $X2=0 $Y2=0
cc_783 N_A_789_316#_c_991_n N_VGND_c_1622_n 0.0129978f $X=7.315 $Y=0.995 $X2=0
+ $Y2=0
cc_784 N_A_789_316#_c_992_n N_VGND_c_1622_n 8.34622e-19 $X=7.735 $Y=0.995 $X2=0
+ $Y2=0
cc_785 N_A_789_316#_c_999_n N_VGND_c_1622_n 0.00961319f $X=7.345 $Y=1.16 $X2=0
+ $Y2=0
cc_786 N_A_789_316#_c_992_n N_VGND_c_1623_n 0.0060234f $X=7.735 $Y=0.995 $X2=0
+ $Y2=0
cc_787 N_A_789_316#_c_993_n N_VGND_c_1623_n 0.00325586f $X=8.16 $Y=1.16 $X2=0
+ $Y2=0
cc_788 N_A_789_316#_c_995_n N_VGND_c_1623_n 0.0113378f $X=8.235 $Y=0.995 $X2=0
+ $Y2=0
cc_789 N_A_789_316#_c_996_n N_VGND_c_1623_n 8.61839e-19 $X=8.655 $Y=0.995 $X2=0
+ $Y2=0
cc_790 N_A_789_316#_c_996_n N_VGND_c_1625_n 0.0161314f $X=8.655 $Y=0.995 $X2=0
+ $Y2=0
cc_791 N_A_789_316#_c_998_n N_VGND_c_1628_n 0.0077748f $X=4.1 $Y=0.51 $X2=0
+ $Y2=0
cc_792 N_A_789_316#_c_991_n N_VGND_c_1630_n 0.0046653f $X=7.315 $Y=0.995 $X2=0
+ $Y2=0
cc_793 N_A_789_316#_c_992_n N_VGND_c_1630_n 0.00420076f $X=7.735 $Y=0.995 $X2=0
+ $Y2=0
cc_794 N_A_789_316#_c_995_n N_VGND_c_1631_n 0.0046653f $X=8.235 $Y=0.995 $X2=0
+ $Y2=0
cc_795 N_A_789_316#_c_996_n N_VGND_c_1631_n 0.00428949f $X=8.655 $Y=0.995 $X2=0
+ $Y2=0
cc_796 N_A_789_316#_M1012_d N_VGND_c_1637_n 0.0052901f $X=3.96 $Y=0.235 $X2=0
+ $Y2=0
cc_797 N_A_789_316#_c_991_n N_VGND_c_1637_n 0.00796766f $X=7.315 $Y=0.995 $X2=0
+ $Y2=0
cc_798 N_A_789_316#_c_992_n N_VGND_c_1637_n 0.00694102f $X=7.735 $Y=0.995 $X2=0
+ $Y2=0
cc_799 N_A_789_316#_c_995_n N_VGND_c_1637_n 0.00796766f $X=8.235 $Y=0.995 $X2=0
+ $Y2=0
cc_800 N_A_789_316#_c_996_n N_VGND_c_1637_n 0.00802461f $X=8.655 $Y=0.995 $X2=0
+ $Y2=0
cc_801 N_A_789_316#_c_998_n N_VGND_c_1637_n 0.00690003f $X=4.1 $Y=0.51 $X2=0
+ $Y2=0
cc_802 N_VPWR_c_1177_n A_193_369# 0.00448763f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_803 N_VPWR_c_1177_n N_A_288_47#_M1025_d 0.00192946f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_804 N_VPWR_c_1178_n N_A_288_47#_c_1337_n 0.00114558f $X=0.68 $Y=2.34 $X2=0
+ $Y2=0
cc_805 N_VPWR_c_1185_n N_A_288_47#_c_1337_n 0.0180901f $X=2.6 $Y=2.72 $X2=0
+ $Y2=0
cc_806 N_VPWR_c_1177_n N_A_288_47#_c_1337_n 0.00858407f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_807 N_VPWR_c_1179_n N_A_288_47#_c_1329_n 0.00423173f $X=2.72 $Y=2.22 $X2=0
+ $Y2=0
cc_808 N_VPWR_c_1185_n N_A_288_47#_c_1329_n 0.00582929f $X=2.6 $Y=2.72 $X2=0
+ $Y2=0
cc_809 N_VPWR_c_1177_n N_A_288_47#_c_1329_n 8.66284e-19 $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_810 N_VPWR_c_1179_n N_A_288_47#_c_1330_n 0.00289411f $X=2.72 $Y=2.22 $X2=0
+ $Y2=0
cc_811 N_VPWR_c_1190_n N_A_288_47#_c_1330_n 0.0172466f $X=4.76 $Y=2.72 $X2=0
+ $Y2=0
cc_812 N_VPWR_c_1177_n N_A_288_47#_c_1330_n 0.00412848f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_813 N_VPWR_M1002_d N_A_288_47#_c_1334_n 5.30843e-19 $X=2.585 $Y=1.725 $X2=0
+ $Y2=0
cc_814 N_VPWR_c_1179_n N_A_288_47#_c_1334_n 0.014737f $X=2.72 $Y=2.22 $X2=0
+ $Y2=0
cc_815 N_VPWR_c_1185_n N_A_288_47#_c_1334_n 0.00180834f $X=2.6 $Y=2.72 $X2=0
+ $Y2=0
cc_816 N_VPWR_c_1190_n N_A_288_47#_c_1334_n 0.00243737f $X=4.76 $Y=2.72 $X2=0
+ $Y2=0
cc_817 N_VPWR_c_1177_n N_A_288_47#_c_1334_n 0.093852f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_818 N_VPWR_c_1179_n N_A_288_47#_c_1374_n 0.00163392f $X=2.72 $Y=2.22 $X2=0
+ $Y2=0
cc_819 N_VPWR_c_1185_n N_A_288_47#_c_1374_n 8.27583e-19 $X=2.6 $Y=2.72 $X2=0
+ $Y2=0
cc_820 N_VPWR_c_1177_n N_A_288_47#_c_1374_n 0.0298306f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_821 N_VPWR_c_1179_n N_A_288_47#_c_1335_n 0.00250319f $X=2.72 $Y=2.22 $X2=0
+ $Y2=0
cc_822 N_VPWR_c_1190_n N_A_288_47#_c_1335_n 8.27838e-19 $X=4.76 $Y=2.72 $X2=0
+ $Y2=0
cc_823 N_VPWR_c_1177_n N_A_288_47#_c_1335_n 0.0296902f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_824 N_VPWR_c_1177_n A_373_413# 0.00300836f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_825 N_VPWR_c_1177_n N_A_873_316#_M1023_d 0.00130544f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_826 N_VPWR_c_1180_n N_A_873_316#_c_1466_n 0.0125871f $X=5.02 $Y=2.17 $X2=0
+ $Y2=0
cc_827 N_VPWR_c_1180_n N_A_873_316#_c_1468_n 3.9298e-19 $X=5.02 $Y=2.17 $X2=0
+ $Y2=0
cc_828 N_VPWR_c_1180_n N_A_873_316#_c_1513_n 0.00347614f $X=5.02 $Y=2.17 $X2=0
+ $Y2=0
cc_829 N_VPWR_c_1187_n N_A_873_316#_c_1513_n 0.00567337f $X=7.02 $Y=2.72 $X2=0
+ $Y2=0
cc_830 N_VPWR_c_1177_n N_A_873_316#_c_1513_n 0.00186252f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_831 N_VPWR_c_1187_n N_A_873_316#_c_1476_n 0.0233641f $X=7.02 $Y=2.72 $X2=0
+ $Y2=0
cc_832 N_VPWR_c_1177_n N_A_873_316#_c_1476_n 0.00706654f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_833 N_VPWR_c_1177_n A_1061_369# 0.00267305f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_834 N_VPWR_c_1177_n A_1280_413# 0.00221859f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_835 N_VPWR_c_1177_n N_X_M1004_s 0.00215535f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_836 N_VPWR_c_1177_n N_X_M1014_s 0.00389051f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_837 N_VPWR_c_1182_n N_X_c_1565_n 0.0735075f $X=8.025 $Y=1.66 $X2=0 $Y2=0
cc_838 N_VPWR_c_1182_n N_X_c_1574_n 0.0158777f $X=8.025 $Y=1.66 $X2=0 $Y2=0
cc_839 N_VPWR_c_1191_n N_X_c_1577_n 0.0228123f $X=7.94 $Y=2.72 $X2=0 $Y2=0
cc_840 N_VPWR_c_1177_n N_X_c_1577_n 0.0148391f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_841 N_VPWR_c_1184_n X 0.0728724f $X=8.94 $Y=1.66 $X2=0 $Y2=0
cc_842 N_VPWR_c_1192_n X 0.0190418f $X=8.855 $Y=2.72 $X2=0 $Y2=0
cc_843 N_VPWR_c_1177_n X 0.0118297f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_844 N_VPWR_c_1184_n N_VGND_c_1625_n 0.0086927f $X=8.94 $Y=1.66 $X2=0 $Y2=0
cc_845 N_A_288_47#_c_1337_n A_373_413# 0.0041168f $X=2.075 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_846 N_A_288_47#_c_1329_n A_373_413# 0.0134763f $X=2.16 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_847 N_A_288_47#_c_1334_n A_373_413# 0.00266219f $X=3.31 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_848 N_A_288_47#_c_1374_n A_373_413# 0.00398835f $X=2.22 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_849 N_A_288_47#_c_1338_n N_VGND_c_1620_n 0.00748073f $X=1.905 $Y=0.45 $X2=0
+ $Y2=0
cc_850 N_A_288_47#_c_1325_n N_VGND_c_1620_n 3.77264e-19 $X=1.99 $Y=1.235 $X2=0
+ $Y2=0
cc_851 N_A_288_47#_c_1338_n N_VGND_c_1627_n 0.020375f $X=1.905 $Y=0.45 $X2=0
+ $Y2=0
cc_852 N_A_288_47#_c_1328_n N_VGND_c_1628_n 0.00895969f $X=3.675 $Y=0.51 $X2=0
+ $Y2=0
cc_853 N_A_288_47#_M1006_d N_VGND_c_1637_n 0.00354687f $X=1.44 $Y=0.235 $X2=0
+ $Y2=0
cc_854 N_A_288_47#_M1012_s N_VGND_c_1637_n 0.00264447f $X=3.55 $Y=0.235 $X2=0
+ $Y2=0
cc_855 N_A_288_47#_c_1338_n N_VGND_c_1637_n 0.0203474f $X=1.905 $Y=0.45 $X2=0
+ $Y2=0
cc_856 N_A_288_47#_c_1328_n N_VGND_c_1637_n 0.00841871f $X=3.675 $Y=0.51 $X2=0
+ $Y2=0
cc_857 N_A_288_47#_c_1338_n A_398_47# 0.00244815f $X=1.905 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_858 N_A_288_47#_c_1325_n A_398_47# 0.00145797f $X=1.99 $Y=1.235 $X2=-0.19
+ $Y2=-0.24
cc_859 N_A_873_316#_c_1468_n A_1061_369# 0.00496775f $X=5.415 $Y=2.155 $X2=-0.19
+ $Y2=-0.24
cc_860 N_A_873_316#_c_1513_n A_1061_369# 0.00306462f $X=5.5 $Y=2.24 $X2=-0.19
+ $Y2=-0.24
cc_861 N_A_873_316#_c_1476_n A_1061_369# 0.00812168f $X=6.115 $Y=2.24 $X2=-0.19
+ $Y2=-0.24
cc_862 N_A_873_316#_c_1514_n N_VGND_c_1621_n 0.0207476f $X=4.52 $Y=0.42 $X2=0
+ $Y2=0
cc_863 N_A_873_316#_c_1514_n N_VGND_c_1628_n 0.0127262f $X=4.52 $Y=0.42 $X2=0
+ $Y2=0
cc_864 N_A_873_316#_c_1540_p N_VGND_c_1629_n 0.0080925f $X=5.5 $Y=0.38 $X2=0
+ $Y2=0
cc_865 N_A_873_316#_c_1475_n N_VGND_c_1629_n 0.0333963f $X=6.06 $Y=0.38 $X2=0
+ $Y2=0
cc_866 N_A_873_316#_M1007_d N_VGND_c_1637_n 0.00403727f $X=4.385 $Y=0.235 $X2=0
+ $Y2=0
cc_867 N_A_873_316#_M1010_d N_VGND_c_1637_n 0.00340843f $X=5.86 $Y=0.235 $X2=0
+ $Y2=0
cc_868 N_A_873_316#_c_1540_p N_VGND_c_1637_n 0.00641762f $X=5.5 $Y=0.38 $X2=0
+ $Y2=0
cc_869 N_A_873_316#_c_1475_n N_VGND_c_1637_n 0.0256442f $X=6.06 $Y=0.38 $X2=0
+ $Y2=0
cc_870 N_A_873_316#_c_1514_n N_VGND_c_1637_n 0.00779458f $X=4.52 $Y=0.42 $X2=0
+ $Y2=0
cc_871 N_A_873_316#_c_1464_n A_1065_47# 0.00347944f $X=5.415 $Y=1.565 $X2=-0.19
+ $Y2=-0.24
cc_872 N_A_873_316#_c_1540_p A_1065_47# 0.00236827f $X=5.5 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_873 N_A_873_316#_c_1475_n A_1065_47# 0.00762432f $X=6.06 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_874 N_X_c_1561_n N_VGND_c_1622_n 0.00390889f $X=7.685 $Y=1.065 $X2=0 $Y2=0
cc_875 N_X_c_1561_n N_VGND_c_1623_n 0.0115783f $X=7.685 $Y=1.065 $X2=0 $Y2=0
cc_876 N_X_c_1574_n N_VGND_c_1623_n 0.0165613f $X=8.36 $Y=1.185 $X2=0 $Y2=0
cc_877 N_X_c_1582_n N_VGND_c_1623_n 0.0349816f $X=7.685 $Y=0.495 $X2=0 $Y2=0
cc_878 X N_VGND_c_1625_n 0.0470634f $X=8.43 $Y=0.425 $X2=0 $Y2=0
cc_879 N_X_c_1582_n N_VGND_c_1630_n 0.0188909f $X=7.685 $Y=0.495 $X2=0 $Y2=0
cc_880 X N_VGND_c_1631_n 0.0190723f $X=8.43 $Y=0.425 $X2=0 $Y2=0
cc_881 N_X_M1003_s N_VGND_c_1637_n 0.00390695f $X=7.39 $Y=0.235 $X2=0 $Y2=0
cc_882 N_X_M1011_s N_VGND_c_1637_n 0.0039413f $X=8.31 $Y=0.235 $X2=0 $Y2=0
cc_883 N_X_c_1582_n N_VGND_c_1637_n 0.0120046f $X=7.685 $Y=0.495 $X2=0 $Y2=0
cc_884 X N_VGND_c_1637_n 0.0119018f $X=8.43 $Y=0.425 $X2=0 $Y2=0
cc_885 N_VGND_c_1637_n A_193_47# 0.00482635f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_886 N_VGND_c_1637_n A_398_47# 0.0089813f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_887 N_VGND_c_1637_n A_1065_47# 0.00329874f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_888 N_VGND_c_1637_n A_1282_47# 0.00726162f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a41o_2.spice.pex
* Created: Thu Aug 27 14:06:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A41O_2%A_79_21# 1 2 3 10 12 15 17 19 22 27 28 29 30
+ 31 32 35 39 41 45 47 49
c101 27 0 1.51504e-19 $X=1.065 $Y=1.16
r102 50 52 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r103 45 47 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=2.545 $Y=0.38
+ $X2=3.88 $Y2=0.38
r104 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=0.465
+ $X2=2.545 $Y2=0.38
r105 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.46 $Y=0.465
+ $X2=2.46 $Y2=0.635
r106 42 49 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.705 $Y=0.72
+ $X2=1.6 $Y2=0.72
r107 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=0.72
+ $X2=2.46 $Y2=0.635
r108 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.375 $Y=0.72
+ $X2=1.705 $Y2=0.72
r109 37 49 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=0.635
+ $X2=1.6 $Y2=0.72
r110 37 39 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.6 $Y=0.635
+ $X2=1.6 $Y2=0.42
r111 33 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=2
r112 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.62 $Y2=1.665
r113 31 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.15 $Y2=1.58
r114 29 49 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.495 $Y=0.72
+ $X2=1.6 $Y2=0.72
r115 29 30 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.495 $Y=0.72
+ $X2=1.15 $Y2=0.72
r116 28 52 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.065 $Y=1.16
+ $X2=0.89 $Y2=1.16
r117 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.065
+ $Y=1.16 $X2=1.065 $Y2=1.16
r118 25 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=1.495
+ $X2=1.15 $Y2=1.58
r119 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.065 $Y=1.495
+ $X2=1.065 $Y2=1.16
r120 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=0.805
+ $X2=1.15 $Y2=0.72
r121 24 27 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.065 $Y=0.805
+ $X2=1.065 $Y2=1.16
r122 20 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r123 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r124 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r125 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r126 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r127 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r128 10 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r129 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r130 3 35 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.485 $X2=1.62 $Y2=2
r131 2 47 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.38
r132 1 39 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%B1 1 3 6 8 14
c32 8 0 1.78912e-19 $X=1.635 $Y=1.19
r33 11 14 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.565 $Y=1.16
+ $X2=1.83 $Y2=1.16
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.16 $X2=1.565 $Y2=1.16
r35 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.16
r36 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.325 $X2=1.83
+ $Y2=1.985
r37 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.995 $X2=1.83
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%A4 1 3 6 8 9 13 14
c37 13 0 2.0811e-19 $X=2.25 $Y=1.16
c38 6 0 1.22839e-19 $X=2.25 $Y=1.985
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r40 8 9 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.167 $Y=1.19
+ $X2=2.167 $Y2=1.53
r41 8 14 1.03204 $w=3.33e-07 $l=3e-08 $layer=LI1_cond $X=2.167 $Y=1.19 $X2=2.167
+ $Y2=1.16
r42 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.325
+ $X2=2.25 $Y2=1.16
r43 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.25 $Y=1.325 $X2=2.25
+ $Y2=1.985
r44 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=0.995
+ $X2=2.25 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.25 $Y=0.995 $X2=2.25
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%A3 3 6 10 11 13 16
c41 10 0 1.22839e-19 $X=2.77 $Y=1.16
r42 13 18 12.8421 $w=1.88e-07 $l=2.2e-07 $layer=LI1_cond $X=2.99 $Y=1.53
+ $X2=2.77 $Y2=1.53
r43 11 17 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.75 $Y2=1.325
r44 11 16 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.75 $Y2=0.995
r45 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.16 $X2=2.77 $Y2=1.16
r46 8 18 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.77 $Y=1.435 $X2=2.77
+ $Y2=1.53
r47 8 10 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.77 $Y=1.435
+ $X2=2.77 $Y2=1.16
r48 6 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.67 $Y=1.985
+ $X2=2.67 $Y2=1.325
r49 3 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.56 $X2=2.67
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%A2 1 3 6 8 9 10 16
r41 17 18 12.5262 $w=1.68e-07 $l=1.92e-07 $layer=LI1_cond $X=3.25 $Y=1.16
+ $X2=3.442 $Y2=1.16
r42 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.16 $X2=3.25 $Y2=1.16
r43 9 18 0.195722 $w=1.68e-07 $l=3e-09 $layer=LI1_cond $X=3.445 $Y=1.16
+ $X2=3.442 $Y2=1.16
r44 9 10 14.4725 $w=2.13e-07 $l=2.7e-07 $layer=LI1_cond $X=3.442 $Y=1.26
+ $X2=3.442 $Y2=1.53
r45 9 18 0.80403 $w=2.13e-07 $l=1.5e-08 $layer=LI1_cond $X=3.442 $Y=1.26
+ $X2=3.442 $Y2=1.245
r46 8 18 12.0604 $w=2.13e-07 $l=2.25e-07 $layer=LI1_cond $X=3.442 $Y=0.85
+ $X2=3.442 $Y2=1.075
r47 4 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.325
+ $X2=3.25 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.25 $Y=1.325 $X2=3.25
+ $Y2=1.985
r49 1 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.25 $Y=0.995 $X2=3.25
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%A1 1 3 6 8 9 10 17
r27 14 17 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=3.67 $Y=1.16 $X2=3.87
+ $Y2=1.16
r28 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.895 $Y=1.16
+ $X2=3.895 $Y2=1.53
r29 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.87
+ $Y=1.16 $X2=3.87 $Y2=1.16
r30 8 9 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=3.895 $Y=0.85 $X2=3.895
+ $Y2=1.16
r31 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r32 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.325 $X2=3.67
+ $Y2=1.985
r33 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.67 $Y=0.995 $X2=3.67
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%VPWR 1 2 3 4 13 15 21 25 29 32 33 34 36 45 51
+ 52 58 61
c68 2 0 1.51504e-19 $X=0.965 $Y=1.485
r69 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 52 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 49 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.46 $Y2=2.72
r74 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 48 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r76 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 45 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=3.46 $Y2=2.72
r78 45 47 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 44 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r80 44 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r81 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r82 41 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.14 $Y2=2.72
r83 41 43 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=2.07 $Y2=2.72
r84 40 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 37 55 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r87 37 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 36 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.14 $Y2=2.72
r89 36 39 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 34 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 34 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r92 32 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r93 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.46 $Y2=2.72
r94 31 47 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.585 $Y=2.72
+ $X2=2.99 $Y2=2.72
r95 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.585 $Y=2.72
+ $X2=2.46 $Y2=2.72
r96 27 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=2.635
+ $X2=3.46 $Y2=2.72
r97 27 29 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.46 $Y=2.635
+ $X2=3.46 $Y2=2.34
r98 23 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.72
r99 23 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.34
r100 19 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.72
r101 19 21 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2
r102 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r103 13 55 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r104 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r105 4 29 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=1.485 $X2=3.46 $Y2=2.34
r106 3 25 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.34
r107 2 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r108 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r109 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%X 1 2 9 11 12 13 14 15 24
r15 15 33 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=2.21
+ $X2=0.69 $Y2=1.96
r16 14 33 5.25359 $w=1.88e-07 $l=9e-08 $layer=LI1_cond $X=0.69 $Y=1.87 $X2=0.69
+ $Y2=1.96
r17 13 14 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.69 $Y=1.53
+ $X2=0.69 $Y2=1.87
r18 12 13 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.69 $Y=1.19
+ $X2=0.69 $Y2=1.53
r19 11 24 2.51005 $w=1.88e-07 $l=4.3e-08 $layer=LI1_cond $X=0.69 $Y=0.807
+ $X2=0.69 $Y2=0.85
r20 11 38 3.1836 $w=1.88e-07 $l=5.2e-08 $layer=LI1_cond $X=0.69 $Y=0.807
+ $X2=0.69 $Y2=0.755
r21 11 12 17.3952 $w=1.88e-07 $l=2.98e-07 $layer=LI1_cond $X=0.69 $Y=0.892
+ $X2=0.69 $Y2=1.19
r22 11 24 2.45167 $w=1.88e-07 $l=4.2e-08 $layer=LI1_cond $X=0.69 $Y=0.892
+ $X2=0.69 $Y2=0.85
r23 9 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.46 $X2=0.68
+ $Y2=0.755
r24 2 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
r25 1 9 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%A_381_297# 1 2 3 12 16 21 23 25
c37 21 0 2.91989e-20 $X=2.04 $Y=1.96
r38 17 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=1.88
+ $X2=2.88 $Y2=1.88
r39 16 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=1.88
+ $X2=3.88 $Y2=1.88
r40 16 17 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.795 $Y=1.88
+ $X2=2.965 $Y2=1.88
r41 13 21 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=1.88
+ $X2=2.04 $Y2=1.88
r42 12 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=1.88
+ $X2=2.88 $Y2=1.88
r43 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.795 $Y=1.88
+ $X2=2.125 $Y2=1.88
r44 3 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=1.96
r45 2 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.96
r46 1 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r62 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r63 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r64 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r65 37 40 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r66 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r67 36 39 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r68 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r69 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r70 34 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.53
+ $Y2=0
r71 33 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r72 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r73 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r75 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r76 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r77 29 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.61
+ $Y2=0
r78 28 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r79 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r80 25 43 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r81 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r82 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r83 24 27 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r84 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r85 22 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r86 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r87 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.38
r88 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r89 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r90 10 43 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r91 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r92 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.38
r93 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r94 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


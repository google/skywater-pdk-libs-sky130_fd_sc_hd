# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o21bai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645000 1.075000 6.810000 1.285000 ;
        RECT 6.585000 1.285000 6.810000 2.455000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.065000 1.075000 4.475000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.555000 1.285000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.455000 4.315000 1.625000 ;
        RECT 1.065000 1.625000 1.275000 2.465000 ;
        RECT 1.420000 0.645000 2.675000 0.815000 ;
        RECT 1.865000 1.625000 2.115000 2.465000 ;
        RECT 2.445000 0.815000 2.675000 1.075000 ;
        RECT 2.445000 1.075000 2.895000 1.445000 ;
        RECT 2.445000 1.445000 4.315000 1.455000 ;
        RECT 3.225000 1.625000 3.475000 2.125000 ;
        RECT 4.065000 1.625000 4.315000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.900000 0.085000 ;
        RECT 0.225000  0.085000 0.395000 0.895000 ;
        RECT 3.265000  0.085000 3.435000 0.555000 ;
        RECT 4.105000  0.085000 4.275000 0.555000 ;
        RECT 4.945000  0.085000 5.115000 0.555000 ;
        RECT 5.785000  0.085000 5.955000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.900000 2.805000 ;
        RECT 0.645000 1.795000 0.855000 2.635000 ;
        RECT 1.445000 1.795000 1.695000 2.635000 ;
        RECT 2.285000 1.795000 2.535000 2.635000 ;
        RECT 4.905000 1.795000 5.155000 2.635000 ;
        RECT 5.745000 1.795000 5.995000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.145000 1.455000 0.895000 1.625000 ;
      RECT 0.145000 1.625000 0.475000 2.435000 ;
      RECT 0.565000 0.290000 0.895000 0.895000 ;
      RECT 0.725000 0.895000 0.895000 1.075000 ;
      RECT 0.725000 1.075000 2.275000 1.285000 ;
      RECT 0.725000 1.285000 0.895000 1.455000 ;
      RECT 1.080000 0.305000 3.095000 0.475000 ;
      RECT 2.775000 1.795000 3.055000 2.295000 ;
      RECT 2.775000 2.295000 4.735000 2.465000 ;
      RECT 2.845000 0.475000 3.095000 0.725000 ;
      RECT 2.845000 0.725000 6.455000 0.905000 ;
      RECT 3.605000 0.255000 3.935000 0.725000 ;
      RECT 3.645000 1.795000 3.895000 2.295000 ;
      RECT 4.445000 0.255000 4.775000 0.725000 ;
      RECT 4.485000 1.455000 6.415000 1.625000 ;
      RECT 4.485000 1.625000 4.735000 2.295000 ;
      RECT 5.285000 0.255000 5.615000 0.725000 ;
      RECT 5.325000 1.625000 5.575000 2.465000 ;
      RECT 6.125000 0.255000 6.455000 0.725000 ;
      RECT 6.165000 1.625000 6.415000 2.465000 ;
  END
END sky130_fd_sc_hd__o21bai_4
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nshort w=650000u l=150000u
+  ad=5.97e+11p pd=5.79e+06u as=3.51e+11p ps=3.68e+06u
M1001 VGND C Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_245_297# C a_161_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u
M1004 VPWR A a_341_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.915e+11p pd=2.67e+06u as=2.7e+11p ps=2.54e+06u
M1005 a_161_297# a_91_199# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.2e+11p ps=3.04e+06u
M1006 Y a_91_199# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_91_199# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1008 a_341_297# B a_245_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_91_199# D_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__nand2b_2.pex.spice
* Created: Thu Aug 27 14:29:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND2B_2%A_N 3 6 8 11 13
r29 11 14 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.16
+ $X2=0.535 $Y2=1.325
r30 11 13 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.16
+ $X2=0.535 $Y2=0.995
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.16 $X2=0.54 $Y2=1.16
r32 8 12 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.54 $Y2=1.16
r33 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.695
+ $X2=0.47 $Y2=1.325
r34 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_2%A_27_93# 1 2 9 13 17 21 23 24 27 30 31 35
+ 39 46
c66 35 0 1.04593e-19 $X=1.195 $Y=1.16
c67 27 0 1.63453e-19 $X=1.9 $Y=1.16
c68 21 0 1.56255e-19 $X=1.9 $Y=0.56
r69 45 46 8.0507 $w=3.63e-07 $l=1.5e-07 $layer=LI1_cond $X=0.26 $Y=1.677
+ $X2=0.41 $Y2=1.677
r70 39 41 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.227 $Y=0.675
+ $X2=0.227 $Y2=0.84
r71 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.16 $X2=1.195 $Y2=1.16
r72 33 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.195 $Y=1.495
+ $X2=1.195 $Y2=1.16
r73 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.03 $Y=1.58
+ $X2=1.195 $Y2=1.495
r74 31 46 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.03 $Y=1.58
+ $X2=0.41 $Y2=1.58
r75 30 45 2.0523 $w=3.63e-07 $l=6.5e-08 $layer=LI1_cond $X=0.195 $Y=1.677
+ $X2=0.26 $Y2=1.677
r76 30 41 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.195 $Y=1.495
+ $X2=0.195 $Y2=0.84
r77 26 27 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.48 $Y=1.16 $X2=1.9
+ $Y2=1.16
r78 25 26 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=1.44 $Y=1.16 $X2=1.48
+ $Y2=1.16
r79 24 36 37.7695 $w=2.7e-07 $l=1.7e-07 $layer=POLY_cond $X=1.365 $Y=1.16
+ $X2=1.195 $Y2=1.16
r80 24 25 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.365 $Y=1.16
+ $X2=1.44 $Y2=1.16
r81 23 36 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.035 $Y=1.16
+ $X2=1.195 $Y2=1.16
r82 19 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.9 $Y=1.025
+ $X2=1.9 $Y2=1.16
r83 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.9 $Y=1.025
+ $X2=1.9 $Y2=0.56
r84 15 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.48 $Y=1.025
+ $X2=1.48 $Y2=1.16
r85 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.48 $Y=1.025
+ $X2=1.48 $Y2=0.56
r86 11 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.44 $Y=1.295
+ $X2=1.44 $Y2=1.16
r87 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.44 $Y=1.295
+ $X2=1.44 $Y2=1.985
r88 7 23 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.96 $Y=1.295
+ $X2=1.035 $Y2=1.16
r89 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.96 $Y=1.295 $X2=0.96
+ $Y2=1.985
r90 2 45 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.695
r91 1 39 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_2%B 3 7 11 15 17 22 23 24 25 32
c58 23 0 1.63453e-19 $X=1.99 $Y=1.445
c59 7 0 8.81896e-20 $X=2.32 $Y=0.56
r60 25 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r61 24 25 23.0136 $w=1.98e-07 $l=4.15e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.95 $Y2=1.175
r62 24 39 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.18 $Y2=1.175
r63 22 39 3.3237 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=2.085 $Y=1.175 $X2=2.18
+ $Y2=1.175
r64 22 23 10.7196 $w=3.58e-07 $l=2.55e-07 $layer=LI1_cond $X=2.085 $Y=1.275
+ $X2=2.085 $Y2=1.53
r65 20 21 10.5164 $w=2.75e-07 $l=6e-08 $layer=POLY_cond $X=2.68 $Y=1.16 $X2=2.74
+ $Y2=1.16
r66 17 32 27.9249 $w=2.9e-07 $l=1.35e-07 $layer=POLY_cond $X=2.815 $Y=1.16
+ $X2=2.95 $Y2=1.16
r67 17 21 12.6442 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=2.815 $Y=1.16
+ $X2=2.74 $Y2=1.16
r68 13 21 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.74 $Y=1.015
+ $X2=2.74 $Y2=1.16
r69 13 15 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.74 $Y=1.015
+ $X2=2.74 $Y2=0.56
r70 9 20 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.68 $Y=1.305
+ $X2=2.68 $Y2=1.16
r71 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.68 $Y=1.305
+ $X2=2.68 $Y2=1.985
r72 5 20 63.0982 $w=2.75e-07 $l=3.6e-07 $layer=POLY_cond $X=2.32 $Y=1.16
+ $X2=2.68 $Y2=1.16
r73 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.32 $Y=1.025
+ $X2=2.32 $Y2=0.56
r74 1 5 10.5164 $w=2.75e-07 $l=6e-08 $layer=POLY_cond $X=2.26 $Y=1.16 $X2=2.32
+ $Y2=1.16
r75 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.26 $Y=1.295 $X2=2.26
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_2%VPWR 1 2 3 12 16 18 22 24 29 35 40 43 46
r45 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 42 43 9.49736 $w=6.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.99 $Y=2.49
+ $X2=2.11 $Y2=2.49
r47 38 42 7.21444 $w=6.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.61 $Y=2.49
+ $X2=1.99 $Y2=2.49
r48 38 40 8.64302 $w=6.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.61 $Y=2.49
+ $X2=1.535 $Y2=2.49
r49 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 33 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 32 43 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.11 $Y2=2.72
r55 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 29 45 4.81317 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=2.805 $Y=2.72
+ $X2=3.012 $Y2=2.72
r57 29 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.805 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 24 35 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.58 $Y=2.72
+ $X2=0.707 $Y2=2.72
r59 24 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.58 $Y=2.72
+ $X2=0.23 $Y2=2.72
r60 22 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r62 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.97 $Y=1.66
+ $X2=2.97 $Y2=2.34
r63 16 45 2.95301 $w=3.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=3.012 $Y2=2.72
r64 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2.34
r65 15 35 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=0.707 $Y2=2.72
r66 15 40 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=1.535 $Y2=2.72
r67 10 35 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=2.635
+ $X2=0.707 $Y2=2.72
r68 10 12 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.707 $Y=2.635
+ $X2=0.707 $Y2=2
r69 3 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.485 $X2=2.89 $Y2=2.34
r70 3 18 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.485 $X2=2.89 $Y2=1.66
r71 2 42 300 $w=1.7e-07 $l=1.06637e-06 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=1.485 $X2=1.99 $Y2=2.34
r72 1 12 300 $w=1.7e-07 $l=6.08933e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_2%Y 1 2 3 12 13 18 21 22 23 24 25 32 41 50
c49 32 0 8.81896e-20 $X=1.67 $Y=0.905
c50 2 0 4.63282e-20 $X=1.035 $Y=1.485
r51 32 50 2.34165 $w=3.28e-07 $l=6.42262e-08 $layer=LI1_cond $X=1.67 $Y=0.905
+ $X2=1.69 $Y2=0.85
r52 25 50 0.557927 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.69 $Y=0.835
+ $X2=1.69 $Y2=0.85
r53 25 47 4.27744 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.69 $Y=0.835
+ $X2=1.69 $Y2=0.72
r54 25 32 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.67 $Y=0.92
+ $X2=1.67 $Y2=0.905
r55 24 33 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.615 $Y=1.92
+ $X2=1.67 $Y2=1.92
r56 24 41 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.615 $Y=1.92
+ $X2=1.2 $Y2=1.92
r57 24 33 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=1.67 $Y=1.81
+ $X2=1.67 $Y2=1.835
r58 23 24 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=1.67 $Y=1.53
+ $X2=1.67 $Y2=1.81
r59 22 23 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.67 $Y=1.19 $X2=1.67
+ $Y2=1.53
r60 22 25 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=1.67 $Y=1.19
+ $X2=1.67 $Y2=0.92
r61 16 21 3.01263 $w=3.15e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.497 $Y=1.835
+ $X2=2.457 $Y2=1.92
r62 16 18 7.33373 $w=2.73e-07 $l=1.75e-07 $layer=LI1_cond $X=2.497 $Y=1.835
+ $X2=2.497 $Y2=1.66
r63 13 33 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.81 $Y=1.92
+ $X2=1.67 $Y2=1.92
r64 12 21 3.63293 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.28 $Y=1.92
+ $X2=2.457 $Y2=1.92
r65 12 13 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.28 $Y=1.92
+ $X2=1.81 $Y2=1.92
r66 3 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.335
+ $Y=1.485 $X2=2.47 $Y2=2
r67 3 18 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.47 $Y2=1.66
r68 2 41 300 $w=1.7e-07 $l=5.91777e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.485 $X2=1.2 $Y2=2
r69 1 47 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r46 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r47 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r49 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r50 30 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.53
+ $Y2=0
r51 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.99
+ $Y2=0
r52 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r53 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r54 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r55 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r56 25 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r57 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r59 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r60 22 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.53
+ $Y2=0
r61 22 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.07
+ $Y2=0
r62 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r63 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r64 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r65 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 11 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0
r67 11 13 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0.36
r68 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r69 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r70 2 13 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.53 $Y2=0.36
r71 1 9 91 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.465 $X2=0.745 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_2%A_229_47# 1 2 3 10 12 14 16 17 18 22
c48 17 0 1.56255e-19 $X=2.15 $Y=0.695
r49 20 22 10.372 $w=3.48e-07 $l=3.15e-07 $layer=LI1_cond $X=2.96 $Y=0.695
+ $X2=2.96 $Y2=0.38
r50 19 29 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.275 $Y=0.8
+ $X2=2.15 $Y2=0.8
r51 18 20 7.38573 $w=2.1e-07 $l=2.21359e-07 $layer=LI1_cond $X=2.785 $Y=0.8
+ $X2=2.96 $Y2=0.695
r52 18 19 26.9351 $w=2.08e-07 $l=5.1e-07 $layer=LI1_cond $X=2.785 $Y=0.8
+ $X2=2.275 $Y2=0.8
r53 17 29 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.15 $Y=0.695
+ $X2=2.15 $Y2=0.8
r54 16 27 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.15 $Y=0.465
+ $X2=2.15 $Y2=0.36
r55 16 17 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=2.15 $Y=0.465
+ $X2=2.15 $Y2=0.695
r56 15 25 3.96222 $w=2.1e-07 $l=1.38e-07 $layer=LI1_cond $X=1.355 $Y=0.36
+ $X2=1.217 $Y2=0.36
r57 14 27 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=0.36
+ $X2=2.15 $Y2=0.36
r58 14 15 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=0.36
+ $X2=1.355 $Y2=0.36
r59 10 25 3.01473 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=1.217 $Y=0.465
+ $X2=1.217 $Y2=0.36
r60 10 12 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=1.217 $Y=0.465
+ $X2=1.217 $Y2=0.72
r61 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.815
+ $Y=0.235 $X2=2.95 $Y2=0.38
r62 2 29 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.72
r63 2 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.38
r64 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.235 $X2=1.27 $Y2=0.38
r65 1 12 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.235 $X2=1.27 $Y2=0.72
.ends


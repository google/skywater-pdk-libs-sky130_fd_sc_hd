* File: sky130_fd_sc_hd__a221o_4.pex.spice
* Created: Tue Sep  1 18:52:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A221O_4%A_79_21# 1 2 3 4 5 16 18 21 23 25 28 30 32
+ 35 37 39 42 44 53 54 55 56 60 61 62 64 65 67 70 77 82 89
c186 89 0 1.68975e-19 $X=1.73 $Y=1.16
c187 82 0 1.79953e-19 $X=4.98 $Y=0.73
c188 61 0 3.07602e-19 $X=4.18 $Y=0.725
c189 55 0 1.64628e-19 $X=1.985 $Y=1.54
c190 54 0 6.31497e-20 $X=4.405 $Y=1.54
c191 53 0 1.74554e-19 $X=1.9 $Y=1.455
c192 1 0 1.19717e-19 $X=3.175 $Y=0.235
r193 86 87 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r194 77 78 23.819 $w=2.1e-07 $l=4.1e-07 $layer=LI1_cond $X=4.57 $Y=1.58 $X2=4.98
+ $Y2=1.58
r195 68 80 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.065 $Y=0.365
+ $X2=4.94 $Y2=0.365
r196 68 70 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=5.065 $Y=0.365
+ $X2=5.82 $Y2=0.365
r197 67 78 1.9771 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.98 $Y=1.455
+ $X2=4.98 $Y2=1.58
r198 66 82 4.53567 $w=2.1e-07 $l=1.08167e-07 $layer=LI1_cond $X=4.98 $Y=0.905
+ $X2=4.94 $Y2=0.815
r199 66 67 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.98 $Y=0.905
+ $X2=4.98 $Y2=1.455
r200 65 82 4.53567 $w=2.1e-07 $l=9e-08 $layer=LI1_cond $X=4.94 $Y=0.725 $X2=4.94
+ $Y2=0.815
r201 64 80 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=4.94 $Y=0.475
+ $X2=4.94 $Y2=0.365
r202 64 65 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=4.94 $Y=0.475
+ $X2=4.94 $Y2=0.725
r203 63 75 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.305 $Y=0.815
+ $X2=4.18 $Y2=0.815
r204 62 82 1.9031 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.815 $Y=0.815
+ $X2=4.94 $Y2=0.815
r205 62 63 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.815 $Y=0.815
+ $X2=4.305 $Y2=0.815
r206 61 75 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=4.18 $Y=0.725 $X2=4.18
+ $Y2=0.815
r207 60 73 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=0.475
+ $X2=4.18 $Y2=0.39
r208 60 61 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=4.18 $Y=0.475
+ $X2=4.18 $Y2=0.725
r209 56 73 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.055 $Y=0.39
+ $X2=4.18 $Y2=0.39
r210 56 58 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.055 $Y=0.39
+ $X2=3.3 $Y2=0.39
r211 54 77 10.0641 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=4.405 $Y=1.54
+ $X2=4.57 $Y2=1.58
r212 54 55 157.882 $w=1.68e-07 $l=2.42e-06 $layer=LI1_cond $X=4.405 $Y=1.54
+ $X2=1.985 $Y2=1.54
r213 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.9 $Y=1.455
+ $X2=1.985 $Y2=1.54
r214 52 53 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.9 $Y=1.285
+ $X2=1.9 $Y2=1.455
r215 51 89 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.68 $Y=1.16 $X2=1.73
+ $Y2=1.16
r216 51 87 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.68 $Y=1.16
+ $X2=1.31 $Y2=1.16
r217 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.16 $X2=1.68 $Y2=1.16
r218 47 86 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.66 $Y=1.16
+ $X2=0.89 $Y2=1.16
r219 47 83 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.66 $Y=1.16
+ $X2=0.47 $Y2=1.16
r220 46 50 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=0.66 $Y=1.18
+ $X2=1.68 $Y2=1.18
r221 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.66
+ $Y=1.16 $X2=0.66 $Y2=1.16
r222 44 52 6.6395 $w=1.97e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.815 $Y=1.18
+ $X2=1.9 $Y2=1.285
r223 44 50 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=1.18
+ $X2=1.68 $Y2=1.18
r224 40 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r225 40 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r226 37 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r227 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r228 33 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r229 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r230 30 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r231 30 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r232 26 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r233 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r234 23 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r235 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r236 19 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r237 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r238 16 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r239 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r240 5 77 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.435
+ $Y=1.485 $X2=4.57 $Y2=1.62
r241 4 70 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.38
r242 3 82 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.73
r243 3 80 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.39
r244 2 75 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.73
r245 2 73 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.39
r246 1 58 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.3 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%A2 1 3 6 8 10 13 15 22
c48 15 0 1.68975e-19 $X=2.54 $Y=1.19
c49 1 0 1.55941e-19 $X=2.15 $Y=0.995
r50 20 22 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.43 $Y=1.16
+ $X2=2.57 $Y2=1.16
r51 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=1.16 $X2=2.43 $Y2=1.16
r52 17 20 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.43 $Y2=1.16
r53 15 21 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=2.54 $Y=1.18
+ $X2=2.43 $Y2=1.18
r54 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r55 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r56 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r57 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r58 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r59 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
r60 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995 $X2=2.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%A1 3 7 9 11 12 14 17 18 31 36 38
c59 31 0 1.27649e-19 $X=3.93 $Y=1.16
c60 12 0 1.79953e-19 $X=3.93 $Y=0.995
r61 36 38 32.0404 $w=1.78e-07 $l=5.2e-07 $layer=LI1_cond $X=3.19 $Y=1.195
+ $X2=3.71 $Y2=1.195
r62 29 31 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.875 $Y=1.16
+ $X2=3.93 $Y2=1.16
r63 27 29 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=3.51 $Y=1.16
+ $X2=3.875 $Y2=1.16
r64 26 27 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=3.415 $Y=1.16
+ $X2=3.51 $Y2=1.16
r65 24 26 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=3.02 $Y=1.16
+ $X2=3.415 $Y2=1.16
r66 21 24 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=2.99 $Y=1.16 $X2=3.02
+ $Y2=1.16
r67 18 38 8.97179 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=1.18
+ $X2=3.71 $Y2=1.18
r68 18 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.875
+ $Y=1.16 $X2=3.875 $Y2=1.16
r69 17 36 10.2921 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=3 $Y=1.18 $X2=3.19
+ $Y2=1.18
r70 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.16 $X2=3.02 $Y2=1.16
r71 12 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.16
r72 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=0.56
r73 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.16
r74 9 11 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
r75 5 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.325
+ $X2=3.415 $Y2=1.16
r76 5 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.415 $Y=1.325
+ $X2=3.415 $Y2=1.985
r77 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r78 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325 $X2=2.99
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%C1 1 3 6 8 10 13 15 21 22 25
c53 22 0 6.31497e-20 $X=4.77 $Y=1.16
c54 13 0 1.29399e-19 $X=4.78 $Y=1.985
c55 8 0 8.27827e-20 $X=4.77 $Y=0.995
c56 1 0 8.33213e-20 $X=4.35 $Y=0.995
r57 22 23 1.48308 $w=3.25e-07 $l=1e-08 $layer=POLY_cond $X=4.77 $Y=1.16 $X2=4.78
+ $Y2=1.16
r58 20 22 35.5938 $w=3.25e-07 $l=2.4e-07 $layer=POLY_cond $X=4.53 $Y=1.16
+ $X2=4.77 $Y2=1.16
r59 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.16 $X2=4.53 $Y2=1.16
r60 18 20 25.2123 $w=3.25e-07 $l=1.7e-07 $layer=POLY_cond $X=4.36 $Y=1.16
+ $X2=4.53 $Y2=1.16
r61 17 18 1.48308 $w=3.25e-07 $l=1e-08 $layer=POLY_cond $X=4.35 $Y=1.16 $X2=4.36
+ $Y2=1.16
r62 15 21 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=4.41 $Y=1.18
+ $X2=4.53 $Y2=1.18
r63 15 25 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=4.41 $Y=1.18
+ $X2=4.405 $Y2=1.18
r64 11 23 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.78 $Y=1.325
+ $X2=4.78 $Y2=1.16
r65 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.78 $Y=1.325
+ $X2=4.78 $Y2=1.985
r66 8 22 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.995 $X2=4.77
+ $Y2=1.16
r67 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r68 4 18 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=1.325 $X2=4.36
+ $Y2=1.16
r69 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.36 $Y=1.325 $X2=4.36
+ $Y2=1.985
r70 1 17 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=0.995 $X2=4.35
+ $Y2=1.16
r71 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995 $X2=4.35
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%B1 1 3 6 8 10 13 15 20 23 24
c49 1 0 1.79953e-19 $X=5.19 $Y=0.995
r50 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.87
+ $Y=1.16 $X2=5.87 $Y2=1.16
r51 20 24 28.5195 $w=2.08e-07 $l=5.4e-07 $layer=LI1_cond $X=5.33 $Y=1.18
+ $X2=5.87 $Y2=1.18
r52 18 19 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=5.61 $Y=1.16 $X2=5.62
+ $Y2=1.16
r53 17 18 60.25 $w=3.28e-07 $l=4.1e-07 $layer=POLY_cond $X=5.2 $Y=1.16 $X2=5.61
+ $Y2=1.16
r54 16 17 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=5.19 $Y=1.16 $X2=5.2
+ $Y2=1.16
r55 15 23 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.695 $Y=1.16
+ $X2=5.87 $Y2=1.16
r56 15 19 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.695 $Y=1.16
+ $X2=5.62 $Y2=1.16
r57 11 19 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.62 $Y=1.325
+ $X2=5.62 $Y2=1.16
r58 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.62 $Y=1.325
+ $X2=5.62 $Y2=1.985
r59 8 18 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.16
r60 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r61 4 17 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.2 $Y=1.325 $X2=5.2
+ $Y2=1.16
r62 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.2 $Y=1.325 $X2=5.2
+ $Y2=1.985
r63 1 16 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.16
r64 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995 $X2=5.19
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%B2 3 5 7 10 12 14 15 22 24
r43 23 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.88 $Y=1.16 $X2=6.97
+ $Y2=1.16
r44 21 23 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.845 $Y=1.16
+ $X2=6.88 $Y2=1.16
r45 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.845
+ $Y=1.16 $X2=6.845 $Y2=1.16
r46 19 21 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=6.55 $Y=1.16
+ $X2=6.845 $Y2=1.16
r47 17 19 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.46 $Y=1.16 $X2=6.55
+ $Y2=1.16
r48 15 22 0.362376 $w=1.008e-06 $l=3e-08 $layer=LI1_cond $X=6.775 $Y=1.19
+ $X2=6.775 $Y2=1.16
r49 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=1.16
r50 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=0.56
r51 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.88 $Y=1.325
+ $X2=6.88 $Y2=1.16
r52 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.88 $Y=1.325
+ $X2=6.88 $Y2=1.985
r53 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=0.995
+ $X2=6.55 $Y2=1.16
r54 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.55 $Y=0.995 $X2=6.55
+ $Y2=0.56
r55 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.46 $Y=1.325
+ $X2=6.46 $Y2=1.16
r56 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.46 $Y=1.325 $X2=6.46
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 67 68
c99 1 0 1.27562e-19 $X=0.135 $Y=1.485
r100 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r101 65 68 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=7.59 $Y2=2.72
r102 64 67 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=7.59 $Y2=2.72
r103 64 65 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r104 62 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r105 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r106 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r108 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r109 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r110 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r111 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r112 50 71 3.80464 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r113 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 48 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 48 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r116 46 61 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.5 $Y=2.72 $X2=3.45
+ $Y2=2.72
r117 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.5 $Y=2.72
+ $X2=3.625 $Y2=2.72
r118 45 64 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.75 $Y=2.72
+ $X2=3.625 $Y2=2.72
r120 43 58 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.53 $Y2=2.72
r121 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.78 $Y2=2.72
r122 42 61 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.905 $Y=2.72
+ $X2=3.45 $Y2=2.72
r123 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.905 $Y=2.72
+ $X2=2.78 $Y2=2.72
r124 40 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.61 $Y2=2.72
r125 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.94 $Y2=2.72
r126 39 58 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.53 $Y2=2.72
r127 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=1.94 $Y2=2.72
r128 37 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=0.69 $Y2=2.72
r129 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=1.1 $Y2=2.72
r130 36 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.225 $Y=2.72
+ $X2=1.61 $Y2=2.72
r131 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=2.72
+ $X2=1.1 $Y2=2.72
r132 32 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.635
+ $X2=3.625 $Y2=2.72
r133 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.625 $Y=2.635
+ $X2=3.625 $Y2=2.3
r134 28 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r135 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.3
r136 24 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r137 24 26 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=1.96
r138 20 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2.72
r139 20 22 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=1.96
r140 16 71 3.21325 $w=2.3e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.192 $Y2=2.72
r141 16 18 33.8217 $w=2.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=1.96
r142 5 34 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.485 $X2=3.625 $Y2=2.3
r143 4 30 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2.3
r144 3 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r145 2 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r146 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%X 1 2 3 4 15 19 21 23 27 29 31 33 34 35 37
+ 40 41 42 50 51
c76 35 0 1.27562e-19 $X=0.555 $Y=1.54
c77 33 0 1.27553e-19 $X=0.515 $Y=0.82
c78 23 0 1.55941e-19 $X=1.355 $Y=0.815
r79 42 51 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=1.54 $X2=0.21
+ $Y2=1.455
r80 42 51 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=0.21 $Y=1.45 $X2=0.21
+ $Y2=1.455
r81 41 42 13.0276 $w=2.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.21 $Y=1.19
+ $X2=0.21 $Y2=1.45
r82 40 50 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=0.82 $X2=0.21
+ $Y2=0.905
r83 40 41 13.5287 $w=2.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.21 $Y=0.92
+ $X2=0.21 $Y2=1.19
r84 40 50 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.21 $Y=0.92
+ $X2=0.21 $Y2=0.905
r85 35 42 9.42571 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.555 $Y=1.54
+ $X2=0.325 $Y2=1.54
r86 35 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=1.54
+ $X2=0.68 $Y2=1.54
r87 33 40 8.37002 $w=3.08e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0.82
+ $X2=0.325 $Y2=0.82
r88 33 34 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.515 $Y=0.82
+ $X2=0.68 $Y2=0.815
r89 29 39 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.625
+ $X2=1.52 $Y2=1.54
r90 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.625
+ $X2=1.52 $Y2=2.3
r91 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=0.725
+ $X2=1.52 $Y2=0.39
r92 24 34 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0.815
+ $X2=0.68 $Y2=0.815
r93 23 25 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=1.52 $Y2=0.725
r94 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=0.845 $Y2=0.815
r95 22 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=1.54
+ $X2=0.68 $Y2=1.54
r96 21 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.395 $Y=1.54
+ $X2=1.52 $Y2=1.54
r97 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.395 $Y=1.54
+ $X2=0.805 $Y2=1.54
r98 17 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.625
+ $X2=0.68 $Y2=1.54
r99 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.625
+ $X2=0.68 $Y2=2.3
r100 13 34 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.68 $Y2=0.815
r101 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.68 $Y2=0.39
r102 4 39 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.62
r103 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.3
r104 3 37 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.62
r105 3 19 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.3
r106 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r107 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%A_445_297# 1 2 3 4 15 21 23 24 25 30 32 33
+ 34 38
c72 23 0 1.29399e-19 $X=5.41 $Y=1.625
r73 33 34 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=4.06 $Y=1.92
+ $X2=4.23 $Y2=1.92
r74 26 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.575 $Y=1.54
+ $X2=5.41 $Y2=1.54
r75 25 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.555 $Y=1.54
+ $X2=6.68 $Y2=1.54
r76 25 26 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.555 $Y=1.54
+ $X2=5.575 $Y2=1.54
r77 23 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=1.625 $X2=5.41
+ $Y2=1.54
r78 23 24 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.41 $Y=1.625
+ $X2=5.41 $Y2=1.875
r79 21 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.245 $Y=1.96
+ $X2=5.41 $Y2=1.875
r80 21 34 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=5.245 $Y=1.96
+ $X2=4.23 $Y2=1.96
r81 20 32 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=3.33 $Y=1.88
+ $X2=3.202 $Y2=1.88
r82 20 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.33 $Y=1.88
+ $X2=4.06 $Y2=1.88
r83 16 30 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.485 $Y=1.88
+ $X2=2.36 $Y2=1.88
r84 15 32 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.075 $Y=1.88
+ $X2=3.202 $Y2=1.88
r85 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.075 $Y=1.88
+ $X2=2.485 $Y2=1.88
r86 4 38 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.535
+ $Y=1.485 $X2=6.67 $Y2=1.62
r87 3 36 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.275
+ $Y=1.485 $X2=5.41 $Y2=1.62
r88 2 32 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.205 $Y2=1.96
r89 1 30 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%A_804_297# 1 2 3 4 19 23 27 28
r35 26 28 10.0761 $w=6.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.25 $Y=2.13
+ $X2=6.385 $Y2=2.13
r36 26 27 13.9388 $w=6.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.25 $Y=2.13
+ $X2=5.745 $Y2=2.13
r37 21 23 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.1 $Y=2.295
+ $X2=7.1 $Y2=1.96
r38 19 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.975 $Y=2.38
+ $X2=7.1 $Y2=2.295
r39 19 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.975 $Y=2.38
+ $X2=6.385 $Y2=2.38
r40 18 27 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=4.99 $Y=2.34
+ $X2=5.745 $Y2=2.34
r41 15 18 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=4.145 $Y=2.34
+ $X2=4.99 $Y2=2.34
r42 4 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.955
+ $Y=1.485 $X2=7.09 $Y2=1.96
r43 3 26 150 $w=1.7e-07 $l=7.56075e-07 $layer=licon1_PDIFF $count=4 $X=5.695
+ $Y=1.485 $X2=6.25 $Y2=1.96
r44 2 18 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.485 $X2=4.99 $Y2=2.3
r45 1 15 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.485 $X2=4.145 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 56 57 58 83 84
c127 33 0 1.79013e-19 $X=2.78 $Y=0.73
c128 1 0 1.27553e-19 $X=0.135 $Y=0.235
r129 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r130 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r131 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r132 78 81 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.67 $Y2=0
r133 77 80 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.67
+ $Y2=0
r134 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r135 75 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r136 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r137 72 75 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=4.37 $Y2=0
r138 71 74 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.37
+ $Y2=0
r139 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r140 69 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r141 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r142 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r143 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r144 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r145 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r146 60 87 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r147 60 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r148 58 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r149 58 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r150 56 80 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.67
+ $Y2=0
r151 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.76
+ $Y2=0
r152 55 83 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=6.845 $Y=0
+ $X2=7.59 $Y2=0
r153 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=0 $X2=6.76
+ $Y2=0
r154 53 74 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r155 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.56
+ $Y2=0
r156 52 77 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.645 $Y=0
+ $X2=4.83 $Y2=0
r157 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=0 $X2=4.56
+ $Y2=0
r158 50 68 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=2.53 $Y2=0
r159 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.78
+ $Y2=0
r160 49 71 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.99 $Y2=0
r161 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.78
+ $Y2=0
r162 47 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r163 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.94
+ $Y2=0
r164 46 68 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.53 $Y2=0
r165 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.94
+ $Y2=0
r166 44 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r167 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r168 43 65 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r169 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r170 39 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=0.085
+ $X2=6.76 $Y2=0
r171 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.76 $Y=0.085
+ $X2=6.76 $Y2=0.39
r172 35 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0
r173 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0.39
r174 31 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r175 31 33 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.73
r176 27 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r177 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.39
r178 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r179 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.39
r180 19 87 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r181 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r182 6 41 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.235 $X2=6.76 $Y2=0.39
r183 5 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.39
r184 4 33 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.73
r185 3 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.39
r186 2 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r187 1 21 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%A_445_47# 1 2 9 11 13 15 16 19 22
c72 16 0 1.79013e-19 $X=2.225 $Y=0.85
c73 15 0 1.19717e-19 $X=3.34 $Y=0.85
c74 13 0 8.33213e-20 $X=3.72 $Y=0.73
r75 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.485 $Y=0.85
+ $X2=3.485 $Y2=0.85
r76 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.08 $Y=0.85
+ $X2=2.08 $Y2=0.85
r77 16 18 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.225 $Y=0.85
+ $X2=2.08 $Y2=0.85
r78 15 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.34 $Y=0.85
+ $X2=3.485 $Y2=0.85
r79 15 16 1.37995 $w=1.4e-07 $l=1.115e-06 $layer=MET1_cond $X=3.34 $Y=0.85
+ $X2=2.225 $Y2=0.85
r80 11 23 6.48473 $w=2.6e-07 $l=1.32288e-07 $layer=LI1_cond $X=3.61 $Y=0.775
+ $X2=3.485 $Y2=0.79
r81 11 13 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=3.61 $Y=0.775
+ $X2=3.72 $Y2=0.775
r82 7 19 19.0838 $w=1.79e-07 $l=2.8e-07 $layer=LI1_cond $X=2.36 $Y=0.835
+ $X2=2.08 $Y2=0.835
r83 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.36 $Y=0.735
+ $X2=2.36 $Y2=0.39
r84 2 13 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.73
r85 1 9 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_4%A_1053_47# 1 2 3 10 16 20 22
c35 10 0 8.27827e-20 $X=6.375 $Y=0.775
r36 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.18 $Y=0.725
+ $X2=7.18 $Y2=0.39
r37 16 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=7.015 $Y=0.815
+ $X2=7.18 $Y2=0.725
r38 16 22 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.015 $Y=0.815
+ $X2=6.505 $Y2=0.815
r39 12 15 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=5.4 $Y=0.775
+ $X2=6.34 $Y2=0.775
r40 10 22 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=6.375 $Y=0.775
+ $X2=6.505 $Y2=0.775
r41 10 15 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=6.375 $Y=0.775
+ $X2=6.34 $Y2=0.775
r42 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.045
+ $Y=0.235 $X2=7.18 $Y2=0.39
r43 2 15 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=6.215
+ $Y=0.235 $X2=6.34 $Y2=0.74
r44 1 12 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.73
.ends


* File: sky130_fd_sc_hd__o221a_1.pxi.spice
* Created: Tue Sep  1 19:22:27 2020
* 
x_PM_SKY130_FD_SC_HD__O221A_1%C1 N_C1_c_71_n N_C1_M1011_g N_C1_M1009_g
+ N_C1_c_72_n N_C1_c_73_n C1 PM_SKY130_FD_SC_HD__O221A_1%C1
x_PM_SKY130_FD_SC_HD__O221A_1%B1 N_B1_M1007_g N_B1_M1005_g B1 N_B1_c_101_n
+ N_B1_c_102_n PM_SKY130_FD_SC_HD__O221A_1%B1
x_PM_SKY130_FD_SC_HD__O221A_1%B2 N_B2_M1001_g N_B2_M1006_g B2 B2 N_B2_c_138_n
+ N_B2_c_139_n PM_SKY130_FD_SC_HD__O221A_1%B2
x_PM_SKY130_FD_SC_HD__O221A_1%A2 N_A2_M1002_g N_A2_M1010_g A2 A2 N_A2_c_178_n
+ N_A2_c_179_n N_A2_c_180_n PM_SKY130_FD_SC_HD__O221A_1%A2
x_PM_SKY130_FD_SC_HD__O221A_1%A1 N_A1_M1000_g N_A1_c_213_n N_A1_M1004_g A1
+ N_A1_c_215_n PM_SKY130_FD_SC_HD__O221A_1%A1
x_PM_SKY130_FD_SC_HD__O221A_1%A_51_297# N_A_51_297#_M1011_s N_A_51_297#_M1009_s
+ N_A_51_297#_M1001_d N_A_51_297#_M1003_g N_A_51_297#_M1008_g
+ N_A_51_297#_c_254_n N_A_51_297#_c_247_n N_A_51_297#_c_248_n
+ N_A_51_297#_c_256_n N_A_51_297#_c_257_n N_A_51_297#_c_270_n
+ N_A_51_297#_c_289_n N_A_51_297#_c_282_n N_A_51_297#_c_296_n
+ N_A_51_297#_c_258_n N_A_51_297#_c_259_n N_A_51_297#_c_260_n
+ N_A_51_297#_c_249_n N_A_51_297#_c_283_n N_A_51_297#_c_250_n
+ N_A_51_297#_c_251_n N_A_51_297#_c_252_n PM_SKY130_FD_SC_HD__O221A_1%A_51_297#
x_PM_SKY130_FD_SC_HD__O221A_1%VPWR N_VPWR_M1009_d N_VPWR_M1000_d N_VPWR_c_367_n
+ N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n VPWR N_VPWR_c_371_n
+ N_VPWR_c_372_n N_VPWR_c_366_n N_VPWR_c_374_n PM_SKY130_FD_SC_HD__O221A_1%VPWR
x_PM_SKY130_FD_SC_HD__O221A_1%X N_X_M1003_d N_X_M1008_d N_X_c_421_n X X
+ N_X_c_424_n PM_SKY130_FD_SC_HD__O221A_1%X
x_PM_SKY130_FD_SC_HD__O221A_1%A_149_47# N_A_149_47#_M1011_d N_A_149_47#_M1006_d
+ N_A_149_47#_c_446_n PM_SKY130_FD_SC_HD__O221A_1%A_149_47#
x_PM_SKY130_FD_SC_HD__O221A_1%A_240_47# N_A_240_47#_M1007_d N_A_240_47#_M1002_d
+ N_A_240_47#_c_460_n N_A_240_47#_c_474_n N_A_240_47#_c_461_n
+ PM_SKY130_FD_SC_HD__O221A_1%A_240_47#
x_PM_SKY130_FD_SC_HD__O221A_1%VGND N_VGND_M1002_s N_VGND_M1004_d N_VGND_c_496_n
+ N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n
+ VGND N_VGND_c_502_n N_VGND_c_503_n PM_SKY130_FD_SC_HD__O221A_1%VGND
cc_1 VNB N_C1_c_71_n 0.019852f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=0.995
cc_2 VNB N_C1_c_72_n 0.0380332f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_3 VNB N_C1_c_73_n 0.00807297f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.16
cc_4 VNB C1 0.0192649f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_5 VNB B1 0.00386436f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_6 VNB N_B1_c_101_n 0.0200744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B1_c_102_n 0.0166686f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_8 VNB B2 0.00189141f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_9 VNB N_B2_c_138_n 0.0274101f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_10 VNB N_B2_c_139_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_178_n 0.0284295f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_12 VNB N_A2_c_179_n 0.00311861f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_13 VNB N_A2_c_180_n 0.0217006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_213_n 0.0163355f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.985
cc_15 VNB A1 0.00584225f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_16 VNB N_A1_c_215_n 0.0208013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_51_297#_c_247_n 0.0154614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_51_297#_c_248_n 0.00713281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_51_297#_c_249_n 0.00759302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_51_297#_c_250_n 0.00268099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_51_297#_c_251_n 0.0300871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_51_297#_c_252_n 0.0199436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_366_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_421_n 0.0467716f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_25 VNB X 0.0221562f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_26 VNB N_A_149_47#_c_446_n 0.00264414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_240_47#_c_460_n 0.019203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_240_47#_c_461_n 0.00567857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_496_n 0.00416643f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.16
cc_30 VNB N_VGND_c_497_n 0.00635813f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_31 VNB N_VGND_c_498_n 0.0569573f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_499_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_500_n 0.0176326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_501_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_502_n 0.0257487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_503_n 0.231119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_C1_M1009_g 0.0228639f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.985
cc_38 VPB N_C1_c_72_n 0.0168812f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_39 VPB N_C1_c_73_n 5.21492e-19 $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.16
cc_40 VPB N_B1_M1005_g 0.0186506f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.985
cc_41 VPB N_B1_c_101_n 0.00412261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B2_M1001_g 0.0226161f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=0.56
cc_43 VPB B2 0.00124626f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.16
cc_44 VPB N_B2_c_138_n 0.00714808f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_45 VPB N_A2_M1010_g 0.0212788f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.985
cc_46 VPB A2 0.00276845f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.16
cc_47 VPB N_A2_c_178_n 0.00785953f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_48 VPB N_A1_M1000_g 0.0184008f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=0.56
cc_49 VPB N_A1_c_215_n 0.00419373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_51_297#_M1008_g 0.0237823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_51_297#_c_254_n 0.031508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_51_297#_c_248_n 0.00612519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_51_297#_c_256_n 0.00834438f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_51_297#_c_257_n 0.00961884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_51_297#_c_258_n 0.00515488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_51_297#_c_259_n 0.00224647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_51_297#_c_260_n 0.00154651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_51_297#_c_251_n 0.00786464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_367_n 0.0024829f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.16
cc_60 VPB N_VPWR_c_368_n 0.00275526f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_61 VPB N_VPWR_c_369_n 0.0216822f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_370_n 0.0036584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_371_n 0.0486921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_372_n 0.0250663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_366_n 0.0532282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_374_n 0.0050755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB X 0.0321768f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_68 VPB N_X_c_424_n 0.0405094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 N_C1_M1009_g N_B1_M1005_g 0.0203192f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_70 N_C1_c_73_n B1 6.65977e-19 $X=0.67 $Y=1.16 $X2=0 $Y2=0
cc_71 N_C1_c_73_n N_B1_c_101_n 0.0211059f $X=0.67 $Y=1.16 $X2=0 $Y2=0
cc_72 N_C1_c_71_n N_B1_c_102_n 0.0214815f $X=0.67 $Y=0.995 $X2=0 $Y2=0
cc_73 N_C1_c_71_n N_A_51_297#_c_248_n 0.00498556f $X=0.67 $Y=0.995 $X2=0 $Y2=0
cc_74 N_C1_M1009_g N_A_51_297#_c_248_n 0.00464446f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_75 N_C1_c_72_n N_A_51_297#_c_248_n 0.00615756f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_76 N_C1_c_73_n N_A_51_297#_c_248_n 0.00511985f $X=0.67 $Y=1.16 $X2=0 $Y2=0
cc_77 C1 N_A_51_297#_c_248_n 0.0207096f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_78 N_C1_M1009_g N_A_51_297#_c_257_n 0.0119713f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_79 N_C1_c_72_n N_A_51_297#_c_257_n 0.00902338f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_80 C1 N_A_51_297#_c_257_n 0.0130132f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_81 N_C1_M1009_g N_A_51_297#_c_270_n 4.98187e-19 $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_82 N_C1_c_71_n N_A_51_297#_c_249_n 0.00708682f $X=0.67 $Y=0.995 $X2=0 $Y2=0
cc_83 N_C1_c_72_n N_A_51_297#_c_249_n 0.00552858f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_84 C1 N_A_51_297#_c_249_n 0.0125238f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_85 N_C1_M1009_g N_VPWR_c_367_n 0.01187f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_86 N_C1_M1009_g N_VPWR_c_369_n 0.00544582f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_87 N_C1_M1009_g N_VPWR_c_366_n 0.0102189f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_88 N_C1_c_71_n N_A_240_47#_c_461_n 2.76599e-19 $X=0.67 $Y=0.995 $X2=0 $Y2=0
cc_89 N_C1_c_71_n N_VGND_c_498_n 0.00426565f $X=0.67 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C1_c_71_n N_VGND_c_503_n 0.00702451f $X=0.67 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B1_M1005_g N_B2_M1001_g 0.0495813f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_92 B1 B2 0.0160063f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B1_c_101_n B2 5.32225e-19 $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B1_M1005_g B2 9.81323e-19 $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_95 B1 N_B2_c_138_n 0.00118606f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_96 N_B1_c_101_n N_B2_c_138_n 0.0495813f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B1_c_102_n N_B2_c_139_n 0.0272763f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B1_M1005_g N_A_51_297#_c_248_n 0.00229717f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_99 B1 N_A_51_297#_c_248_n 0.016562f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_100 N_B1_c_101_n N_A_51_297#_c_248_n 0.00295107f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B1_c_102_n N_A_51_297#_c_248_n 0.00192903f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_M1005_g N_A_51_297#_c_256_n 0.0109308f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_103 B1 N_A_51_297#_c_256_n 0.02438f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_104 N_B1_c_101_n N_A_51_297#_c_256_n 0.00292298f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B1_M1005_g N_A_51_297#_c_270_n 0.00586523f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B1_M1005_g N_A_51_297#_c_282_n 0.00547192f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B1_M1005_g N_A_51_297#_c_283_n 0.00117881f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B1_M1005_g N_VPWR_c_367_n 0.00717065f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_109 N_B1_M1005_g N_VPWR_c_371_n 0.00513223f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_110 N_B1_M1005_g N_VPWR_c_366_n 0.00848813f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_111 B1 N_A_149_47#_c_446_n 0.00527792f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B1_c_101_n N_A_149_47#_c_446_n 0.00146804f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B1_c_102_n N_A_149_47#_c_446_n 0.00939545f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_114 B1 N_A_240_47#_c_461_n 0.00709717f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_115 N_B1_c_101_n N_A_240_47#_c_461_n 7.30268e-19 $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B1_c_102_n N_A_240_47#_c_461_n 0.00550561f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B1_c_102_n N_VGND_c_498_n 0.00368123f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_c_102_n N_VGND_c_503_n 0.00538566f $X=1.09 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B2_M1001_g A2 0.00171316f $X=1.51 $Y=1.985 $X2=0 $Y2=0
cc_120 B2 A2 0.0243348f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_121 B2 N_A2_c_178_n 6.66734e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B2_c_138_n N_A2_c_178_n 0.0101681f $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_123 B2 N_A2_c_179_n 0.0243348f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B2_c_138_n N_A2_c_179_n 9.64103e-19 $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_125 B2 N_A_51_297#_M1001_d 0.00472395f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_126 N_B2_M1001_g N_A_51_297#_c_256_n 0.00107932f $X=1.51 $Y=1.985 $X2=0 $Y2=0
cc_127 B2 N_A_51_297#_c_256_n 0.0140608f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_128 N_B2_M1001_g N_A_51_297#_c_270_n 0.00404889f $X=1.51 $Y=1.985 $X2=0 $Y2=0
cc_129 B2 N_A_51_297#_c_270_n 0.00585651f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_130 N_B2_M1001_g N_A_51_297#_c_289_n 0.00964365f $X=1.51 $Y=1.985 $X2=0 $Y2=0
cc_131 B2 N_A_51_297#_c_289_n 0.00157524f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_132 B2 N_A_51_297#_c_289_n 0.00594534f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_133 N_B2_M1001_g N_A_51_297#_c_283_n 0.00749973f $X=1.51 $Y=1.985 $X2=0 $Y2=0
cc_134 B2 N_A_51_297#_c_283_n 0.0160501f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_135 N_B2_c_138_n N_A_51_297#_c_283_n 6.24447e-19 $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B2_M1001_g N_VPWR_c_371_n 0.00426014f $X=1.51 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B2_M1001_g N_VPWR_c_366_n 0.00707977f $X=1.51 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B2_c_139_n N_A_149_47#_c_446_n 0.00817144f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B2_c_138_n N_A_240_47#_c_460_n 0.00406449f $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B2_c_139_n N_A_240_47#_c_460_n 0.00748768f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_141 B2 N_A_240_47#_c_461_n 0.0294941f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_142 N_B2_c_138_n N_A_240_47#_c_461_n 0.00103987f $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_143 N_B2_c_139_n N_A_240_47#_c_461_n 0.00773828f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B2_c_139_n N_VGND_c_496_n 0.00252945f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B2_c_139_n N_VGND_c_498_n 0.00368123f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B2_c_139_n N_VGND_c_503_n 0.00660066f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A2_M1010_g N_A1_M1000_g 0.0497122f $X=2.485 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A2_c_180_n N_A1_c_213_n 0.0124239f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_178_n A1 0.00142612f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_179_n A1 0.0160278f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A2_c_178_n N_A1_c_215_n 0.0497122f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_152 A2 N_A_51_297#_M1001_d 0.00977963f $X=2.005 $Y=1.445 $X2=0 $Y2=0
cc_153 N_A2_M1010_g N_A_51_297#_c_296_n 0.00883733f $X=2.485 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A2_M1010_g N_A_51_297#_c_259_n 0.00345654f $X=2.485 $Y=1.985 $X2=0
+ $Y2=0
cc_155 A2 N_A_51_297#_c_259_n 0.00839634f $X=2.005 $Y=1.445 $X2=0 $Y2=0
cc_156 N_A2_M1010_g N_A_51_297#_c_283_n 0.0117718f $X=2.485 $Y=1.985 $X2=0 $Y2=0
cc_157 A2 N_A_51_297#_c_283_n 0.030784f $X=2.005 $Y=1.445 $X2=0 $Y2=0
cc_158 N_A2_c_178_n N_A_51_297#_c_283_n 6.31723e-19 $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_c_179_n N_A_51_297#_c_283_n 0.00232255f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A2_M1010_g N_VPWR_c_368_n 0.0026105f $X=2.485 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A2_M1010_g N_VPWR_c_371_n 0.00430753f $X=2.485 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A2_M1010_g N_VPWR_c_366_n 0.00711996f $X=2.485 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_c_178_n N_A_240_47#_c_460_n 0.00541932f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A2_c_179_n N_A_240_47#_c_460_n 0.0381966f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A2_c_180_n N_A_240_47#_c_460_n 0.0137594f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A2_c_180_n N_A_240_47#_c_474_n 0.011223f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_c_180_n N_VGND_c_496_n 0.00316354f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_c_180_n N_VGND_c_500_n 0.00425021f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A2_c_180_n N_VGND_c_503_n 0.00709f $X=2.375 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_M1000_g N_A_51_297#_M1008_g 0.0216527f $X=2.845 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A1_M1000_g N_A_51_297#_c_258_n 0.0139164f $X=2.845 $Y=1.985 $X2=0 $Y2=0
cc_172 A1 N_A_51_297#_c_258_n 0.0297283f $X=2.925 $Y=1.105 $X2=0 $Y2=0
cc_173 N_A1_c_215_n N_A_51_297#_c_258_n 0.00306699f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_174 A1 N_A_51_297#_c_259_n 0.00338836f $X=2.925 $Y=1.105 $X2=0 $Y2=0
cc_175 N_A1_M1000_g N_A_51_297#_c_260_n 7.09459e-19 $X=2.845 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A1_c_215_n N_A_51_297#_c_260_n 2.50987e-19 $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_177 A1 N_A_51_297#_c_250_n 0.0170576f $X=2.925 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A1_c_215_n N_A_51_297#_c_250_n 2.00717e-19 $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_179 A1 N_A_51_297#_c_251_n 0.00134784f $X=2.925 $Y=1.105 $X2=0 $Y2=0
cc_180 N_A1_c_215_n N_A_51_297#_c_251_n 0.0217109f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A1_c_213_n N_A_51_297#_c_252_n 0.012217f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_M1000_g N_VPWR_c_368_n 0.0153942f $X=2.845 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A1_M1000_g N_VPWR_c_371_n 0.0046653f $X=2.845 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A1_M1000_g N_VPWR_c_366_n 0.00783311f $X=2.845 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A1_c_213_n N_A_240_47#_c_460_n 0.00240887f $X=2.905 $Y=0.995 $X2=0
+ $Y2=0
cc_186 A1 N_A_240_47#_c_460_n 0.0148551f $X=2.925 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A1_c_215_n N_A_240_47#_c_460_n 0.00179264f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A1_c_213_n N_A_240_47#_c_474_n 0.00509815f $X=2.905 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A1_c_213_n N_VGND_c_497_n 0.00159991f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_190 A1 N_VGND_c_497_n 0.00844867f $X=2.925 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A1_c_215_n N_VGND_c_497_n 2.31083e-19 $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A1_c_213_n N_VGND_c_500_n 0.00541964f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_213_n N_VGND_c_503_n 0.00955661f $X=2.905 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_51_297#_c_256_n N_VPWR_M1009_d 0.00323198f $X=1.155 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_195 N_A_51_297#_c_258_n N_VPWR_M1000_d 0.00229612f $X=3.3 $Y=1.54 $X2=0 $Y2=0
cc_196 N_A_51_297#_c_257_n N_VPWR_c_367_n 0.0154507f $X=0.755 $Y=1.54 $X2=0
+ $Y2=0
cc_197 N_A_51_297#_c_270_n N_VPWR_c_367_n 0.0057552f $X=1.24 $Y=1.875 $X2=0
+ $Y2=0
cc_198 N_A_51_297#_c_282_n N_VPWR_c_367_n 0.0137304f $X=1.325 $Y=1.96 $X2=0
+ $Y2=0
cc_199 N_A_51_297#_c_283_n N_VPWR_c_367_n 0.0126441f $X=2.275 $Y=1.96 $X2=0
+ $Y2=0
cc_200 N_A_51_297#_M1008_g N_VPWR_c_368_n 0.00308386f $X=3.325 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_51_297#_c_258_n N_VPWR_c_368_n 0.0197404f $X=3.3 $Y=1.54 $X2=0 $Y2=0
cc_202 N_A_51_297#_c_254_n N_VPWR_c_369_n 0.02094f $X=0.455 $Y=2.3 $X2=0 $Y2=0
cc_203 N_A_51_297#_c_289_n N_VPWR_c_371_n 0.00343127f $X=1.575 $Y=1.96 $X2=0
+ $Y2=0
cc_204 N_A_51_297#_c_282_n N_VPWR_c_371_n 0.00239782f $X=1.325 $Y=1.96 $X2=0
+ $Y2=0
cc_205 N_A_51_297#_c_283_n N_VPWR_c_371_n 0.0578769f $X=2.275 $Y=1.96 $X2=0
+ $Y2=0
cc_206 N_A_51_297#_M1008_g N_VPWR_c_372_n 0.00570217f $X=3.325 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_51_297#_M1009_s N_VPWR_c_366_n 0.00465839f $X=0.255 $Y=1.485 $X2=0
+ $Y2=0
cc_208 N_A_51_297#_M1001_d N_VPWR_c_366_n 0.00680903f $X=1.585 $Y=1.485 $X2=0
+ $Y2=0
cc_209 N_A_51_297#_M1008_g N_VPWR_c_366_n 0.0116479f $X=3.325 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_51_297#_c_254_n N_VPWR_c_366_n 0.0114713f $X=0.455 $Y=2.3 $X2=0 $Y2=0
cc_211 N_A_51_297#_c_289_n N_VPWR_c_366_n 0.00615797f $X=1.575 $Y=1.96 $X2=0
+ $Y2=0
cc_212 N_A_51_297#_c_282_n N_VPWR_c_366_n 0.0045742f $X=1.325 $Y=1.96 $X2=0
+ $Y2=0
cc_213 N_A_51_297#_c_283_n N_VPWR_c_366_n 0.0395775f $X=2.275 $Y=1.96 $X2=0
+ $Y2=0
cc_214 N_A_51_297#_c_256_n A_245_297# 0.00119842f $X=1.155 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_215 N_A_51_297#_c_270_n A_245_297# 0.00254363f $X=1.24 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_216 N_A_51_297#_c_289_n A_245_297# 0.00293242f $X=1.575 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_217 N_A_51_297#_c_282_n A_245_297# 8.18448e-19 $X=1.325 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A_51_297#_c_283_n A_512_297# 0.00182723f $X=2.275 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_51_297#_c_258_n N_X_M1008_d 0.0022945f $X=3.3 $Y=1.54 $X2=0 $Y2=0
cc_220 N_A_51_297#_c_250_n N_X_c_421_n 0.0214469f $X=3.47 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_51_297#_c_251_n N_X_c_421_n 0.00524099f $X=3.47 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_51_297#_c_252_n N_X_c_421_n 0.00777615f $X=3.427 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_51_297#_M1008_g X 0.00642397f $X=3.325 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_51_297#_c_258_n X 0.00893296f $X=3.3 $Y=1.54 $X2=0 $Y2=0
cc_225 N_A_51_297#_c_260_n X 0.00806556f $X=3.385 $Y=1.455 $X2=0 $Y2=0
cc_226 N_A_51_297#_c_250_n X 0.0170593f $X=3.47 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_51_297#_c_251_n X 0.00548511f $X=3.47 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_51_297#_c_252_n X 0.0025028f $X=3.427 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_51_297#_M1008_g N_X_c_424_n 0.00564711f $X=3.325 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_51_297#_c_258_n N_X_c_424_n 0.00137824f $X=3.3 $Y=1.54 $X2=0 $Y2=0
cc_231 N_A_51_297#_c_250_n N_X_c_424_n 0.00504355f $X=3.47 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_51_297#_c_251_n N_X_c_424_n 0.00262516f $X=3.47 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_51_297#_c_259_n N_A_240_47#_c_460_n 0.00519125f $X=2.72 $Y=1.54 $X2=0
+ $Y2=0
cc_234 N_A_51_297#_c_248_n N_A_240_47#_c_461_n 0.00202031f $X=0.67 $Y=1.455
+ $X2=0 $Y2=0
cc_235 N_A_51_297#_c_256_n N_A_240_47#_c_461_n 0.00265948f $X=1.155 $Y=1.54
+ $X2=0 $Y2=0
cc_236 N_A_51_297#_c_258_n N_VGND_c_497_n 0.00257474f $X=3.3 $Y=1.54 $X2=0 $Y2=0
cc_237 N_A_51_297#_c_252_n N_VGND_c_497_n 0.00283964f $X=3.427 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_51_297#_c_247_n N_VGND_c_498_n 0.0210537f $X=0.41 $Y=0.39 $X2=0 $Y2=0
cc_239 N_A_51_297#_c_249_n N_VGND_c_498_n 0.00261859f $X=0.67 $Y=0.735 $X2=0
+ $Y2=0
cc_240 N_A_51_297#_c_252_n N_VGND_c_502_n 0.00540301f $X=3.427 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_51_297#_M1011_s N_VGND_c_503_n 0.00257894f $X=0.285 $Y=0.235 $X2=0
+ $Y2=0
cc_242 N_A_51_297#_c_247_n N_VGND_c_503_n 0.0124562f $X=0.41 $Y=0.39 $X2=0 $Y2=0
cc_243 N_A_51_297#_c_249_n N_VGND_c_503_n 0.00404964f $X=0.67 $Y=0.735 $X2=0
+ $Y2=0
cc_244 N_A_51_297#_c_252_n N_VGND_c_503_n 0.0108183f $X=3.427 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_366_n A_245_297# 0.00257328f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_246 N_VPWR_c_366_n A_512_297# 0.00409664f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_247 N_VPWR_c_366_n N_X_M1008_d 0.00225742f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_248 N_VPWR_c_372_n N_X_c_424_n 0.0444565f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_c_366_n N_X_c_424_n 0.0253782f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_250 N_X_c_421_n N_VGND_c_497_n 0.0275853f $X=3.93 $Y=0.585 $X2=0 $Y2=0
cc_251 N_X_c_421_n N_VGND_c_502_n 0.0433666f $X=3.93 $Y=0.585 $X2=0 $Y2=0
cc_252 N_X_M1003_d N_VGND_c_503_n 0.00226107f $X=3.4 $Y=0.235 $X2=0 $Y2=0
cc_253 N_X_c_421_n N_VGND_c_503_n 0.0259874f $X=3.93 $Y=0.585 $X2=0 $Y2=0
cc_254 N_A_149_47#_c_446_n N_A_240_47#_M1007_d 0.00329099f $X=1.755 $Y=0.39
+ $X2=-0.19 $Y2=-0.24
cc_255 N_A_149_47#_M1006_d N_A_240_47#_c_460_n 0.00319946f $X=1.62 $Y=0.235
+ $X2=0 $Y2=0
cc_256 N_A_149_47#_c_446_n N_A_240_47#_c_460_n 0.0156303f $X=1.755 $Y=0.39 $X2=0
+ $Y2=0
cc_257 N_A_149_47#_c_446_n N_A_240_47#_c_461_n 0.0186894f $X=1.755 $Y=0.39 $X2=0
+ $Y2=0
cc_258 N_A_149_47#_c_446_n N_VGND_c_496_n 0.0102966f $X=1.755 $Y=0.39 $X2=0
+ $Y2=0
cc_259 N_A_149_47#_c_446_n N_VGND_c_498_n 0.0506122f $X=1.755 $Y=0.39 $X2=0
+ $Y2=0
cc_260 N_A_149_47#_M1011_d N_VGND_c_503_n 0.00246352f $X=0.745 $Y=0.235 $X2=0
+ $Y2=0
cc_261 N_A_149_47#_M1006_d N_VGND_c_503_n 0.0021262f $X=1.62 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_149_47#_c_446_n N_VGND_c_503_n 0.0412133f $X=1.755 $Y=0.39 $X2=0
+ $Y2=0
cc_263 N_A_240_47#_c_460_n N_VGND_M1002_s 0.00315719f $X=2.53 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_264 N_A_240_47#_c_460_n N_VGND_c_496_n 0.012101f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_265 N_A_240_47#_c_460_n N_VGND_c_497_n 0.00787895f $X=2.53 $Y=0.82 $X2=0
+ $Y2=0
cc_266 N_A_240_47#_c_460_n N_VGND_c_498_n 0.00384963f $X=2.53 $Y=0.82 $X2=0
+ $Y2=0
cc_267 N_A_240_47#_c_460_n N_VGND_c_500_n 0.00193763f $X=2.53 $Y=0.82 $X2=0
+ $Y2=0
cc_268 N_A_240_47#_c_474_n N_VGND_c_500_n 0.0171957f $X=2.695 $Y=0.39 $X2=0
+ $Y2=0
cc_269 N_A_240_47#_M1007_d N_VGND_c_503_n 0.00220248f $X=1.2 $Y=0.235 $X2=0
+ $Y2=0
cc_270 N_A_240_47#_M1002_d N_VGND_c_503_n 0.00215764f $X=2.56 $Y=0.235 $X2=0
+ $Y2=0
cc_271 N_A_240_47#_c_460_n N_VGND_c_503_n 0.0122175f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_272 N_A_240_47#_c_474_n N_VGND_c_503_n 0.0121066f $X=2.695 $Y=0.39 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__o2111a_4.spice
* Created: Tue Sep  1 19:20:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2111a_4.pex.spice"
.subckt sky130_fd_sc_hd__o2111a_4  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1009 N_A_27_47#_M1009_d N_D1_M1009_g N_A_27_297#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1024 N_A_27_47#_M1024_d N_D1_M1024_g N_A_27_297#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1011 A_445_47# N_C1_M1011_g N_A_27_47#_M1024_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1020 N_A_361_47#_M1020_d N_B1_M1020_g A_445_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75001.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1012 N_A_361_47#_M1020_d N_B1_M1012_g A_277_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.06825 PD=0.92 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.9
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1014 A_277_47# N_C1_M1014_g N_A_27_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.169 PD=0.86 PS=1.82 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A2_M1018_g N_A_361_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.102375 PD=1.82 PS=0.965 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75000.2
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_361_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.102375 PD=0.92 PS=0.965 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1001_d N_A1_M1005_g N_A_361_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A2_M1021_g N_A_361_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.144625 AS=0.12025 PD=1.095 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_27_297#_M1006_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.144625 PD=1.005 PS=1.095 NRD=14.76 NRS=22.152 M=1 R=4.33333
+ SA=75002.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1006_d N_A_27_297#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.092625 PD=1.005 PS=0.935 NRD=0 NRS=0.912 M=1 R=4.33333
+ SA=75002.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1025 N_X_M1025_d N_A_27_297#_M1025_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.092625 PD=0.945 PS=0.935 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1027 N_X_M1025_d N_A_27_297#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.182 PD=0.945 PS=1.86 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_297#_M1002_d N_D1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1015 N_A_27_297#_M1015_d N_D1_M1015_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_A_27_297#_M1015_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1000_d N_B1_M1016_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1022_d N_B1_M1022_g N_A_27_297#_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1022_d N_C1_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.305 PD=1.27 PS=1.61 NRD=0 NRS=32.4853 M=1 R=6.66667 SA=75002.3
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1008 N_A_27_297#_M1003_s N_A2_M1008_g A_681_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.305 AS=0.1375 PD=1.61 PS=1.275 NRD=0 NRS=16.2328 M=1 R=6.66667 SA=75003
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 A_681_297# N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.1375
+ AS=0.14 PD=1.275 PS=1.28 NRD=16.2328 NRS=0 M=1 R=6.66667 SA=75003.5 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1019 A_852_297# N_A1_M1019_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.1775
+ AS=0.14 PD=1.355 PS=1.28 NRD=24.1128 NRS=0 M=1 R=6.66667 SA=75003.9 SB=75000.7
+ A=0.15 P=2.3 MULT=1
MM1026 N_A_27_297#_M1026_d N_A2_M1026_g A_852_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1775 PD=2.52 PS=1.355 NRD=0 NRS=24.1128 M=1 R=6.66667 SA=75004.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_27_297#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1007_d N_A_27_297#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1017 N_X_M1017_d N_A_27_297#_M1017_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1023 N_X_M1017_d N_A_27_297#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=12.4227 P=18.69
c_62 VNB 0 6.66153e-20 $X=0.145 $Y=-0.085
c_121 VPB 0 1.45e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__o2111a_4.pxi.spice"
*
.ends
*
*

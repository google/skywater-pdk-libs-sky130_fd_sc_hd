* File: sky130_fd_sc_hd__buf_8.spice.SKY130_FD_SC_HD__BUF_8.pxi
* Created: Thu Aug 27 14:10:05 2020
* 
x_PM_SKY130_FD_SC_HD__BUF_8%A N_A_M1007_g N_A_M1002_g N_A_M1012_g N_A_M1004_g
+ N_A_c_107_n N_A_M1021_g N_A_M1013_g A A A PM_SKY130_FD_SC_HD__BUF_8%A
x_PM_SKY130_FD_SC_HD__BUF_8%A_27_47# N_A_27_47#_M1007_d N_A_27_47#_M1012_d
+ N_A_27_47#_M1002_s N_A_27_47#_M1004_s N_A_27_47#_M1000_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1003_g N_A_27_47#_M1005_g N_A_27_47#_M1009_g N_A_27_47#_M1006_g
+ N_A_27_47#_M1010_g N_A_27_47#_M1008_g N_A_27_47#_M1014_g N_A_27_47#_M1011_g
+ N_A_27_47#_M1016_g N_A_27_47#_M1015_g N_A_27_47#_M1017_g N_A_27_47#_M1019_g
+ N_A_27_47#_M1018_g N_A_27_47#_M1020_g N_A_27_47#_c_201_n N_A_27_47#_c_355_p
+ N_A_27_47#_c_184_n N_A_27_47#_c_185_n N_A_27_47#_c_202_n N_A_27_47#_c_203_n
+ N_A_27_47#_c_223_n N_A_27_47#_c_349_p N_A_27_47#_c_186_n N_A_27_47#_c_187_n
+ N_A_27_47#_c_188_n N_A_27_47#_c_189_n N_A_27_47#_c_205_n N_A_27_47#_c_190_n
+ N_A_27_47#_c_191_n N_A_27_47#_c_192_n PM_SKY130_FD_SC_HD__BUF_8%A_27_47#
x_PM_SKY130_FD_SC_HD__BUF_8%VPWR N_VPWR_M1002_d N_VPWR_M1013_d N_VPWR_M1005_d
+ N_VPWR_M1008_d N_VPWR_M1015_d N_VPWR_M1020_d N_VPWR_c_374_n N_VPWR_c_375_n
+ N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n
+ N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n
+ N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n VPWR VPWR N_VPWR_c_389_n
+ N_VPWR_c_390_n N_VPWR_c_373_n N_VPWR_c_392_n N_VPWR_c_393_n
+ PM_SKY130_FD_SC_HD__BUF_8%VPWR
x_PM_SKY130_FD_SC_HD__BUF_8%X N_X_M1000_d N_X_M1009_d N_X_M1014_d N_X_M1017_d
+ N_X_M1001_s N_X_M1006_s N_X_M1011_s N_X_M1019_s N_X_c_548_p N_X_c_525_n
+ N_X_c_463_n N_X_c_464_n N_X_c_469_n N_X_c_470_n N_X_c_551_p N_X_c_529_n
+ N_X_c_465_n N_X_c_471_n N_X_c_545_p N_X_c_533_n N_X_c_553_p N_X_c_466_n
+ N_X_c_472_n N_X_c_467_n N_X_c_473_n X X X N_X_c_537_n
+ PM_SKY130_FD_SC_HD__BUF_8%X
x_PM_SKY130_FD_SC_HD__BUF_8%VGND N_VGND_M1007_s N_VGND_M1021_s N_VGND_M1003_s
+ N_VGND_M1010_s N_VGND_M1016_s N_VGND_M1018_s N_VGND_c_566_n N_VGND_c_567_n
+ N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n
+ N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n N_VGND_c_576_n N_VGND_c_577_n
+ N_VGND_c_578_n VGND VGND N_VGND_c_579_n VGND N_VGND_c_580_n N_VGND_c_581_n
+ N_VGND_c_582_n N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n
+ PM_SKY130_FD_SC_HD__BUF_8%VGND
cc_1 VNB N_A_M1007_g 0.0228678f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_M1012_g 0.0170552f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_A_M1004_g 4.49778e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_4 VNB N_A_c_107_n 0.0679847f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_5 VNB N_A_M1021_g 0.0172396f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_6 VNB N_A_M1013_g 4.62826e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_7 VNB A 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_8 VNB N_A_27_47#_M1000_g 0.0174794f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_9 VNB N_A_27_47#_M1001_g 4.62903e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_10 VNB N_A_27_47#_M1003_g 0.0170561f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_11 VNB N_A_27_47#_M1005_g 4.49847e-19 $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_12 VNB N_A_27_47#_M1009_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_13 VNB N_A_27_47#_M1006_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_14 VNB N_A_27_47#_M1010_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_15 VNB N_A_27_47#_M1008_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_16 VNB N_A_27_47#_M1014_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_M1011_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_M1016_g 0.0170518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_M1015_g 4.49527e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_M1017_g 0.0165623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_M1019_g 4.12504e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_M1018_g 0.0233974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_M1020_g 7.17862e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_184_n 0.00292127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_185_n 0.00183779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_186_n 0.00104171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_187_n 0.00305801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_188_n 0.00102395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_189_n 0.00274061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_190_n 0.00127298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_191_n 0.00134032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_192_n 0.137816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_373_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_463_n 0.00308383f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_35 VNB N_X_c_464_n 0.00141134f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_36 VNB N_X_c_465_n 0.00308383f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.175
cc_37 VNB N_X_c_466_n 0.00127314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_467_n 0.00127314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB X 0.00451082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_566_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.295
cc_41 VNB N_VGND_c_567_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_42 VNB N_VGND_c_568_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_569_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_44 VNB N_VGND_c_570_n 0.0112357f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_45 VNB N_VGND_c_571_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_46 VNB N_VGND_c_572_n 0.0317254f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_47 VNB N_VGND_c_573_n 0.0112511f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.175
cc_48 VNB N_VGND_c_574_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_575_n 0.0118636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_576_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_577_n 0.0112357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_578_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_579_n 0.0152765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_580_n 0.011863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_581_n 0.0172587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_582_n 0.292703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_583_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_584_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_585_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VPB N_A_M1002_g 0.0266267f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_A_M1004_g 0.0191647f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_A_c_107_n 0.00598216f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_63 VPB N_A_M1013_g 0.0194261f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_64 VPB N_A_27_47#_M1001_g 0.0198358f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_65 VPB N_A_27_47#_M1005_g 0.0189386f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_66 VPB N_A_27_47#_M1006_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_67 VPB N_A_27_47#_M1008_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_68 VPB N_A_27_47#_M1011_g 0.0189613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_M1015_g 0.0189336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_M1019_g 0.0183577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_M1020_g 0.0266676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_201_n 0.0331497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_202_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_203_n 0.0106324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_188_n 0.00306481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_205_n 0.00345546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_374_n 0.00410835f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.295
cc_78 VPB N_VPWR_c_375_n 0.00354062f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_79 VPB N_VPWR_c_376_n 3.15634e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_377_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.16
cc_81 VPB N_VPWR_c_378_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_82 VPB N_VPWR_c_379_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_83 VPB N_VPWR_c_380_n 0.0452743f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_84 VPB N_VPWR_c_381_n 0.0178658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_382_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_383_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_384_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_385_n 0.0160841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_386_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_387_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_388_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_389_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_390_n 0.0172587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_373_n 0.0596433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_392_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_393_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_X_c_469_n 0.00326551f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_98 VPB N_X_c_470_n 0.00168851f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.16
cc_99 VPB N_X_c_471_n 0.00326551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_X_c_472_n 0.00137166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_X_c_473_n 0.00137166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB X 0.00132527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB X 0.00360398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 N_A_M1021_g N_A_27_47#_M1000_g 0.0213484f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_105 N_A_M1013_g N_A_27_47#_M1001_g 0.0213484f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_M1002_g N_A_27_47#_c_201_n 0.0106215f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_M1004_g N_A_27_47#_c_201_n 7.66249e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_M1007_g N_A_27_47#_c_184_n 0.0126041f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_M1012_g N_A_27_47#_c_184_n 0.0114493f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A_c_107_n N_A_27_47#_c_184_n 0.00322376f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_111 A N_A_27_47#_c_184_n 0.0473007f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_112 N_A_c_107_n N_A_27_47#_c_185_n 0.00413894f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_113 A N_A_27_47#_c_185_n 0.0138086f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_114 N_A_M1002_g N_A_27_47#_c_202_n 0.0107189f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_M1004_g N_A_27_47#_c_202_n 0.0107189f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_c_107_n N_A_27_47#_c_202_n 0.00198252f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_117 A N_A_27_47#_c_202_n 0.0578998f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A_M1002_g N_A_27_47#_c_203_n 0.00168781f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_c_107_n N_A_27_47#_c_203_n 0.00600433f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_120 A N_A_27_47#_c_203_n 0.0231044f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A_M1002_g N_A_27_47#_c_223_n 7.67038e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_M1004_g N_A_27_47#_c_223_n 0.0107272f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_M1013_g N_A_27_47#_c_223_n 0.0109954f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_M1021_g N_A_27_47#_c_186_n 0.0126765f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_125 A N_A_27_47#_c_186_n 0.00392548f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_126 N_A_M1021_g N_A_27_47#_c_187_n 0.00420813f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_127 N_A_c_107_n N_A_27_47#_c_188_n 0.00448196f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_128 A N_A_27_47#_c_188_n 0.00218678f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_129 N_A_M1004_g N_A_27_47#_c_205_n 0.00139111f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_c_107_n N_A_27_47#_c_205_n 0.00198252f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_131 N_A_M1013_g N_A_27_47#_c_205_n 0.0133819f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_c_107_n N_A_27_47#_c_190_n 0.00213376f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_133 A N_A_27_47#_c_190_n 0.0138019f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_c_107_n N_A_27_47#_c_191_n 0.00177712f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_135 A N_A_27_47#_c_191_n 0.0144236f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_c_107_n N_A_27_47#_c_192_n 0.0213484f $X=1.31 $Y=1.025 $X2=0 $Y2=0
cc_137 N_A_M1002_g N_VPWR_c_374_n 0.00268723f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_M1004_g N_VPWR_c_374_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_M1013_g N_VPWR_c_375_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1002_g N_VPWR_c_381_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1004_g N_VPWR_c_383_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1013_g N_VPWR_c_383_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1002_g N_VPWR_c_373_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1004_g N_VPWR_c_373_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1013_g N_VPWR_c_373_n 0.00952874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1007_g N_VGND_c_566_n 0.0094499f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_147 N_A_M1012_g N_VGND_c_566_n 0.00772492f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_148 N_A_M1021_g N_VGND_c_566_n 5.9099e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_M1012_g N_VGND_c_567_n 5.9099e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_150 N_A_M1021_g N_VGND_c_567_n 0.00769102f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_M1012_g N_VGND_c_573_n 0.00350562f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_M1021_g N_VGND_c_573_n 0.00350562f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_153 N_A_M1007_g N_VGND_c_579_n 0.00350562f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A_M1007_g N_VGND_c_582_n 0.00517665f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A_M1012_g N_VGND_c_582_n 0.00418574f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_M1021_g N_VGND_c_582_n 0.00418574f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_202_n N_VPWR_M1002_d 0.00185611f $X=0.935 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_27_47#_c_205_n N_VPWR_M1013_d 0.00332925f $X=1.507 $Y=1.53 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_202_n N_VPWR_c_374_n 0.0104788f $X=0.935 $Y=1.53 $X2=0 $Y2=0
cc_160 N_A_27_47#_M1001_g N_VPWR_c_375_n 0.00137415f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_205_n N_VPWR_c_375_n 0.0102773f $X=1.507 $Y=1.53 $X2=0 $Y2=0
cc_162 N_A_27_47#_M1001_g N_VPWR_c_376_n 7.05049e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_M1005_g N_VPWR_c_376_n 0.0112732f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_27_47#_M1006_g N_VPWR_c_376_n 0.0110878f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_27_47#_M1008_g N_VPWR_c_376_n 6.72101e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_M1006_g N_VPWR_c_377_n 6.72101e-19 $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_M1008_g N_VPWR_c_377_n 0.0110878f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_27_47#_M1011_g N_VPWR_c_377_n 0.0110878f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_27_47#_M1015_g N_VPWR_c_377_n 6.72101e-19 $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_M1011_g N_VPWR_c_378_n 0.0046653f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_27_47#_M1015_g N_VPWR_c_378_n 0.0046653f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1011_g N_VPWR_c_379_n 6.72101e-19 $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1015_g N_VPWR_c_379_n 0.0110878f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1019_g N_VPWR_c_379_n 0.0110878f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1020_g N_VPWR_c_379_n 6.72101e-19 $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1019_g N_VPWR_c_380_n 8.09353e-19 $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_M1020_g N_VPWR_c_380_n 0.0161769f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_201_n N_VPWR_c_381_n 0.0210382f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_223_n N_VPWR_c_383_n 0.0189039f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1001_g N_VPWR_c_385_n 0.00585385f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1005_g N_VPWR_c_385_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1006_g N_VPWR_c_387_n 0.0046653f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_27_47#_M1008_g N_VPWR_c_387_n 0.0046653f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1019_g N_VPWR_c_389_n 0.0046653f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1020_g N_VPWR_c_389_n 0.0046653f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_27_47#_M1002_s N_VPWR_c_373_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_M1004_s N_VPWR_c_373_n 0.00215201f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1001_g N_VPWR_c_373_n 0.0106402f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_27_47#_M1005_g N_VPWR_c_373_n 0.00796766f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1006_g N_VPWR_c_373_n 0.00796766f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1008_g N_VPWR_c_373_n 0.00796766f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1011_g N_VPWR_c_373_n 0.00796766f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1015_g N_VPWR_c_373_n 0.00796766f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1019_g N_VPWR_c_373_n 0.00796766f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1020_g N_VPWR_c_373_n 0.00796766f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_201_n N_VPWR_c_373_n 0.0124268f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_223_n N_VPWR_c_373_n 0.0122217f $X=1.1 $Y=1.63 $X2=0 $Y2=0
cc_198 N_A_27_47#_M1003_g N_X_c_463_n 0.0111101f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_27_47#_M1009_g N_X_c_463_n 0.0114884f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_189_n N_X_c_463_n 0.0467269f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_192_n N_X_c_463_n 0.00205431f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1000_g N_X_c_464_n 7.27465e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_186_n N_X_c_464_n 0.00628034f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_189_n N_X_c_464_n 0.0136643f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_192_n N_X_c_464_n 0.00213429f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_27_47#_M1005_g N_X_c_469_n 0.013304f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_27_47#_M1006_g N_X_c_469_n 0.0135832f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_189_n N_X_c_469_n 0.0412229f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_192_n N_X_c_469_n 0.00201555f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1001_g N_X_c_470_n 7.19058e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_189_n N_X_c_470_n 0.0121473f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_205_n N_X_c_470_n 0.00690855f $X=1.507 $Y=1.53 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_192_n N_X_c_470_n 0.00211055f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_27_47#_M1010_g N_X_c_465_n 0.0115326f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_215 N_A_27_47#_M1014_g N_X_c_465_n 0.0115326f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_189_n N_X_c_465_n 0.0467269f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_192_n N_X_c_465_n 0.00205431f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_27_47#_M1008_g N_X_c_471_n 0.0136273f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_27_47#_M1011_g N_X_c_471_n 0.0136273f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_189_n N_X_c_471_n 0.0412229f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_192_n N_X_c_471_n 0.00201555f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_189_n N_X_c_466_n 0.0136643f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_192_n N_X_c_466_n 0.00213429f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_189_n N_X_c_472_n 0.0121473f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_192_n N_X_c_472_n 0.00211055f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_189_n N_X_c_467_n 0.0136643f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_192_n N_X_c_467_n 0.00213429f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_189_n N_X_c_473_n 0.0121473f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_192_n N_X_c_473_n 0.00211055f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_27_47#_M1016_g X 0.0120816f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A_27_47#_M1015_g X 7.43505e-19 $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A_27_47#_M1017_g X 0.0150937f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A_27_47#_M1019_g X 0.00402798f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_27_47#_M1018_g X 0.00421537f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_235 N_A_27_47#_M1020_g X 0.00384694f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_189_n X 0.0335381f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_192_n X 0.0316594f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_27_47#_M1015_g X 0.0135832f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A_27_47#_M1019_g X 0.0140861f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_27_47#_M1020_g X 0.0015501f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_189_n X 0.0209281f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_192_n X 0.00215943f $X=4.67 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_184_n N_VGND_M1007_s 0.00162006f $X=1.015 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_27_47#_c_186_n N_VGND_M1021_s 0.00337318f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_184_n N_VGND_c_566_n 0.016419f $X=1.015 $Y=0.82 $X2=0 $Y2=0
cc_246 N_A_27_47#_M1000_g N_VGND_c_567_n 0.00799556f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A_27_47#_M1003_g N_VGND_c_567_n 5.77787e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_186_n N_VGND_c_567_n 0.0153948f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_189_n N_VGND_c_567_n 0.00197677f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_27_47#_M1000_g N_VGND_c_568_n 5.77787e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_251 N_A_27_47#_M1003_g N_VGND_c_568_n 0.00769005f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A_27_47#_M1009_g N_VGND_c_568_n 0.00769005f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1010_g N_VGND_c_568_n 5.77787e-19 $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A_27_47#_M1009_g N_VGND_c_569_n 5.77787e-19 $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A_27_47#_M1010_g N_VGND_c_569_n 0.00769005f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_256 N_A_27_47#_M1014_g N_VGND_c_569_n 0.00769005f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_257 N_A_27_47#_M1016_g N_VGND_c_569_n 5.77787e-19 $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A_27_47#_M1014_g N_VGND_c_570_n 0.00350562f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A_27_47#_M1016_g N_VGND_c_570_n 0.00350562f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_27_47#_M1014_g N_VGND_c_571_n 5.77787e-19 $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A_27_47#_M1016_g N_VGND_c_571_n 0.00769005f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A_27_47#_M1017_g N_VGND_c_571_n 0.00769005f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_263 N_A_27_47#_M1018_g N_VGND_c_571_n 5.77787e-19 $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_264 N_A_27_47#_M1017_g N_VGND_c_572_n 7.31324e-19 $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_265 N_A_27_47#_M1018_g N_VGND_c_572_n 0.0125262f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_184_n N_VGND_c_573_n 0.00193763f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_349_p N_VGND_c_573_n 0.0110017f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_186_n N_VGND_c_573_n 0.00193763f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1000_g N_VGND_c_575_n 0.0046653f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_270 N_A_27_47#_M1003_g N_VGND_c_575_n 0.00350562f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_271 N_A_27_47#_M1009_g N_VGND_c_577_n 0.00350562f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_272 N_A_27_47#_M1010_g N_VGND_c_577_n 0.00350562f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_355_p N_VGND_c_579_n 0.0115672f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_184_n N_VGND_c_579_n 0.00193763f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1017_g N_VGND_c_580_n 0.0035053f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_276 N_A_27_47#_M1018_g N_VGND_c_580_n 0.0046653f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_277 N_A_27_47#_M1007_d N_VGND_c_582_n 0.00377256f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1012_d N_VGND_c_582_n 0.00266498f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1000_g N_VGND_c_582_n 0.00796766f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_280 N_A_27_47#_M1003_g N_VGND_c_582_n 0.00418574f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A_27_47#_M1009_g N_VGND_c_582_n 0.00418574f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_27_47#_M1010_g N_VGND_c_582_n 0.00418574f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_27_47#_M1014_g N_VGND_c_582_n 0.00418574f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A_27_47#_M1016_g N_VGND_c_582_n 0.00418574f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A_27_47#_M1017_g N_VGND_c_582_n 0.00418516f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_27_47#_M1018_g N_VGND_c_582_n 0.00796766f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_355_p N_VGND_c_582_n 0.0064623f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_184_n N_VGND_c_582_n 0.00895872f $X=1.015 $Y=0.82 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_349_p N_VGND_c_582_n 0.00644569f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_186_n N_VGND_c_582_n 0.00485047f $X=1.42 $Y=0.82 $X2=0 $Y2=0
cc_291 N_VPWR_c_373_n N_X_M1001_s 0.00570907f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_373_n N_X_M1006_s 0.00570907f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_373_n N_X_M1011_s 0.00570907f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_c_373_n N_X_M1019_s 0.00570907f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_295 N_VPWR_c_385_n N_X_c_525_n 0.0113958f $X=2.195 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_c_373_n N_X_c_525_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_M1005_d N_X_c_469_n 0.00185611f $X=2.225 $Y=1.485 $X2=0 $Y2=0
cc_298 N_VPWR_c_376_n N_X_c_469_n 0.0140015f $X=2.36 $Y=2 $X2=0 $Y2=0
cc_299 N_VPWR_c_387_n N_X_c_529_n 0.0113958f $X=3.035 $Y=2.72 $X2=0 $Y2=0
cc_300 N_VPWR_c_373_n N_X_c_529_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_M1008_d N_X_c_471_n 0.00185611f $X=3.065 $Y=1.485 $X2=0 $Y2=0
cc_302 N_VPWR_c_377_n N_X_c_471_n 0.0140015f $X=3.2 $Y=2 $X2=0 $Y2=0
cc_303 N_VPWR_c_378_n N_X_c_533_n 0.0113958f $X=3.875 $Y=2.72 $X2=0 $Y2=0
cc_304 N_VPWR_c_373_n N_X_c_533_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_305 N_VPWR_M1015_d X 0.00185611f $X=3.905 $Y=1.485 $X2=0 $Y2=0
cc_306 N_VPWR_c_379_n X 0.0140015f $X=4.04 $Y=2 $X2=0 $Y2=0
cc_307 N_VPWR_c_389_n N_X_c_537_n 0.0113958f $X=4.715 $Y=2.72 $X2=0 $Y2=0
cc_308 N_VPWR_c_373_n N_X_c_537_n 0.00646998f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_309 N_VPWR_c_380_n N_VGND_c_572_n 0.00942828f $X=4.88 $Y=1.66 $X2=0 $Y2=0
cc_310 N_X_c_463_n N_VGND_M1003_s 0.00162006f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_311 N_X_c_465_n N_VGND_M1010_s 0.00162006f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_312 X N_VGND_M1016_s 0.00162006f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_313 N_X_c_463_n N_VGND_c_568_n 0.016419f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_314 N_X_c_465_n N_VGND_c_569_n 0.016419f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_315 N_X_c_465_n N_VGND_c_570_n 0.00193763f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_316 N_X_c_545_p N_VGND_c_570_n 0.0113595f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_317 X N_VGND_c_570_n 0.00193763f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_318 X N_VGND_c_571_n 0.016419f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_319 N_X_c_548_p N_VGND_c_575_n 0.0113595f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_320 N_X_c_463_n N_VGND_c_575_n 0.00193763f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_321 N_X_c_463_n N_VGND_c_577_n 0.00193763f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_322 N_X_c_551_p N_VGND_c_577_n 0.0113595f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_323 N_X_c_465_n N_VGND_c_577_n 0.00193763f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_324 N_X_c_553_p N_VGND_c_580_n 0.0113958f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_325 X N_VGND_c_580_n 0.00197879f $X=4.29 $Y=0.765 $X2=0 $Y2=0
cc_326 N_X_M1000_d N_VGND_c_582_n 0.00418657f $X=1.805 $Y=0.235 $X2=0 $Y2=0
cc_327 N_X_M1009_d N_VGND_c_582_n 0.00266406f $X=2.645 $Y=0.235 $X2=0 $Y2=0
cc_328 N_X_M1014_d N_VGND_c_582_n 0.00266406f $X=3.485 $Y=0.235 $X2=0 $Y2=0
cc_329 N_X_M1017_d N_VGND_c_582_n 0.00418582f $X=4.325 $Y=0.235 $X2=0 $Y2=0
cc_330 N_X_c_548_p N_VGND_c_582_n 0.0064623f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_331 N_X_c_463_n N_VGND_c_582_n 0.00895872f $X=2.695 $Y=0.82 $X2=0 $Y2=0
cc_332 N_X_c_551_p N_VGND_c_582_n 0.0064623f $X=2.78 $Y=0.56 $X2=0 $Y2=0
cc_333 N_X_c_465_n N_VGND_c_582_n 0.00895872f $X=3.535 $Y=0.82 $X2=0 $Y2=0
cc_334 N_X_c_545_p N_VGND_c_582_n 0.0064623f $X=3.62 $Y=0.56 $X2=0 $Y2=0
cc_335 N_X_c_553_p N_VGND_c_582_n 0.00646998f $X=4.46 $Y=0.56 $X2=0 $Y2=0
cc_336 X N_VGND_c_582_n 0.00909756f $X=4.29 $Y=0.765 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nand3b_1.spice
* Created: Thu Aug 27 14:29:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand3b_1.spice.pex"
.subckt sky130_fd_sc_hd__nand3b_1  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_N_M1004_g N_A_53_93#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=37.812 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 A_232_47# N_C_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.121799 PD=0.92 PS=1.19673 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1000 A_316_47# N_B_M1000_g A_232_47# VNB NSHORT L=0.15 W=0.65 AD=0.125125
+ AS=0.08775 PD=1.035 PS=0.92 NRD=25.38 NRS=14.76 M=1 R=4.33333 SA=75000.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_A_53_93#_M1006_g A_316_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.125125 PD=1.86 PS=1.035 NRD=0 NRS=25.38 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_53_93#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.1092 PD=0.789718 PS=1.36 NRD=28.1316 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_C_M1007_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.205282 PD=1.27 PS=1.88028 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.4 SB=75001.2
+ A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=1 AD=0.1925
+ AS=0.135 PD=1.385 PS=1.27 NRD=10.8153 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1005_d N_A_53_93#_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.1925 PD=2.56 PS=1.385 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75001.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__nand3b_1.spice.SKY130_FD_SC_HD__NAND3B_1.pxi"
*
.ends
*
*

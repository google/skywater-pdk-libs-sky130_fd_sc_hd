* File: sky130_fd_sc_hd__a221oi_4.spice.pex
* Created: Thu Aug 27 14:02:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A221OI_4%C1 1 3 6 8 10 13 15 17 20 22 24 27 29 40
r80 39 40 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.75 $Y2=1.16
r81 37 39 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.33 $Y2=1.16
r82 35 37 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.17 $Y2=1.16
r83 33 35 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.91 $Y2=1.16
r84 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r85 29 34 36.8773 $w=1.98e-07 $l=6.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=0.49 $Y2=1.175
r86 29 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r87 25 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r88 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r89 22 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r91 18 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r92 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r93 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r94 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r95 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r96 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r97 8 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r98 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r99 4 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r100 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.985
r101 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r102 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%B2 1 3 4 6 9 11 13 16 20 22 24 27 31 32 35
+ 39 40 49
c124 32 0 1.68801e-19 $X=5.63 $Y=1.16
c125 11 0 1.5152e-19 $X=3.03 $Y=0.995
c126 4 0 1.49368e-19 $X=2.61 $Y=0.995
c127 1 0 3.01892e-19 $X=2.19 $Y=0.995
r128 46 47 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.03 $Y=1.16 $X2=3.11
+ $Y2=1.16
r129 45 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=3.03 $Y2=1.16
r130 44 45 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.61 $Y=1.16 $X2=2.69
+ $Y2=1.16
r131 42 44 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.19 $Y=1.16
+ $X2=2.61 $Y2=1.16
r132 39 40 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=5.465 $Y=1.53
+ $X2=3.935 $Y2=1.53
r133 38 40 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.765 $Y=1.53
+ $X2=3.935 $Y2=1.53
r134 36 49 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.5 $Y=1.16 $X2=3.53
+ $Y2=1.16
r135 36 47 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=3.5 $Y=1.16
+ $X2=3.11 $Y2=1.16
r136 35 38 17.034 $w=2.65e-07 $l=4.49055e-07 $layer=LI1_cond $X=3.59 $Y=1.16
+ $X2=3.765 $Y2=1.53
r137 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.5
+ $Y=1.16 $X2=3.5 $Y2=1.16
r138 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=1.16 $X2=5.63 $Y2=1.16
r139 29 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.63 $Y=1.445
+ $X2=5.465 $Y2=1.53
r140 29 31 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.63 $Y=1.445
+ $X2=5.63 $Y2=1.16
r141 25 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.16
r142 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.985
r143 22 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=1.16
r144 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=0.56
r145 18 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.16
r146 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.985
r147 14 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r148 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.985
r149 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.03 $Y=0.995
+ $X2=3.03 $Y2=1.16
r150 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.03 $Y=0.995
+ $X2=3.03 $Y2=0.56
r151 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.16
r152 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.985
r153 4 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=0.995
+ $X2=2.61 $Y2=1.16
r154 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.61 $Y=0.995
+ $X2=2.61 $Y2=0.56
r155 1 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=0.995
+ $X2=2.19 $Y2=1.16
r156 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.19 $Y=0.995
+ $X2=2.19 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r64 39 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.12 $Y=1.16 $X2=5.21
+ $Y2=1.16
r65 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.12
+ $Y=1.16 $X2=5.12 $Y2=1.16
r66 37 39 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=5.12 $Y2=1.16
r67 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.37 $Y=1.16
+ $X2=4.79 $Y2=1.16
r68 34 36 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.1 $Y=1.16 $X2=4.37
+ $Y2=1.16
r69 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.1 $Y=1.16
+ $X2=4.1 $Y2=1.16
r70 31 34 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.95 $Y=1.16 $X2=4.1
+ $Y2=1.16
r71 29 40 29.84 $w=2.78e-07 $l=7.25e-07 $layer=LI1_cond $X=4.395 $Y=1.135
+ $X2=5.12 $Y2=1.135
r72 29 35 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.395 $Y=1.135
+ $X2=4.1 $Y2=1.135
r73 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.16
r74 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.985
r75 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=1.16
r76 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=0.56
r77 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.16
r78 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.985
r79 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=1.16
r80 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=0.56
r81 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.325
+ $X2=4.37 $Y2=1.16
r82 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.37 $Y=1.325
+ $X2=4.37 $Y2=1.985
r83 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=1.16
r84 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=0.56
r85 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.325
+ $X2=3.95 $Y2=1.16
r86 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.95 $Y=1.325 $X2=3.95
+ $Y2=1.985
r87 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.95 $Y2=1.16
r88 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.95 $Y=0.995 $X2=3.95
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 31 32 34
+ 35 37 38 39 50 51
c126 32 0 1.80815e-19 $X=6.13 $Y=1.16
r127 49 51 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9 $Y=1.16 $X2=9.07
+ $Y2=1.16
r128 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9
+ $Y=1.16 $X2=9 $Y2=1.16
r129 47 49 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=8.65 $Y=1.16 $X2=9
+ $Y2=1.16
r130 45 47 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=8.32 $Y=1.16
+ $X2=8.65 $Y2=1.16
r131 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.32
+ $Y=1.16 $X2=8.32 $Y2=1.16
r132 42 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.23 $Y=1.16 $X2=8.32
+ $Y2=1.16
r133 39 50 25.7864 $w=1.98e-07 $l=4.65e-07 $layer=LI1_cond $X=8.535 $Y=1.175
+ $X2=9 $Y2=1.175
r134 39 46 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=8.535 $Y=1.175
+ $X2=8.32 $Y2=1.175
r135 38 46 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=8.265 $Y=1.175
+ $X2=8.32 $Y2=1.175
r136 36 38 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=8.18 $Y=1.275
+ $X2=8.265 $Y2=1.175
r137 36 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.18 $Y=1.275
+ $X2=8.18 $Y2=1.445
r138 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.095 $Y=1.53
+ $X2=8.18 $Y2=1.445
r139 34 35 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=8.095 $Y=1.53
+ $X2=6.295 $Y2=1.53
r140 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.13
+ $Y=1.16 $X2=6.13 $Y2=1.16
r141 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.13 $Y=1.445
+ $X2=6.295 $Y2=1.53
r142 29 31 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.13 $Y=1.445
+ $X2=6.13 $Y2=1.16
r143 25 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.07 $Y=1.325
+ $X2=9.07 $Y2=1.16
r144 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.07 $Y=1.325
+ $X2=9.07 $Y2=1.985
r145 22 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.07 $Y=0.995
+ $X2=9.07 $Y2=1.16
r146 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.07 $Y=0.995
+ $X2=9.07 $Y2=0.56
r147 18 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.65 $Y=1.325
+ $X2=8.65 $Y2=1.16
r148 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.65 $Y=1.325
+ $X2=8.65 $Y2=1.985
r149 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.65 $Y=0.995
+ $X2=8.65 $Y2=1.16
r150 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.65 $Y=0.995
+ $X2=8.65 $Y2=0.56
r151 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.16
r152 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.985
r153 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=1.16
r154 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=0.56
r155 4 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=1.325
+ $X2=6.13 $Y2=1.16
r156 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.13 $Y=1.325
+ $X2=6.13 $Y2=1.985
r157 1 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=1.16
r158 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 35 41
r58 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=1.16
+ $X2=7.81 $Y2=1.16
r59 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=7.39 $Y=1.16
+ $X2=7.66 $Y2=1.16
r60 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.97 $Y=1.16
+ $X2=7.39 $Y2=1.16
r61 35 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.66
+ $Y=1.16 $X2=7.66 $Y2=1.16
r62 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=6.64 $Y=1.16
+ $X2=6.97 $Y2=1.16
r63 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.64
+ $Y=1.16 $X2=6.64 $Y2=1.16
r64 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=1.16 $X2=6.64
+ $Y2=1.16
r65 29 35 0.259574 $w=1.408e-06 $l=3e-08 $layer=LI1_cond $X=7.18 $Y=1.19
+ $X2=7.18 $Y2=1.16
r66 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.81 $Y=1.325
+ $X2=7.81 $Y2=1.16
r67 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.81 $Y=1.325
+ $X2=7.81 $Y2=1.985
r68 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.81 $Y=0.995
+ $X2=7.81 $Y2=1.16
r69 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.81 $Y=0.995
+ $X2=7.81 $Y2=0.56
r70 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=1.325
+ $X2=7.39 $Y2=1.16
r71 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.39 $Y=1.325
+ $X2=7.39 $Y2=1.985
r72 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=0.995
+ $X2=7.39 $Y2=1.16
r73 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.39 $Y=0.995
+ $X2=7.39 $Y2=0.56
r74 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=1.325
+ $X2=6.97 $Y2=1.16
r75 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.97 $Y=1.325
+ $X2=6.97 $Y2=1.985
r76 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=1.16
r77 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=0.56
r78 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=1.325
+ $X2=6.55 $Y2=1.16
r79 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.55 $Y=1.325 $X2=6.55
+ $Y2=1.985
r80 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=0.995
+ $X2=6.55 $Y2=1.16
r81 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.55 $Y=0.995 $X2=6.55
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%A_27_297# 1 2 3 4 5 6 7 22 24 26 30 32 35
+ 37 38 39 41 43 50 54
c79 50 0 1.39053e-19 $X=5.42 $Y=1.96
r80 48 50 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=4.58 $Y=1.94
+ $X2=5.42 $Y2=1.94
r81 46 48 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=3.74 $Y=1.94
+ $X2=4.58 $Y2=1.94
r82 44 58 4.13622 $w=2.1e-07 $l=1.48e-07 $layer=LI1_cond $X=3.03 $Y=1.94
+ $X2=2.882 $Y2=1.94
r83 44 46 37.4978 $w=2.08e-07 $l=7.1e-07 $layer=LI1_cond $X=3.03 $Y=1.94
+ $X2=3.74 $Y2=1.94
r84 41 58 2.93448 $w=2.95e-07 $l=1.05e-07 $layer=LI1_cond $X=2.882 $Y=1.835
+ $X2=2.882 $Y2=1.94
r85 41 43 8.39916 $w=2.93e-07 $l=2.15e-07 $layer=LI1_cond $X=2.882 $Y=1.835
+ $X2=2.882 $Y2=1.62
r86 40 43 0.195329 $w=2.93e-07 $l=5e-09 $layer=LI1_cond $X=2.882 $Y=1.615
+ $X2=2.882 $Y2=1.62
r87 38 40 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=2.735 $Y=1.53
+ $X2=2.882 $Y2=1.615
r88 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.735 $Y=1.53
+ $X2=2.125 $Y2=1.53
r89 35 56 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=2.295 $X2=2
+ $Y2=2.38
r90 35 37 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=2 $Y=2.295 $X2=2
+ $Y2=1.63
r91 34 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2 $Y=1.615
+ $X2=2.125 $Y2=1.53
r92 34 37 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=2 $Y=1.615 $X2=2
+ $Y2=1.63
r93 33 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.38
+ $X2=1.12 $Y2=2.38
r94 32 56 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.875 $Y=2.38 $X2=2
+ $Y2=2.38
r95 32 33 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.875 $Y=2.38
+ $X2=1.245 $Y2=2.38
r96 28 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.295
+ $X2=1.12 $Y2=2.38
r97 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.12 $Y=2.295
+ $X2=1.12 $Y2=1.96
r98 27 53 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=2.38
+ $X2=0.247 $Y2=2.38
r99 26 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=2.38
+ $X2=1.12 $Y2=2.38
r100 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=2.38
+ $X2=0.405 $Y2=2.38
r101 22 53 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=2.295
+ $X2=0.247 $Y2=2.38
r102 22 24 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.247 $Y=2.295
+ $X2=0.247 $Y2=1.62
r103 7 50 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.42 $Y2=1.96
r104 6 48 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.485 $X2=4.58 $Y2=1.96
r105 5 46 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.485 $X2=3.74 $Y2=1.96
r106 4 58 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.485 $X2=2.9 $Y2=1.96
r107 4 43 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.485 $X2=2.9 $Y2=1.62
r108 3 56 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.31
r109 3 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.63
r110 2 30 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.96
r111 1 53 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r112 1 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%Y 1 2 3 4 5 6 7 8 27 31 33 34 35 36 39 43
+ 46 47 50 52 63 65 66 67 68 69 70 71 72
c150 65 0 1.32347e-19 $X=1.54 $Y=0.815
c151 39 0 1.69544e-19 $X=1.54 $Y=0.39
r152 70 71 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=6.29 $Y=0.775
+ $X2=6.46 $Y2=0.775
r153 69 70 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.68 $Y=0.82
+ $X2=6.29 $Y2=0.82
r154 68 69 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=5.51 $Y=0.775
+ $X2=5.68 $Y2=0.775
r155 66 72 6.57889 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.605 $Y=1.445
+ $X2=1.605 $Y2=1.275
r156 66 67 4.06715 $w=2.25e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.605 $Y=1.445
+ $X2=1.56 $Y2=1.53
r157 61 63 53.2364 $w=1.73e-07 $l=8.4e-07 $layer=LI1_cond $X=6.76 $Y=0.732
+ $X2=7.6 $Y2=0.732
r158 61 71 19.013 $w=1.73e-07 $l=3e-07 $layer=LI1_cond $X=6.76 $Y=0.732 $X2=6.46
+ $Y2=0.732
r159 56 68 32.3221 $w=1.73e-07 $l=5.1e-07 $layer=LI1_cond $X=5 $Y=0.732 $X2=5.51
+ $Y2=0.732
r160 54 56 53.2364 $w=1.73e-07 $l=8.4e-07 $layer=LI1_cond $X=4.16 $Y=0.732 $X2=5
+ $Y2=0.732
r161 52 54 57.9896 $w=1.73e-07 $l=9.15e-07 $layer=LI1_cond $X=3.245 $Y=0.732
+ $X2=4.16 $Y2=0.732
r162 49 52 6.81835 $w=1.75e-07 $l=1.23386e-07 $layer=LI1_cond $X=3.16 $Y=0.82
+ $X2=3.245 $Y2=0.732
r163 49 50 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.16 $Y=0.82
+ $X2=3.16 $Y2=1.095
r164 48 72 1.72457 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=1.705 $Y=1.185
+ $X2=1.605 $Y2=1.185
r165 47 50 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.075 $Y=1.185
+ $X2=3.16 $Y2=1.095
r166 47 48 84.4141 $w=1.78e-07 $l=1.37e-06 $layer=LI1_cond $X=3.075 $Y=1.185
+ $X2=1.705 $Y2=1.185
r167 46 72 4.72821 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=1.605 $Y=1.095 $X2=1.605
+ $Y2=1.185
r168 45 65 3.70371 $w=2.65e-07 $l=1.1811e-07 $layer=LI1_cond $X=1.605 $Y=0.905
+ $X2=1.54 $Y2=0.815
r169 45 46 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=1.605 $Y=0.905
+ $X2=1.605 $Y2=1.095
r170 41 67 4.06715 $w=2.25e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.54 $Y=1.615
+ $X2=1.56 $Y2=1.53
r171 41 43 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.54 $Y=1.615
+ $X2=1.54 $Y2=1.62
r172 37 65 3.70371 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.815
r173 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r174 35 65 2.76582 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r175 35 36 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r176 33 67 2.36881 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.415 $Y=1.53
+ $X2=1.56 $Y2=1.53
r177 33 34 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.415 $Y=1.53
+ $X2=0.825 $Y2=1.53
r178 29 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.7 $Y=1.615
+ $X2=0.825 $Y2=1.53
r179 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.7 $Y=1.615 $X2=0.7
+ $Y2=1.62
r180 25 36 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r181 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.7 $Y2=0.39
r182 8 43 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.62
r183 7 31 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.62
r184 6 63 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=7.465
+ $Y=0.235 $X2=7.6 $Y2=0.73
r185 5 61 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.235 $X2=6.76 $Y2=0.73
r186 4 56 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5 $Y2=0.73
r187 3 54 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.235 $X2=4.16 $Y2=0.73
r188 2 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r189 1 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%A_471_297# 1 2 3 4 5 6 7 8 9 28 30 32 40 41
+ 42 50 53 54 55 58 69
c90 42 0 1.51067e-19 $X=8.355 $Y=1.915
c91 40 0 5.9496e-20 $X=5.88 $Y=2.045
r92 58 60 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=9.28 $Y=1.62
+ $X2=9.28 $Y2=2.3
r93 56 58 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=9.28 $Y=1.615
+ $X2=9.28 $Y2=1.62
r94 54 56 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.155 $Y=1.53
+ $X2=9.28 $Y2=1.615
r95 54 55 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=9.155 $Y=1.53
+ $X2=8.605 $Y2=1.53
r96 53 69 7.24004 $w=1.7e-07 $l=1.48661e-07 $layer=LI1_cond $X=8.52 $Y=1.785
+ $X2=8.48 $Y2=1.915
r97 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.52 $Y=1.615
+ $X2=8.605 $Y2=1.53
r98 52 53 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.52 $Y=1.615
+ $X2=8.52 $Y2=1.785
r99 48 69 7.24004 $w=1.7e-07 $l=1.48661e-07 $layer=LI1_cond $X=8.44 $Y=2.045
+ $X2=8.48 $Y2=1.915
r100 48 50 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.44 $Y=2.045
+ $X2=8.44 $Y2=2.3
r101 45 47 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=6.76 $Y=1.915
+ $X2=7.6 $Y2=1.915
r102 43 65 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=6.005 $Y=1.915
+ $X2=5.88 $Y2=1.915
r103 43 45 33.4652 $w=2.58e-07 $l=7.55e-07 $layer=LI1_cond $X=6.005 $Y=1.915
+ $X2=6.76 $Y2=1.915
r104 42 69 0.132371 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=8.355 $Y=1.915
+ $X2=8.48 $Y2=1.915
r105 42 47 33.4652 $w=2.58e-07 $l=7.55e-07 $layer=LI1_cond $X=8.355 $Y=1.915
+ $X2=7.6 $Y2=1.915
r106 41 67 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.88 $Y=2.215
+ $X2=5.88 $Y2=2.34
r107 40 65 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=5.88 $Y=2.045
+ $X2=5.88 $Y2=1.915
r108 40 41 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.88 $Y=2.045
+ $X2=5.88 $Y2=2.215
r109 37 39 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=4.16 $Y=2.34 $X2=5
+ $Y2=2.34
r110 35 37 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=3.32 $Y=2.34
+ $X2=4.16 $Y2=2.34
r111 33 63 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=2.565 $Y=2.34
+ $X2=2.44 $Y2=2.34
r112 33 35 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=2.565 $Y=2.34
+ $X2=3.32 $Y2=2.34
r113 32 67 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.755 $Y=2.34
+ $X2=5.88 $Y2=2.34
r114 32 39 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=5.755 $Y=2.34
+ $X2=5 $Y2=2.34
r115 28 63 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=2.44 $Y=2.215
+ $X2=2.44 $Y2=2.34
r116 28 30 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.44 $Y=2.215
+ $X2=2.44 $Y2=1.96
r117 9 60 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.28 $Y2=2.3
r118 9 58 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.28 $Y2=1.62
r119 8 69 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=1.96
r120 8 50 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=2.3
r121 7 47 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=7.465
+ $Y=1.485 $X2=7.6 $Y2=1.96
r122 6 45 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.485 $X2=6.76 $Y2=1.96
r123 5 67 600 $w=1.7e-07 $l=8.98248e-07 $layer=licon1_PDIFF $count=1 $X=5.705
+ $Y=1.485 $X2=5.88 $Y2=2.3
r124 5 65 600 $w=1.7e-07 $l=5.55653e-07 $layer=licon1_PDIFF $count=1 $X=5.705
+ $Y=1.485 $X2=5.88 $Y2=1.96
r125 4 39 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5 $Y2=2.3
r126 3 37 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.485 $X2=4.16 $Y2=2.3
r127 2 35 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.485 $X2=3.32 $Y2=2.3
r128 1 63 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.355
+ $Y=1.485 $X2=2.48 $Y2=2.3
r129 1 30 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=2.355
+ $Y=1.485 $X2=2.48 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%VPWR 1 2 3 4 15 18 19 20 27 28 39 40 45 53
r105 51 53 9.48275 $w=5.88e-07 $l=1.35e-07 $layer=LI1_cond $X=8.05 $Y=2.51
+ $X2=8.185 $Y2=2.51
r106 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r107 49 51 0.608175 $w=5.88e-07 $l=3e-08 $layer=LI1_cond $X=8.02 $Y=2.51
+ $X2=8.05 $Y2=2.51
r108 43 47 2.63543 $w=5.88e-07 $l=1.3e-07 $layer=LI1_cond $X=6.21 $Y=2.51
+ $X2=6.34 $Y2=2.51
r109 43 45 7.4555 $w=5.88e-07 $l=3.5e-08 $layer=LI1_cond $X=6.21 $Y=2.51
+ $X2=6.175 $Y2=2.51
r110 43 44 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r112 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r113 37 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r114 36 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.51 $Y=2.72
+ $X2=8.185 $Y2=2.72
r115 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r116 31 52 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.05 $Y2=2.72
r117 31 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r118 30 33 10.339 $w=5.88e-07 $l=5.1e-07 $layer=LI1_cond $X=6.67 $Y=2.51
+ $X2=7.18 $Y2=2.51
r119 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r120 28 47 2.63543 $w=5.88e-07 $l=1.3e-07 $layer=LI1_cond $X=6.47 $Y=2.51
+ $X2=6.34 $Y2=2.51
r121 28 30 4.0545 $w=5.88e-07 $l=2e-07 $layer=LI1_cond $X=6.47 $Y=2.51 $X2=6.67
+ $Y2=2.51
r122 27 49 2.63543 $w=5.88e-07 $l=1.3e-07 $layer=LI1_cond $X=7.89 $Y=2.51
+ $X2=8.02 $Y2=2.51
r123 27 33 14.3935 $w=5.88e-07 $l=7.1e-07 $layer=LI1_cond $X=7.89 $Y=2.51
+ $X2=7.18 $Y2=2.51
r124 24 45 387.856 $w=1.68e-07 $l=5.945e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=6.175 $Y2=2.72
r125 20 44 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=6.21 $Y2=2.72
r126 20 24 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r127 18 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.775 $Y=2.72
+ $X2=8.51 $Y2=2.72
r128 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.775 $Y=2.72
+ $X2=8.86 $Y2=2.72
r129 17 39 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.945 $Y=2.72
+ $X2=9.43 $Y2=2.72
r130 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.945 $Y=2.72
+ $X2=8.86 $Y2=2.72
r131 13 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=2.635
+ $X2=8.86 $Y2=2.72
r132 13 15 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=8.86 $Y=2.635
+ $X2=8.86 $Y2=1.96
r133 4 15 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.725
+ $Y=1.485 $X2=8.86 $Y2=1.96
r134 3 49 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=2.3
r135 2 33 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=1.485 $X2=7.18 $Y2=2.3
r136 1 47 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%VGND 1 2 3 4 5 6 7 22 24 28 33 35 38 42 46
+ 49 50 52 53 55 56 59 60 62 63 65 66 67 92 93
r138 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r139 90 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.43
+ $Y2=0
r140 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r141 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r142 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r143 84 87 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=8.05 $Y2=0
r144 83 86 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=8.05
+ $Y2=0
r145 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r146 81 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r147 80 81 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r148 78 81 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=5.75
+ $Y2=0
r149 77 80 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=5.75
+ $Y2=0
r150 77 78 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r151 75 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r152 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r153 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r154 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r155 69 96 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r156 69 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.69 $Y2=0
r157 67 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r158 67 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r159 65 89 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=8.97 $Y2=0
r160 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.195 $Y=0 $X2=9.28
+ $Y2=0
r161 64 92 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.365 $Y=0 $X2=9.43
+ $Y2=0
r162 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.365 $Y=0 $X2=9.28
+ $Y2=0
r163 62 86 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.355 $Y=0
+ $X2=8.05 $Y2=0
r164 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=0 $X2=8.44
+ $Y2=0
r165 61 89 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.525 $Y=0
+ $X2=8.97 $Y2=0
r166 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=0 $X2=8.44
+ $Y2=0
r167 59 80 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.75
+ $Y2=0
r168 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.92
+ $Y2=0
r169 58 83 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.005 $Y=0
+ $X2=6.21 $Y2=0
r170 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0 $X2=5.92
+ $Y2=0
r171 55 56 3.26614 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=0.76
+ $X2=2.735 $Y2=0.76
r172 52 74 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r173 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r174 51 77 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.07
+ $Y2=0
r175 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r176 49 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r177 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r178 48 74 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.61 $Y2=0
r179 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r180 44 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=0.085
+ $X2=9.28 $Y2=0
r181 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.28 $Y=0.085
+ $X2=9.28 $Y2=0.39
r182 40 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0
r183 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0.39
r184 36 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r185 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.39
r186 35 56 28.3995 $w=2.78e-07 $l=6.9e-07 $layer=LI1_cond $X=2.045 $Y=0.785
+ $X2=2.735 $Y2=0.785
r187 31 35 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.96 $Y=0.645
+ $X2=2.045 $Y2=0.785
r188 31 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.96 $Y=0.645
+ $X2=1.96 $Y2=0.39
r189 30 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r190 30 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r191 26 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r192 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r193 22 96 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r194 22 24 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.39
r195 7 46 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.145
+ $Y=0.235 $X2=9.28 $Y2=0.39
r196 6 42 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.305
+ $Y=0.235 $X2=8.44 $Y2=0.39
r197 5 38 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.92 $Y2=0.39
r198 4 55 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.685
+ $Y=0.235 $X2=2.82 $Y2=0.76
r199 3 33 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r200 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r201 1 24 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%A_453_47# 1 2 3 4 15 21 26 27
c36 26 0 1.5152e-19 $X=2.61 $Y=0.365
c37 15 0 1.49368e-19 $X=3.255 $Y=0.365
r38 26 27 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.61 $Y=0.34
+ $X2=3.035 $Y2=0.34
r39 24 26 11.6259 $w=2.18e-07 $l=2.1e-07 $layer=LI1_cond $X=2.4 $Y=0.365
+ $X2=2.61 $Y2=0.365
r40 19 21 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=4.58 $Y=0.365
+ $X2=5.42 $Y2=0.365
r41 17 19 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=3.74 $Y=0.365
+ $X2=4.58 $Y2=0.365
r42 15 27 12.1497 $w=2.18e-07 $l=2.2e-07 $layer=LI1_cond $X=3.255 $Y=0.365
+ $X2=3.035 $Y2=0.365
r43 15 17 25.4061 $w=2.18e-07 $l=4.85e-07 $layer=LI1_cond $X=3.255 $Y=0.365
+ $X2=3.74 $Y2=0.365
r44 4 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.235 $X2=5.42 $Y2=0.39
r45 3 19 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.58 $Y2=0.39
r46 2 17 91 $w=1.7e-07 $l=7.08273e-07 $layer=licon1_NDIFF $count=2 $X=3.105
+ $Y=0.235 $X2=3.74 $Y2=0.39
r47 1 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_4%A_1241_47# 1 2 3 4 13 19 20 21 25
r46 23 25 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.86 $Y=0.725
+ $X2=8.86 $Y2=0.39
r47 22 30 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=8.185 $Y=0.815
+ $X2=8.06 $Y2=0.815
r48 21 23 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=8.695 $Y=0.815
+ $X2=8.86 $Y2=0.725
r49 21 22 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=8.695 $Y=0.815
+ $X2=8.185 $Y2=0.815
r50 20 30 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=8.06 $Y=0.725 $X2=8.06
+ $Y2=0.815
r51 19 28 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.06 $Y=0.475
+ $X2=8.06 $Y2=0.365
r52 19 20 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=8.06 $Y=0.475
+ $X2=8.06 $Y2=0.725
r53 15 18 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=6.34 $Y=0.365
+ $X2=7.18 $Y2=0.365
r54 13 28 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=7.935 $Y=0.365
+ $X2=8.06 $Y2=0.365
r55 13 18 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=7.935 $Y=0.365
+ $X2=7.18 $Y2=0.365
r56 4 25 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.725
+ $Y=0.235 $X2=8.86 $Y2=0.39
r57 3 30 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.73
r58 3 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.39
r59 2 18 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.045
+ $Y=0.235 $X2=7.18 $Y2=0.39
r60 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.205
+ $Y=0.235 $X2=6.34 $Y2=0.39
.ends


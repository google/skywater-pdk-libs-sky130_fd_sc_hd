* File: sky130_fd_sc_hd__a2111oi_0.pex.spice
* Created: Tue Sep  1 18:50:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2111OI_0%D1 1 2 3 5 6 8 12 15 16 17 22
c36 15 0 1.12786e-19 $X=0.23 $Y=0.85
c37 12 0 3.19383e-20 $X=0.7 $Y=0.805
r38 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.35
+ $Y=0.93 $X2=0.35 $Y2=0.93
r39 16 17 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r40 16 23 8.56101 $w=3.48e-07 $l=2.6e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=0.93
r41 15 23 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=0.85 $X2=0.26
+ $Y2=0.93
r42 14 22 153.3 $w=2.7e-07 $l=6.9e-07 $layer=POLY_cond $X=0.35 $Y=1.62 $X2=0.35
+ $Y2=0.93
r43 10 22 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=0.35 $Y=0.88 $X2=0.35
+ $Y2=0.93
r44 10 12 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.35 $Y=0.805
+ $X2=0.7 $Y2=0.805
r45 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.77 $Y=1.77 $X2=0.77
+ $Y2=2.165
r46 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.7 $Y=0.73 $X2=0.7
+ $Y2=0.805
r47 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.7 $Y=0.73 $X2=0.7
+ $Y2=0.445
r48 2 14 29.8935 $w=1.5e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.485 $Y=1.695
+ $X2=0.35 $Y2=1.62
r49 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.695 $Y=1.695
+ $X2=0.77 $Y2=1.77
r50 1 2 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.695 $Y=1.695
+ $X2=0.485 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%C1 3 7 9 10 11 12 18
c38 18 0 1.03836e-19 $X=1.04 $Y=1.22
c39 7 0 1.52116e-19 $X=1.13 $Y=2.165
c40 3 0 1.12786e-19 $X=1.13 $Y=0.445
r41 18 21 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.04 $Y=1.22 $X2=1.04
+ $Y2=1.41
r42 18 20 44.4629 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=1.04 $Y=1.22
+ $X2=1.04 $Y2=1.065
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.22 $X2=1.04 $Y2=1.22
r44 11 12 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.14 $Y=1.87 $X2=1.14
+ $Y2=2.21
r45 10 11 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.14 $Y=1.53 $X2=1.14
+ $Y2=1.87
r46 10 19 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.14 $Y=1.53 $X2=1.14
+ $Y2=1.22
r47 9 19 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=1.14 $Y=1.19 $X2=1.14
+ $Y2=1.22
r48 7 21 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.13 $Y=2.165
+ $X2=1.13 $Y2=1.41
r49 3 20 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.13 $Y=0.445
+ $X2=1.13 $Y2=1.065
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%B1 3 7 9 10 14
r33 14 17 48.1856 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=1.595 $Y=1.22
+ $X2=1.595 $Y2=1.395
r34 14 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.22
+ $X2=1.595 $Y2=1.055
r35 9 10 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.67 $Y=1.19 $X2=1.67
+ $Y2=1.53
r36 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.22 $X2=1.61 $Y2=1.22
r37 7 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.63 $Y=0.445
+ $X2=1.63 $Y2=1.055
r38 3 17 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.49 $Y=2.165 $X2=1.49
+ $Y2=1.395
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%A1 1 3 6 9 15 16 17 18 23
c63 17 0 2.20172e-19 $X=2.53 $Y=1.19
r64 30 36 1.91462 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.49 $Y=1.4 $X2=2.49
+ $Y2=1.235
r65 26 36 1.91462 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.49 $Y=1.07
+ $X2=2.49 $Y2=1.235
r66 24 36 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=2.46 $Y=1.235 $X2=2.49
+ $Y2=1.235
r67 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.46
+ $Y=1.235 $X2=2.46 $Y2=1.235
r68 18 30 5.5488 $w=2.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.49 $Y=1.53 $X2=2.49
+ $Y2=1.4
r69 17 36 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.53 $Y=1.235 $X2=2.49
+ $Y2=1.235
r70 16 26 9.39028 $w=2.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.49 $Y=0.85
+ $X2=2.49 $Y2=1.07
r71 14 23 53.1961 $w=3.2e-07 $l=2.95e-07 $layer=POLY_cond $X=2.165 $Y=1.25
+ $X2=2.46 $Y2=1.25
r72 14 15 3.5291 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=2.165 $Y=1.25 $X2=2.075
+ $Y2=1.25
r73 9 10 61.9714 $w=1.75e-07 $l=1.55e-07 $layer=POLY_cond $X=2.075 $Y=1.682
+ $X2=1.92 $Y2=1.682
r74 8 15 33.9972 $w=1.65e-07 $l=1.6e-07 $layer=POLY_cond $X=2.075 $Y=1.41
+ $X2=2.075 $Y2=1.25
r75 8 9 71.9113 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=2.075 $Y=1.41
+ $X2=2.075 $Y2=1.595
r76 4 15 33.9972 $w=1.65e-07 $l=1.67332e-07 $layer=POLY_cond $X=2.06 $Y=1.09
+ $X2=2.075 $Y2=1.25
r77 4 6 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.06 $Y=1.09 $X2=2.06
+ $Y2=0.445
r78 1 10 6.48137 $w=1.5e-07 $l=8.8e-08 $layer=POLY_cond $X=1.92 $Y=1.77 $X2=1.92
+ $Y2=1.682
r79 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.92 $Y=1.77 $X2=1.92
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%A2 1 3 4 6 7 8 9 10 13 14 15 20
c48 10 0 1.507e-19 $X=2.525 $Y=1.695
r49 14 15 12.7108 $w=3.38e-07 $l=3.75e-07 $layer=LI1_cond $X=2.965 $Y=1.155
+ $X2=2.965 $Y2=1.53
r50 14 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.98
+ $Y=1.155 $X2=2.98 $Y2=1.155
r51 13 14 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=2.965 $Y=0.85
+ $X2=2.965 $Y2=1.155
r52 12 20 99.6211 $w=2.8e-07 $l=4.65e-07 $layer=POLY_cond $X=2.975 $Y=1.62
+ $X2=2.975 $Y2=1.155
r53 11 20 58.9157 $w=2.8e-07 $l=2.75e-07 $layer=POLY_cond $X=2.975 $Y=0.88
+ $X2=2.975 $Y2=1.155
r54 9 12 30.2628 $w=1.5e-07 $l=1.73494e-07 $layer=POLY_cond $X=2.835 $Y=1.695
+ $X2=2.975 $Y2=1.62
r55 9 10 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.835 $Y=1.695
+ $X2=2.525 $Y2=1.695
r56 7 11 30.2628 $w=1.5e-07 $l=1.73494e-07 $layer=POLY_cond $X=2.835 $Y=0.805
+ $X2=2.975 $Y2=0.88
r57 7 8 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.835 $Y=0.805
+ $X2=2.495 $Y2=0.805
r58 4 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.45 $Y=1.77
+ $X2=2.525 $Y2=1.695
r59 4 6 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.45 $Y=1.77 $X2=2.45
+ $Y2=2.165
r60 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.42 $Y=0.73
+ $X2=2.495 $Y2=0.805
r61 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.42 $Y=0.73 $X2=2.42
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%Y 1 2 3 12 14 15 18 20 21 22 23 24 49
c52 14 0 1.03836e-19 $X=1.71 $Y=0.75
r53 49 50 5.13628 $w=4.23e-07 $l=4.5e-08 $layer=LI1_cond $X=0.572 $Y=1.87
+ $X2=0.572 $Y2=1.825
r54 46 47 10.1433 $w=2.61e-07 $l=2.17e-07 $layer=LI1_cond $X=0.695 $Y=0.75
+ $X2=0.912 $Y2=0.75
r55 40 53 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=0.572 $Y=2.037
+ $X2=0.572 $Y2=1.99
r56 32 46 2.91302 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=0.695 $Y=0.885
+ $X2=0.695 $Y2=0.75
r57 24 40 4.69112 $w=4.23e-07 $l=1.73e-07 $layer=LI1_cond $X=0.572 $Y=2.21
+ $X2=0.572 $Y2=2.037
r58 23 53 2.71163 $w=4.23e-07 $l=1e-07 $layer=LI1_cond $X=0.572 $Y=1.89
+ $X2=0.572 $Y2=1.99
r59 23 49 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=0.572 $Y=1.89
+ $X2=0.572 $Y2=1.87
r60 23 50 1.23232 $w=1.78e-07 $l=2e-08 $layer=LI1_cond $X=0.695 $Y=1.805
+ $X2=0.695 $Y2=1.825
r61 22 23 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.805
r62 21 22 20.9495 $w=1.78e-07 $l=3.4e-07 $layer=LI1_cond $X=0.695 $Y=1.19
+ $X2=0.695 $Y2=1.53
r63 20 46 0.233716 $w=2.61e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=0.75
+ $X2=0.695 $Y2=0.75
r64 20 21 17.2525 $w=1.78e-07 $l=2.8e-07 $layer=LI1_cond $X=0.695 $Y=0.91
+ $X2=0.695 $Y2=1.19
r65 20 32 1.5404 $w=1.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.695 $Y=0.91
+ $X2=0.695 $Y2=0.885
r66 16 18 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.875 $Y=0.615
+ $X2=1.875 $Y2=0.445
r67 15 47 5.7837 $w=2.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.04 $Y=0.75
+ $X2=0.912 $Y2=0.75
r68 14 16 6.90553 $w=2.7e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.71 $Y=0.75
+ $X2=1.875 $Y2=0.615
r69 14 15 28.5977 $w=2.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.71 $Y=0.75
+ $X2=1.04 $Y2=0.75
r70 10 47 0.881292 $w=2.55e-07 $l=1.35e-07 $layer=LI1_cond $X=0.912 $Y=0.615
+ $X2=0.912 $Y2=0.75
r71 10 12 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=0.912 $Y=0.615
+ $X2=0.912 $Y2=0.42
r72 3 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.4
+ $Y=1.845 $X2=0.525 $Y2=1.99
r73 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.235 $X2=1.845 $Y2=0.445
r74 1 12 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.235 $X2=0.915 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%A_313_369# 1 2 9 11 13 16
c29 16 0 1.52116e-19 $X=1.705 $Y=1.99
c30 11 0 3.47928e-20 $X=2.705 $Y=2.085
r31 11 18 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.705 $Y=2.085
+ $X2=2.705 $Y2=1.995
r32 11 13 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.705 $Y=2.085
+ $X2=2.705 $Y2=2.33
r33 10 16 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=1.995
+ $X2=1.705 $Y2=1.995
r34 9 18 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=1.995
+ $X2=2.705 $Y2=1.995
r35 9 10 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.54 $Y=1.995
+ $X2=1.87 $Y2=1.995
r36 2 18 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.845 $X2=2.705 $Y2=1.99
r37 2 13 600 $w=1.7e-07 $l=5.67913e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.845 $X2=2.705 $Y2=2.33
r38 1 16 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.845 $X2=1.705 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%VPWR 1 6 8 10 17 18 21
r36 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r39 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=2.72
+ $X2=2.205 $Y2=2.72
r40 15 17 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.37 $Y=2.72
+ $X2=2.99 $Y2=2.72
r41 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=2.72
+ $X2=2.205 $Y2=2.72
r42 10 12 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.04 $Y=2.72
+ $X2=0.23 $Y2=2.72
r43 8 22 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 8 12 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r45 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2.72
r46 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.205 $Y=2.635
+ $X2=2.205 $Y2=2.34
r47 1 6 600 $w=1.7e-07 $l=5.90741e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.845 $X2=2.205 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_0%VGND 1 2 3 12 16 20 23 24 26 27 28 36 42
+ 43 46
c53 26 0 3.19383e-20 $X=1.21 $Y=0
c54 20 0 3.46791e-20 $X=2.635 $Y=0.36
r55 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r56 43 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r57 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r58 40 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.635
+ $Y2=0
r59 40 42 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.99
+ $Y2=0
r60 39 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r61 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r62 36 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.635
+ $Y2=0
r63 36 38 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=1.61
+ $Y2=0
r64 35 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r65 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r66 28 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r67 28 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r68 26 34 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.21 $Y=0 $X2=1.15
+ $Y2=0
r69 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=0 $X2=1.375
+ $Y2=0
r70 25 38 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.54 $Y=0 $X2=1.61
+ $Y2=0
r71 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=1.375
+ $Y2=0
r72 23 31 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.23
+ $Y2=0
r73 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.45
+ $Y2=0
r74 22 34 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=1.15
+ $Y2=0
r75 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.45
+ $Y2=0
r76 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0
r77 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0.36
r78 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0
r79 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0.36
r80 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.45 $Y=0.085
+ $X2=0.45 $Y2=0
r81 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.45 $Y=0.085
+ $X2=0.45 $Y2=0.38
r82 3 20 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.635 $Y2=0.36
r83 2 16 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=1.205
+ $Y=0.235 $X2=1.375 $Y2=0.36
r84 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.235 $X2=0.45 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__fah_1.spice
* Created: Thu Aug 27 14:21:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__fah_1.spice.pex"
.subckt sky130_fd_sc_hd__fah_1  VNB VPB A B CI VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1029 N_VGND_M1029_d N_A_67_199#_M1029_g N_A_27_47#_M1029_s VNB NSHORT L=0.15
+ W=0.65 AD=0.106066 AS=0.169 PD=0.982558 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1031 N_A_67_199#_M1031_d N_A_M1031_g N_VGND_M1029_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1664 AS=0.104434 PD=1.8 PS=0.967442 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_310_49#_M1018_s VNB NSHORT L=0.15 W=0.64
+ AD=0.169947 AS=0.1664 PD=1.17085 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1000 N_A_508_297#_M1000_d N_B_M1000_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17 AS=0.172603 PD=1.86 PS=1.18915 NRD=0 NRS=47.076 M=1 R=4.33333
+ SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1027 N_A_719_47#_M1027_d N_B_M1027_g N_A_310_49#_M1027_s VNB NSHORT L=0.15
+ W=0.64 AD=0.088 AS=0.16285 PD=0.915 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_27_47#_M1013_d N_A_508_297#_M1013_g N_A_719_47#_M1027_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2176 AS=0.088 PD=1.96 PS=0.915 NRD=14.052 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1002 N_A_1008_47#_M1002_d N_A_508_297#_M1002_g N_A_310_49#_M1002_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.189675 AS=0.1664 PD=1.24 PS=1.8 NRD=47.808 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1014 N_A_27_47#_M1014_d N_B_M1014_g N_A_1008_47#_M1002_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1664 AS=0.189675 PD=1.8 PS=1.24 NRD=0 NRS=10.308 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_1332_297#_M1004_d N_A_719_47#_M1004_g N_A_1262_49#_M1004_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.088 AS=0.1664 PD=0.915 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_508_297#_M1021_d N_A_1008_47#_M1021_g N_A_1332_297#_M1004_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1664 AS=0.088 PD=1.8 PS=0.915 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_1617_49#_M1009_d N_A_1008_47#_M1009_g N_A_1262_49#_M1009_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0928 AS=0.1664 PD=0.93 PS=1.8 NRD=2.808 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_1640_380#_M1003_d N_A_719_47#_M1003_g N_A_1617_49#_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1792 AS=0.0928 PD=1.84 PS=0.93 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_VGND_M1024_d N_CI_M1024_g N_A_1262_49#_M1024_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.1728 PD=0.91 PS=1.82 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1028 N_A_1640_380#_M1028_d N_A_1262_49#_M1028_g N_VGND_M1024_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_A_1332_297#_M1011_g N_COUT_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.1755 PD=0.92 PS=1.84 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1017 N_SUM_M1017_d N_A_1617_49#_M1017_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.65 AD=0.221 AS=0.08775 PD=1.98 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_67_199#_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.28 PD=1.3 PS=2.56 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1007 N_A_67_199#_M1007_d N_A_M1007_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.15 PD=2.52 PS=1.3 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7 SB=75000.2
+ A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_310_49#_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2075 AS=0.275 PD=1.415 PS=2.55 NRD=22.6353 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1012 N_A_508_297#_M1012_d N_B_M1012_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.2075 PD=2.52 PS=1.415 NRD=0 NRS=3.9203 M=1 R=6.66667 SA=75000.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1023 N_A_719_47#_M1023_d N_B_M1023_g N_A_27_47#_M1023_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1155 AS=0.3594 PD=1.115 PS=2.8 NRD=0 NRS=87.4286 M=1 R=5.6
+ SA=75000.3 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_A_310_49#_M1010_d N_A_508_297#_M1010_g N_A_719_47#_M1023_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2184 AS=0.1155 PD=2.2 PS=1.115 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 N_A_1008_47#_M1022_d N_A_508_297#_M1022_g N_A_27_47#_M1022_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.152262 AS=0.323 PD=1.3 PS=2.73 NRD=0 NRS=7.0329 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1020 N_A_310_49#_M1020_d N_B_M1020_g N_A_1008_47#_M1022_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2184 AS=0.152262 PD=2.2 PS=1.3 NRD=0 NRS=14.0658 M=1 R=5.6
+ SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1026 N_A_1332_297#_M1026_d N_A_719_47#_M1026_g N_A_508_297#_M1026_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1134 AS=0.2562 PD=1.11 PS=2.29 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_1262_49#_M1008_d N_A_1008_47#_M1008_g N_A_1332_297#_M1026_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.711425 AS=0.1134 PD=3.4 PS=1.11 NRD=139.535 NRS=0
+ M=1 R=5.6 SA=75000.6 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1019 N_A_1617_49#_M1019_d N_A_1008_47#_M1019_g N_A_1640_380#_M1019_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1134 AS=0.21515 PD=1.11 PS=2.2 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1016 N_A_1262_49#_M1016_d N_A_719_47#_M1016_g N_A_1617_49#_M1019_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.310686 AS=0.1134 PD=1.57957 PS=1.11 NRD=75.6283 NRS=0 M=1
+ R=5.6 SA=75000.6 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1025 N_VPWR_M1025_d N_CI_M1025_g N_A_1262_49#_M1016_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.369864 PD=1.27 PS=1.88043 NRD=0 NRS=18.2225 M=1 R=6.66667
+ SA=75001.3 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_1640_380#_M1005_d N_A_1262_49#_M1005_g N_VPWR_M1025_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_1332_297#_M1001_g N_COUT_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1030 N_SUM_M1030_d N_A_1617_49#_M1030_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.135 PD=2.57 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.544 P=28.81
pX33_noxref noxref_20 B B PROBETYPE=1
c_118 VNB 0 2.31345e-19 $X=0.145 $Y=-0.085
c_235 VPB 0 6.77358e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__fah_1.spice.SKY130_FD_SC_HD__FAH_1.pxi"
*
.ends
*
*

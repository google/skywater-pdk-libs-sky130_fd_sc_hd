* File: sky130_fd_sc_hd__maj3_4.spice
* Created: Thu Aug 27 14:27:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__maj3_4.spice.pex"
.subckt sky130_fd_sc_hd__maj3_4  VNB VPB C A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C	C
* VPB	VPB
* VNB	VNB
MM1002 A_151_47# N_C_M1002_g N_A_47_297#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.079625 AS=0.182 PD=0.895 PS=1.86 NRD=12.456 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g A_151_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.079625 PD=0.92 PS=0.895 NRD=0 NRS=12.456 M=1 R=4.33333 SA=75000.6
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1012 A_314_47# N_A_M1012_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001 SB=75003.3
+ A=0.0975 P=1.6 MULT=1
MM1015 N_A_47_297#_M1015_d N_B_M1015_g A_314_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75001.4
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1014 A_482_47# N_B_M1014_g N_A_47_297#_M1015_d VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.08775 PD=0.86 PS=0.92 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_C_M1016_g A_482_47# VNB NSHORT L=0.15 W=0.65 AD=0.157625
+ AS=0.06825 PD=1.135 PS=0.86 NRD=21.228 NRS=9.228 M=1 R=4.33333 SA=75002.2
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1016_d N_A_47_297#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.157625 AS=0.08775 PD=1.135 PS=0.92 NRD=16.608 NRS=0 M=1 R=4.33333
+ SA=75002.9 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_47_297#_M1005_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1005_d N_A_47_297#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A_47_297#_M1018_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 A_151_297# N_C_M1011_g N_A_47_297#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1225 AS=0.37 PD=1.245 PS=2.74 NRD=13.2778 NRS=16.7253 M=1 R=6.66667
+ SA=75000.3 SB=75004.1 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g A_151_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.1225 PD=1.27 PS=1.245 NRD=0 NRS=13.2778 M=1 R=6.66667 SA=75000.7
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1008 A_314_297# N_A_M1008_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75001.1 SB=75003.3
+ A=0.15 P=2.3 MULT=1
MM1004 N_A_47_297#_M1004_d N_B_M1004_g A_314_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75001.5
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1019 A_482_297# N_B_M1019_g N_A_47_297#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.135 PD=1.21 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g A_482_297# VPB PHIGHVT L=0.15 W=1 AD=0.2425
+ AS=0.105 PD=1.485 PS=1.21 NRD=19.6803 NRS=9.8303 M=1 R=6.66667 SA=75002.3
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1001_d N_A_47_297#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2425 AS=0.135 PD=1.485 PS=1.27 NRD=20.685 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_47_297#_M1006_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1006_d N_A_47_297#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_47_297#_M1010_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=8.7312 P=14.09
c_44 VNB 0 1.11508e-19 $X=0.14 $Y=-0.085
c_528 A_314_297# 0 1.01236e-19 $X=1.57 $Y=1.485
*
.include "sky130_fd_sc_hd__maj3_4.spice.SKY130_FD_SC_HD__MAJ3_4.pxi"
*
.ends
*
*

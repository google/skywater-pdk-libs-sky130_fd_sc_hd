* File: sky130_fd_sc_hd__lpflow_decapkapwr_6.pex.spice
* Created: Tue Sep  1 19:11:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%VGND 1 7 9 12 15 23 26 29
r22 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r23 26 28 0.445255 $w=8.22e-07 $l=3e-08 $layer=LI1_cond $X=2.5 $Y=0.385 $X2=2.53
+ $Y2=0.385
r24 21 23 0.900738 $w=1.219e-06 $l=9e-08 $layer=LI1_cond $X=0.647 $Y=0.385
+ $X2=0.647 $Y2=0.475
r25 20 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r26 17 21 3.85316 $w=1.219e-06 $l=3.85e-07 $layer=LI1_cond $X=0.647 $Y=0
+ $X2=0.647 $Y2=0.385
r27 17 20 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r28 13 23 8.15669 $w=1.219e-06 $l=8.15e-07 $layer=LI1_cond $X=0.647 $Y=1.29
+ $X2=0.647 $Y2=0.475
r29 12 15 21.4725 $w=1.706e-06 $l=8.8476e-07 $layer=POLY_cond $X=1.11 $Y=1.29
+ $X2=1.38 $Y2=2.05
r30 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.11
+ $Y=1.29 $X2=1.11 $Y2=1.29
r31 9 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r32 9 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r33 8 21 2.26174 $w=9.4e-07 $l=6.48e-07 $layer=LI1_cond $X=1.295 $Y=0.385
+ $X2=0.647 $Y2=0.385
r34 7 26 4.05283 $w=9.4e-07 $l=2.95e-07 $layer=LI1_cond $X=2.205 $Y=0.385
+ $X2=2.5 $Y2=0.385
r35 7 8 11.8106 $w=9.38e-07 $l=9.1e-07 $layer=LI1_cond $X=2.205 $Y=0.385
+ $X2=1.295 $Y2=0.385
r36 1 26 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=2.365 $Y=0.235
+ $X2=2.5 $Y2=0.475
r37 1 23 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%KAPWR 1 9 12 16 17 18 20 34 36
+ 38
r28 36 38 0.0085136 $w=2.6e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=2.21
+ $X2=0.23 $Y2=2.21
r29 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.21
+ $X2=2.53 $Y2=2.21
r30 31 33 2.06694 $w=1.208e-06 $l=2.05e-07 $layer=LI1_cond $X=2.07 $Y=2.005
+ $X2=2.07 $Y2=2.21
r31 30 31 1.76446 $w=1.208e-06 $l=1.75e-07 $layer=LI1_cond $X=2.07 $Y=1.83
+ $X2=2.07 $Y2=2.005
r32 22 26 0.397826 $w=9.18e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=2.005
+ $X2=0.26 $Y2=2.005
r33 22 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.21
+ $X2=0.23 $Y2=2.21
r34 20 31 2.34412 $w=9.2e-07 $l=6.05e-07 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=2.07 $Y2=2.005
r35 20 26 15.9793 $w=9.18e-07 $l=1.205e-06 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=0.26 $Y2=2.005
r36 17 30 7.2595 $w=1.208e-06 $l=7.2e-07 $layer=LI1_cond $X=2.07 $Y=1.11
+ $X2=2.07 $Y2=1.83
r37 16 18 36.3375 $w=1.17e-06 $l=7.15e-07 $layer=POLY_cond $X=2.2 $Y=0.69
+ $X2=1.485 $Y2=0.69
r38 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.2 $Y=1.11
+ $X2=2.2 $Y2=1.11
r39 12 36 0.0120192 $w=2.6e-07 $l=2.5e-08 $layer=MET1_cond $X=0.19 $Y=2.21
+ $X2=0.215 $Y2=2.21
r40 12 34 1.27874 $w=2.6e-07 $l=2.253e-06 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=2.53 $Y2=2.21
r41 12 38 0.0266759 $w=2.6e-07 $l=4.7e-08 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=0.23 $Y2=2.21
r42 9 18 6.24815 $w=8.1e-07 $l=1.05e-07 $layer=POLY_cond $X=1.38 $Y=0.51
+ $X2=1.485 $Y2=0.51
r43 1 30 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.615 $X2=2.5 $Y2=1.83
r44 1 26 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_6%VPWR 1 8 9
r13 8 9 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72 $X2=2.53
+ $Y2=2.72
r14 4 8 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r15 1 9 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r16 1 4 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends


* File: sky130_fd_sc_hd__clkdlybuf4s50_2.pex.spice
* Created: Tue Sep  1 19:01:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A 3 7 9 15
r30 12 15 34.1305 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.315 $Y=1.16
+ $X2=0.48 $Y2=1.16
r31 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=1.16 $X2=0.315 $Y2=1.16
r32 5 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.48 $Y=1.305
+ $X2=0.48 $Y2=1.16
r33 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.48 $Y=1.305 $X2=0.48
+ $Y2=1.985
r34 1 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.48 $Y=1.015
+ $X2=0.48 $Y2=1.16
r35 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.48 $Y=1.015 $X2=0.48
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_27_47# 1 2 9 13 17 21 23 24 25 26
+ 29 30
c66 30 0 3.32424e-19 $X=1.27 $Y=1.16
c67 29 0 2.17216e-19 $X=1.27 $Y=1.16
c68 13 0 1.48431e-19 $X=1.165 $Y=2.075
c69 9 0 1.48431e-19 $X=1.165 $Y=0.56
r70 30 34 14.3413 $w=6.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.1
+ $Y2=1.295
r71 30 33 14.3413 $w=6.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.1
+ $Y2=1.025
r72 29 31 9.97944 $w=4.67e-07 $l=3.82e-07 $layer=LI1_cond $X=1.1 $Y=1.16 $X2=1.1
+ $Y2=1.542
r73 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r74 27 29 8.88223 $w=4.67e-07 $l=3.4e-07 $layer=LI1_cond $X=1.1 $Y=0.82 $X2=1.1
+ $Y2=1.16
r75 25 31 6.56345 $w=1.75e-07 $l=2.5e-07 $layer=LI1_cond $X=0.85 $Y=1.542
+ $X2=1.1 $Y2=1.542
r76 25 26 26.6182 $w=1.73e-07 $l=4.2e-07 $layer=LI1_cond $X=0.85 $Y=1.542
+ $X2=0.43 $Y2=1.542
r77 23 27 6.73017 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.85 $Y=0.82 $X2=1.1
+ $Y2=0.82
r78 23 24 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.85 $Y=0.82
+ $X2=0.415 $Y2=0.82
r79 19 26 7.80978 $w=1.75e-07 $l=2.12492e-07 $layer=LI1_cond $X=0.257 $Y=1.63
+ $X2=0.43 $Y2=1.542
r80 19 21 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=1.63
+ $X2=0.257 $Y2=1.965
r81 15 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.25 $Y=0.735
+ $X2=0.415 $Y2=0.82
r82 15 17 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.25 $Y=0.735
+ $X2=0.25 $Y2=0.47
r83 13 34 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.165 $Y=2.075
+ $X2=1.165 $Y2=1.295
r84 9 33 49.7577 $w=5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.165 $Y=0.56
+ $X2=1.165 $Y2=1.025
r85 2 21 300 $w=1.7e-07 $l=5.4111e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.265 $Y2=1.965
r86 1 17 182 $w=1.7e-07 $l=2.92874e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_283_47# 1 2 9 13 19 22 27 28 31 32
+ 33 34
c66 28 0 5.23118e-19 $X=2.14 $Y=1.16
r67 31 32 9.09563 $w=4.03e-07 $l=1.8e-07 $layer=LI1_cond $X=1.592 $Y=1.965
+ $X2=1.592 $Y2=1.785
r68 28 37 15.4315 $w=7.35e-07 $l=1.45e-07 $layer=POLY_cond $X=2.342 $Y=1.16
+ $X2=2.342 $Y2=1.305
r69 28 36 15.4315 $w=7.35e-07 $l=1.45e-07 $layer=POLY_cond $X=2.342 $Y=1.16
+ $X2=2.342 $Y2=1.015
r70 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r71 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=1.16
+ $X2=1.71 $Y2=1.16
r72 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.795 $Y=1.16
+ $X2=2.14 $Y2=1.16
r73 23 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.245
+ $X2=1.71 $Y2=1.16
r74 23 32 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.71 $Y=1.245
+ $X2=1.71 $Y2=1.785
r75 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.075
+ $X2=1.71 $Y2=1.16
r76 22 33 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.71 $Y=1.075
+ $X2=1.71 $Y2=0.9
r77 17 33 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=1.617 $Y=0.723
+ $X2=1.617 $Y2=0.9
r78 17 19 9.3494 $w=3.53e-07 $l=2.88e-07 $layer=LI1_cond $X=1.617 $Y=0.723
+ $X2=1.617 $Y2=0.435
r79 13 37 82.3945 $w=5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.46 $Y=2.075 $X2=2.46
+ $Y2=1.305
r80 9 36 48.6877 $w=5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.46 $Y=0.56 $X2=2.46
+ $Y2=1.015
r81 2 31 300 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.665 $X2=1.555 $Y2=1.965
r82 1 19 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%A_390_47# 1 2 9 13 15 16 19 23 25 28
+ 32 34 35 36 37 40 43
r84 41 50 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.055 $Y=1.16
+ $X2=3.115 $Y2=1.16
r85 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.055
+ $Y=1.16 $X2=3.055 $Y2=1.16
r86 38 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.56 $Y=1.16
+ $X2=2.56 $Y2=1.545
r87 38 43 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.56 $Y=1.16
+ $X2=2.56 $Y2=0.82
r88 38 40 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.645 $Y=1.16
+ $X2=3.055 $Y2=1.16
r89 36 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=1.545
+ $X2=2.56 $Y2=1.545
r90 36 37 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.475 $Y=1.545
+ $X2=2.235 $Y2=1.545
r91 34 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.82
+ $X2=2.56 $Y2=0.82
r92 34 35 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.475 $Y=0.82
+ $X2=2.235 $Y2=0.82
r93 30 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.11 $Y=1.63
+ $X2=2.235 $Y2=1.545
r94 30 32 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=2.11 $Y=1.63
+ $X2=2.11 $Y2=1.96
r95 26 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.11 $Y=0.735
+ $X2=2.235 $Y2=0.82
r96 26 28 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.11 $Y=0.735
+ $X2=2.11 $Y2=0.47
r97 21 25 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.54 $Y=1.295
+ $X2=3.54 $Y2=1.16
r98 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.54 $Y=1.295
+ $X2=3.54 $Y2=1.985
r99 17 25 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.54 $Y=1.025
+ $X2=3.54 $Y2=1.16
r100 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.54 $Y=1.025
+ $X2=3.54 $Y2=0.445
r101 16 50 15.1926 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.19 $Y=1.16
+ $X2=3.115 $Y2=1.16
r102 15 25 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.465 $Y=1.16
+ $X2=3.54 $Y2=1.16
r103 15 16 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=3.465 $Y=1.16
+ $X2=3.19 $Y2=1.16
r104 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.325
+ $X2=3.115 $Y2=1.16
r105 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.115 $Y=1.325
+ $X2=3.115 $Y2=1.985
r106 7 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=0.995
+ $X2=3.115 $Y2=1.16
r107 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.115 $Y=0.995
+ $X2=3.115 $Y2=0.445
r108 2 32 300 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=2 $X=1.95
+ $Y=1.665 $X2=2.075 $Y2=1.96
r109 1 28 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.235 $X2=2.075 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%VPWR 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
c45 12 0 1.60901e-19 $X=0.765 $Y=1.965
r46 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r47 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r49 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r50 39 47 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.795 $Y=2.72
+ $X2=3.967 $Y2=2.72
r51 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.795 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.765 $Y2=2.72
r59 32 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.765 $Y2=2.72
r61 27 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r62 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 23 37 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.685 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=2.72
+ $X2=2.85 $Y2=2.72
r66 22 41 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.015 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.72
+ $X2=2.85 $Y2=2.72
r68 18 47 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.925 $Y=2.635
+ $X2=3.967 $Y2=2.72
r69 18 20 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=3.925 $Y=2.635
+ $X2=3.925 $Y2=1.965
r70 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=2.635
+ $X2=2.85 $Y2=2.72
r71 14 16 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.85 $Y=2.635
+ $X2=2.85 $Y2=1.965
r72 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2.72
r73 10 12 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=1.965
r74 3 20 300 $w=1.7e-07 $l=5.97997e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=1.485 $X2=3.88 $Y2=1.965
r75 2 16 300 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=2 $X=2.71
+ $Y=1.665 $X2=2.85 $Y2=1.965
r76 1 12 300 $w=1.7e-07 $l=5.755e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.765 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%X 1 2 7 8 9 10 11 12 28 42
c26 8 0 9.5523e-20 $X=3.475 $Y=0.85
r27 20 42 2.37163 $w=2.8e-07 $l=1.85e-07 $layer=LI1_cond $X=3.485 $Y=0.64
+ $X2=3.485 $Y2=0.455
r28 12 33 6.54797 $w=4.38e-07 $l=2.5e-07 $layer=LI1_cond $X=3.405 $Y=2.21
+ $X2=3.405 $Y2=1.96
r29 11 33 2.35727 $w=4.38e-07 $l=9e-08 $layer=LI1_cond $X=3.405 $Y=1.87
+ $X2=3.405 $Y2=1.96
r30 11 29 3.14303 $w=4.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.405 $Y=1.87
+ $X2=3.405 $Y2=1.75
r31 10 29 4.66216 $w=4.38e-07 $l=1.78e-07 $layer=LI1_cond $X=3.405 $Y=1.572
+ $X2=3.405 $Y2=1.75
r32 10 28 1.10006 $w=4.38e-07 $l=4.2e-08 $layer=LI1_cond $X=3.405 $Y=1.572
+ $X2=3.405 $Y2=1.53
r33 10 28 1.76982 $w=2.78e-07 $l=4.3e-08 $layer=LI1_cond $X=3.485 $Y=1.487
+ $X2=3.485 $Y2=1.53
r34 9 10 12.2241 $w=2.78e-07 $l=2.97e-07 $layer=LI1_cond $X=3.485 $Y=1.19
+ $X2=3.485 $Y2=1.487
r35 8 9 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.485 $Y=0.85 $X2=3.485
+ $Y2=1.19
r36 8 20 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=3.485 $Y=0.85
+ $X2=3.485 $Y2=0.64
r37 7 42 0.311471 $w=3.68e-07 $l=1e-08 $layer=LI1_cond $X=3.475 $Y=0.455
+ $X2=3.485 $Y2=0.455
r38 7 38 4.51633 $w=3.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.475 $Y=0.455
+ $X2=3.33 $Y2=0.455
r39 2 33 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=3.19
+ $Y=1.485 $X2=3.33 $Y2=1.96
r40 1 38 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.235 $X2=3.33 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S50_2%VGND 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
c51 12 0 1.71523e-19 $X=0.75 $Y=0.425
c52 1 0 8.64836e-20 $X=0.555 $Y=0.235
r53 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r54 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r55 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r56 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r57 39 47 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.967
+ $Y2=0
r58 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.45
+ $Y2=0
r59 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r60 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r61 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r62 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r63 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r64 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r65 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r66 32 34 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.15
+ $Y2=0
r67 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r68 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.23
+ $Y2=0
r69 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r70 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 23 37 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.53
+ $Y2=0
r72 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.85
+ $Y2=0
r73 22 41 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.45
+ $Y2=0
r74 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.85
+ $Y2=0
r75 18 47 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.967 $Y2=0
r76 18 20 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.47
r77 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=0.085
+ $X2=2.85 $Y2=0
r78 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.85 $Y=0.085
+ $X2=2.85 $Y2=0.4
r79 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r80 10 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.425
r81 3 20 182 $w=1.7e-07 $l=3.64005e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.235 $X2=3.88 $Y2=0.47
r82 2 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.235 $X2=2.85 $Y2=0.4
r83 1 12 182 $w=1.7e-07 $l=2.73998e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.75 $Y2=0.425
.ends


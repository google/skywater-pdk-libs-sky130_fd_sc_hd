* File: sky130_fd_sc_hd__or4_4.pex.spice
* Created: Tue Sep  1 19:28:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4_4%D 1 3 6 8 9 16
r33 13 16 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.285 $Y=1.16
+ $X2=0.495 $Y2=1.16
r34 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.285
+ $Y=1.16 $X2=0.285 $Y2=1.16
r35 8 9 12.5353 $w=2.83e-07 $l=3.1e-07 $layer=LI1_cond $X=0.227 $Y=0.85
+ $X2=0.227 $Y2=1.16
r36 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r37 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.985
r38 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_4%C 3 6 10 11 13 14 19 23
r48 21 23 2.46952 $w=3.48e-07 $l=7.5e-08 $layer=LI1_cond $X=1.055 $Y=1.795
+ $X2=1.055 $Y2=1.87
r49 13 21 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=1.055 $Y=1.79
+ $X2=1.055 $Y2=1.795
r50 13 29 8.65312 $w=3.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.055 $Y=1.79
+ $X2=1.055 $Y2=1.62
r51 13 14 11.0305 $w=3.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=1.875
+ $X2=1.055 $Y2=2.21
r52 13 23 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=1.055 $Y=1.875
+ $X2=1.055 $Y2=1.87
r53 11 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=0.965 $Y2=1.325
r54 11 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=0.965 $Y2=0.995
r55 10 29 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.965 $Y=1.16
+ $X2=0.965 $Y2=1.62
r56 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.16 $X2=0.965 $Y2=1.16
r57 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.025 $Y=1.985
+ $X2=1.025 $Y2=1.325
r58 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.025 $Y=0.56
+ $X2=1.025 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_4%B 1 3 6 10 11 14 15 31
c40 11 0 5.72837e-20 $X=1.445 $Y=1.16
c41 6 0 2.99791e-19 $X=1.445 $Y=1.985
r42 21 31 2.70104 $w=3.18e-07 $l=7.5e-08 $layer=LI1_cond $X=1.56 $Y=1.945
+ $X2=1.56 $Y2=1.87
r43 14 31 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=1.56 $Y=1.865
+ $X2=1.56 $Y2=1.87
r44 14 15 9.3636 $w=3.18e-07 $l=2.6e-07 $layer=LI1_cond $X=1.56 $Y=1.95 $X2=1.56
+ $Y2=2.21
r45 14 21 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=1.56 $Y=1.95 $X2=1.56
+ $Y2=1.945
r46 13 14 13.9192 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=1.505 $Y=1.45
+ $X2=1.505 $Y2=1.785
r47 10 13 11.6456 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.445 $Y=1.16
+ $X2=1.445 $Y2=1.45
r48 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=1.16 $X2=1.445 $Y2=1.16
r49 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.325
+ $X2=1.445 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.445 $Y=1.325
+ $X2=1.445 $Y2=1.985
r51 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.445 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.445 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_4%A 3 6 8 12 13 14
c41 13 0 1.24234e-19 $X=1.925 $Y=1.16
c42 8 0 1.75557e-19 $X=2.065 $Y=1.53
r43 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.16
+ $X2=1.925 $Y2=1.325
r44 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.16
+ $X2=1.925 $Y2=0.995
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.16 $X2=1.925 $Y2=1.16
r46 8 20 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.065 $Y=1.53
+ $X2=1.925 $Y2=1.53
r47 8 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.925 $Y=1.445
+ $X2=1.925 $Y2=1.53
r48 8 13 16.0859 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=1.925 $Y=1.445
+ $X2=1.925 $Y2=1.16
r49 6 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.865 $Y=1.985
+ $X2=1.865 $Y2=1.325
r50 3 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.865 $Y=0.56
+ $X2=1.865 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_4%A_32_297# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 40 43 46 48 49 52 54 57 58 63 69 74 81
c139 74 0 5.72837e-20 $X=1.655 $Y=0.74
c140 54 0 1.60701e-19 $X=2.18 $Y=0.74
r141 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.815 $Y=1.16
+ $X2=3.235 $Y2=1.16
r142 71 73 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.625 $Y=0.74
+ $X2=0.785 $Y2=0.74
r143 64 81 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.475 $Y=1.16
+ $X2=3.655 $Y2=1.16
r144 64 79 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.475 $Y=1.16
+ $X2=3.235 $Y2=1.16
r145 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.475
+ $Y=1.16 $X2=3.475 $Y2=1.16
r146 61 78 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.455 $Y=1.16
+ $X2=2.815 $Y2=1.16
r147 61 75 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.455 $Y=1.16
+ $X2=2.395 $Y2=1.16
r148 60 63 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.455 $Y=1.16
+ $X2=3.475 $Y2=1.16
r149 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.455
+ $Y=1.16 $X2=2.455 $Y2=1.16
r150 58 60 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.35 $Y=1.16
+ $X2=2.455 $Y2=1.16
r151 57 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=1.075
+ $X2=2.35 $Y2=1.16
r152 56 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.265 $Y=0.825
+ $X2=2.265 $Y2=1.075
r153 55 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.74
+ $X2=1.655 $Y2=0.74
r154 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.18 $Y=0.74
+ $X2=2.265 $Y2=0.825
r155 54 55 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.18 $Y=0.74
+ $X2=1.74 $Y2=0.74
r156 50 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.655
+ $X2=1.655 $Y2=0.74
r157 50 52 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=0.655
+ $X2=1.655 $Y2=0.49
r158 49 73 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=0.74
+ $X2=0.785 $Y2=0.74
r159 48 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.74
+ $X2=1.655 $Y2=0.74
r160 48 49 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.57 $Y=0.74 $X2=0.87
+ $Y2=0.74
r161 44 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.655
+ $X2=0.785 $Y2=0.74
r162 44 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=0.655
+ $X2=0.785 $Y2=0.49
r163 43 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.625 $Y=1.495
+ $X2=0.625 $Y2=1.58
r164 42 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.625 $Y=0.825
+ $X2=0.625 $Y2=0.74
r165 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.625 $Y=0.825
+ $X2=0.625 $Y2=1.495
r166 38 69 22.3775 $w=1.68e-07 $l=3.43e-07 $layer=LI1_cond $X=0.282 $Y=1.58
+ $X2=0.625 $Y2=1.58
r167 38 40 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=2.34
r168 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.325
+ $X2=3.655 $Y2=1.16
r169 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.655 $Y=1.325
+ $X2=3.655 $Y2=1.985
r170 31 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=0.995
+ $X2=3.655 $Y2=1.16
r171 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.655 $Y=0.995
+ $X2=3.655 $Y2=0.56
r172 27 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.325
+ $X2=3.235 $Y2=1.16
r173 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.235 $Y=1.325
+ $X2=3.235 $Y2=1.985
r174 24 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=0.995
+ $X2=3.235 $Y2=1.16
r175 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.235 $Y=0.995
+ $X2=3.235 $Y2=0.56
r176 20 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.325
+ $X2=2.815 $Y2=1.16
r177 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.815 $Y=1.325
+ $X2=2.815 $Y2=1.985
r178 17 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=0.995
+ $X2=2.815 $Y2=1.16
r179 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.815 $Y=0.995
+ $X2=2.815 $Y2=0.56
r180 13 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.325
+ $X2=2.395 $Y2=1.16
r181 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.395 $Y=1.325
+ $X2=2.395 $Y2=1.985
r182 10 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.395 $Y2=1.16
r183 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.395 $Y=0.995
+ $X2=2.395 $Y2=0.56
r184 3 38 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.485 $X2=0.285 $Y2=1.66
r185 3 40 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.485 $X2=0.285 $Y2=2.34
r186 2 52 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.235 $X2=1.655 $Y2=0.49
r187 1 46 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.785 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_4%VPWR 1 2 3 12 16 18 20 22 24 29 34 40 43 47 51
r55 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 41 51 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r61 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 35 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.15 $Y=2.72
+ $X2=3.025 $Y2=2.72
r63 35 37 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.15 $Y=2.72 $X2=3.45
+ $Y2=2.72
r64 34 46 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.74 $Y=2.72 $X2=3.94
+ $Y2=2.72
r65 34 37 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 30 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.13 $Y2=2.72
r70 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 29 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.9 $Y=2.72
+ $X2=3.025 $Y2=2.72
r72 29 32 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.9 $Y=2.72 $X2=2.53
+ $Y2=2.72
r73 26 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 24 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.13 $Y2=2.72
r75 24 26 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 22 51 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 18 46 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.865 $Y=2.635
+ $X2=3.94 $Y2=2.72
r78 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.865 $Y=2.635
+ $X2=3.865 $Y2=1.96
r79 14 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=2.635
+ $X2=3.025 $Y2=2.72
r80 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.025 $Y=2.635
+ $X2=3.025 $Y2=1.96
r81 10 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=2.635
+ $X2=2.13 $Y2=2.72
r82 10 12 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.13 $Y=2.635
+ $X2=2.13 $Y2=1.96
r83 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.73
+ $Y=1.485 $X2=3.865 $Y2=1.96
r84 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.89
+ $Y=1.485 $X2=3.025 $Y2=1.96
r85 1 12 300 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=1.485 $X2=2.13 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_4%X 1 2 3 4 13 15 19 21 23 24 27 31 33 35 39 41
+ 43 46
r74 43 46 2.98271 $w=2.45e-07 $l=9e-08 $layer=LI1_cond $X=3.932 $Y=0.815
+ $X2=3.932 $Y2=0.905
r75 43 46 0.705577 $w=2.43e-07 $l=1.5e-08 $layer=LI1_cond $X=3.932 $Y=0.92
+ $X2=3.932 $Y2=0.905
r76 42 43 25.1656 $w=2.43e-07 $l=5.35e-07 $layer=LI1_cond $X=3.932 $Y=1.455
+ $X2=3.932 $Y2=0.92
r77 36 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.61 $Y=0.815
+ $X2=3.445 $Y2=0.815
r78 35 43 4.04323 $w=1.8e-07 $l=1.22e-07 $layer=LI1_cond $X=3.81 $Y=0.815
+ $X2=3.932 $Y2=0.815
r79 35 36 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=3.81 $Y=0.815 $X2=3.61
+ $Y2=0.815
r80 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.57 $Y=1.54
+ $X2=3.445 $Y2=1.54
r81 33 42 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.81 $Y=1.54
+ $X2=3.932 $Y2=1.455
r82 33 34 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.81 $Y=1.54
+ $X2=3.57 $Y2=1.54
r83 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=1.625
+ $X2=3.445 $Y2=1.54
r84 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.445 $Y=1.625
+ $X2=3.445 $Y2=2.3
r85 25 39 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.445 $Y=0.725
+ $X2=3.445 $Y2=0.815
r86 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.445 $Y=0.725
+ $X2=3.445 $Y2=0.39
r87 23 39 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=0.815
+ $X2=3.445 $Y2=0.815
r88 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.28 $Y=0.815
+ $X2=2.77 $Y2=0.815
r89 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.73 $Y=1.54
+ $X2=2.605 $Y2=1.54
r90 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.32 $Y=1.54
+ $X2=3.445 $Y2=1.54
r91 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.32 $Y=1.54 $X2=2.73
+ $Y2=1.54
r92 17 24 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.645 $Y=0.725
+ $X2=2.77 $Y2=0.815
r93 17 19 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=2.645 $Y=0.725
+ $X2=2.645 $Y2=0.485
r94 13 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=1.625
+ $X2=2.605 $Y2=1.54
r95 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.605 $Y=1.625
+ $X2=2.605 $Y2=2.3
r96 4 41 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.485 $X2=3.445 $Y2=1.62
r97 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.485 $X2=3.445 $Y2=2.3
r98 3 38 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.485 $X2=2.605 $Y2=1.62
r99 3 15 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.485 $X2=2.605 $Y2=2.3
r100 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.31
+ $Y=0.235 $X2=3.445 $Y2=0.39
r101 1 19 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.605 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__OR4_4%VGND 1 2 3 4 5 16 18 20 24 28 30 34 36 38 40
+ 42 47 56 59 62 66 70
c84 30 0 1.60701e-19 $X=2.94 $Y=0
r85 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r86 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r87 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r88 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r89 57 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.23
+ $Y2=0
r90 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r91 53 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r92 51 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r93 51 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r94 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r95 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=0 $X2=3.025
+ $Y2=0
r96 48 50 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.11 $Y=0 $X2=3.45
+ $Y2=0
r97 47 65 3.40825 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=3.96
+ $Y2=0
r98 47 50 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=3.45
+ $Y2=0
r99 46 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r100 46 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r101 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r102 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.235
+ $Y2=0
r103 43 45 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.61
+ $Y2=0
r104 42 59 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=2.15
+ $Y2=0
r105 42 45 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.96 $Y=0 $X2=1.61
+ $Y2=0
r106 40 70 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0
+ $X2=0.23 $Y2=0
r107 36 65 3.40825 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.96 $Y2=0
r108 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.865 $Y=0.085
+ $X2=3.865 $Y2=0.39
r109 32 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=0.085
+ $X2=3.025 $Y2=0
r110 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.025 $Y=0.085
+ $X2=3.025 $Y2=0.39
r111 31 59 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.15
+ $Y2=0
r112 30 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0 $X2=3.025
+ $Y2=0
r113 30 31 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=2.34
+ $Y2=0
r114 26 59 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r115 26 28 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.4
r116 22 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r117 22 24 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.4
r118 21 53 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=0 $X2=0.185
+ $Y2=0
r119 20 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.235
+ $Y2=0
r120 20 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.37
+ $Y2=0
r121 16 53 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.185 $Y2=0
r122 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.42
r123 5 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.865 $Y2=0.39
r124 4 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.235 $X2=3.025 $Y2=0.39
r125 3 28 182 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.235 $X2=2.175 $Y2=0.4
r126 2 24 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.235 $Y2=0.4
r127 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.42
.ends


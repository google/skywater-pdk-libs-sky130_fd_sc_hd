* File: sky130_fd_sc_hd__a32o_4.spice.pex
* Created: Thu Aug 27 14:05:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A32O_4%A_79_21# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 41 50 51 52 53 58 60 62 67 71 73 74 75 82
c166 82 0 1.75139e-19 $X=1.73 $Y=1.16
c167 71 0 1.30021e-19 $X=6.255 $Y=0.72
c168 50 0 1.00633e-19 $X=1.885 $Y=1.495
r169 79 80 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r170 74 75 4.00505 $w=1.78e-07 $l=6.5e-08 $layer=LI1_cond $X=6.135 $Y=1.995
+ $X2=6.2 $Y2=1.995
r171 69 71 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=5.365 $Y=0.72
+ $X2=6.255 $Y2=0.72
r172 65 67 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.3 $Y=2 $X2=7.14
+ $Y2=2
r173 65 75 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.3 $Y=2 $X2=6.2
+ $Y2=2
r174 62 74 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.45 $Y=1.99
+ $X2=6.135 $Y2=1.99
r175 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.365 $Y=1.905
+ $X2=5.45 $Y2=1.99
r176 59 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=1.665
+ $X2=5.365 $Y2=1.58
r177 59 60 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.365 $Y=1.665
+ $X2=5.365 $Y2=1.905
r178 58 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=1.495
+ $X2=5.365 $Y2=1.58
r179 57 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=0.805
+ $X2=5.365 $Y2=0.72
r180 57 58 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.365 $Y=0.805
+ $X2=5.365 $Y2=1.495
r181 53 69 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.28 $Y=0.72
+ $X2=5.365 $Y2=0.72
r182 53 55 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.28 $Y=0.72
+ $X2=4.56 $Y2=0.72
r183 51 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.28 $Y=1.58
+ $X2=5.365 $Y2=1.58
r184 51 52 215.947 $w=1.68e-07 $l=3.31e-06 $layer=LI1_cond $X=5.28 $Y=1.58
+ $X2=1.97 $Y2=1.58
r185 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.885 $Y=1.495
+ $X2=1.97 $Y2=1.58
r186 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.885 $Y=1.325
+ $X2=1.885 $Y2=1.495
r187 48 82 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.73 $Y2=1.16
r188 48 80 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.395 $Y=1.16
+ $X2=1.31 $Y2=1.16
r189 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.395
+ $Y=1.16 $X2=1.395 $Y2=1.16
r190 44 79 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.89 $Y2=1.16
r191 44 76 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.47 $Y2=1.16
r192 43 47 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=0.655 $Y=1.16
+ $X2=1.395 $Y2=1.16
r193 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.655
+ $Y=1.16 $X2=0.655 $Y2=1.16
r194 41 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.8 $Y=1.16
+ $X2=1.885 $Y2=1.325
r195 41 47 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.8 $Y=1.16
+ $X2=1.395 $Y2=1.16
r196 37 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r197 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r198 34 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r199 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r200 30 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r201 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r202 27 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r203 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r204 23 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r205 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r206 20 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r207 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r208 16 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r209 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r210 13 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r211 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r212 4 67 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=7.005
+ $Y=1.485 $X2=7.14 $Y2=2
r213 3 65 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=6.165
+ $Y=1.485 $X2=6.3 $Y2=2
r214 2 71 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.235 $X2=6.255 $Y2=0.72
r215 1 55 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%A3 1 3 6 8 10 13 15 16 20
c44 16 0 1.75139e-19 $X=2.995 $Y=1.19
r45 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.715
+ $Y=1.16 $X2=2.715 $Y2=1.16
r46 20 22 21.7726 $w=3.21e-07 $l=1.45e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.715 $Y2=1.16
r47 19 20 63.0654 $w=3.21e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r48 16 23 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=2.995 $Y=1.185
+ $X2=2.715 $Y2=1.185
r49 15 23 9.42908 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=2.535 $Y=1.185
+ $X2=2.715 $Y2=1.185
r50 11 20 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r52 8 20 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r54 4 19 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
r56 1 19 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995 $X2=2.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%A2 1 3 6 8 10 13 15 16 26
r45 24 26 12.8343 $w=3.38e-07 $l=9e-08 $layer=POLY_cond $X=3.84 $Y=1.17 $X2=3.93
+ $Y2=1.17
r46 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.16 $X2=3.84 $Y2=1.16
r47 22 24 47.0592 $w=3.38e-07 $l=3.3e-07 $layer=POLY_cond $X=3.51 $Y=1.17
+ $X2=3.84 $Y2=1.17
r48 20 22 1.42604 $w=3.38e-07 $l=1e-08 $layer=POLY_cond $X=3.5 $Y=1.17 $X2=3.51
+ $Y2=1.17
r49 16 25 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=3.935 $Y=1.2
+ $X2=3.84 $Y2=1.2
r50 15 25 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=3.475 $Y=1.2
+ $X2=3.84 $Y2=1.2
r51 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.5
+ $Y=1.16 $X2=3.5 $Y2=1.16
r52 11 26 21.7938 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.93 $Y=1.345
+ $X2=3.93 $Y2=1.17
r53 11 13 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.93 $Y=1.345
+ $X2=3.93 $Y2=1.985
r54 8 26 21.7938 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.17
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=0.56
r56 4 22 21.7938 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.51 $Y=1.345
+ $X2=3.51 $Y2=1.17
r57 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.51 $Y=1.345 $X2=3.51
+ $Y2=1.985
r58 1 22 21.7938 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.17
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995 $X2=3.51
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%A1 3 7 11 15 17 18 25
r44 25 27 21.5591 $w=3.13e-07 $l=1.4e-07 $layer=POLY_cond $X=4.77 $Y=1.18
+ $X2=4.91 $Y2=1.18
r45 23 25 30.7987 $w=3.13e-07 $l=2e-07 $layer=POLY_cond $X=4.57 $Y=1.18 $X2=4.77
+ $Y2=1.18
r46 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.57
+ $Y=1.16 $X2=4.57 $Y2=1.16
r47 18 24 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.855 $Y=1.2
+ $X2=4.57 $Y2=1.2
r48 18 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.91
+ $Y=1.16 $X2=4.91 $Y2=1.16
r49 17 24 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=4.395 $Y=1.2
+ $X2=4.57 $Y2=1.2
r50 13 25 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.345
+ $X2=4.77 $Y2=1.18
r51 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.77 $Y=1.345
+ $X2=4.77 $Y2=1.985
r52 9 25 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.015
+ $X2=4.77 $Y2=1.18
r53 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.77 $Y=1.015
+ $X2=4.77 $Y2=0.56
r54 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.35 $Y=1.345 $X2=4.35
+ $Y2=1.985
r55 1 23 33.8786 $w=3.13e-07 $l=2.2e-07 $layer=POLY_cond $X=4.35 $Y=1.18
+ $X2=4.57 $Y2=1.18
r56 1 5 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.18 $X2=4.35
+ $Y2=1.345
r57 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%B1 3 7 11 15 17 19 21 37
c51 37 0 1.83668e-19 $X=6.465 $Y=1.175
r52 37 38 7.35254 $w=2.95e-07 $l=4.5e-08 $layer=POLY_cond $X=6.465 $Y=1.175
+ $X2=6.51 $Y2=1.175
r53 35 37 7.35254 $w=2.95e-07 $l=4.5e-08 $layer=POLY_cond $X=6.42 $Y=1.175
+ $X2=6.465 $Y2=1.175
r54 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.42
+ $Y=1.16 $X2=6.42 $Y2=1.16
r55 33 35 53.9186 $w=2.95e-07 $l=3.3e-07 $layer=POLY_cond $X=6.09 $Y=1.175
+ $X2=6.42 $Y2=1.175
r56 31 33 1.6339 $w=2.95e-07 $l=1e-08 $layer=POLY_cond $X=6.08 $Y=1.175 $X2=6.09
+ $Y2=1.175
r57 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.08
+ $Y=1.16 $X2=6.08 $Y2=1.16
r58 29 31 5.71864 $w=2.95e-07 $l=3.5e-08 $layer=POLY_cond $X=6.045 $Y=1.175
+ $X2=6.08 $Y2=1.175
r59 21 36 5.32799 $w=5.48e-07 $l=2.45e-07 $layer=LI1_cond $X=6.665 $Y=1.35
+ $X2=6.42 $Y2=1.35
r60 19 36 4.67558 $w=5.48e-07 $l=2.15e-07 $layer=LI1_cond $X=6.205 $Y=1.35
+ $X2=6.42 $Y2=1.35
r61 19 32 2.71836 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.205 $Y=1.35
+ $X2=6.08 $Y2=1.35
r62 17 32 7.2852 $w=5.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.745 $Y=1.35
+ $X2=6.08 $Y2=1.35
r63 13 38 18.5736 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.51 $Y=1.325
+ $X2=6.51 $Y2=1.175
r64 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.51 $Y=1.325
+ $X2=6.51 $Y2=1.985
r65 9 37 18.5736 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.465 $Y=1.025
+ $X2=6.465 $Y2=1.175
r66 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.465 $Y=1.025
+ $X2=6.465 $Y2=0.56
r67 5 33 18.5736 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.09 $Y=1.325
+ $X2=6.09 $Y2=1.175
r68 5 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.09 $Y=1.325 $X2=6.09
+ $Y2=1.985
r69 1 29 18.5736 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.045 $Y=1.025
+ $X2=6.045 $Y2=1.175
r70 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.045 $Y=1.025
+ $X2=6.045 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%B2 3 7 11 15 17 18 19 24 28
c39 28 0 1.61536e-19 $X=7.127 $Y=1.295
c40 18 0 2.21319e-20 $X=7.125 $Y=1.53
c41 3 0 1.30021e-19 $X=6.93 $Y=0.56
r42 24 26 31.5403 $w=2.98e-07 $l=1.95e-07 $layer=POLY_cond $X=7.35 $Y=1.17
+ $X2=7.545 $Y2=1.17
r43 19 32 16.7628 $w=2.18e-07 $l=3.2e-07 $layer=LI1_cond $X=7.545 $Y=1.185
+ $X2=7.225 $Y2=1.185
r44 19 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.545
+ $Y=1.16 $X2=7.545 $Y2=1.16
r45 18 28 13.366 $w=1.93e-07 $l=2.35e-07 $layer=LI1_cond $X=7.127 $Y=1.53
+ $X2=7.127 $Y2=1.295
r46 17 28 3.62192 $w=1.95e-07 $l=1.1e-07 $layer=LI1_cond $X=7.127 $Y=1.185
+ $X2=7.127 $Y2=1.295
r47 17 32 3.2268 $w=2.2e-07 $l=9.8e-08 $layer=LI1_cond $X=7.127 $Y=1.185
+ $X2=7.225 $Y2=1.185
r48 13 24 18.8112 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=7.35 $Y=1.325
+ $X2=7.35 $Y2=1.17
r49 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.35 $Y=1.325
+ $X2=7.35 $Y2=1.985
r50 9 24 18.8112 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=7.35 $Y=1.015
+ $X2=7.35 $Y2=1.17
r51 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.35 $Y=1.015
+ $X2=7.35 $Y2=0.56
r52 5 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.93 $Y=1.325 $X2=6.93
+ $Y2=1.985
r53 1 24 67.9329 $w=2.98e-07 $l=4.2e-07 $layer=POLY_cond $X=6.93 $Y=1.17
+ $X2=7.35 $Y2=1.17
r54 1 5 18.8112 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=6.93 $Y=1.17 $X2=6.93
+ $Y2=1.325
r55 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.93 $Y=1.025
+ $X2=6.93 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%VPWR 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 55 57 79 80 86
c122 3 0 1.00633e-19 $X=1.805 $Y=1.485
c123 1 0 3.98522e-20 $X=0.135 $Y=1.485
r124 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r125 79 80 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r126 77 80 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=7.59 $Y2=2.72
r127 76 79 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=7.59 $Y2=2.72
r128 76 77 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r129 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r130 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r131 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r134 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r135 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r136 65 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r137 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r138 62 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.1 $Y2=2.72
r139 62 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 61 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r141 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r142 58 83 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r143 58 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r144 57 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.1 $Y2=2.72
r145 57 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 55 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r147 55 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r148 53 73 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.395 $Y=2.72
+ $X2=4.37 $Y2=2.72
r149 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=2.72
+ $X2=4.56 $Y2=2.72
r150 52 76 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.725 $Y=2.72
+ $X2=4.83 $Y2=2.72
r151 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=2.72
+ $X2=4.56 $Y2=2.72
r152 50 70 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=2.72
+ $X2=3.45 $Y2=2.72
r153 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=2.72
+ $X2=3.72 $Y2=2.72
r154 49 73 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.37 $Y2=2.72
r155 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=3.72 $Y2=2.72
r156 47 67 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.53 $Y2=2.72
r157 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.78 $Y2=2.72
r158 46 70 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.45 $Y2=2.72
r159 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.78 $Y2=2.72
r160 44 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.61 $Y2=2.72
r161 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.94 $Y2=2.72
r162 43 67 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.53 $Y2=2.72
r163 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=1.94 $Y2=2.72
r164 39 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2.72
r165 39 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2.34
r166 35 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2.72
r167 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2.34
r168 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r169 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.34
r170 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r171 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r172 23 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r173 23 25 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r174 19 83 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r175 19 21 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2
r176 6 41 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2.34
r177 5 37 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2.34
r178 4 33 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2.34
r179 3 29 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r180 2 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r181 1 21 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%X 1 2 3 4 13 15 19 23 25 27 31 35 37 38 39 40
+ 41 47 48 50
c49 50 0 3.98522e-20 $X=0.235 $Y=0.85
r50 47 50 2.35727 $w=2.18e-07 $l=4.5e-08 $layer=LI1_cond $X=0.23 $Y=0.805
+ $X2=0.23 $Y2=0.85
r51 41 48 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=1.58 $X2=0.23
+ $Y2=1.495
r52 41 48 1.30959 $w=2.18e-07 $l=2.5e-08 $layer=LI1_cond $X=0.23 $Y=1.47
+ $X2=0.23 $Y2=1.495
r53 40 41 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.23 $Y2=1.47
r54 39 47 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=0.72 $X2=0.23
+ $Y2=0.805
r55 39 40 16.7628 $w=2.18e-07 $l=3.2e-07 $layer=LI1_cond $X=0.23 $Y=0.87
+ $X2=0.23 $Y2=1.19
r56 39 50 1.04768 $w=2.18e-07 $l=2e-08 $layer=LI1_cond $X=0.23 $Y=0.87 $X2=0.23
+ $Y2=0.85
r57 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.96
r58 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.52 $Y=0.635
+ $X2=1.52 $Y2=0.42
r59 28 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.58
+ $X2=0.68 $Y2=1.58
r60 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=1.58
+ $X2=1.52 $Y2=1.665
r61 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=1.58
+ $X2=0.765 $Y2=1.58
r62 26 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.72
+ $X2=0.68 $Y2=0.72
r63 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=1.52 $Y2=0.635
r64 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=0.765 $Y2=0.72
r65 21 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.58
r66 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.96
r67 17 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.68 $Y2=0.72
r68 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.68 $Y2=0.42
r69 16 41 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.34 $Y=1.58 $X2=0.23
+ $Y2=1.58
r70 15 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=1.58
+ $X2=0.68 $Y2=1.58
r71 15 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.595 $Y=1.58
+ $X2=0.34 $Y2=1.58
r72 14 39 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.34 $Y=0.72 $X2=0.23
+ $Y2=0.72
r73 13 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0.72
+ $X2=0.68 $Y2=0.72
r74 13 14 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.595 $Y=0.72
+ $X2=0.34 $Y2=0.72
r75 4 35 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r76 3 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
r77 2 31 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.42
r78 1 19 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%A_445_297# 1 2 3 4 5 6 21 23 24 27 29 33 35
+ 39 40 45 47 49 50
r74 45 52 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=2.255 $X2=7.6
+ $Y2=2.34
r75 45 47 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.6 $Y=2.255
+ $X2=7.6 $Y2=1.92
r76 42 44 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.88 $Y=2.34
+ $X2=6.72 $Y2=2.34
r77 40 42 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=5.065 $Y=2.34
+ $X2=5.88 $Y2=2.34
r78 39 52 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.475 $Y=2.34
+ $X2=7.6 $Y2=2.34
r79 39 44 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.475 $Y=2.34
+ $X2=6.72 $Y2=2.34
r80 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.98 $Y=2.255
+ $X2=5.065 $Y2=2.34
r81 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.98 $Y=2.085
+ $X2=4.98 $Y2=2.255
r82 36 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=2 $X2=4.14
+ $Y2=2
r83 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.895 $Y=2
+ $X2=4.98 $Y2=2.085
r84 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.895 $Y=2 $X2=4.225
+ $Y2=2
r85 31 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.085
+ $X2=4.14 $Y2=2
r86 31 33 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.14 $Y=2.085
+ $X2=4.14 $Y2=2.3
r87 30 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=2 $X2=3.3
+ $Y2=2
r88 29 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=2 $X2=4.14
+ $Y2=2
r89 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.055 $Y=2 $X2=3.385
+ $Y2=2
r90 25 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.085 $X2=3.3
+ $Y2=2
r91 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.3 $Y=2.085
+ $X2=3.3 $Y2=2.3
r92 23 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2 $X2=3.3
+ $Y2=2
r93 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.215 $Y=2 $X2=2.445
+ $Y2=2
r94 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=2.085
+ $X2=2.445 $Y2=2
r95 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.36 $Y=2.085
+ $X2=2.36 $Y2=2.3
r96 6 52 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.425
+ $Y=1.485 $X2=7.56 $Y2=2.34
r97 6 47 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=7.425
+ $Y=1.485 $X2=7.56 $Y2=1.92
r98 5 44 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.585
+ $Y=1.485 $X2=6.72 $Y2=2.34
r99 4 42 600 $w=1.7e-07 $l=1.39862e-06 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.485 $X2=5.88 $Y2=2.34
r100 3 33 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2.3
r101 2 27 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=1.485 $X2=3.3 $Y2=2.3
r102 1 21 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 42 44 56 65 66 72 75
r112 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r113 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r114 66 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r115 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r116 63 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=7.14
+ $Y2=0
r117 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.305 $Y=0
+ $X2=7.59 $Y2=0
r118 62 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r119 61 62 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r120 59 62 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=6.67
+ $Y2=0
r121 58 61 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=6.67
+ $Y2=0
r122 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r123 56 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=0 $X2=7.14
+ $Y2=0
r124 56 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=6.67 $Y2=0
r125 55 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r126 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r127 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r128 52 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r129 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r130 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r131 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r132 48 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r133 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r134 45 69 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r135 45 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r136 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r137 44 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r138 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r139 42 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r140 40 54 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.53
+ $Y2=0
r141 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.78
+ $Y2=0
r142 39 58 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.99
+ $Y2=0
r143 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.78
+ $Y2=0
r144 37 51 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.61 $Y2=0
r145 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.94
+ $Y2=0
r146 36 54 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.105 $Y=0
+ $X2=2.53 $Y2=0
r147 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=1.94
+ $Y2=0
r148 32 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0
r149 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0.38
r150 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r151 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.38
r152 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r153 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.38
r154 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r155 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r156 16 69 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r157 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r158 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.005
+ $Y=0.235 $X2=7.14 $Y2=0.38
r159 4 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.38
r160 3 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r161 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r162 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%A_445_47# 1 2 9 11 13
r25 11 13 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=2.445 $Y=0.74
+ $X2=3.72 $Y2=0.74
r26 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=0.655
+ $X2=2.445 $Y2=0.74
r27 7 9 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.36 $Y=0.655
+ $X2=2.36 $Y2=0.42
r28 2 13 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.74
r29 1 9 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%A_635_47# 1 2 3 16
r20 14 16 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.38
+ $X2=4.98 $Y2=0.38
r21 11 14 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.3 $Y=0.38 $X2=4.14
+ $Y2=0.38
r22 3 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.38
r23 2 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.38
r24 1 11 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.3 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A32O_4%A_1142_47# 1 2 3 10 14 15 16 17 20
r32 18 20 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.56 $Y=0.645
+ $X2=7.56 $Y2=0.42
r33 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.475 $Y=0.73
+ $X2=7.56 $Y2=0.645
r34 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.475 $Y=0.73
+ $X2=6.805 $Y2=0.73
r35 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.72 $Y=0.645
+ $X2=6.805 $Y2=0.73
r36 14 23 3.40825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.72 $Y=0.465
+ $X2=6.72 $Y2=0.36
r37 14 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.72 $Y=0.465
+ $X2=6.72 $Y2=0.645
r38 10 23 3.40825 $w=1.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=6.635 $Y=0.38
+ $X2=6.72 $Y2=0.36
r39 10 12 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.635 $Y=0.38
+ $X2=5.835 $Y2=0.38
r40 3 20 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.56 $Y2=0.42
r41 2 23 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=6.54
+ $Y=0.235 $X2=6.72 $Y2=0.42
r42 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.71
+ $Y=0.235 $X2=5.835 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a32oi_2.spice
* Created: Tue Sep  1 18:55:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a32oi_2.pex.spice"
.subckt sky130_fd_sc_hd__a32oi_2  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1006 N_A_27_47#_M1006_d N_B2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1016 N_A_27_47#_M1016_d N_B2_M1016_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1008 N_A_27_47#_M1016_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_27_47#_M1009_d N_B1_M1009_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1012_d N_A1_M1012_g N_A_478_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1012_d N_A1_M1019_g N_A_478_47#_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.091 PD=0.92 PS=0.93 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1001 N_A_478_47#_M1019_s N_A2_M1001_g N_A_730_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.08775 PD=0.93 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1005 N_A_478_47#_M1005_d N_A2_M1005_g N_A_730_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_730_47#_M1004_d N_A3_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.20475 PD=1.02 PS=1.93 NRD=3.684 NRS=9.228 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_A_730_47#_M1004_d N_A3_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=12.912 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_297#_M1002_d N_B2_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1010 N_A_27_297#_M1010_d N_B2_M1010_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_A_27_297#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1000_d N_B1_M1015_g N_A_27_297#_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1011 N_A_27_297#_M1015_s N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.3775 PD=1.27 PS=1.755 NRD=0 NRS=13.7703 M=1 R=6.66667 SA=75001.9
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1013 N_A_27_297#_M1013_d N_A1_M1013_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.3775 PD=1.3 PS=1.755 NRD=0 NRS=12.7853 M=1 R=6.66667 SA=75002.8
+ SB=75002.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_27_297#_M1013_d N_A2_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.305 PD=1.3 PS=1.61 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1017 N_A_27_297#_M1017_d N_A2_M1017_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.305 PD=1.275 PS=1.61 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1007 N_A_27_297#_M1017_d N_A3_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1375 AS=0.335 PD=1.275 PS=1.67 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75004.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1018 N_A_27_297#_M1018_d N_A3_M1018_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.335 PD=2.52 PS=1.67 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75005.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__a32oi_2.pxi.spice"
*
.ends
*
*

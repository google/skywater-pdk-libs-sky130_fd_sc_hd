* File: sky130_fd_sc_hd__a221o_1.pex.spice
* Created: Thu Aug 27 14:01:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A221O_1%C1 1 3 6 8 14
r28 11 14 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r30 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r31 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r32 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r33 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%B2 3 7 8 11 12 13
c32 3 0 1.14647e-19 $X=0.89 $Y=1.985
r33 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.995
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r35 8 12 10.8136 $w=1.98e-07 $l=1.95e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.89 $Y2=1.175
r36 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.95 $Y=0.56 $X2=0.95
+ $Y2=0.995
r37 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r38 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%B1 3 6 8 9 13 15
r44 14 17 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.39 $Y=1.175
+ $X2=1.56 $Y2=1.175
r45 13 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.16
+ $X2=1.38 $Y2=1.325
r46 13 15 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.16
+ $X2=1.38 $Y2=0.995
r47 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.39
+ $Y=1.16 $X2=1.39 $Y2=1.16
r48 9 17 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=1.615 $Y=1.175 $X2=1.56
+ $Y2=1.175
r49 8 17 9.2607 $w=2.78e-07 $l=2.25e-07 $layer=LI1_cond $X=1.56 $Y=0.85 $X2=1.56
+ $Y2=1.075
r50 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.985
+ $X2=1.31 $Y2=1.325
r51 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.56 $X2=1.31
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%A1 3 6 8 9 13 15
r41 13 16 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.162 $Y=1.16
+ $X2=2.162 $Y2=1.325
r42 13 15 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=2.162 $Y=1.16
+ $X2=2.162 $Y2=0.995
r43 9 22 3.21434 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=1.16
+ $X2=2.135 $Y2=1.075
r44 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.16 $X2=2.135 $Y2=1.16
r45 8 22 9.09823 $w=2.83e-07 $l=2.25e-07 $layer=LI1_cond $X=2.112 $Y=0.85
+ $X2=2.112 $Y2=1.075
r46 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.25 $Y=1.985
+ $X2=2.25 $Y2=1.325
r47 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.25 $Y=0.56 $X2=2.25
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%A2 3 6 8 11 12 13
r36 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.67 $Y2=1.325
r37 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.67 $Y2=0.995
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.16 $X2=2.67 $Y2=1.16
r39 8 12 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=2.67 $Y2=1.175
r40 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.73 $Y=1.985
+ $X2=2.73 $Y2=1.325
r41 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.73 $Y=0.56 $X2=2.73
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%A_27_47# 1 2 3 4 15 18 22 26 28 29 30 31 33
+ 34 35 41 42 43 47 48 50
c120 48 0 2.21533e-19 $X=3.15 $Y=1.16
r121 48 51 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.16
+ $X2=3.15 $Y2=1.325
r122 48 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.16
+ $X2=3.15 $Y2=0.995
r123 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.16 $X2=3.15 $Y2=1.16
r124 45 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.15 $Y=1.455
+ $X2=3.15 $Y2=1.16
r125 44 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.15 $Y=0.905
+ $X2=3.15 $Y2=1.16
r126 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.065 $Y=0.82
+ $X2=3.15 $Y2=0.905
r127 42 43 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.065 $Y=0.82
+ $X2=2.605 $Y2=0.82
r128 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.52 $Y=0.735
+ $X2=2.605 $Y2=0.82
r129 40 41 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.52 $Y=0.505
+ $X2=2.52 $Y2=0.735
r130 37 39 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=1.52 $Y=0.38
+ $X2=2.04 $Y2=0.38
r131 35 37 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.24 $Y=0.38
+ $X2=1.52 $Y2=0.38
r132 34 40 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.435 $Y=0.38
+ $X2=2.52 $Y2=0.505
r133 34 39 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=2.435 $Y=0.38
+ $X2=2.04 $Y2=0.38
r134 32 35 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.155 $Y=0.505
+ $X2=1.24 $Y2=0.38
r135 32 33 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.155 $Y=0.505
+ $X2=1.155 $Y2=0.735
r136 30 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.065 $Y=1.54
+ $X2=3.15 $Y2=1.455
r137 30 31 177.455 $w=1.68e-07 $l=2.72e-06 $layer=LI1_cond $X=3.065 $Y=1.54
+ $X2=0.345 $Y2=1.54
r138 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=0.82
+ $X2=1.155 $Y2=0.735
r139 28 29 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.07 $Y=0.82
+ $X2=0.345 $Y2=0.82
r140 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.345 $Y2=1.54
r141 24 26 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.65
r142 20 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.345 $Y2=0.82
r143 20 22 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.56
r144 18 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.195 $Y=1.985
+ $X2=3.195 $Y2=1.325
r145 15 50 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.195 $Y=0.56
+ $X2=3.195 $Y2=0.995
r146 4 26 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
r147 3 39 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.235 $X2=2.04 $Y2=0.42
r148 2 37 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.42
r149 1 22 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%A_109_297# 1 2 9 12 14 15
c25 14 0 1.14647e-19 $X=1.52 $Y=2.34
r26 14 15 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=2.36
+ $X2=1.355 $Y2=2.36
r27 12 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.845 $Y=2.38
+ $X2=1.355 $Y2=2.38
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.68 $Y=2.295
+ $X2=0.845 $Y2=2.38
r29 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=2.295 $X2=0.68
+ $Y2=1.96
r30 2 14 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r31 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%A_193_297# 1 2 7 9 11 16
r23 14 16 5.94149 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.1 $Y=1.96
+ $X2=1.245 $Y2=1.96
r24 9 18 3.3405 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=2.525 $Y=2.035
+ $X2=2.525 $Y2=1.915
r25 9 11 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.525 $Y=2.035
+ $X2=2.525 $Y2=2.3
r26 7 18 3.47969 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=2.4 $Y=1.915
+ $X2=2.525 $Y2=1.915
r27 7 16 55.4613 $w=2.38e-07 $l=1.155e-06 $layer=LI1_cond $X=2.4 $Y=1.915
+ $X2=1.245 $Y2=1.915
r28 2 18 600 $w=1.7e-07 $l=5.39096e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.485 $Y2=1.95
r29 2 11 600 $w=1.7e-07 $l=8.91417e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.485 $Y2=2.3
r30 1 14 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%VPWR 1 2 9 13 15 17 19 29 36 37 40 43
c52 13 0 1.18411e-19 $X=2.985 $Y=1.96
r53 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 37 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 34 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=2.72
+ $X2=2.985 $Y2=2.72
r58 34 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.15 $Y=2.72 $X2=3.45
+ $Y2=2.72
r59 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r62 30 40 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=2.23 $Y=2.72
+ $X2=2.052 $Y2=2.72
r63 30 32 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r64 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=2.72
+ $X2=2.985 $Y2=2.72
r65 29 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.82 $Y=2.72
+ $X2=2.53 $Y2=2.72
r66 28 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 19 40 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=2.052 $Y2=2.72
r69 19 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=1.61 $Y2=2.72
r70 17 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r71 17 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 15 27 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 15 21 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 11 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=2.635
+ $X2=2.985 $Y2=2.72
r75 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.985 $Y=2.635
+ $X2=2.985 $Y2=1.96
r76 7 40 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.052 $Y=2.635
+ $X2=2.052 $Y2=2.72
r77 7 9 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=2.052 $Y=2.635
+ $X2=2.052 $Y2=2.3
r78 2 13 300 $w=1.7e-07 $l=5.57786e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=2.985 $Y2=1.96
r79 1 9 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.485 $X2=2.04 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%X 1 2 7 9 10 11 12 16
r18 12 16 11.2985 $w=2.53e-07 $l=2.5e-07 $layer=LI1_cond $X=3.447 $Y=2.21
+ $X2=3.447 $Y2=1.96
r19 11 21 4.55602 $w=2.41e-07 $l=9e-08 $layer=LI1_cond $X=3.447 $Y=0.51
+ $X2=3.447 $Y2=0.42
r20 9 16 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=3.447 $Y=1.922
+ $X2=3.447 $Y2=1.96
r21 9 10 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=3.447 $Y=1.922
+ $X2=3.447 $Y2=1.795
r22 7 11 8.92078 $w=2.41e-07 $l=1.75186e-07 $layer=LI1_cond $X=3.49 $Y=0.665
+ $X2=3.447 $Y2=0.51
r23 7 10 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=3.49 $Y=0.665
+ $X2=3.49 $Y2=1.795
r24 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.27
+ $Y=1.485 $X2=3.405 $Y2=1.96
r25 1 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.27
+ $Y=0.235 $X2=3.405 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A221O_1%VGND 1 2 9 11 14 16 21 31 32 40 43
c49 9 0 1.03121e-19 $X=2.94 $Y=0.4
r50 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r51 32 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r52 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r53 29 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.94
+ $Y2=0
r54 29 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.45
+ $Y2=0
r55 28 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r56 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r57 25 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r58 25 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r59 24 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r60 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r62 21 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.94
+ $Y2=0
r63 21 27 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.53
+ $Y2=0
r64 16 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r65 14 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r66 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r67 11 43 9.87585 $w=4.98e-07 $l=3.55e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.44
r68 11 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r69 11 16 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0 $X2=0.515
+ $Y2=0
r70 11 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0 $X2=0.845
+ $Y2=0
r71 7 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085 $X2=2.94
+ $Y2=0
r72 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.4
r73 2 9 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.235 $X2=2.94 $Y2=0.4
r74 1 43 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.44
.ends


* File: sky130_fd_sc_hd__decap_4.spice.SKY130_FD_SC_HD__DECAP_4.pxi
* Created: Thu Aug 27 14:13:38 2020
* 
x_PM_SKY130_FD_SC_HD__DECAP_4%VGND N_VGND_M1001_s VGND N_VGND_c_11_n
+ N_VGND_M1000_g N_VGND_c_12_n N_VGND_c_13_n PM_SKY130_FD_SC_HD__DECAP_4%VGND
x_PM_SKY130_FD_SC_HD__DECAP_4%VPWR N_VPWR_M1000_s VPWR N_VPWR_M1001_g
+ N_VPWR_c_21_n N_VPWR_c_22_n PM_SKY130_FD_SC_HD__DECAP_4%VPWR
cc_1 VNB N_VGND_c_11_n 0.0336337f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.29
cc_2 VNB N_VGND_c_12_n 0.115583f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=0.51
cc_3 VNB N_VGND_c_13_n 0.121884f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=0
cc_4 VNB N_VPWR_M1001_g 0.151224f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.29
cc_5 VNB N_VPWR_c_21_n 0.0137616f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=0.645
cc_6 VNB N_VPWR_c_22_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0
cc_7 VPB N_VGND_c_11_n 0.11759f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.29
cc_8 VPB N_VGND_c_12_n 0.00381416f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=0.51
cc_9 VPB N_VPWR_c_21_n 0.132884f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=0.645
cc_10 VPB N_VPWR_c_22_n 0.0419189f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=0
cc_11 N_VGND_c_11_n N_VPWR_M1001_g 0.0689775f $X=0.27 $Y=1.29 $X2=0 $Y2=0
cc_12 N_VGND_c_12_n N_VPWR_M1001_g 0.142049f $X=1.58 $Y=0.51 $X2=0 $Y2=0
cc_13 N_VGND_c_11_n N_VPWR_c_21_n 0.172773f $X=0.27 $Y=1.29 $X2=0 $Y2=0
cc_14 N_VGND_c_12_n N_VPWR_c_21_n 0.16291f $X=1.58 $Y=0.51 $X2=0 $Y2=0

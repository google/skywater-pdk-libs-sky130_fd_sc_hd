* File: sky130_fd_sc_hd__a31o_2.pex.spice
* Created: Tue Sep  1 18:55:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A31O_2%A_79_21# 1 2 7 9 12 14 16 19 22 23 24 26 29
+ 33 37 39 44
c88 33 0 1.5053e-19 $X=0.72 $Y=1.16
c89 26 0 1.88247e-19 $X=2.62 $Y=1.495
c90 22 0 1.62889e-19 $X=0.64 $Y=1.495
c91 1 0 1.71438e-19 $X=2.285 $Y=0.235
r92 38 39 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.62 $Y=1.58
+ $X2=2.96 $Y2=1.58
r93 34 44 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.72 $Y=1.16
+ $X2=0.89 $Y2=1.16
r94 34 41 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.72 $Y=1.16
+ $X2=0.47 $Y2=1.16
r95 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.16 $X2=0.72 $Y2=1.16
r96 27 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=1.665
+ $X2=2.96 $Y2=1.58
r97 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=1.665
+ $X2=2.96 $Y2=1.96
r98 26 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.495
+ $X2=2.62 $Y2=1.58
r99 25 37 2.48377 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=2.62 $Y=0.505
+ $X2=2.54 $Y2=0.38
r100 25 26 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.62 $Y=0.505
+ $X2=2.62 $Y2=1.495
r101 23 38 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=1.58
+ $X2=2.62 $Y2=1.58
r102 23 24 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.535 $Y=1.58
+ $X2=0.725 $Y2=1.58
r103 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.64 $Y=1.495
+ $X2=0.725 $Y2=1.58
r104 21 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=1.245
+ $X2=0.64 $Y2=1.16
r105 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.64 $Y=1.245
+ $X2=0.64 $Y2=1.495
r106 17 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r107 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r108 14 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r109 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r110 10 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r111 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r112 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r113 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r114 2 29 300 $w=1.7e-07 $l=5.64137e-07 $layer=licon1_PDIFF $count=2 $X=2.765
+ $Y=1.485 $X2=2.96 $Y2=1.96
r115 1 37 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=2.285
+ $Y=0.235 $X2=2.54 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%A3 1 3 6 8 9 13
c39 13 0 2.44922e-19 $X=1.31 $Y=1.16
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.16 $X2=1.31 $Y2=1.16
r41 9 14 1.31655 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=1.23 $Y=1.19 $X2=1.23
+ $Y2=1.16
r42 8 14 13.6043 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.23 $Y=0.85 $X2=1.23
+ $Y2=1.16
r43 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r44 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r45 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%A2 3 6 9 13 16 17 18 21
c52 13 0 1.58449e-19 $X=1.71 $Y=0.78
r53 17 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.16
+ $X2=1.79 $Y2=1.325
r54 17 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.16
+ $X2=1.79 $Y2=0.995
r55 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.16 $X2=1.79 $Y2=1.16
r56 11 18 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.615 $Y=0.695
+ $X2=1.615 $Y2=0.51
r57 10 13 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=0.78
+ $X2=1.71 $Y2=0.78
r58 10 11 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.78
+ $X2=1.615 $Y2=0.695
r59 9 16 0.961343 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=1.71 $Y=1.075
+ $X2=1.71 $Y2=1.167
r60 8 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.865
+ $X2=1.71 $Y2=0.78
r61 8 9 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.71 $Y=0.865 $X2=1.71
+ $Y2=1.075
r62 6 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=1.325
r63 3 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.56 $X2=1.73
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%A1 3 6 10 11 16 18 21
c52 21 0 1.58449e-19 $X=2.27 $Y=0.995
c53 18 0 1.51344e-19 $X=2.075 $Y=0.51
c54 10 0 1.71438e-19 $X=2.27 $Y=1.16
r55 14 18 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=2.07 $Y=0.7 $X2=2.07
+ $Y2=0.51
r56 14 16 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.07 $Y=0.785 $X2=2.27
+ $Y2=0.785
r57 11 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.16
+ $X2=2.27 $Y2=1.325
r58 11 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.16
+ $X2=2.27 $Y2=0.995
r59 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.27
+ $Y=1.16 $X2=2.27 $Y2=1.16
r60 8 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.27 $Y=0.87 $X2=2.27
+ $Y2=0.785
r61 8 10 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.27 $Y=0.87 $X2=2.27
+ $Y2=1.16
r62 6 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.21 $Y=1.985
+ $X2=2.21 $Y2=1.325
r63 3 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.21 $Y=0.56 $X2=2.21
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%B1 3 5 7 8 9 16
c32 5 0 1.51344e-19 $X=2.75 $Y=0.995
r33 14 16 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.98 $Y2=1.16
r34 12 14 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.69 $Y=1.16 $X2=2.75
+ $Y2=1.16
r35 8 9 17.6317 $w=1.93e-07 $l=3.1e-07 $layer=LI1_cond $X=2.992 $Y=1.16
+ $X2=2.992 $Y2=0.85
r36 8 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=1.16 $X2=2.98 $Y2=1.16
r37 5 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=0.995
+ $X2=2.75 $Y2=1.16
r38 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.995 $X2=2.75
+ $Y2=0.56
r39 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.16
r40 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.69 $Y=1.325 $X2=2.69
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%VPWR 1 2 3 10 12 16 20 23 24 25 31 37 38 44
r59 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 38 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 35 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=1.98 $Y2=2.72
r63 35 37 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 34 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.98 $Y2=2.72
r67 31 33 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 30 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r69 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 27 41 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r71 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 25 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 25 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 23 29 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.06 $Y2=2.72
r76 22 33 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.06 $Y2=2.72
r78 18 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.72
r79 18 20 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.26
r80 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=2.635
+ $X2=1.06 $Y2=2.72
r81 14 16 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.06 $Y=2.635
+ $X2=1.06 $Y2=2
r82 10 41 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.192 $Y2=2.72
r83 10 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r84 3 20 600 $w=1.7e-07 $l=8.5805e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.98 $Y2=2.26
r85 2 16 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r86 1 12 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%X 1 2 7 9 13 17 19 20 21 22 29 30
c35 2 0 9.99956e-20 $X=0.545 $Y=1.485
r36 22 30 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=1.92
+ $X2=0.217 $Y2=1.835
r37 22 30 1.12985 $w=2.53e-07 $l=2.5e-08 $layer=LI1_cond $X=0.217 $Y=1.81
+ $X2=0.217 $Y2=1.835
r38 21 22 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=0.217 $Y=1.53
+ $X2=0.217 $Y2=1.81
r39 20 21 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.217 $Y=1.19
+ $X2=0.217 $Y2=1.53
r40 19 29 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=0.8
+ $X2=0.217 $Y2=0.885
r41 19 20 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=0.217 $Y=0.91
+ $X2=0.217 $Y2=1.19
r42 19 29 1.12985 $w=2.53e-07 $l=2.5e-08 $layer=LI1_cond $X=0.217 $Y=0.91
+ $X2=0.217 $Y2=0.885
r43 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.005
+ $X2=0.68 $Y2=2.3
r44 11 13 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.715
+ $X2=0.68 $Y2=0.42
r45 10 22 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.92
+ $X2=0.217 $Y2=1.92
r46 9 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.595 $Y=1.92
+ $X2=0.68 $Y2=2.005
r47 9 10 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.595 $Y=1.92
+ $X2=0.345 $Y2=1.92
r48 8 19 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.8
+ $X2=0.217 $Y2=0.8
r49 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.595 $Y=0.8
+ $X2=0.68 $Y2=0.715
r50 7 8 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.595 $Y=0.8 $X2=0.345
+ $Y2=0.8
r51 2 17 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.3
r52 1 13 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%A_277_297# 1 2 7 9 11 13 15
c25 2 0 1.88247e-19 $X=2.285 $Y=1.485
r26 13 20 3.04246 $w=2.5e-07 $l=9.88686e-08 $layer=LI1_cond $X=2.46 $Y=2.005
+ $X2=2.49 $Y2=1.92
r27 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.46 $Y=2.005
+ $X2=2.46 $Y2=2.26
r28 12 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.605 $Y=1.92
+ $X2=1.48 $Y2=1.92
r29 11 20 4.1007 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.335 $Y=1.92
+ $X2=2.49 $Y2=1.92
r30 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.335 $Y=1.92
+ $X2=1.605 $Y2=1.92
r31 7 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=2.005 $X2=1.48
+ $Y2=1.92
r32 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.48 $Y=2.005
+ $X2=1.48 $Y2=2.26
r33 2 20 600 $w=1.7e-07 $l=5.23498e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.485 $X2=2.48 $Y2=1.92
r34 2 15 600 $w=1.7e-07 $l=8.67035e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.485 $X2=2.48 $Y2=2.26
r35 1 18 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.92
r36 1 9 600 $w=1.7e-07 $l=8.39792e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_HD__A31O_2%VGND 1 2 3 10 12 15 16 18 22 24 29 41 45
c56 15 0 3.14973e-20 $X=1.12 $Y=0.3
r57 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r58 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r59 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r60 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r61 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r62 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r63 32 35 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r64 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r65 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r66 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.61
+ $Y2=0
r67 29 44 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=3.047
+ $Y2=0
r68 29 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.53
+ $Y2=0
r69 28 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r70 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r71 25 38 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r72 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r73 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r74 24 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.69
+ $Y2=0
r75 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r76 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r77 16 44 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.005 $Y=0.085
+ $X2=3.047 $Y2=0
r78 16 18 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.005 $Y=0.085
+ $X2=3.005 $Y2=0.4
r79 15 21 3.30798 $w=3.3e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=0.3 $X2=1.12
+ $Y2=0.38
r80 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r81 14 15 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.3
r82 10 38 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r83 10 12 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.38
r84 3 18 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.4
r85 2 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r86 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__xnor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
M1000 VPWR a_47_47# Y VPB phighvt w=1e+06u l=150000u
+  ad=1.39e+12p pd=8.78e+06u as=3.3e+11p ps=2.66e+06u
M1001 a_285_47# A VGND VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=3.445e+11p ps=3.66e+06u
M1002 a_377_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1003 VPWR A a_47_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1004 Y B a_377_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_129_47# B a_47_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=1.69e+11p ps=1.82e+06u
M1006 a_285_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_129_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_47_47# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_47_47# a_285_47# VNB nshort w=650000u l=150000u
+  ad=1.95e+11p pd=1.9e+06u as=0p ps=0u
.ends


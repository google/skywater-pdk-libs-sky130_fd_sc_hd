* File: sky130_fd_sc_hd__and3_2.pex.spice
* Created: Tue Sep  1 18:57:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND3_2%A 3 7 9 16
r27 15 16 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.48 $Y=1.16
+ $X2=0.485 $Y2=1.16
r28 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.48 $Y2=1.16
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r30 9 13 9.27941 $w=3.83e-07 $l=3.1e-07 $layer=LI1_cond $X=0.277 $Y=0.85
+ $X2=0.277 $Y2=1.16
r31 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.16
r32 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.475
r33 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r34 1 3 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.48 $Y=1.325 $X2=0.48
+ $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_2%B 1 3 8 9 12
r42 12 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=2.3
+ $X2=0.97 $Y2=2.135
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=2.3 $X2=0.98 $Y2=2.3
r44 9 13 5.76222 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.15 $Y=2.295
+ $X2=0.98 $Y2=2.295
r45 8 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.9 $Y=1.765 $X2=0.9
+ $Y2=2.135
r46 5 8 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.9 $Y=1.48 $X2=0.9
+ $Y2=1.765
r47 1 5 54.102 $w=1.96e-07 $l=2.45967e-07 $layer=POLY_cond $X=0.845 $Y=1.26
+ $X2=0.9 $Y2=1.48
r48 1 3 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.845 $Y=1.26
+ $X2=0.845 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_2%C 3 7 9 10 14
r49 14 17 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.317 $Y=1.16
+ $X2=1.317 $Y2=1.325
r50 14 16 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.317 $Y=1.16
+ $X2=1.317 $Y2=0.995
r51 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.16 $X2=1.31 $Y2=1.16
r52 10 15 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=1.27 $Y=0.85
+ $X2=1.27 $Y2=1.16
r53 10 22 5.01423 $w=4.08e-07 $l=1e-07 $layer=LI1_cond $X=1.27 $Y=0.85 $X2=1.27
+ $Y2=0.75
r54 9 22 12.0255 $w=2.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.18 $Y=0.51 $X2=1.18
+ $Y2=0.75
r55 7 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.375 $Y=1.695
+ $X2=1.375 $Y2=1.325
r56 3 16 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.25 $Y=0.475
+ $X2=1.25 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_2%A_29_311# 1 2 3 10 12 15 17 19 22 26 28 32 33
+ 35 36 40 42 46 49 50 56
r115 55 56 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.275 $Y=1.16
+ $X2=2.29 $Y2=1.16
r116 54 55 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.87 $Y=1.16
+ $X2=2.275 $Y2=1.16
r117 53 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.87 $Y2=1.16
r118 47 53 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.805 $Y=1.16
+ $X2=1.855 $Y2=1.16
r119 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=1.16 $X2=1.805 $Y2=1.16
r120 44 46 13.2781 $w=2.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.775 $Y=1.425
+ $X2=1.775 $Y2=1.16
r121 43 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.33 $Y=1.51
+ $X2=1.205 $Y2=1.51
r122 42 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.66 $Y=1.51
+ $X2=1.775 $Y2=1.425
r123 42 43 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.66 $Y=1.51
+ $X2=1.33 $Y2=1.51
r124 38 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.595
+ $X2=1.205 $Y2=1.51
r125 38 40 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.205 $Y=1.595
+ $X2=1.205 $Y2=1.725
r126 37 49 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.895 $Y=1.51
+ $X2=0.767 $Y2=1.51
r127 36 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.08 $Y=1.51
+ $X2=1.205 $Y2=1.51
r128 36 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.08 $Y=1.51
+ $X2=0.895 $Y2=1.51
r129 35 49 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.767 $Y=1.425
+ $X2=0.767 $Y2=1.51
r130 34 35 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=0.767 $Y=0.57
+ $X2=0.767 $Y2=1.425
r131 32 49 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.64 $Y=1.51
+ $X2=0.767 $Y2=1.51
r132 32 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.64 $Y=1.51
+ $X2=0.355 $Y2=1.51
r133 28 34 6.81977 $w=2.65e-07 $l=1.85957e-07 $layer=LI1_cond $X=0.64 $Y=0.437
+ $X2=0.767 $Y2=0.57
r134 28 30 15.8733 $w=2.63e-07 $l=3.65e-07 $layer=LI1_cond $X=0.64 $Y=0.437
+ $X2=0.275 $Y2=0.437
r135 24 33 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.227 $Y=1.595
+ $X2=0.355 $Y2=1.51
r136 24 26 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.227 $Y=1.595
+ $X2=0.227 $Y2=1.76
r137 20 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.325
+ $X2=2.29 $Y2=1.16
r138 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.29 $Y=1.325
+ $X2=2.29 $Y2=1.985
r139 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=1.16
r140 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=0.56
r141 13 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.325
+ $X2=1.87 $Y2=1.16
r142 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.87 $Y=1.325
+ $X2=1.87 $Y2=1.985
r143 10 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=1.16
r144 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=0.56
r145 3 40 600 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.555 $X2=1.165 $Y2=1.725
r146 2 26 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.555 $X2=0.27 $Y2=1.76
r147 1 30 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.265 $X2=0.275 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_2%VPWR 1 2 3 11 12 16 18 20 25 27 29 35 40 44
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r51 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 35 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 30 40 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.77 $Y=2.72
+ $X2=1.662 $Y2=2.72
r58 30 32 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.77 $Y=2.72 $X2=2.07
+ $Y2=2.72
r59 29 43 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.587 $Y2=2.72
r60 29 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 27 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 27 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 22 25 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=0.62 $Y=1.86 $X2=0.69
+ $Y2=1.86
r64 18 43 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.545 $Y=2.635
+ $X2=2.587 $Y2=2.72
r65 18 20 29.9192 $w=2.58e-07 $l=6.75e-07 $layer=LI1_cond $X=2.545 $Y=2.635
+ $X2=2.545 $Y2=1.96
r66 14 40 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.662 $Y=2.635
+ $X2=1.662 $Y2=2.72
r67 14 16 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=1.662 $Y=2.635
+ $X2=1.662 $Y2=1.955
r68 13 35 8.84583 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=0.715 $Y=2.72
+ $X2=0.357 $Y2=2.72
r69 12 40 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.662 $Y2=2.72
r70 12 13 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=0.715 $Y2=2.72
r71 11 35 17.8437 $w=6.51e-07 $l=7.09415e-07 $layer=LI1_cond $X=0.62 $Y=2.13
+ $X2=0.357 $Y2=2.72
r72 10 22 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.62 $Y=1.955
+ $X2=0.62 $Y2=1.86
r73 10 11 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=0.62 $Y=1.955
+ $X2=0.62 $Y2=2.13
r74 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.485 $X2=2.5 $Y2=1.96
r75 2 16 300 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_PDIFF $count=2 $X=1.45
+ $Y=1.485 $X2=1.66 $Y2=1.955
r76 1 25 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=0.555
+ $Y=1.555 $X2=0.69 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_2%X 1 2 8 11 12 13 14 15 20 23 26
r34 32 34 0.345023 $w=5.18e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=1.185
+ $X2=2.16 $Y2=1.185
r35 20 23 3.904 $w=2.5e-07 $l=8e-08 $layer=LI1_cond $X=2.105 $Y=0.59 $X2=2.105
+ $Y2=0.51
r36 15 34 8.51056 $w=5.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.53 $Y=1.185
+ $X2=2.16 $Y2=1.185
r37 14 26 10.4768 $w=2.73e-07 $l=2.5e-07 $layer=LI1_cond $X=2.107 $Y=2.21
+ $X2=2.107 $Y2=1.96
r38 13 31 6.85717 $w=2.48e-07 $l=1.23e-07 $layer=LI1_cond $X=2.105 $Y=0.592
+ $X2=2.105 $Y2=0.715
r39 13 20 0.0921954 $w=2.48e-07 $l=2e-09 $layer=LI1_cond $X=2.105 $Y=0.592
+ $X2=2.105 $Y2=0.59
r40 13 23 0.1464 $w=2.5e-07 $l=3e-09 $layer=LI1_cond $X=2.105 $Y=0.507 $X2=2.105
+ $Y2=0.51
r41 11 26 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=2.107 $Y=1.932
+ $X2=2.107 $Y2=1.96
r42 11 12 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.107 $Y=1.932
+ $X2=2.107 $Y2=1.795
r43 9 34 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.16 $Y=1.445 $X2=2.16
+ $Y2=1.185
r44 9 12 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.16 $Y=1.445
+ $X2=2.16 $Y2=1.795
r45 8 32 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.145 $Y=0.925
+ $X2=2.145 $Y2=1.185
r46 8 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.145 $Y=0.925
+ $X2=2.145 $Y2=0.715
r47 2 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.485 $X2=2.08 $Y2=1.96
r48 1 23 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.235 $X2=2.065 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_2%VGND 1 2 9 11 13 15 17 25 31 35
r35 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r37 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r38 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r39 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r40 26 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.64
+ $Y2=0
r41 26 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=2.07
+ $Y2=0
r42 25 34 4.27912 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.58
+ $Y2=0
r43 25 28 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.07
+ $Y2=0
r44 24 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r45 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r46 19 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r47 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.64
+ $Y2=0
r48 17 23 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.15
+ $Y2=0
r49 15 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r50 15 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 11 34 3.04293 $w=2.75e-07 $l=1.04307e-07 $layer=LI1_cond $X=2.537 $Y=0.085
+ $X2=2.58 $Y2=0
r52 11 13 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=2.537 $Y=0.085
+ $X2=2.537 $Y2=0.515
r53 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.085 $X2=1.64
+ $Y2=0
r54 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.64 $Y=0.085 $X2=1.64
+ $Y2=0.495
r55 2 13 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.485 $Y2=0.515
r56 1 9 182 $w=1.7e-07 $l=4.14337e-07 $layer=licon1_NDIFF $count=1 $X=1.325
+ $Y=0.265 $X2=1.64 $Y2=0.495
.ends


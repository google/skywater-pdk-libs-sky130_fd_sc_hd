* File: sky130_fd_sc_hd__and3_2.spice
* Created: Thu Aug 27 14:07:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and3_2.pex.spice"
.subckt sky130_fd_sc_hd__and3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_112_53# N_A_M1001_g N_A_29_311#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1007 A_184_53# N_B_M1007_g A_112_53# VNB NSHORT L=0.15 W=0.42 AD=0.05355
+ AS=0.0441 PD=0.675 PS=0.63 NRD=20.712 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_C_M1008_g A_184_53# VNB NSHORT L=0.15 W=0.42 AD=0.10237
+ AS=0.05355 PD=0.867477 PS=0.675 NRD=49.992 NRS=20.712 M=1 R=2.8 SA=75000.9
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1008_d N_A_29_311#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.15843 AS=0.08775 PD=1.34252 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_29_311#_M1004_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.08775 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_29_311#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 N_A_29_311#_M1006_d N_B_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.074375 AS=0.0567 PD=0.815 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_C_M1005_g N_A_29_311#_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0891761 AS=0.074375 PD=0.795634 PS=0.815 NRD=73.7765 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_29_311#_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.212324 PD=1.27 PS=1.89437 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1002_d N_A_29_311#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__and3_2.pxi.spice"
*
.ends
*
*

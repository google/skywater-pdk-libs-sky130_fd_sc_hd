* File: sky130_fd_sc_hd__dlrbp_1.spice.pex
* Created: Thu Aug 27 14:16:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRBP_1%GATE 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39587e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r47 19 20 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.205 $Y=1.19
+ $X2=0.205 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r49 15 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%A_27_47# 1 2 9 13 17 19 20 23 27 30 34 35 36
+ 41 44 46 49 50 53 56 57 60 64
c146 57 0 1.8552e-19 $X=2.555 $Y=1.53
c147 13 0 2.69793e-20 $X=0.89 $Y=2.135
c148 9 0 2.69793e-20 $X=0.89 $Y=0.445
r149 57 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r150 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.53
+ $X2=2.555 $Y2=1.53
r151 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r152 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r153 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.53
+ $X2=2.555 $Y2=1.53
r154 49 50 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.41 $Y=1.53
+ $X2=0.84 $Y2=1.53
r155 48 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r156 47 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r157 45 64 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r158 44 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r159 44 46 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r160 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r161 38 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r162 37 41 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r163 36 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r164 36 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r165 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r166 34 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r167 28 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r168 28 30 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r169 26 60 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r170 26 27 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r171 25 60 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r172 21 23 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.215 $Y=1.245
+ $X2=3.215 $Y2=0.415
r173 20 25 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r174 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.14 $Y=1.32
+ $X2=3.215 $Y2=1.245
r175 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.14 $Y=1.32
+ $X2=2.805 $Y2=1.32
r176 17 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.73 $Y=2.275
+ $X2=2.73 $Y2=1.685
r177 11 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r178 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r179 7 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r180 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r181 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r182 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%A_299_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c84 32 0 1.12109e-19 $X=2.255 $Y=0.93
c85 18 0 7.13094e-20 $X=1.97 $Y=0.7
r86 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=1.095
r87 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=0.765
r88 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r89 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r90 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.155 $Y2=0.93
r91 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.055 $Y2=1.495
r92 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=2.055 $Y2=1.495
r93 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=1.785 $Y2=1.58
r94 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r95 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=2.155 $Y2=0.93
r96 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=1.705 $Y2=0.7
r97 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r98 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r99 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=2.165
+ $X2=2.25 $Y2=1.095
r100 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.765
r101 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r102 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%A_193_47# 1 2 7 9 12 16 18 24 25 27 28 31 34
+ 39 40
c117 39 0 2.54761e-19 $X=3.18 $Y=1.74
c118 24 0 2.84791e-19 $X=3.01 $Y=1.575
r119 39 42 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.18 $Y2=1.875
r120 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r121 34 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.01 $Y=1.87
+ $X2=3.01 $Y2=1.87
r122 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r123 28 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r124 27 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.865 $Y=1.87
+ $X2=3.01 $Y2=1.87
r125 27 28 1.93688 $w=1.4e-07 $l=1.565e-06 $layer=MET1_cond $X=2.865 $Y=1.87
+ $X2=1.3 $Y2=1.87
r126 25 31 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r127 25 26 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r128 24 40 8.96243 $w=3.11e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.01 $Y=1.575
+ $X2=3.095 $Y2=1.74
r129 23 24 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=1.575
r130 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=0.9 $X2=2.765 $Y2=0.9
r131 18 23 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.925 $Y=0.9
+ $X2=3.01 $Y2=1.035
r132 18 20 6.82929 $w=2.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.925 $Y=0.9
+ $X2=2.765 $Y2=0.9
r133 16 26 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r134 12 42 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.15 $Y=2.275
+ $X2=3.15 $Y2=1.875
r135 7 21 43.0683 $w=3.2e-07 $l=2.14068e-07 $layer=POLY_cond $X=2.725 $Y=0.705
+ $X2=2.765 $Y2=0.9
r136 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.725 $Y=0.705
+ $X2=2.725 $Y2=0.415
r137 2 31 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r138 1 16 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%A_711_307# 1 2 9 13 15 17 20 22 23 26 30 32
+ 33 36 38 41 42 45 47 52 55
c114 36 0 1.91094e-19 $X=3.925 $Y=1.7
c115 13 0 2.20671e-19 $X=3.69 $Y=0.445
r116 56 58 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.63 $Y=1.7 $X2=3.69
+ $Y2=1.7
r117 53 63 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.805 $Y=1.16
+ $X2=5.935 $Y2=1.16
r118 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.805
+ $Y=1.16 $X2=5.805 $Y2=1.16
r119 50 52 18.39 $w=2.33e-07 $l=3.75e-07 $layer=LI1_cond $X=5.772 $Y=1.535
+ $X2=5.772 $Y2=1.16
r120 49 52 16.4284 $w=2.33e-07 $l=3.35e-07 $layer=LI1_cond $X=5.772 $Y=0.825
+ $X2=5.772 $Y2=1.16
r121 48 55 3.351 $w=2.8e-07 $l=1.07121e-07 $layer=LI1_cond $X=4.95 $Y=1.65
+ $X2=4.865 $Y2=1.7
r122 47 50 6.81752 $w=2.3e-07 $l=1.64754e-07 $layer=LI1_cond $X=5.655 $Y=1.65
+ $X2=5.772 $Y2=1.535
r123 47 48 35.3249 $w=2.28e-07 $l=7.05e-07 $layer=LI1_cond $X=5.655 $Y=1.65
+ $X2=4.95 $Y2=1.65
r124 43 55 3.18746 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=1.865
+ $X2=4.865 $Y2=1.7
r125 43 45 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.865 $Y=1.865
+ $X2=4.865 $Y2=2.27
r126 41 49 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=5.655 $Y=0.74
+ $X2=5.772 $Y2=0.825
r127 41 42 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.655 $Y=0.74
+ $X2=4.54 $Y2=0.74
r128 38 42 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.39 $Y=0.655
+ $X2=4.54 $Y2=0.74
r129 38 40 3.86333 $w=3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.39 $Y=0.655 $X2=4.39
+ $Y2=0.56
r130 36 58 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.69 $Y2=1.7
r131 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r132 33 55 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=1.7 $X2=4.865
+ $Y2=1.7
r133 33 35 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=4.78 $Y=1.7
+ $X2=3.925 $Y2=1.7
r134 28 32 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.875 $Y=1.325
+ $X2=6.875 $Y2=1.16
r135 28 30 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.875 $Y=1.325
+ $X2=6.875 $Y2=2.165
r136 24 32 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.875 $Y=0.995
+ $X2=6.875 $Y2=1.16
r137 24 26 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.875 $Y=0.995
+ $X2=6.875 $Y2=0.445
r138 23 63 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.01 $Y=1.16
+ $X2=5.935 $Y2=1.16
r139 22 32 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.8 $Y=1.16
+ $X2=6.875 $Y2=1.16
r140 22 23 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=6.8 $Y=1.16 $X2=6.01
+ $Y2=1.16
r141 18 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=1.325
+ $X2=5.935 $Y2=1.16
r142 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.935 $Y=1.325
+ $X2=5.935 $Y2=1.985
r143 15 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=0.995
+ $X2=5.935 $Y2=1.16
r144 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.935 $Y=0.995
+ $X2=5.935 $Y2=0.56
r145 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.69 $Y=1.535
+ $X2=3.69 $Y2=1.7
r146 11 13 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.69 $Y=1.535
+ $X2=3.69 $Y2=0.445
r147 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=1.7
r148 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=2.275
r149 2 55 600 $w=1.7e-07 $l=3.46627e-07 $layer=licon1_PDIFF $count=1 $X=4.69
+ $Y=1.485 $X2=4.865 $Y2=1.755
r150 2 45 600 $w=1.7e-07 $l=8.68101e-07 $layer=licon1_PDIFF $count=1 $X=4.69
+ $Y=1.485 $X2=4.865 $Y2=2.27
r151 1 40 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=4.295
+ $Y=0.235 $X2=4.42 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%A_560_47# 1 2 9 11 13 14 15 16 20 25 27 30
+ 34
c80 34 0 1.54454e-19 $X=3.33 $Y=0.995
c81 16 0 2.87957e-19 $X=3.27 $Y=2.34
r82 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.16 $X2=4.115 $Y2=1.16
r83 28 34 0.89609 $w=3.3e-07 $l=3.47851e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=3.33 $Y2=0.995
r84 28 30 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=4.115 $Y2=1.16
r85 27 33 18.4264 $w=2.8e-07 $l=4.19452e-07 $layer=LI1_cond $X=3.52 $Y=1.96
+ $X2=3.437 $Y2=2.34
r86 26 34 8.61065 $w=1.7e-07 $l=4.14246e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.33 $Y2=0.995
r87 26 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.96
r88 25 34 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=0.995
+ $X2=3.33 $Y2=0.995
r89 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=0.995
r90 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r91 20 22 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=2.935 $Y2=0.45
r92 16 33 3.65648 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.27 $Y=2.34
+ $X2=3.437 $Y2=2.34
r93 16 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.27 $Y=2.34
+ $X2=2.94 $Y2=2.34
r94 14 31 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=4.54 $Y=1.16
+ $X2=4.115 $Y2=1.16
r95 14 15 5.03009 $w=3.3e-07 $l=8.2e-08 $layer=POLY_cond $X=4.54 $Y=1.16
+ $X2=4.622 $Y2=1.16
r96 11 15 37.0704 $w=1.5e-07 $l=1.68953e-07 $layer=POLY_cond $X=4.63 $Y=0.995
+ $X2=4.622 $Y2=1.16
r97 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.63 $Y=0.995
+ $X2=4.63 $Y2=0.56
r98 7 15 37.0704 $w=1.5e-07 $l=1.68464e-07 $layer=POLY_cond $X=4.615 $Y=1.325
+ $X2=4.622 $Y2=1.16
r99 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.615 $Y=1.325
+ $X2=4.615 $Y2=1.985
r100 2 18 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.065 $X2=2.94 $Y2=2.34
r101 1 22 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.935 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%RESET_B 3 6 8 9 13 15 22
c36 9 0 1.26975e-19 $X=5.23 $Y=1.105
r37 14 22 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.05 $Y=1.16 $X2=5.29
+ $Y2=1.16
r38 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.16
+ $X2=5.05 $Y2=1.325
r39 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.16
+ $X2=5.05 $Y2=0.995
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=1.16 $X2=5.05 $Y2=1.16
r41 9 22 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=1.16
+ $X2=5.29 $Y2=1.16
r42 8 14 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.855 $Y=1.16
+ $X2=5.05 $Y2=1.16
r43 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.075 $Y=1.985
+ $X2=5.075 $Y2=1.325
r44 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.075 $Y=0.56
+ $X2=5.075 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%A_1308_47# 1 2 9 12 16 20 24 25 27 29
r40 25 30 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=1.16
+ $X2=7.325 $Y2=1.325
r41 25 29 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=1.16
+ $X2=7.325 $Y2=0.995
r42 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.16 $X2=7.31 $Y2=1.16
r43 22 27 0.189605 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=6.83 $Y=1.16
+ $X2=6.705 $Y2=1.16
r44 22 24 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.83 $Y=1.16
+ $X2=7.31 $Y2=1.16
r45 18 27 6.72893 $w=2.37e-07 $l=1.65e-07 $layer=LI1_cond $X=6.705 $Y=1.325
+ $X2=6.705 $Y2=1.16
r46 18 20 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=6.705 $Y=1.325
+ $X2=6.705 $Y2=2.165
r47 14 27 6.72893 $w=2.37e-07 $l=1.71377e-07 $layer=LI1_cond $X=6.692 $Y=0.995
+ $X2=6.705 $Y2=1.16
r48 14 16 24.8415 $w=2.23e-07 $l=4.85e-07 $layer=LI1_cond $X=6.692 $Y=0.995
+ $X2=6.692 $Y2=0.51
r49 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.35 $Y=1.985
+ $X2=7.35 $Y2=1.325
r50 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.35 $Y=0.56 $X2=7.35
+ $Y2=0.995
r51 2 20 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=6.54
+ $Y=1.845 $X2=6.665 $Y2=2.165
r52 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.54
+ $Y=0.235 $X2=6.665 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%VPWR 1 2 3 4 5 6 21 25 29 31 33 38 51 56 63
+ 64 67 70 74 80 82 89
r110 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r111 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r112 82 85 10.8734 $w=7.68e-07 $l=7e-07 $layer=LI1_cond $X=5.505 $Y=2.02
+ $X2=5.505 $Y2=2.72
r113 79 80 10.9687 $w=6.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.405 $Y=2.47
+ $X2=4.59 $Y2=2.47
r114 76 79 0.624817 $w=6.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.37 $Y=2.47
+ $X2=4.405 $Y2=2.47
r115 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r116 73 76 9.46152 $w=6.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.84 $Y=2.47
+ $X2=4.37 $Y2=2.47
r117 73 74 9.18355 $w=6.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=2.47
+ $X2=3.755 $Y2=2.47
r118 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 64 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r121 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r122 61 89 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.305 $Y=2.72
+ $X2=7.157 $Y2=2.72
r123 61 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.305 $Y=2.72
+ $X2=7.59 $Y2=2.72
r124 60 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r125 60 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r126 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r127 57 85 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=5.89 $Y=2.72
+ $X2=5.505 $Y2=2.72
r128 57 59 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.89 $Y=2.72
+ $X2=6.67 $Y2=2.72
r129 56 89 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=7.157 $Y2=2.72
r130 56 59 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=6.67 $Y2=2.72
r131 55 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r132 55 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 54 80 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=4.59 $Y2=2.72
r134 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r135 51 85 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=5.505 $Y2=2.72
r136 51 54 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=4.83 $Y2=2.72
r137 50 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r138 49 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.755 $Y2=2.72
r139 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r140 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r141 47 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 46 49 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r143 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r144 44 70 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r145 44 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r146 42 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r147 42 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r149 39 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r150 39 41 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r151 38 70 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r152 38 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r153 33 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r154 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 31 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r156 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r157 27 89 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.157 $Y=2.635
+ $X2=7.157 $Y2=2.72
r158 27 29 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=7.157 $Y=2.635
+ $X2=7.157 $Y2=2
r159 23 70 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r160 23 25 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r161 19 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r162 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r163 6 29 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=6.95
+ $Y=1.845 $X2=7.14 $Y2=2
r164 5 82 150 $w=1.7e-07 $l=7.98906e-07 $layer=licon1_PDIFF $count=4 $X=5.15
+ $Y=1.485 $X2=5.725 $Y2=2.02
r165 4 79 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.485 $X2=4.405 $Y2=2.34
r166 3 73 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.705
+ $Y=2.065 $X2=3.84 $Y2=2.3
r167 2 25 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r168 1 21 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%Q 1 2 7 8 9 10 11 12
r17 12 32 8.23174 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=6.235 $Y=2.21
+ $X2=6.235 $Y2=1.96
r18 11 32 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=6.235 $Y=1.87
+ $X2=6.235 $Y2=1.96
r19 10 11 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=6.235 $Y=1.53
+ $X2=6.235 $Y2=1.87
r20 9 10 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=6.235 $Y=1.19
+ $X2=6.235 $Y2=1.53
r21 8 9 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=6.235 $Y=0.85
+ $X2=6.235 $Y2=1.19
r22 7 8 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=6.235 $Y=0.51
+ $X2=6.235 $Y2=0.85
r23 2 32 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.01
+ $Y=1.485 $X2=6.145 $Y2=1.96
r24 1 7 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=6.01
+ $Y=0.235 $X2=6.145 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%Q_N 1 2 7 8 9 30 35
r13 16 35 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=7.605 $Y=1.915
+ $X2=7.605 $Y2=1.87
r14 8 35 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=7.605 $Y=1.85
+ $X2=7.605 $Y2=1.87
r15 8 9 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=7.605 $Y=1.935
+ $X2=7.605 $Y2=2.21
r16 8 16 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=7.605 $Y=1.935
+ $X2=7.605 $Y2=1.915
r17 7 30 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=7.56 $Y=0.425 $X2=7.65
+ $Y2=0.425
r18 7 30 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.65 $Y=0.595 $X2=7.65
+ $Y2=0.425
r19 7 8 47.9934 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=7.65 $Y=0.595
+ $X2=7.65 $Y2=1.785
r20 2 8 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.425
+ $Y=1.485 $X2=7.56 $Y2=1.96
r21 1 7 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.56 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_1%VGND 1 2 3 4 5 18 22 26 30 32 34 39 44 57 64
+ 65 68 71 74 79 85 87
c110 65 0 2.71124e-20 $X=7.59 $Y=0
c111 2 0 7.13094e-20 $X=1.905 $Y=0.235
r112 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r113 83 85 9.43642 $w=5.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.75 $Y=0.2
+ $X2=5.89 $Y2=0.2
r114 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r115 81 83 0.524596 $w=5.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.725 $Y=0.2
+ $X2=5.75 $Y2=0.2
r116 78 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r117 77 81 9.12797 $w=5.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.29 $Y=0.2
+ $X2=5.725 $Y2=0.2
r118 77 79 10.0659 $w=5.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.29 $Y=0.2
+ $X2=5.12 $Y2=0.2
r119 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r120 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r121 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r122 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r123 65 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r124 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r125 62 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=7.14
+ $Y2=0
r126 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.305 $Y=0
+ $X2=7.59 $Y2=0
r127 61 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r128 61 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=5.75
+ $Y2=0
r129 60 85 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=5.89
+ $Y2=0
r130 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r131 57 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=0 $X2=7.14
+ $Y2=0
r132 57 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=6.67 $Y2=0
r133 56 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r134 56 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r135 55 79 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.12
+ $Y2=0
r136 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r137 53 74 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.902
+ $Y2=0
r138 53 55 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.83
+ $Y2=0
r139 51 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r140 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r141 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r142 48 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r143 47 50 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r144 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r145 45 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r146 45 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r147 44 74 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=3.902 $Y2=0
r148 44 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=3.45 $Y2=0
r149 43 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r150 43 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r151 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r152 40 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r153 40 42 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r154 39 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r155 39 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r156 34 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r157 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r158 32 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r159 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r160 28 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0
r161 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0.38
r162 24 74 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.902 $Y=0.085
+ $X2=3.902 $Y2=0
r163 24 26 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=3.902 $Y=0.085
+ $X2=3.902 $Y2=0.445
r164 20 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r165 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r166 16 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r167 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r168 5 30 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=6.95
+ $Y=0.235 $X2=7.14 $Y2=0.38
r169 4 81 91 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_NDIFF $count=2 $X=5.15
+ $Y=0.235 $X2=5.725 $Y2=0.36
r170 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.235 $X2=3.9 $Y2=0.445
r171 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r172 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


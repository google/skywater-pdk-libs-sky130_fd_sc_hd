* File: sky130_fd_sc_hd__nand3b_4.spice.SKY130_FD_SC_HD__NAND3B_4.pxi
* Created: Thu Aug 27 14:29:59 2020
* 
x_PM_SKY130_FD_SC_HD__NAND3B_4%A_N N_A_N_M1023_g N_A_N_M1018_g A_N N_A_N_c_116_n
+ PM_SKY130_FD_SC_HD__NAND3B_4%A_N
x_PM_SKY130_FD_SC_HD__NAND3B_4%A_27_47# N_A_27_47#_M1023_s N_A_27_47#_M1018_s
+ N_A_27_47#_M1004_g N_A_27_47#_M1001_g N_A_27_47#_M1006_g N_A_27_47#_M1015_g
+ N_A_27_47#_M1008_g N_A_27_47#_M1019_g N_A_27_47#_M1014_g N_A_27_47#_M1020_g
+ N_A_27_47#_c_150_n N_A_27_47#_c_161_n N_A_27_47#_c_162_n N_A_27_47#_c_151_n
+ N_A_27_47#_c_152_n N_A_27_47#_c_206_p N_A_27_47#_c_153_n N_A_27_47#_c_154_n
+ N_A_27_47#_c_155_n N_A_27_47#_c_156_n PM_SKY130_FD_SC_HD__NAND3B_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND3B_4%B N_B_M1007_g N_B_M1010_g N_B_M1009_g N_B_M1011_g
+ N_B_M1012_g N_B_M1016_g N_B_M1013_g N_B_M1021_g B B B N_B_c_264_n
+ PM_SKY130_FD_SC_HD__NAND3B_4%B
x_PM_SKY130_FD_SC_HD__NAND3B_4%C N_C_M1000_g N_C_M1002_g N_C_M1003_g N_C_M1017_g
+ N_C_M1005_g N_C_M1022_g N_C_M1025_g N_C_M1024_g C C C C N_C_c_342_n
+ N_C_c_343_n PM_SKY130_FD_SC_HD__NAND3B_4%C
x_PM_SKY130_FD_SC_HD__NAND3B_4%VPWR N_VPWR_M1018_d N_VPWR_M1001_s N_VPWR_M1015_s
+ N_VPWR_M1020_s N_VPWR_M1011_s N_VPWR_M1021_s N_VPWR_M1002_d N_VPWR_M1017_d
+ N_VPWR_M1024_d N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n
+ N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n
+ N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_430_n
+ N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n VPWR N_VPWR_c_434_n
+ N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_416_n N_VPWR_c_438_n N_VPWR_c_439_n
+ PM_SKY130_FD_SC_HD__NAND3B_4%VPWR
x_PM_SKY130_FD_SC_HD__NAND3B_4%Y N_Y_M1004_s N_Y_M1008_s N_Y_M1001_d N_Y_M1019_d
+ N_Y_M1010_d N_Y_M1016_d N_Y_M1002_s N_Y_M1022_s N_Y_c_523_n N_Y_c_526_n
+ N_Y_c_547_n N_Y_c_550_n N_Y_c_552_n N_Y_c_527_n N_Y_c_572_n N_Y_c_528_n
+ N_Y_c_594_n N_Y_c_529_n N_Y_c_530_n N_Y_c_605_n N_Y_c_531_n N_Y_c_532_n Y Y
+ N_Y_c_525_n Y N_Y_c_534_n N_Y_c_535_n PM_SKY130_FD_SC_HD__NAND3B_4%Y
x_PM_SKY130_FD_SC_HD__NAND3B_4%VGND N_VGND_M1023_d N_VGND_M1000_d N_VGND_M1003_d
+ N_VGND_M1025_d N_VGND_c_657_n N_VGND_c_658_n N_VGND_c_659_n N_VGND_c_660_n
+ N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n
+ N_VGND_c_666_n VGND N_VGND_c_667_n N_VGND_c_668_n N_VGND_c_669_n
+ N_VGND_c_670_n PM_SKY130_FD_SC_HD__NAND3B_4%VGND
x_PM_SKY130_FD_SC_HD__NAND3B_4%A_215_47# N_A_215_47#_M1004_d N_A_215_47#_M1006_d
+ N_A_215_47#_M1014_d N_A_215_47#_M1009_s N_A_215_47#_M1013_s
+ N_A_215_47#_c_743_n PM_SKY130_FD_SC_HD__NAND3B_4%A_215_47#
x_PM_SKY130_FD_SC_HD__NAND3B_4%A_633_47# N_A_633_47#_M1007_d N_A_633_47#_M1012_d
+ N_A_633_47#_M1000_s N_A_633_47#_M1005_s N_A_633_47#_c_777_n
+ N_A_633_47#_c_778_n N_A_633_47#_c_791_n N_A_633_47#_c_779_n
+ N_A_633_47#_c_799_n N_A_633_47#_c_780_n N_A_633_47#_c_781_n
+ PM_SKY130_FD_SC_HD__NAND3B_4%A_633_47#
cc_1 VNB N_A_N_M1023_g 0.0256913f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB A_N 0.00171637f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_3 VNB N_A_N_c_116_n 0.0273695f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_4 VNB N_A_27_47#_M1004_g 0.0207485f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_5 VNB N_A_27_47#_M1001_g 5.53572e-19 $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_6 VNB N_A_27_47#_M1006_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1015_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1008_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1019_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1014_g 0.0175122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1020_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_150_n 0.0183576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_151_n 0.00970788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_152_n 0.00406828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_153_n 0.00993195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_154_n 0.0188025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_155_n 0.03161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_156_n 0.0581706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B_M1007_g 0.017661f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_B_M1010_g 4.13233e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_21 VNB N_B_M1009_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=1.16
cc_22 VNB N_B_M1011_g 4.49286e-19 $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=1.305
cc_23 VNB N_B_M1012_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_B_M1016_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_B_M1013_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B_M1021_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB B 0.00271316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_B_c_264_n 0.0624411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_C_M1000_g 0.0238914f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_30 VNB N_C_M1002_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_31 VNB N_C_M1003_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=1.16
cc_32 VNB N_C_M1017_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=1.305
cc_33 VNB N_C_M1005_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_C_M1022_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_C_M1025_g 0.0237664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_C_M1024_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB C 0.00341134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_C_c_342_n 0.0304355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_C_c_343_n 0.0678784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_416_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_523_n 0.00736934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB Y 0.00246646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_525_n 0.00304777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_657_n 0.00885089f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=1.305
cc_45 VNB N_VGND_c_658_n 0.0082423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_659_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_660_n 0.035793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_661_n 0.092353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_662_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_663_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_664_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_665_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_666_n 0.00634414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_667_n 0.0171188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_668_n 0.0134401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_669_n 0.367788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_670_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_215_47#_c_743_n 0.00503226f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_633_47#_c_777_n 0.00935305f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_60 VNB N_A_633_47#_c_778_n 0.00835607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_633_47#_c_779_n 0.004418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_633_47#_c_780_n 0.0036494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_633_47#_c_781_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VPB N_A_N_M1018_g 0.0316181f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_65 VPB N_A_N_c_116_n 0.00641609f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_66 VPB N_A_27_47#_M1001_g 0.0264483f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_67 VPB N_A_27_47#_M1015_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_M1019_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_M1020_g 0.0194268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_161_n 0.0085685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_162_n 0.0336524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_154_n 0.00660992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B_M1010_g 0.0186547f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_74 VPB N_B_M1011_g 0.0191571f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=1.305
cc_75 VPB N_B_M1016_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_B_M1021_g 0.026721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_C_M1002_g 0.026721f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_78 VPB N_C_M1017_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=1.305
cc_79 VPB N_C_M1022_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_C_M1024_g 0.0264483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_417_n 0.0245646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_418_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_419_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_420_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_421_n 0.0153464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_422_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_423_n 0.0501811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_424_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_425_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_426_n 0.0172923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_427_n 0.00323604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_428_n 0.0172923f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_429_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_430_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_431_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_432_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_433_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_434_n 0.0177718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_435_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_436_n 0.0134401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_416_n 0.054605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_438_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_439_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_Y_c_526_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_Y_c_527_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_Y_c_528_n 0.0128506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_Y_c_529_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_Y_c_530_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_Y_c_531_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_Y_c_532_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB Y 0.00198971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_Y_c_534_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_Y_c_535_n 0.00635302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 N_A_N_c_116_n N_A_27_47#_M1001_g 2.68352e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_N_M1023_g N_A_27_47#_c_150_n 0.0108374f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_N_M1018_g N_A_27_47#_c_161_n 0.00338942f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_N_M1018_g N_A_27_47#_c_162_n 0.0095746f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_N_M1023_g N_A_27_47#_c_151_n 0.0112031f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_119 A_N N_A_27_47#_c_151_n 0.0251973f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_120 N_A_N_c_116_n N_A_27_47#_c_151_n 0.00505312f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_N_M1023_g N_A_27_47#_c_152_n 0.00291964f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_122 A_N N_A_27_47#_c_152_n 0.0135639f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_123 N_A_N_c_116_n N_A_27_47#_c_152_n 8.35206e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_N_M1023_g N_A_27_47#_c_153_n 0.00163224f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_125 N_A_N_M1023_g N_A_27_47#_c_154_n 0.0136859f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_126 A_N N_A_27_47#_c_154_n 0.015054f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_127 A_N N_A_27_47#_c_155_n 7.26316e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_128 N_A_N_c_116_n N_A_27_47#_c_155_n 0.0152652f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_N_M1018_g N_VPWR_c_417_n 0.0057288f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_130 A_N N_VPWR_c_417_n 0.0150811f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_131 N_A_N_c_116_n N_VPWR_c_417_n 0.00386161f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_N_M1018_g N_VPWR_c_434_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_N_M1018_g N_VPWR_c_416_n 0.0117818f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_N_M1023_g N_VGND_c_657_n 0.0044954f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_135 N_A_N_M1023_g N_VGND_c_667_n 0.00422241f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_136 N_A_N_M1023_g N_VGND_c_669_n 0.00797683f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1014_g N_B_M1007_g 0.0279197f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1020_g N_B_M1010_g 0.0279197f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_156_n N_B_c_264_n 0.0279197f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1001_g N_VPWR_c_417_n 0.00427388f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_c_161_n N_VPWR_c_417_n 0.0402242f $X=0.255 $Y=1.615 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_c_151_n N_VPWR_c_417_n 0.00855453f $X=1.005 $Y=0.81 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_c_152_n N_VPWR_c_417_n 0.0244885f $X=1.145 $Y=1.075 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_155_n N_VPWR_c_417_n 0.00639477f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_M1015_g N_VPWR_c_418_n 0.00146448f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_M1019_g N_VPWR_c_418_n 0.00146448f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_M1020_g N_VPWR_c_419_n 0.00146448f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_M1001_g N_VPWR_c_424_n 0.00541359f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_M1015_g N_VPWR_c_424_n 0.00541359f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_27_47#_M1019_g N_VPWR_c_426_n 0.00540367f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_M1020_g N_VPWR_c_426_n 0.00421248f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_162_n N_VPWR_c_434_n 0.0217551f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_153 N_A_27_47#_M1018_s N_VPWR_c_416_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_M1001_g N_VPWR_c_416_n 0.0108276f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_27_47#_M1015_g N_VPWR_c_416_n 0.00950154f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_M1019_g N_VPWR_c_416_n 0.00945548f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_M1020_g N_VPWR_c_416_n 0.00573823f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_c_162_n N_VPWR_c_416_n 0.0128119f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_159 N_A_27_47#_M1004_g N_Y_c_523_n 0.0068614f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A_27_47#_M1006_g N_Y_c_523_n 0.0112239f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_161 N_A_27_47#_M1008_g N_Y_c_523_n 0.0112192f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_27_47#_M1014_g N_Y_c_523_n 0.0117996f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_151_n N_Y_c_523_n 0.0088422f $X=1.005 $Y=0.81 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_206_p N_Y_c_523_n 0.0864637f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_156_n N_Y_c_523_n 0.0062366f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_27_47#_M1001_g N_Y_c_526_n 0.00331821f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_27_47#_M1015_g N_Y_c_526_n 0.00149073f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_206_p N_Y_c_526_n 0.026643f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_156_n N_Y_c_526_n 0.00206439f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_27_47#_M1001_g N_Y_c_547_n 0.00902485f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_27_47#_M1015_g N_Y_c_547_n 0.00974075f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1019_g N_Y_c_547_n 6.1927e-19 $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_27_47#_M1019_g N_Y_c_550_n 0.00512562f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1020_g N_Y_c_550_n 0.00631111f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1020_g N_Y_c_552_n 5.2007e-19 $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_27_47#_M1020_g Y 0.00351106f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_206_p Y 0.0164737f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_156_n Y 0.00351106f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_27_47#_M1014_g N_Y_c_525_n 0.00351106f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1015_g N_Y_c_534_n 0.0120357f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_27_47#_M1019_g N_Y_c_534_n 0.0120357f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_206_p N_Y_c_534_n 0.0627659f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_156_n N_Y_c_534_n 0.0019951f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1015_g N_Y_c_535_n 4.81356e-19 $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1019_g N_Y_c_535_n 0.0063824f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_27_47#_M1020_g N_Y_c_535_n 0.0212342f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_156_n N_Y_c_535_n 0.00204726f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_151_n N_VGND_M1023_d 0.00285834f $X=1.005 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_27_47#_M1004_g N_VGND_c_657_n 0.00231165f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_151_n N_VGND_c_657_n 0.0191474f $X=1.005 $Y=0.81 $X2=0 $Y2=0
cc_191 N_A_27_47#_M1004_g N_VGND_c_661_n 0.00357877f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A_27_47#_M1006_g N_VGND_c_661_n 0.00357877f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A_27_47#_M1008_g N_VGND_c_661_n 0.00357877f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A_27_47#_M1014_g N_VGND_c_661_n 0.00357877f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_151_n N_VGND_c_661_n 0.00300337f $X=1.005 $Y=0.81 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_150_n N_VGND_c_667_n 0.0217307f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_151_n N_VGND_c_667_n 0.00203746f $X=1.005 $Y=0.81 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_M1023_s N_VGND_c_669_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_M1004_g N_VGND_c_669_n 0.00655123f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_27_47#_M1006_g N_VGND_c_669_n 0.00522516f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_27_47#_M1008_g N_VGND_c_669_n 0.00522516f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1014_g N_VGND_c_669_n 0.00525237f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_150_n N_VGND_c_669_n 0.0128045f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_151_n N_VGND_c_669_n 0.0107957f $X=1.005 $Y=0.81 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_151_n N_A_215_47#_M1004_d 0.00401649f $X=1.005 $Y=0.81
+ $X2=-0.19 $Y2=-0.24
cc_206 N_A_27_47#_M1004_g N_A_215_47#_c_743_n 0.0103313f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1006_g N_A_215_47#_c_743_n 0.00866705f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_M1008_g N_A_215_47#_c_743_n 0.00866705f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_M1014_g N_A_215_47#_c_743_n 0.00866705f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_151_n N_A_215_47#_c_743_n 0.0135762f $X=1.005 $Y=0.81 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_206_p N_A_215_47#_c_743_n 0.00347188f $X=2.46 $Y=1.16 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_155_n N_A_215_47#_c_743_n 9.07366e-19 $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_213 B C 0.0121822f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_214 N_B_c_264_n C 8.71733e-19 $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_215 B N_C_c_342_n 8.07044e-19 $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_216 N_B_c_264_n N_C_c_342_n 0.00741568f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B_M1010_g N_VPWR_c_419_n 0.00146448f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B_M1011_g N_VPWR_c_420_n 0.00146448f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B_M1016_g N_VPWR_c_420_n 0.00146448f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B_M1021_g N_VPWR_c_421_n 0.0033532f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B_M1010_g N_VPWR_c_428_n 0.00421248f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_222 N_B_M1011_g N_VPWR_c_428_n 0.00540367f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B_M1016_g N_VPWR_c_435_n 0.00541359f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_224 N_B_M1021_g N_VPWR_c_435_n 0.00541359f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B_M1010_g N_VPWR_c_416_n 0.00573823f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B_M1011_g N_VPWR_c_416_n 0.00945548f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B_M1016_g N_VPWR_c_416_n 0.00950154f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_228 N_B_M1021_g N_VPWR_c_416_n 0.0108276f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B_M1007_g N_Y_c_523_n 0.00121164f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_230 N_B_M1010_g N_Y_c_550_n 5.2007e-19 $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_231 N_B_M1010_g N_Y_c_552_n 0.00631111f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_232 N_B_M1011_g N_Y_c_552_n 0.00512562f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_233 N_B_M1011_g N_Y_c_527_n 0.0120357f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_234 N_B_M1016_g N_Y_c_527_n 0.0120357f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_235 N_B_c_264_n N_Y_c_527_n 0.0019951f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B_M1011_g N_Y_c_572_n 6.1927e-19 $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_237 N_B_M1016_g N_Y_c_572_n 0.00974075f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_238 N_B_M1021_g N_Y_c_572_n 0.0145598f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_239 N_B_M1021_g N_Y_c_528_n 0.0147646f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_240 B N_Y_c_528_n 0.0126419f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_241 N_B_M1016_g N_Y_c_531_n 0.00149073f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_242 N_B_M1021_g N_Y_c_531_n 0.00149073f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_243 B N_Y_c_531_n 0.026643f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_244 N_B_c_264_n N_Y_c_531_n 0.00206439f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B_M1010_g Y 0.00493083f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_246 N_B_M1011_g Y 8.21208e-19 $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_247 B Y 0.0156785f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_248 N_B_c_264_n Y 0.00977999f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_249 N_B_M1007_g N_Y_c_525_n 0.00410511f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_250 N_B_M1010_g N_Y_c_535_n 0.0207f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B_M1011_g N_Y_c_535_n 0.0063824f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_252 N_B_M1016_g N_Y_c_535_n 4.81356e-19 $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_253 B N_Y_c_535_n 0.0521195f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_254 N_B_c_264_n N_Y_c_535_n 0.00212545f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B_M1013_g N_VGND_c_658_n 0.00231165f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_256 N_B_M1007_g N_VGND_c_661_n 0.00357877f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_257 N_B_M1009_g N_VGND_c_661_n 0.00357877f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_258 N_B_M1012_g N_VGND_c_661_n 0.00357877f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_259 N_B_M1013_g N_VGND_c_661_n 0.00357877f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_260 N_B_M1007_g N_VGND_c_669_n 0.00525237f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_261 N_B_M1009_g N_VGND_c_669_n 0.00522516f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_262 N_B_M1012_g N_VGND_c_669_n 0.00522516f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_263 N_B_M1013_g N_VGND_c_669_n 0.00655123f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_264 N_B_M1007_g N_A_215_47#_c_743_n 0.0109603f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_265 N_B_M1009_g N_A_215_47#_c_743_n 0.00866705f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_266 N_B_M1012_g N_A_215_47#_c_743_n 0.00866705f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_267 N_B_M1013_g N_A_215_47#_c_743_n 0.00866705f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_268 N_B_M1007_g N_A_633_47#_c_777_n 0.00420272f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_269 N_B_M1009_g N_A_633_47#_c_777_n 0.0112239f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_270 N_B_M1012_g N_A_633_47#_c_777_n 0.0112239f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_271 N_B_M1013_g N_A_633_47#_c_777_n 0.0142655f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_272 B N_A_633_47#_c_777_n 0.0893207f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_273 N_B_c_264_n N_A_633_47#_c_777_n 0.00630644f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_274 N_C_M1002_g N_VPWR_c_421_n 0.0033532f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_275 N_C_M1017_g N_VPWR_c_422_n 0.00146448f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_276 N_C_M1022_g N_VPWR_c_422_n 0.00146448f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_277 N_C_M1024_g N_VPWR_c_423_n 0.0233944f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_278 N_C_M1002_g N_VPWR_c_430_n 0.00541359f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_279 N_C_M1017_g N_VPWR_c_430_n 0.00541359f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_280 N_C_M1022_g N_VPWR_c_432_n 0.00541359f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_281 N_C_M1024_g N_VPWR_c_432_n 0.00541359f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_282 N_C_M1002_g N_VPWR_c_416_n 0.0108276f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_283 N_C_M1017_g N_VPWR_c_416_n 0.00950154f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_284 N_C_M1022_g N_VPWR_c_416_n 0.00950154f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_285 N_C_M1024_g N_VPWR_c_416_n 0.0109543f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_286 N_C_M1002_g N_Y_c_528_n 0.0147646f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_287 C N_Y_c_528_n 0.0400987f $X=6.17 $Y=1.105 $X2=0 $Y2=0
cc_288 N_C_c_342_n N_Y_c_528_n 0.00729564f $X=5.215 $Y=1.16 $X2=0 $Y2=0
cc_289 N_C_M1002_g N_Y_c_594_n 0.0145598f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_290 N_C_M1017_g N_Y_c_594_n 0.00975139f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_291 N_C_M1022_g N_Y_c_594_n 6.1949e-19 $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_292 N_C_M1017_g N_Y_c_529_n 0.0120357f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_293 N_C_M1022_g N_Y_c_529_n 0.0120357f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_294 C N_Y_c_529_n 0.0366837f $X=6.17 $Y=1.105 $X2=0 $Y2=0
cc_295 N_C_c_343_n N_Y_c_529_n 0.0019951f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_296 N_C_M1022_g N_Y_c_530_n 0.00149073f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_297 N_C_M1024_g N_Y_c_530_n 0.00338303f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_298 C N_Y_c_530_n 0.0262578f $X=6.17 $Y=1.105 $X2=0 $Y2=0
cc_299 N_C_c_343_n N_Y_c_530_n 0.00206439f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_300 N_C_M1017_g N_Y_c_605_n 6.1949e-19 $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_301 N_C_M1022_g N_Y_c_605_n 0.00975139f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_302 N_C_M1024_g N_Y_c_605_n 0.00902485f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_303 N_C_M1002_g N_Y_c_532_n 0.00149073f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_304 N_C_M1017_g N_Y_c_532_n 0.00149073f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_305 C N_Y_c_532_n 0.026643f $X=6.17 $Y=1.105 $X2=0 $Y2=0
cc_306 N_C_c_343_n N_Y_c_532_n 0.00206439f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_307 N_C_M1000_g N_VGND_c_658_n 0.00321269f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_308 N_C_M1003_g N_VGND_c_659_n 0.00146448f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_309 N_C_M1005_g N_VGND_c_659_n 0.00146448f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_310 N_C_M1025_g N_VGND_c_660_n 0.0162028f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_311 N_C_M1000_g N_VGND_c_663_n 0.00422241f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_312 N_C_M1003_g N_VGND_c_663_n 0.00422241f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_313 N_C_M1005_g N_VGND_c_665_n 0.00422241f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_314 N_C_M1025_g N_VGND_c_665_n 0.00541359f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_315 N_C_M1000_g N_VGND_c_669_n 0.00702263f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_316 N_C_M1003_g N_VGND_c_669_n 0.00569656f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_317 N_C_M1005_g N_VGND_c_669_n 0.00569656f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_318 N_C_M1025_g N_VGND_c_669_n 0.0109543f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_319 N_C_M1000_g N_A_633_47#_c_778_n 0.0112581f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_320 C N_A_633_47#_c_778_n 0.039638f $X=6.17 $Y=1.105 $X2=0 $Y2=0
cc_321 N_C_c_342_n N_A_633_47#_c_778_n 0.00753289f $X=5.215 $Y=1.16 $X2=0 $Y2=0
cc_322 N_C_M1000_g N_A_633_47#_c_791_n 0.00907724f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_323 N_C_M1003_g N_A_633_47#_c_791_n 0.00620543f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_324 N_C_M1005_g N_A_633_47#_c_791_n 5.19281e-19 $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_325 N_C_M1003_g N_A_633_47#_c_779_n 0.00890471f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_326 N_C_M1005_g N_A_633_47#_c_779_n 0.0100649f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_327 N_C_M1025_g N_A_633_47#_c_779_n 0.00268058f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_328 C N_A_633_47#_c_779_n 0.0624206f $X=6.17 $Y=1.105 $X2=0 $Y2=0
cc_329 N_C_c_343_n N_A_633_47#_c_779_n 0.00419427f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_330 N_C_M1003_g N_A_633_47#_c_799_n 5.19281e-19 $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_331 N_C_M1005_g N_A_633_47#_c_799_n 0.00620543f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_332 N_C_M1025_g N_A_633_47#_c_799_n 0.00528656f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_333 N_C_M1000_g N_A_633_47#_c_780_n 0.00137399f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_334 N_C_M1000_g N_A_633_47#_c_781_n 0.00116017f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_335 N_C_M1003_g N_A_633_47#_c_781_n 0.00116017f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_336 C N_A_633_47#_c_781_n 0.0265408f $X=6.17 $Y=1.105 $X2=0 $Y2=0
cc_337 N_C_c_343_n N_A_633_47#_c_781_n 0.00213429f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_338 N_VPWR_c_416_n N_Y_M1001_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_339 N_VPWR_c_416_n N_Y_M1019_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_340 N_VPWR_c_416_n N_Y_M1010_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_341 N_VPWR_c_416_n N_Y_M1016_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_342 N_VPWR_c_416_n N_Y_M1002_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_343 N_VPWR_c_416_n N_Y_M1022_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_344 N_VPWR_c_417_n N_Y_c_526_n 0.0110887f $X=0.68 $Y=1.66 $X2=0 $Y2=0
cc_345 N_VPWR_c_424_n N_Y_c_547_n 0.0189039f $X=1.955 $Y=2.72 $X2=0 $Y2=0
cc_346 N_VPWR_c_416_n N_Y_c_547_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_347 N_VPWR_c_426_n N_Y_c_550_n 0.0184921f $X=2.795 $Y=2.72 $X2=0 $Y2=0
cc_348 N_VPWR_c_416_n N_Y_c_550_n 0.012098f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_349 N_VPWR_c_428_n N_Y_c_552_n 0.0184921f $X=3.635 $Y=2.72 $X2=0 $Y2=0
cc_350 N_VPWR_c_416_n N_Y_c_552_n 0.012098f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_351 N_VPWR_M1011_s N_Y_c_527_n 0.00167154f $X=3.585 $Y=1.485 $X2=0 $Y2=0
cc_352 N_VPWR_c_420_n N_Y_c_527_n 0.0129161f $X=3.72 $Y=2 $X2=0 $Y2=0
cc_353 N_VPWR_c_435_n N_Y_c_572_n 0.0189039f $X=4.475 $Y=2.72 $X2=0 $Y2=0
cc_354 N_VPWR_c_416_n N_Y_c_572_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_355 N_VPWR_M1021_s N_Y_c_528_n 0.00296777f $X=4.425 $Y=1.485 $X2=0 $Y2=0
cc_356 N_VPWR_M1002_d N_Y_c_528_n 0.00296777f $X=4.955 $Y=1.485 $X2=0 $Y2=0
cc_357 N_VPWR_c_421_n N_Y_c_528_n 0.0568271f $X=4.56 $Y=2 $X2=0 $Y2=0
cc_358 N_VPWR_c_430_n N_Y_c_594_n 0.0189039f $X=5.835 $Y=2.72 $X2=0 $Y2=0
cc_359 N_VPWR_c_416_n N_Y_c_594_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_360 N_VPWR_M1017_d N_Y_c_529_n 0.00167154f $X=5.785 $Y=1.485 $X2=0 $Y2=0
cc_361 N_VPWR_c_422_n N_Y_c_529_n 0.0129161f $X=5.92 $Y=2 $X2=0 $Y2=0
cc_362 N_VPWR_c_423_n N_Y_c_530_n 0.0108967f $X=6.84 $Y=1.66 $X2=0 $Y2=0
cc_363 N_VPWR_c_432_n N_Y_c_605_n 0.0189039f $X=6.675 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_416_n N_Y_c_605_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_M1015_s N_Y_c_534_n 0.00167154f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_366 N_VPWR_c_418_n N_Y_c_534_n 0.0129161f $X=2.04 $Y=2 $X2=0 $Y2=0
cc_367 N_VPWR_M1020_s N_Y_c_535_n 0.0016762f $X=2.745 $Y=1.485 $X2=0 $Y2=0
cc_368 N_VPWR_c_419_n N_Y_c_535_n 0.0132033f $X=2.88 $Y=2.34 $X2=0 $Y2=0
cc_369 N_VPWR_c_426_n N_Y_c_535_n 0.00219876f $X=2.795 $Y=2.72 $X2=0 $Y2=0
cc_370 N_VPWR_c_428_n N_Y_c_535_n 0.00219876f $X=3.635 $Y=2.72 $X2=0 $Y2=0
cc_371 N_VPWR_c_416_n N_Y_c_535_n 0.00906442f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_c_423_n N_VGND_c_660_n 0.0137178f $X=6.84 $Y=1.66 $X2=0 $Y2=0
cc_373 N_Y_M1004_s N_VGND_c_669_n 0.00216833f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_374 N_Y_M1008_s N_VGND_c_669_n 0.00216833f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_375 N_Y_c_523_n N_A_215_47#_M1006_d 0.00162207f $X=2.795 $Y=0.77 $X2=0 $Y2=0
cc_376 N_Y_c_523_n N_A_215_47#_M1014_d 0.00206479f $X=2.795 $Y=0.77 $X2=0 $Y2=0
cc_377 N_Y_M1004_s N_A_215_47#_c_743_n 0.00305599f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_378 N_Y_M1008_s N_A_215_47#_c_743_n 0.00305599f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_379 N_Y_c_523_n N_A_215_47#_c_743_n 0.0783214f $X=2.795 $Y=0.77 $X2=0 $Y2=0
cc_380 Y N_A_215_47#_c_743_n 0.0029984f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_381 N_Y_c_523_n N_A_633_47#_c_777_n 0.0121859f $X=2.795 $Y=0.77 $X2=0 $Y2=0
cc_382 N_Y_c_528_n N_A_633_47#_c_777_n 0.0109732f $X=5.335 $Y=1.555 $X2=0 $Y2=0
cc_383 N_Y_c_535_n N_A_633_47#_c_777_n 0.00491983f $X=3.465 $Y=1.725 $X2=0 $Y2=0
cc_384 N_VGND_c_669_n N_A_215_47#_M1004_d 0.00209344f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_385 N_VGND_c_669_n N_A_215_47#_M1006_d 0.00215227f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_669_n N_A_215_47#_M1014_d 0.00215227f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_387 N_VGND_c_669_n N_A_215_47#_M1009_s 0.00215227f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_388 N_VGND_c_669_n N_A_215_47#_M1013_s 0.00209344f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_657_n N_A_215_47#_c_743_n 0.0166761f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_390 N_VGND_c_658_n N_A_215_47#_c_743_n 0.0166761f $X=5.08 $Y=0.38 $X2=0 $Y2=0
cc_391 N_VGND_c_661_n N_A_215_47#_c_743_n 0.208356f $X=4.915 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_669_n N_A_215_47#_c_743_n 0.132034f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_669_n N_A_633_47#_M1007_d 0.00216833f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_394 N_VGND_c_669_n N_A_633_47#_M1012_d 0.00216833f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_395 N_VGND_c_669_n N_A_633_47#_M1000_s 0.00215201f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_669_n N_A_633_47#_M1005_s 0.00215201f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_M1000_d N_A_633_47#_c_778_n 0.00285834f $X=4.955 $Y=0.235 $X2=0
+ $Y2=0
cc_398 N_VGND_c_658_n N_A_633_47#_c_778_n 0.0191473f $X=5.08 $Y=0.38 $X2=0 $Y2=0
cc_399 N_VGND_c_661_n N_A_633_47#_c_778_n 0.00296114f $X=4.915 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_663_n N_A_633_47#_c_778_n 0.00203746f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_669_n N_A_633_47#_c_778_n 0.00998562f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_402 N_VGND_c_663_n N_A_633_47#_c_791_n 0.0188551f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_403 N_VGND_c_669_n N_A_633_47#_c_791_n 0.0122069f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_404 N_VGND_M1003_d N_A_633_47#_c_779_n 0.00162148f $X=5.785 $Y=0.235 $X2=0
+ $Y2=0
cc_405 N_VGND_c_659_n N_A_633_47#_c_779_n 0.0122675f $X=5.92 $Y=0.38 $X2=0 $Y2=0
cc_406 N_VGND_c_660_n N_A_633_47#_c_779_n 0.0087974f $X=6.84 $Y=0.38 $X2=0 $Y2=0
cc_407 N_VGND_c_663_n N_A_633_47#_c_779_n 0.00203746f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_665_n N_A_633_47#_c_779_n 0.00203746f $X=6.675 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_669_n N_A_633_47#_c_779_n 0.00845923f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_665_n N_A_633_47#_c_799_n 0.0188551f $X=6.675 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_669_n N_A_633_47#_c_799_n 0.0122069f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_412 N_A_215_47#_c_743_n N_A_633_47#_M1007_d 0.00305599f $X=4.56 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_413 N_A_215_47#_c_743_n N_A_633_47#_M1012_d 0.00305599f $X=4.56 $Y=0.38 $X2=0
+ $Y2=0
cc_414 N_A_215_47#_M1009_s N_A_633_47#_c_777_n 0.00162207f $X=3.585 $Y=0.235
+ $X2=0 $Y2=0
cc_415 N_A_215_47#_M1013_s N_A_633_47#_c_777_n 0.00111257f $X=4.425 $Y=0.235
+ $X2=0 $Y2=0
cc_416 N_A_215_47#_c_743_n N_A_633_47#_c_777_n 0.0838291f $X=4.56 $Y=0.38 $X2=0
+ $Y2=0
cc_417 N_A_215_47#_M1013_s N_A_633_47#_c_780_n 0.00209037f $X=4.425 $Y=0.235
+ $X2=0 $Y2=0

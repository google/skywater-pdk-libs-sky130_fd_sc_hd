* File: sky130_fd_sc_hd__bufinv_16.pex.spice
* Created: Thu Aug 27 14:10:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUFINV_16%A 3 7 11 15 19 23 25 32 33
c66 32 0 1.44067e-19 $X=1.02 $Y=1.16
c67 23 0 1.25206e-19 $X=1.31 $Y=1.985
c68 19 0 1.25206e-19 $X=1.31 $Y=0.56
r69 31 33 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.31 $Y2=1.16
r70 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.02
+ $Y=1.16 $X2=1.02 $Y2=1.16
r71 29 31 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.02 $Y2=1.16
r72 27 29 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.89
+ $Y2=1.16
r73 25 32 43.5318 $w=1.98e-07 $l=7.85e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=1.02 $Y2=1.175
r74 21 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r75 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r76 17 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r77 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r78 13 29 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r79 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r80 9 29 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.16
r81 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r82 5 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r83 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295 $X2=0.47
+ $Y2=1.985
r84 1 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r85 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_16%A_27_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 72 73 74 77 81 86 88 94 98 101 103 112
c198 112 0 1.44067e-19 $X=3.83 $Y=1.16
c199 94 0 1.39258e-19 $X=3.56 $Y=1.16
c200 59 0 1.25206e-19 $X=3.83 $Y=1.985
c201 55 0 1.25206e-19 $X=3.83 $Y=0.56
r202 109 110 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.41 $Y2=1.16
r203 108 109 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r204 107 108 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r205 95 112 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=3.56 $Y=1.16
+ $X2=3.83 $Y2=1.16
r206 95 110 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.56 $Y=1.16
+ $X2=3.41 $Y2=1.16
r207 94 95 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.56
+ $Y=1.16 $X2=3.56 $Y2=1.16
r208 92 107 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=1.86 $Y=1.16
+ $X2=2.15 $Y2=1.16
r209 92 104 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=1.86 $Y=1.16
+ $X2=1.73 $Y2=1.16
r210 91 94 94.2727 $w=1.98e-07 $l=1.7e-06 $layer=LI1_cond $X=1.86 $Y=1.175
+ $X2=3.56 $Y2=1.175
r211 91 92 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.86
+ $Y=1.16 $X2=1.86 $Y2=1.16
r212 89 103 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.175
+ $X2=1.52 $Y2=1.175
r213 89 91 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.605 $Y=1.175
+ $X2=1.86 $Y2=1.175
r214 88 101 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.445
+ $X2=1.52 $Y2=1.53
r215 87 103 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.52 $Y=1.275
+ $X2=1.52 $Y2=1.175
r216 87 88 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.52 $Y=1.275
+ $X2=1.52 $Y2=1.445
r217 86 103 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.52 $Y=1.075
+ $X2=1.52 $Y2=1.175
r218 85 98 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.905
+ $X2=1.52 $Y2=0.82
r219 85 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.52 $Y=0.905
+ $X2=1.52 $Y2=1.075
r220 81 83 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.1 $Y=1.63 $X2=1.1
+ $Y2=2.31
r221 79 101 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.1 $Y=1.53
+ $X2=1.52 $Y2=1.53
r222 79 81 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.1 $Y=1.615
+ $X2=1.1 $Y2=1.63
r223 75 98 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.1 $Y=0.82
+ $X2=1.52 $Y2=0.82
r224 75 77 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=0.735
+ $X2=1.1 $Y2=0.4
r225 73 79 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.53
+ $X2=1.1 $Y2=1.53
r226 73 74 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=1.53
+ $X2=0.425 $Y2=1.53
r227 71 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=1.1 $Y2=0.82
r228 71 72 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.82
+ $X2=0.425 $Y2=0.82
r229 67 69 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r230 65 74 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r231 65 67 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r232 61 72 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.425 $Y2=0.82
r233 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.735
+ $X2=0.26 $Y2=0.4
r234 57 112 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.16
r235 57 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.985
r236 53 112 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=1.16
r237 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=0.56
r238 49 110 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r239 49 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r240 45 110 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r241 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r242 41 109 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r243 41 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r244 37 109 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r245 37 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r246 33 108 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r247 33 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r248 29 108 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r249 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r250 25 107 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r251 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r252 21 107 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r253 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r254 17 104 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r255 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r256 13 104 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r257 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r258 4 83 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.31
r259 4 81 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.63
r260 3 69 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r261 3 67 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r262 2 77 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r263 1 63 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_16%A_361_47# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 153 157 158 159 160 163 167 171 173 177 181 186 188 194 197 198
+ 200 203 205 224
c464 224 0 1.39258e-19 $X=10.55 $Y=1.16
c465 160 0 1.25206e-19 $X=2.105 $Y=1.53
c466 158 0 1.25206e-19 $X=2.105 $Y=0.82
r467 221 222 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.71 $Y=1.16
+ $X2=10.13 $Y2=1.16
r468 220 221 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.29 $Y=1.16
+ $X2=9.71 $Y2=1.16
r469 219 220 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.87 $Y=1.16
+ $X2=9.29 $Y2=1.16
r470 218 219 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.45 $Y=1.16
+ $X2=8.87 $Y2=1.16
r471 217 218 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.03 $Y=1.16
+ $X2=8.45 $Y2=1.16
r472 216 217 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.61 $Y=1.16
+ $X2=8.03 $Y2=1.16
r473 215 216 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.19 $Y=1.16
+ $X2=7.61 $Y2=1.16
r474 214 215 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.77 $Y=1.16
+ $X2=7.19 $Y2=1.16
r475 213 214 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.35 $Y=1.16
+ $X2=6.77 $Y2=1.16
r476 212 213 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.93 $Y=1.16
+ $X2=6.35 $Y2=1.16
r477 211 212 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.51 $Y=1.16
+ $X2=5.93 $Y2=1.16
r478 210 211 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.09 $Y=1.16
+ $X2=5.51 $Y2=1.16
r479 209 210 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.67 $Y=1.16
+ $X2=5.09 $Y2=1.16
r480 195 224 91.0912 $w=2.7e-07 $l=4.1e-07 $layer=POLY_cond $X=10.14 $Y=1.16
+ $X2=10.55 $Y2=1.16
r481 195 222 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=10.14 $Y=1.16
+ $X2=10.13 $Y2=1.16
r482 194 195 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=10.14
+ $Y=1.16 $X2=10.14 $Y2=1.16
r483 192 209 68.8738 $w=2.7e-07 $l=3.1e-07 $layer=POLY_cond $X=4.36 $Y=1.16
+ $X2=4.67 $Y2=1.16
r484 192 206 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=4.36 $Y=1.16
+ $X2=4.25 $Y2=1.16
r485 191 194 320.527 $w=1.98e-07 $l=5.78e-06 $layer=LI1_cond $X=4.36 $Y=1.175
+ $X2=10.14 $Y2=1.175
r486 191 192 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=4.36
+ $Y=1.16 $X2=4.36 $Y2=1.16
r487 189 205 0.866423 $w=2e-07 $l=8.8e-08 $layer=LI1_cond $X=4.125 $Y=1.175
+ $X2=4.037 $Y2=1.175
r488 189 191 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=4.125 $Y=1.175
+ $X2=4.36 $Y2=1.175
r489 188 203 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.037 $Y=1.445
+ $X2=4.037 $Y2=1.53
r490 187 205 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=4.037 $Y=1.275
+ $X2=4.037 $Y2=1.175
r491 187 188 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=4.037 $Y=1.275
+ $X2=4.037 $Y2=1.445
r492 186 205 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=4.037 $Y=1.075
+ $X2=4.037 $Y2=1.175
r493 185 200 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.037 $Y=0.905
+ $X2=4.037 $Y2=0.82
r494 185 186 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=4.037 $Y=0.905
+ $X2=4.037 $Y2=1.075
r495 181 183 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.62 $Y=1.63
+ $X2=3.62 $Y2=2.31
r496 179 203 27.2053 $w=1.68e-07 $l=4.17e-07 $layer=LI1_cond $X=3.62 $Y=1.53
+ $X2=4.037 $Y2=1.53
r497 179 181 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.62 $Y=1.615
+ $X2=3.62 $Y2=1.63
r498 175 200 27.2053 $w=1.68e-07 $l=4.17e-07 $layer=LI1_cond $X=3.62 $Y=0.82
+ $X2=4.037 $Y2=0.82
r499 175 177 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.4
r500 174 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=1.53
+ $X2=2.78 $Y2=1.53
r501 173 179 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=1.53
+ $X2=3.62 $Y2=1.53
r502 173 174 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.455 $Y=1.53
+ $X2=2.945 $Y2=1.53
r503 172 197 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0.82
+ $X2=2.78 $Y2=0.82
r504 171 175 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0.82
+ $X2=3.62 $Y2=0.82
r505 171 172 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.455 $Y=0.82
+ $X2=2.945 $Y2=0.82
r506 167 169 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.78 $Y=1.63
+ $X2=2.78 $Y2=2.31
r507 165 198 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=1.615
+ $X2=2.78 $Y2=1.53
r508 165 167 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.78 $Y=1.615
+ $X2=2.78 $Y2=1.63
r509 161 197 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.82
r510 161 163 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.78 $Y=0.735
+ $X2=2.78 $Y2=0.4
r511 159 198 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=1.53
+ $X2=2.78 $Y2=1.53
r512 159 160 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.615 $Y=1.53
+ $X2=2.105 $Y2=1.53
r513 157 197 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0.82
+ $X2=2.78 $Y2=0.82
r514 157 158 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.615 $Y=0.82
+ $X2=2.105 $Y2=0.82
r515 153 155 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.94 $Y=1.63
+ $X2=1.94 $Y2=2.31
r516 151 160 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=2.105 $Y2=1.53
r517 151 153 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.94 $Y=1.615
+ $X2=1.94 $Y2=1.63
r518 147 158 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=2.105 $Y2=0.82
r519 147 149 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.4
r520 143 224 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.55 $Y=1.295
+ $X2=10.55 $Y2=1.16
r521 143 145 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.55 $Y=1.295
+ $X2=10.55 $Y2=1.985
r522 139 224 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.55 $Y=1.025
+ $X2=10.55 $Y2=1.16
r523 139 141 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.55 $Y=1.025
+ $X2=10.55 $Y2=0.56
r524 135 222 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.13 $Y=1.295
+ $X2=10.13 $Y2=1.16
r525 135 137 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.13 $Y=1.295
+ $X2=10.13 $Y2=1.985
r526 131 222 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.13 $Y=1.025
+ $X2=10.13 $Y2=1.16
r527 131 133 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.13 $Y=1.025
+ $X2=10.13 $Y2=0.56
r528 127 221 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.71 $Y=1.295
+ $X2=9.71 $Y2=1.16
r529 127 129 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.71 $Y=1.295
+ $X2=9.71 $Y2=1.985
r530 123 221 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.71 $Y=1.025
+ $X2=9.71 $Y2=1.16
r531 123 125 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.71 $Y=1.025
+ $X2=9.71 $Y2=0.56
r532 119 220 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.29 $Y=1.295
+ $X2=9.29 $Y2=1.16
r533 119 121 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.29 $Y=1.295
+ $X2=9.29 $Y2=1.985
r534 115 220 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.29 $Y=1.025
+ $X2=9.29 $Y2=1.16
r535 115 117 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.29 $Y=1.025
+ $X2=9.29 $Y2=0.56
r536 111 219 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.87 $Y=1.295
+ $X2=8.87 $Y2=1.16
r537 111 113 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.87 $Y=1.295
+ $X2=8.87 $Y2=1.985
r538 107 219 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.87 $Y=1.025
+ $X2=8.87 $Y2=1.16
r539 107 109 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.87 $Y=1.025
+ $X2=8.87 $Y2=0.56
r540 103 218 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.45 $Y=1.295
+ $X2=8.45 $Y2=1.16
r541 103 105 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.45 $Y=1.295
+ $X2=8.45 $Y2=1.985
r542 99 218 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.45 $Y=1.025
+ $X2=8.45 $Y2=1.16
r543 99 101 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.45 $Y=1.025
+ $X2=8.45 $Y2=0.56
r544 95 217 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.03 $Y=1.295
+ $X2=8.03 $Y2=1.16
r545 95 97 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.03 $Y=1.295
+ $X2=8.03 $Y2=1.985
r546 91 217 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.03 $Y=1.025
+ $X2=8.03 $Y2=1.16
r547 91 93 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.03 $Y=1.025
+ $X2=8.03 $Y2=0.56
r548 87 216 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.61 $Y=1.295
+ $X2=7.61 $Y2=1.16
r549 87 89 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.61 $Y=1.295
+ $X2=7.61 $Y2=1.985
r550 83 216 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.61 $Y=1.025
+ $X2=7.61 $Y2=1.16
r551 83 85 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.61 $Y=1.025
+ $X2=7.61 $Y2=0.56
r552 79 215 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.19 $Y=1.295
+ $X2=7.19 $Y2=1.16
r553 79 81 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.19 $Y=1.295
+ $X2=7.19 $Y2=1.985
r554 75 215 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.19 $Y=1.025
+ $X2=7.19 $Y2=1.16
r555 75 77 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.19 $Y=1.025
+ $X2=7.19 $Y2=0.56
r556 71 214 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.16
r557 71 73 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.985
r558 67 214 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=1.16
r559 67 69 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=0.56
r560 63 213 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.16
r561 63 65 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.985
r562 59 213 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=1.16
r563 59 61 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=0.56
r564 55 212 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.16
r565 55 57 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.985
r566 51 212 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=1.16
r567 51 53 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=0.56
r568 47 211 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.16
r569 47 49 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.985
r570 43 211 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=1.16
r571 43 45 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=0.56
r572 39 210 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.16
r573 39 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.985
r574 35 210 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=1.16
r575 35 37 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=0.56
r576 31 209 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.16
r577 31 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.985
r578 27 209 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=1.16
r579 27 29 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=0.56
r580 23 206 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.16
r581 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.985
r582 19 206 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=1.16
r583 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=0.56
r584 6 183 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2.31
r585 6 181 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.63
r586 5 169 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2.31
r587 5 167 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.63
r588 4 155 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.31
r589 4 153 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.63
r590 3 177 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.4
r591 2 163 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.4
r592 1 149 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 42 46
+ 50 54 58 60 64 68 72 76 80 84 86 90 92 94 97 98 100 101 103 104 106 107 108
+ 109 111 112 114 115 117 118 120 121 122 123 124 158 164 167 171
r181 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r182 167 168 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r183 164 165 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r184 162 171 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r185 162 168 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.89 $Y2=2.72
r186 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r187 159 167 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.005 $Y=2.72
+ $X2=9.92 $Y2=2.72
r188 159 161 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.005 $Y=2.72
+ $X2=10.35 $Y2=2.72
r189 158 170 3.40825 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=2.72
+ $X2=10.857 $Y2=2.72
r190 158 161 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.675 $Y=2.72
+ $X2=10.35 $Y2=2.72
r191 157 168 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r192 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r193 154 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r194 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r195 151 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r196 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r197 148 151 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r198 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r199 145 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r200 145 165 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r201 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r202 142 164 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=4.88 $Y2=2.72
r203 142 144 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=5.29 $Y2=2.72
r204 141 165 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r205 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r206 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r207 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r208 135 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r209 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r210 132 135 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r211 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r212 124 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r213 124 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r214 122 156 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=8.995 $Y=2.72
+ $X2=8.97 $Y2=2.72
r215 122 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.995 $Y=2.72
+ $X2=9.08 $Y2=2.72
r216 120 153 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.155 $Y=2.72
+ $X2=8.05 $Y2=2.72
r217 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.155 $Y=2.72
+ $X2=8.24 $Y2=2.72
r218 119 156 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=8.325 $Y=2.72
+ $X2=8.97 $Y2=2.72
r219 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.325 $Y=2.72
+ $X2=8.24 $Y2=2.72
r220 117 150 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.315 $Y=2.72
+ $X2=7.13 $Y2=2.72
r221 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.315 $Y=2.72
+ $X2=7.4 $Y2=2.72
r222 116 153 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=8.05 $Y2=2.72
r223 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=7.4 $Y2=2.72
r224 114 147 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.475 $Y=2.72
+ $X2=6.21 $Y2=2.72
r225 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=2.72
+ $X2=6.56 $Y2=2.72
r226 113 150 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.645 $Y=2.72
+ $X2=7.13 $Y2=2.72
r227 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=2.72
+ $X2=6.56 $Y2=2.72
r228 111 144 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.29 $Y2=2.72
r229 111 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=2.72
+ $X2=5.72 $Y2=2.72
r230 110 147 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.805 $Y=2.72
+ $X2=6.21 $Y2=2.72
r231 110 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=2.72
+ $X2=5.72 $Y2=2.72
r232 108 140 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=3.91 $Y2=2.72
r233 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=4.04 $Y2=2.72
r234 106 137 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=2.72
+ $X2=2.99 $Y2=2.72
r235 106 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.72
+ $X2=3.2 $Y2=2.72
r236 105 140 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=3.91 $Y2=2.72
r237 105 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=3.2 $Y2=2.72
r238 103 134 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.07 $Y2=2.72
r239 103 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.36 $Y2=2.72
r240 102 137 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.445 $Y=2.72
+ $X2=2.99 $Y2=2.72
r241 102 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=2.72
+ $X2=2.36 $Y2=2.72
r242 100 131 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r243 100 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.52 $Y2=2.72
r244 99 134 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=2.07 $Y2=2.72
r245 99 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.52 $Y2=2.72
r246 97 127 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r247 97 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.68 $Y2=2.72
r248 96 131 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=1.15 $Y2=2.72
r249 96 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.68 $Y2=2.72
r250 92 170 3.40825 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=10.76 $Y=2.635
+ $X2=10.857 $Y2=2.72
r251 92 94 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.76 $Y=2.635
+ $X2=10.76 $Y2=2
r252 88 167 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.92 $Y=2.635
+ $X2=9.92 $Y2=2.72
r253 88 90 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.92 $Y=2.635
+ $X2=9.92 $Y2=2
r254 87 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.165 $Y=2.72
+ $X2=9.08 $Y2=2.72
r255 86 167 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.835 $Y=2.72
+ $X2=9.92 $Y2=2.72
r256 86 87 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.835 $Y=2.72
+ $X2=9.165 $Y2=2.72
r257 82 123 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.08 $Y=2.635
+ $X2=9.08 $Y2=2.72
r258 82 84 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.08 $Y=2.635
+ $X2=9.08 $Y2=2
r259 78 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=2.635
+ $X2=8.24 $Y2=2.72
r260 78 80 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.24 $Y=2.635
+ $X2=8.24 $Y2=2
r261 74 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=2.635
+ $X2=7.4 $Y2=2.72
r262 74 76 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.4 $Y=2.635
+ $X2=7.4 $Y2=2
r263 70 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=2.635
+ $X2=6.56 $Y2=2.72
r264 70 72 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.56 $Y=2.635
+ $X2=6.56 $Y2=2
r265 66 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=2.635
+ $X2=5.72 $Y2=2.72
r266 66 68 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.72 $Y=2.635
+ $X2=5.72 $Y2=2
r267 62 164 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2.72
r268 62 64 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.88 $Y=2.635
+ $X2=4.88 $Y2=2
r269 61 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=2.72
+ $X2=4.04 $Y2=2.72
r270 60 164 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.88 $Y2=2.72
r271 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.125 $Y2=2.72
r272 56 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.635
+ $X2=4.04 $Y2=2.72
r273 56 58 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.04 $Y=2.635
+ $X2=4.04 $Y2=2
r274 52 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2.72
r275 52 54 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2
r276 48 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r277 48 50 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2
r278 44 101 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r279 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2
r280 40 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r281 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2
r282 13 94 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=10.625
+ $Y=1.485 $X2=10.76 $Y2=2
r283 12 90 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.785
+ $Y=1.485 $X2=9.92 $Y2=2
r284 11 84 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.945
+ $Y=1.485 $X2=9.08 $Y2=2
r285 10 80 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.105
+ $Y=1.485 $X2=8.24 $Y2=2
r286 9 76 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.265
+ $Y=1.485 $X2=7.4 $Y2=2
r287 8 72 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.425
+ $Y=1.485 $X2=6.56 $Y2=2
r288 7 68 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=2
r289 6 64 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=2
r290 5 58 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=2
r291 4 54 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2
r292 3 50 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2
r293 2 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2
r294 1 42 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 49 50 53 57 58 59 60 61 62 65 69 71 73 74 77 81 83 87 91 95 97 101 105 109 111
+ 115 119 123 125 129 133 137 139 143 147 151 153 159 160 163 164 165 166 167
+ 168 169 170 171 172 173 174 176 177
c337 60 0 1.25206e-19 $X=4.625 $Y=1.53
c338 58 0 1.25206e-19 $X=4.625 $Y=0.82
r339 176 177 8.27522 $w=4.43e-07 $l=2.55e-07 $layer=LI1_cond $X=10.817 $Y=1.19
+ $X2=10.817 $Y2=1.445
r340 175 176 11.9435 $w=2.73e-07 $l=2.85e-07 $layer=LI1_cond $X=10.817 $Y=0.905
+ $X2=10.817 $Y2=1.19
r341 154 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.505 $Y=1.53
+ $X2=10.34 $Y2=1.53
r342 153 177 4.51856 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=10.68 $Y=1.53
+ $X2=10.817 $Y2=1.53
r343 153 154 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.68 $Y=1.53
+ $X2=10.505 $Y2=1.53
r344 152 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.505 $Y=0.82
+ $X2=10.34 $Y2=0.82
r345 151 175 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=10.68 $Y=0.82
+ $X2=10.817 $Y2=0.905
r346 151 152 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.68 $Y=0.82
+ $X2=10.505 $Y2=0.82
r347 147 149 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.34 $Y=1.63
+ $X2=10.34 $Y2=2.31
r348 145 174 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.34 $Y=1.615
+ $X2=10.34 $Y2=1.53
r349 145 147 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=10.34 $Y=1.615
+ $X2=10.34 $Y2=1.63
r350 141 173 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.34 $Y=0.735
+ $X2=10.34 $Y2=0.82
r351 141 143 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.34 $Y=0.735
+ $X2=10.34 $Y2=0.4
r352 140 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=1.53
+ $X2=9.5 $Y2=1.53
r353 139 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.175 $Y=1.53
+ $X2=10.34 $Y2=1.53
r354 139 140 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.175 $Y=1.53
+ $X2=9.665 $Y2=1.53
r355 138 171 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=0.82
+ $X2=9.5 $Y2=0.82
r356 137 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.175 $Y=0.82
+ $X2=10.34 $Y2=0.82
r357 137 138 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.175 $Y=0.82
+ $X2=9.665 $Y2=0.82
r358 133 135 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.5 $Y=1.63
+ $X2=9.5 $Y2=2.31
r359 131 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.5 $Y=1.615
+ $X2=9.5 $Y2=1.53
r360 131 133 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=9.5 $Y=1.615
+ $X2=9.5 $Y2=1.63
r361 127 171 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.5 $Y=0.735
+ $X2=9.5 $Y2=0.82
r362 127 129 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.5 $Y=0.735
+ $X2=9.5 $Y2=0.4
r363 126 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.825 $Y=1.53
+ $X2=8.66 $Y2=1.53
r364 125 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.335 $Y=1.53
+ $X2=9.5 $Y2=1.53
r365 125 126 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.335 $Y=1.53
+ $X2=8.825 $Y2=1.53
r366 124 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.825 $Y=0.82
+ $X2=8.66 $Y2=0.82
r367 123 171 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.335 $Y=0.82
+ $X2=9.5 $Y2=0.82
r368 123 124 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.335 $Y=0.82
+ $X2=8.825 $Y2=0.82
r369 119 121 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.66 $Y=1.63
+ $X2=8.66 $Y2=2.31
r370 117 170 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.66 $Y=1.615
+ $X2=8.66 $Y2=1.53
r371 117 119 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.66 $Y=1.615
+ $X2=8.66 $Y2=1.63
r372 113 169 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.66 $Y=0.735
+ $X2=8.66 $Y2=0.82
r373 113 115 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.66 $Y=0.735
+ $X2=8.66 $Y2=0.4
r374 112 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.985 $Y=1.53
+ $X2=7.82 $Y2=1.53
r375 111 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.495 $Y=1.53
+ $X2=8.66 $Y2=1.53
r376 111 112 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=1.53
+ $X2=7.985 $Y2=1.53
r377 110 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.985 $Y=0.82
+ $X2=7.82 $Y2=0.82
r378 109 169 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.495 $Y=0.82
+ $X2=8.66 $Y2=0.82
r379 109 110 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.495 $Y=0.82
+ $X2=7.985 $Y2=0.82
r380 105 107 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.82 $Y=1.63
+ $X2=7.82 $Y2=2.31
r381 103 168 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.82 $Y=1.615
+ $X2=7.82 $Y2=1.53
r382 103 105 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.82 $Y=1.615
+ $X2=7.82 $Y2=1.63
r383 99 167 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.82 $Y=0.735
+ $X2=7.82 $Y2=0.82
r384 99 101 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.82 $Y=0.735
+ $X2=7.82 $Y2=0.4
r385 98 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=1.53
+ $X2=6.98 $Y2=1.53
r386 97 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=1.53
+ $X2=7.82 $Y2=1.53
r387 97 98 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.655 $Y=1.53
+ $X2=7.145 $Y2=1.53
r388 96 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=0.82
+ $X2=6.98 $Y2=0.82
r389 95 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=0.82
+ $X2=7.82 $Y2=0.82
r390 95 96 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.655 $Y=0.82
+ $X2=7.145 $Y2=0.82
r391 91 93 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.98 $Y=1.63
+ $X2=6.98 $Y2=2.31
r392 89 166 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=1.615
+ $X2=6.98 $Y2=1.53
r393 89 91 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.98 $Y=1.615
+ $X2=6.98 $Y2=1.63
r394 85 165 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=0.735
+ $X2=6.98 $Y2=0.82
r395 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.98 $Y=0.735
+ $X2=6.98 $Y2=0.4
r396 84 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=1.53
+ $X2=6.14 $Y2=1.53
r397 83 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.815 $Y=1.53
+ $X2=6.98 $Y2=1.53
r398 83 84 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.815 $Y=1.53
+ $X2=6.305 $Y2=1.53
r399 82 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0.82
+ $X2=6.14 $Y2=0.82
r400 81 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.815 $Y=0.82
+ $X2=6.98 $Y2=0.82
r401 81 82 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.815 $Y=0.82
+ $X2=6.305 $Y2=0.82
r402 77 79 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.14 $Y=1.63
+ $X2=6.14 $Y2=2.31
r403 75 164 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=1.615
+ $X2=6.14 $Y2=1.53
r404 75 77 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.14 $Y=1.615
+ $X2=6.14 $Y2=1.63
r405 74 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=0.735
+ $X2=6.14 $Y2=0.82
r406 73 162 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=6.14 $Y=0.425
+ $X2=6.14 $Y2=0.4
r407 73 74 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.14 $Y=0.425
+ $X2=6.14 $Y2=0.735
r408 72 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=1.53
+ $X2=5.3 $Y2=1.53
r409 71 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=1.53
+ $X2=6.14 $Y2=1.53
r410 71 72 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.975 $Y=1.53
+ $X2=5.465 $Y2=1.53
r411 70 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=0.82
+ $X2=5.3 $Y2=0.82
r412 69 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=0.82
+ $X2=6.14 $Y2=0.82
r413 69 70 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.975 $Y=0.82
+ $X2=5.465 $Y2=0.82
r414 65 67 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.3 $Y=1.63 $X2=5.3
+ $Y2=2.31
r415 63 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=1.615
+ $X2=5.3 $Y2=1.53
r416 63 65 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.3 $Y=1.615
+ $X2=5.3 $Y2=1.63
r417 62 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=0.735
+ $X2=5.3 $Y2=0.82
r418 61 158 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=5.3 $Y=0.425
+ $X2=5.3 $Y2=0.4
r419 61 62 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=5.3 $Y=0.425 $X2=5.3
+ $Y2=0.735
r420 59 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=1.53
+ $X2=5.3 $Y2=1.53
r421 59 60 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.135 $Y=1.53
+ $X2=4.625 $Y2=1.53
r422 57 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=0.82
+ $X2=5.3 $Y2=0.82
r423 57 58 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.135 $Y=0.82
+ $X2=4.625 $Y2=0.82
r424 53 55 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.46 $Y=1.63
+ $X2=4.46 $Y2=2.31
r425 51 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.46 $Y=1.615
+ $X2=4.625 $Y2=1.53
r426 51 53 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.46 $Y=1.615
+ $X2=4.46 $Y2=1.63
r427 50 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.46 $Y=0.735
+ $X2=4.625 $Y2=0.82
r428 49 156 0.924242 $w=3.3e-07 $l=2.5e-08 $layer=LI1_cond $X=4.46 $Y=0.425
+ $X2=4.46 $Y2=0.4
r429 49 50 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=4.46 $Y=0.425
+ $X2=4.46 $Y2=0.735
r430 16 149 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=10.205
+ $Y=1.485 $X2=10.34 $Y2=2.31
r431 16 147 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.205
+ $Y=1.485 $X2=10.34 $Y2=1.63
r432 15 135 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=9.365
+ $Y=1.485 $X2=9.5 $Y2=2.31
r433 15 133 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.365
+ $Y=1.485 $X2=9.5 $Y2=1.63
r434 14 121 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=1.485 $X2=8.66 $Y2=2.31
r435 14 119 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=1.485 $X2=8.66 $Y2=1.63
r436 13 107 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.485 $X2=7.82 $Y2=2.31
r437 13 105 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.485 $X2=7.82 $Y2=1.63
r438 12 93 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=6.98 $Y2=2.31
r439 12 91 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=6.98 $Y2=1.63
r440 11 79 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=6.005
+ $Y=1.485 $X2=6.14 $Y2=2.31
r441 11 77 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.005
+ $Y=1.485 $X2=6.14 $Y2=1.63
r442 10 67 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=2.31
r443 10 65 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=1.63
r444 9 55 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=2.31
r445 9 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=1.63
r446 8 143 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=10.205
+ $Y=0.235 $X2=10.34 $Y2=0.4
r447 7 129 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=9.365
+ $Y=0.235 $X2=9.5 $Y2=0.4
r448 6 115 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.525
+ $Y=0.235 $X2=8.66 $Y2=0.4
r449 5 101 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=7.685
+ $Y=0.235 $X2=7.82 $Y2=0.4
r450 4 87 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.235 $X2=6.98 $Y2=0.4
r451 3 162 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=6.005
+ $Y=0.235 $X2=6.14 $Y2=0.4
r452 2 158 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.165
+ $Y=0.235 $X2=5.3 $Y2=0.4
r453 1 156 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 42 46
+ 50 54 58 60 64 68 72 76 80 84 86 90 92 94 97 98 100 101 103 104 106 107 108
+ 109 111 112 114 115 117 118 120 121 122 123 124 158 164 167 171
r215 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r216 167 168 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r217 164 165 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r218 162 171 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r219 162 168 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=9.89 $Y2=0
r220 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r221 159 167 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.005 $Y=0
+ $X2=9.92 $Y2=0
r222 159 161 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.005 $Y=0
+ $X2=10.35 $Y2=0
r223 158 170 3.40825 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.857 $Y2=0
r224 158 161 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.35 $Y2=0
r225 157 168 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r226 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r227 154 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r228 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r229 151 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r230 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r231 148 151 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r232 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r233 145 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r234 145 165 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r235 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r236 142 164 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=0
+ $X2=4.88 $Y2=0
r237 142 144 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.965 $Y=0
+ $X2=5.29 $Y2=0
r238 141 165 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r239 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r240 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r241 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r242 135 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r243 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r244 132 135 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r245 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r246 124 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r247 124 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r248 122 156 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=8.995 $Y=0
+ $X2=8.97 $Y2=0
r249 122 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.995 $Y=0
+ $X2=9.08 $Y2=0
r250 120 153 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.155 $Y=0
+ $X2=8.05 $Y2=0
r251 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.155 $Y=0
+ $X2=8.24 $Y2=0
r252 119 156 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.97 $Y2=0
r253 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.24 $Y2=0
r254 117 150 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=7.13 $Y2=0
r255 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.315 $Y=0 $X2=7.4
+ $Y2=0
r256 116 153 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=7.485 $Y=0
+ $X2=8.05 $Y2=0
r257 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=0 $X2=7.4
+ $Y2=0
r258 114 147 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.475 $Y=0
+ $X2=6.21 $Y2=0
r259 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=0
+ $X2=6.56 $Y2=0
r260 113 150 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.645 $Y=0
+ $X2=7.13 $Y2=0
r261 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=0
+ $X2=6.56 $Y2=0
r262 111 144 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.635 $Y=0
+ $X2=5.29 $Y2=0
r263 111 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=0
+ $X2=5.72 $Y2=0
r264 110 147 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.805 $Y=0
+ $X2=6.21 $Y2=0
r265 110 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=0
+ $X2=5.72 $Y2=0
r266 108 140 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=3.91 $Y2=0
r267 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=4.04 $Y2=0
r268 106 137 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=0
+ $X2=2.99 $Y2=0
r269 106 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.2
+ $Y2=0
r270 105 140 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.285 $Y=0
+ $X2=3.91 $Y2=0
r271 105 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.2
+ $Y2=0
r272 103 134 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.275 $Y=0
+ $X2=2.07 $Y2=0
r273 103 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0
+ $X2=2.36 $Y2=0
r274 102 137 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.99 $Y2=0
r275 102 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.36 $Y2=0
r276 100 131 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0
+ $X2=1.15 $Y2=0
r277 100 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0
+ $X2=1.52 $Y2=0
r278 99 134 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=2.07 $Y2=0
r279 99 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.52
+ $Y2=0
r280 97 127 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r281 97 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r282 96 131 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=1.15 $Y2=0
r283 96 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r284 92 170 3.40825 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.857 $Y2=0
r285 92 94 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.76 $Y2=0.4
r286 88 167 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.92 $Y=0.085
+ $X2=9.92 $Y2=0
r287 88 90 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.92 $Y=0.085
+ $X2=9.92 $Y2=0.4
r288 87 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.165 $Y=0 $X2=9.08
+ $Y2=0
r289 86 167 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.835 $Y=0 $X2=9.92
+ $Y2=0
r290 86 87 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.835 $Y=0
+ $X2=9.165 $Y2=0
r291 82 123 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.08 $Y=0.085
+ $X2=9.08 $Y2=0
r292 82 84 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.08 $Y=0.085
+ $X2=9.08 $Y2=0.4
r293 78 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=0.085
+ $X2=8.24 $Y2=0
r294 78 80 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.24 $Y=0.085
+ $X2=8.24 $Y2=0.4
r295 74 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0.085
+ $X2=7.4 $Y2=0
r296 74 76 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.4 $Y=0.085
+ $X2=7.4 $Y2=0.4
r297 70 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=0.085
+ $X2=6.56 $Y2=0
r298 70 72 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.56 $Y=0.085
+ $X2=6.56 $Y2=0.4
r299 66 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=0.085
+ $X2=5.72 $Y2=0
r300 66 68 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.72 $Y=0.085
+ $X2=5.72 $Y2=0.4
r301 62 164 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r302 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.4
r303 61 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.04
+ $Y2=0
r304 60 164 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.88
+ $Y2=0
r305 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=4.125 $Y2=0
r306 56 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r307 56 58 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.4
r308 52 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.085
+ $X2=3.2 $Y2=0
r309 52 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.2 $Y=0.085
+ $X2=3.2 $Y2=0.4
r310 48 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0
r311 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.36 $Y=0.085
+ $X2=2.36 $Y2=0.4
r312 44 101 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r313 44 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.4
r314 40 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r315 40 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r316 13 94 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=10.625
+ $Y=0.235 $X2=10.76 $Y2=0.4
r317 12 90 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=9.785
+ $Y=0.235 $X2=9.92 $Y2=0.4
r318 11 84 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.945
+ $Y=0.235 $X2=9.08 $Y2=0.4
r319 10 80 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.105
+ $Y=0.235 $X2=8.24 $Y2=0.4
r320 9 76 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.265
+ $Y=0.235 $X2=7.4 $Y2=0.4
r321 8 72 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.425
+ $Y=0.235 $X2=6.56 $Y2=0.4
r322 7 68 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.4
r323 6 64 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.4
r324 5 58 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.4
r325 4 54 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.4
r326 3 50 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.4
r327 2 46 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r328 1 42 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends


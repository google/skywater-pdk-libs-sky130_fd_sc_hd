* File: sky130_fd_sc_hd__a311o_1.spice.pex
* Created: Thu Aug 27 14:03:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A311O_1%A_75_199# 1 2 3 12 15 20 21 22 23 24 26 27
+ 28 29 30 31 32 35 39 42 43 44 49
c110 43 0 1.87367e-19 $X=0.51 $Y=1.16
c111 42 0 1.12853e-19 $X=0.51 $Y=1.16
c112 20 0 1.0136e-19 $X=0.65 $Y=1.495
r113 43 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r114 43 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r115 42 45 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=1.16
+ $X2=0.58 $Y2=1.325
r116 42 44 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=1.16
+ $X2=0.58 $Y2=0.995
r117 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r118 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.42 $Y=1.665
+ $X2=3.42 $Y2=1.96
r119 33 35 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.42 $Y=0.655
+ $X2=3.42 $Y2=0.42
r120 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.74
+ $X2=3.42 $Y2=0.655
r121 31 32 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.335 $Y=0.74
+ $X2=2.495 $Y2=0.74
r122 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=0.655
+ $X2=2.495 $Y2=0.74
r123 29 47 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.425
+ $X2=2.41 $Y2=0.34
r124 29 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=0.425
+ $X2=2.41 $Y2=0.655
r125 27 47 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=0.34
+ $X2=2.41 $Y2=0.34
r126 27 28 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=2.325 $Y=0.34
+ $X2=1.26 $Y2=0.34
r127 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.26 $Y2=0.34
r128 25 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.175 $Y2=0.655
r129 23 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=1.58
+ $X2=3.42 $Y2=1.665
r130 23 24 169.626 $w=1.68e-07 $l=2.6e-06 $layer=LI1_cond $X=3.335 $Y=1.58
+ $X2=0.735 $Y2=1.58
r131 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=0.74
+ $X2=1.175 $Y2=0.655
r132 21 22 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.09 $Y=0.74
+ $X2=0.735 $Y2=0.74
r133 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.65 $Y=1.495
+ $X2=0.735 $Y2=1.58
r134 20 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=1.495
+ $X2=0.65 $Y2=1.325
r135 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.65 $Y=0.825
+ $X2=0.735 $Y2=0.74
r136 17 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=0.825
+ $X2=0.65 $Y2=0.995
r137 15 50 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.985
+ $X2=0.495 $Y2=1.325
r138 12 49 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
r139 3 39 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.96
r140 2 35 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.42
r141 1 47 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.41 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%A3 3 7 8 11 13
r35 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.16
+ $X2=0.99 $Y2=1.325
r36 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.16
+ $X2=0.99 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=1.16 $X2=0.99 $Y2=1.16
r38 8 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=0.99
+ $Y2=1.16
r39 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.965 $Y=0.56
+ $X2=0.965 $Y2=0.995
r40 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.93 $Y=1.985
+ $X2=0.93 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%A2 3 5 7 8 9 16
r39 14 16 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.5 $Y=1.16 $X2=1.62
+ $Y2=1.16
r40 12 14 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.41 $Y=1.16 $X2=1.5
+ $Y2=1.16
r41 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.16 $X2=1.62 $Y2=1.16
r42 8 9 17.6317 $w=1.93e-07 $l=3.1e-07 $layer=LI1_cond $X=1.607 $Y=0.85
+ $X2=1.607 $Y2=1.16
r43 5 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=0.995 $X2=1.5
+ $Y2=1.16
r44 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.5 $Y=0.995 $X2=1.5
+ $Y2=0.56
r45 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r46 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325 $X2=1.41
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%A1 3 6 8 9 13 15
r38 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.225 $Y2=1.325
r39 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.225 $Y2=0.995
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=1.16 $X2=2.225 $Y2=1.16
r41 9 14 1.30249 $w=2.81e-07 $l=3e-08 $layer=LI1_cond $X=2.137 $Y=1.19 $X2=2.137
+ $Y2=1.16
r42 8 14 13.4591 $w=2.81e-07 $l=3.1e-07 $layer=LI1_cond $X=2.137 $Y=0.85
+ $X2=2.137 $Y2=1.16
r43 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.985
+ $X2=2.17 $Y2=1.325
r44 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.56 $X2=2.17
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%B1 3 6 8 11 13
r34 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.16
+ $X2=2.705 $Y2=1.325
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.16
+ $X2=2.705 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.16 $X2=2.705 $Y2=1.16
r37 8 12 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.99 $Y=1.16
+ $X2=2.705 $Y2=1.16
r38 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.645 $Y=1.985
+ $X2=2.645 $Y2=1.325
r39 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.645 $Y=0.56
+ $X2=2.645 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%C1 1 3 6 8 13
r25 10 13 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.21 $Y=1.16
+ $X2=3.435 $Y2=1.16
r26 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.435
+ $Y=1.16 $X2=3.435 $Y2=1.16
r27 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.325
+ $X2=3.21 $Y2=1.16
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.325 $X2=3.21
+ $Y2=1.985
r29 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.995 $X2=3.21
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%X 1 2 9 12 13 20
r19 13 20 7.11803 $w=3.38e-07 $l=2.1e-07 $layer=LI1_cond $X=0.255 $Y=2.21
+ $X2=0.255 $Y2=2
r20 12 20 2.38745 $w=5.08e-07 $l=4.5e-08 $layer=LI1_cond $X=0.255 $Y=1.955
+ $X2=0.255 $Y2=2
r21 11 12 47.9353 $w=2.73e-07 $l=1.115e-06 $layer=LI1_cond $X=0.17 $Y=0.67
+ $X2=0.17 $Y2=1.785
r22 9 11 11.6272 $w=3.08e-07 $l=2.5e-07 $layer=LI1_cond $X=0.24 $Y=0.42 $X2=0.24
+ $Y2=0.67
r23 2 20 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
r24 1 9 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%VPWR 1 2 9 11 13 25 26 29 34 40
c51 1 0 1.0136e-19 $X=0.57 $Y=1.485
r52 38 40 7.43982 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=2.07 $Y=2.53
+ $X2=2.125 $Y2=2.53
r53 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 36 38 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.96 $Y=2.53
+ $X2=2.07 $Y2=2.53
r55 33 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 32 36 7.61141 $w=5.48e-07 $l=3.5e-07 $layer=LI1_cond $X=1.61 $Y=2.53
+ $X2=1.96 $Y2=2.53
r57 32 34 9.61451 $w=5.48e-07 $l=1.55e-07 $layer=LI1_cond $X=1.61 $Y=2.53
+ $X2=1.455 $Y2=2.53
r58 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 26 39 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 25 40 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=2.125 $Y2=2.72
r62 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r63 22 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 22 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 21 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=1.455 $Y2=2.72
r66 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 19 29 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.84 $Y=2.72
+ $X2=0.717 $Y2=2.72
r68 19 21 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.84 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 13 29 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.717 $Y2=2.72
r70 13 15 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 11 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 7 29 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.717 $Y=2.635
+ $X2=0.717 $Y2=2.72
r74 7 9 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.717 $Y=2.635
+ $X2=0.717 $Y2=2.34
r75 2 36 300 $w=1.7e-07 $l=1.06637e-06 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.485 $X2=1.96 $Y2=2.34
r76 1 9 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.485 $X2=0.705 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%A_201_297# 1 2 7 9 11 13 15
r24 13 20 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=2.005
+ $X2=2.45 $Y2=1.92
r25 13 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.45 $Y=2.005
+ $X2=2.45 $Y2=2.3
r26 12 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=1.92
+ $X2=1.14 $Y2=1.92
r27 11 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=1.92
+ $X2=2.45 $Y2=1.92
r28 11 12 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=2.325 $Y=1.92
+ $X2=1.265 $Y2=1.92
r29 7 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.005 $X2=1.14
+ $Y2=1.92
r30 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=2.005
+ $X2=1.14 $Y2=2.3
r31 2 20 600 $w=1.7e-07 $l=5.10882e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.41 $Y2=1.92
r32 2 15 600 $w=1.7e-07 $l=8.937e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.41 $Y2=2.3
r33 1 18 600 $w=1.7e-07 $l=5.15121e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.485 $X2=1.18 $Y2=1.92
r34 1 9 600 $w=1.7e-07 $l=8.98248e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.485 $X2=1.18 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_1%VGND 1 2 9 13 15 17 22 32 33 36 39
c53 9 0 1.87367e-19 $X=0.755 $Y=0.38
r54 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r56 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r57 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r58 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=2.93
+ $Y2=0
r59 30 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=3.45
+ $Y2=0
r60 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r61 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r62 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r63 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r64 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r65 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r66 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=0.755
+ $Y2=0
r67 23 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=1.15
+ $Y2=0
r68 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.765 $Y=0 $X2=2.93
+ $Y2=0
r69 22 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.765 $Y=0 $X2=2.53
+ $Y2=0
r70 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.755
+ $Y2=0
r71 17 19 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.23
+ $Y2=0
r72 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r73 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r74 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=0.085
+ $X2=2.93 $Y2=0
r75 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.93 $Y=0.085
+ $X2=2.93 $Y2=0.4
r76 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r77 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.38
r78 2 13 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.235 $X2=2.93 $Y2=0.4
r79 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.755 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__maj3_1.spice
* Created: Thu Aug 27 14:27:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__maj3_1.spice.pex"
.subckt sky130_fd_sc_hd__maj3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1013 A_109_47# N_C_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g A_109_47# VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1007 A_265_47# N_A_M1007_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_27_47#_M1008_d N_B_M1008_g A_265_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 A_421_47# N_B_M1001_g N_A_27_47#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_C_M1002_g A_421_47# VNB NSHORT L=0.15 W=0.42 AD=0.115716
+ AS=0.0441 PD=0.953832 PS=0.63 NRD=30 NRS=14.28 M=1 R=2.8 SA=75002.1 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_27_47#_M1009_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.23725 AS=0.179084 PD=2.03 PS=1.47617 NRD=18.456 NRS=33.228 M=1 R=4.33333
+ SA=75001.9 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1010 A_109_341# N_C_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_109_341# VPB PHIGHVT L=0.15 W=0.42 AD=0.0567
+ AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.5 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1003 A_265_341# N_A_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_27_47#_M1004_d N_B_M1004_g A_265_341# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.3
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1011 A_421_341# N_B_M1011_g N_A_27_47#_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_C_M1012_g A_421_341# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.147414 AS=0.0441 PD=0.925775 PS=0.63 NRD=53.9386 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_27_47#_M1000_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.365 AS=0.350986 PD=2.73 PS=2.20423 NRD=19.6803 NRS=33.4703 M=1 R=6.66667
+ SA=75001.4 SB=75000.3 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_67 VPB 0 1.84181e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__maj3_1.spice.SKY130_FD_SC_HD__MAJ3_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a22oi_4.pxi.spice
* Created: Tue Sep  1 18:53:45 2020
* 
x_PM_SKY130_FD_SC_HD__A22OI_4%B2 N_B2_c_108_n N_B2_M1013_g N_B2_M1003_g
+ N_B2_c_109_n N_B2_M1016_g N_B2_M1005_g N_B2_c_110_n N_B2_M1020_g N_B2_M1021_g
+ N_B2_c_111_n N_B2_M1031_g N_B2_M1028_g B2 N_B2_c_112_n N_B2_c_113_n
+ PM_SKY130_FD_SC_HD__A22OI_4%B2
x_PM_SKY130_FD_SC_HD__A22OI_4%B1 N_B1_c_189_n N_B1_M1017_g N_B1_M1000_g
+ N_B1_c_190_n N_B1_M1022_g N_B1_M1006_g N_B1_c_191_n N_B1_M1026_g N_B1_M1024_g
+ N_B1_c_192_n N_B1_M1027_g N_B1_M1029_g B1 N_B1_c_193_n N_B1_c_194_n
+ PM_SKY130_FD_SC_HD__A22OI_4%B1
x_PM_SKY130_FD_SC_HD__A22OI_4%A1 N_A1_c_257_n N_A1_M1010_g N_A1_M1001_g
+ N_A1_c_258_n N_A1_M1014_g N_A1_M1009_g N_A1_c_259_n N_A1_M1018_g N_A1_M1012_g
+ N_A1_c_260_n N_A1_M1023_g N_A1_M1030_g A1 N_A1_c_261_n N_A1_c_262_n
+ PM_SKY130_FD_SC_HD__A22OI_4%A1
x_PM_SKY130_FD_SC_HD__A22OI_4%A2 N_A2_c_320_n N_A2_M1008_g N_A2_M1002_g
+ N_A2_c_321_n N_A2_M1011_g N_A2_M1004_g N_A2_c_322_n N_A2_M1015_g N_A2_M1007_g
+ N_A2_c_323_n N_A2_M1019_g N_A2_M1025_g A2 N_A2_c_324_n N_A2_c_325_n
+ PM_SKY130_FD_SC_HD__A22OI_4%A2
x_PM_SKY130_FD_SC_HD__A22OI_4%A_27_297# N_A_27_297#_M1003_s N_A_27_297#_M1005_s
+ N_A_27_297#_M1028_s N_A_27_297#_M1006_s N_A_27_297#_M1029_s
+ N_A_27_297#_M1009_s N_A_27_297#_M1030_s N_A_27_297#_M1004_s
+ N_A_27_297#_M1025_s N_A_27_297#_c_395_n N_A_27_297#_c_396_n
+ N_A_27_297#_c_410_n N_A_27_297#_c_458_p N_A_27_297#_c_412_n
+ N_A_27_297#_c_449_p N_A_27_297#_c_414_n N_A_27_297#_c_454_p
+ N_A_27_297#_c_416_n N_A_27_297#_c_397_n N_A_27_297#_c_480_p
+ N_A_27_297#_c_398_n N_A_27_297#_c_471_p N_A_27_297#_c_399_n
+ N_A_27_297#_c_485_p N_A_27_297#_c_400_n N_A_27_297#_c_484_p
+ N_A_27_297#_c_401_n N_A_27_297#_c_402_n N_A_27_297#_c_486_p
+ N_A_27_297#_c_481_p N_A_27_297#_c_482_p N_A_27_297#_c_483_p
+ N_A_27_297#_c_403_n N_A_27_297#_c_404_n N_A_27_297#_c_405_n
+ PM_SKY130_FD_SC_HD__A22OI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A22OI_4%Y N_Y_M1017_d N_Y_M1026_d N_Y_M1010_d N_Y_M1018_d
+ N_Y_M1003_d N_Y_M1021_d N_Y_M1000_d N_Y_M1024_d N_Y_c_512_n N_Y_c_535_n
+ N_Y_c_510_n N_Y_c_511_n N_Y_c_514_n N_Y_c_515_n N_Y_c_516_n N_Y_c_517_n
+ N_Y_c_518_n Y Y PM_SKY130_FD_SC_HD__A22OI_4%Y
x_PM_SKY130_FD_SC_HD__A22OI_4%VPWR N_VPWR_M1001_d N_VPWR_M1012_d N_VPWR_M1002_d
+ N_VPWR_M1007_d N_VPWR_c_608_n N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n
+ N_VPWR_c_612_n N_VPWR_c_613_n N_VPWR_c_614_n N_VPWR_c_615_n N_VPWR_c_616_n
+ VPWR N_VPWR_c_617_n N_VPWR_c_618_n N_VPWR_c_607_n N_VPWR_c_620_n
+ N_VPWR_c_621_n PM_SKY130_FD_SC_HD__A22OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A22OI_4%A_27_47# N_A_27_47#_M1013_d N_A_27_47#_M1016_d
+ N_A_27_47#_M1031_d N_A_27_47#_M1022_s N_A_27_47#_M1027_s N_A_27_47#_c_709_n
+ N_A_27_47#_c_710_n N_A_27_47#_c_711_n N_A_27_47#_c_724_n N_A_27_47#_c_712_n
+ N_A_27_47#_c_732_n N_A_27_47#_c_713_n N_A_27_47#_c_714_n N_A_27_47#_c_715_n
+ PM_SKY130_FD_SC_HD__A22OI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__A22OI_4%VGND N_VGND_M1013_s N_VGND_M1020_s N_VGND_M1008_d
+ N_VGND_M1015_d N_VGND_c_777_n N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n
+ N_VGND_c_781_n N_VGND_c_782_n N_VGND_c_783_n N_VGND_c_784_n N_VGND_c_785_n
+ N_VGND_c_786_n VGND N_VGND_c_787_n N_VGND_c_788_n N_VGND_c_789_n
+ N_VGND_c_790_n PM_SKY130_FD_SC_HD__A22OI_4%VGND
x_PM_SKY130_FD_SC_HD__A22OI_4%A_803_47# N_A_803_47#_M1010_s N_A_803_47#_M1014_s
+ N_A_803_47#_M1023_s N_A_803_47#_M1011_s N_A_803_47#_M1019_s
+ N_A_803_47#_c_883_n N_A_803_47#_c_895_n N_A_803_47#_c_884_n
+ N_A_803_47#_c_885_n N_A_803_47#_c_903_n N_A_803_47#_c_886_n
+ N_A_803_47#_c_887_n N_A_803_47#_c_888_n PM_SKY130_FD_SC_HD__A22OI_4%A_803_47#
cc_1 VNB N_B2_c_108_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B2_c_109_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_B2_c_110_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_B2_c_111_n 0.016004f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_B2_c_112_n 0.0177948f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_6 VNB N_B2_c_113_n 0.0691925f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_7 VNB N_B1_c_189_n 0.01577f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_B1_c_190_n 0.0159234f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_9 VNB N_B1_c_191_n 0.0159506f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_10 VNB N_B1_c_192_n 0.0219013f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_11 VNB N_B1_c_193_n 0.0770067f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=1.16
cc_12 VNB N_B1_c_194_n 0.0100559f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_13 VNB N_A1_c_257_n 0.0219013f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_A1_c_258_n 0.0159553f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_15 VNB N_A1_c_259_n 0.0159544f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_16 VNB N_A1_c_260_n 0.0162225f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_17 VNB N_A1_c_261_n 0.00333731f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=1.16
cc_18 VNB N_A1_c_262_n 0.0652416f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_19 VNB N_A2_c_320_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_A2_c_321_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_21 VNB N_A2_c_322_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_22 VNB N_A2_c_323_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_23 VNB N_A2_c_324_n 0.0236945f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=1.16
cc_24 VNB N_A2_c_325_n 0.0689339f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_25 VNB N_Y_c_510_n 0.00103672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_511_n 0.00813346f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_27 VNB N_VPWR_c_607_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_709_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_29 VNB N_A_27_47#_c_710_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_30 VNB N_A_27_47#_c_711_n 0.0104565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_712_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_32 VNB N_A_27_47#_c_713_n 0.00299845f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_33 VNB N_A_27_47#_c_714_n 0.00262034f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_34 VNB N_A_27_47#_c_715_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_35 VNB N_VGND_c_777_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_36 VNB N_VGND_c_778_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_37 VNB N_VGND_c_779_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_38 VNB N_VGND_c_780_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_39 VNB N_VGND_c_781_n 0.0172255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_782_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_41 VNB N_VGND_c_783_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_42 VNB N_VGND_c_784_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_43 VNB N_VGND_c_785_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_44 VNB N_VGND_c_786_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_45 VNB N_VGND_c_787_n 0.103644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_788_n 0.0191348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_789_n 0.377151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_790_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_803_47#_c_883_n 0.00262034f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_50 VNB N_A_803_47#_c_884_n 0.00337422f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_51 VNB N_A_803_47#_c_885_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_52 VNB N_A_803_47#_c_886_n 0.0126428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_803_47#_c_887_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_54 VNB N_A_803_47#_c_888_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=1.16
cc_55 VPB N_B2_M1003_g 0.0253871f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_56 VPB N_B2_M1005_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_57 VPB N_B2_M1021_g 0.018138f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_58 VPB N_B2_M1028_g 0.0183758f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_59 VPB N_B2_c_113_n 0.0108493f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_60 VPB N_B1_M1000_g 0.0178886f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_B1_M1006_g 0.0180858f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_B1_M1024_g 0.0181158f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_63 VPB N_B1_M1029_g 0.0251939f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_64 VPB N_B1_c_193_n 0.0156051f $X=-0.19 $Y=1.305 $X2=1.64 $Y2=1.16
cc_65 VPB N_A1_M1001_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_66 VPB N_A1_M1009_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_67 VPB N_A1_M1012_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_68 VPB N_A1_M1030_g 0.0185045f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_69 VPB N_A1_c_262_n 0.0103962f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_70 VPB N_A2_M1002_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_71 VPB N_A2_M1004_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_72 VPB N_A2_M1007_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_73 VPB N_A2_M1025_g 0.0252703f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_74 VPB N_A2_c_325_n 0.0108808f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_75 VPB N_A_27_297#_c_395_n 0.00753428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_297#_c_396_n 0.0356473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_297#_c_397_n 0.00907639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_297#_c_398_n 0.00240741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_297#_c_399_n 0.00257732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_297#_c_400_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_297#_c_401_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_297#_c_402_n 0.00365821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_297#_c_403_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_297#_c_404_n 0.00469599f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_297#_c_405_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_Y_c_512_n 0.00460272f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_87 VPB N_Y_c_510_n 0.00113183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_Y_c_514_n 0.00239046f $X=-0.19 $Y=1.305 $X2=0.992 $Y2=1.16
cc_89 VPB N_Y_c_515_n 0.00234676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_Y_c_516_n 0.00202148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_Y_c_517_n 5.28005e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_Y_c_518_n 0.00239278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB Y 0.00195997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_608_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_95 VPB N_VPWR_c_609_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_96 VPB N_VPWR_c_610_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_611_n 0.00393015f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_98 VPB N_VPWR_c_612_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_99 VPB N_VPWR_c_613_n 0.103005f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_100 VPB N_VPWR_c_614_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_615_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_102 VPB N_VPWR_c_616_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_103 VPB N_VPWR_c_617_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.992 $Y2=1.19
cc_104 VPB N_VPWR_c_618_n 0.0193807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_607_n 0.0474036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_620_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_621_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 N_B2_c_111_n N_B1_c_189_n 0.018739f $X=1.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_109 N_B2_M1028_g N_B1_M1000_g 0.018739f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_110 N_B2_c_112_n N_B1_c_193_n 0.00190901f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_111 N_B2_c_113_n N_B1_c_193_n 0.018739f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B2_M1003_g N_A_27_297#_c_395_n 7.12665e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B2_M1003_g N_A_27_297#_c_396_n 0.011048f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B2_M1005_g N_A_27_297#_c_396_n 6.53272e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B2_c_112_n N_A_27_297#_c_396_n 0.0271922f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B2_M1003_g N_A_27_297#_c_410_n 0.0101149f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B2_M1005_g N_A_27_297#_c_410_n 0.00988743f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_118 N_B2_M1021_g N_A_27_297#_c_412_n 0.00988743f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B2_M1028_g N_A_27_297#_c_412_n 0.00988743f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B2_M1028_g N_Y_c_512_n 0.0113206f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B2_c_112_n N_Y_c_512_n 0.0179392f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B2_c_111_n N_Y_c_510_n 9.27367e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B2_c_112_n N_Y_c_510_n 0.0108226f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_124 N_B2_c_113_n N_Y_c_510_n 0.0010701f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B2_M1005_g N_Y_c_515_n 0.0112596f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B2_M1021_g N_Y_c_515_n 0.0113206f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B2_c_112_n N_Y_c_515_n 0.0419177f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_128 N_B2_c_113_n N_Y_c_515_n 0.00214201f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_129 N_B2_c_112_n N_Y_c_516_n 0.0204933f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B2_c_113_n N_Y_c_516_n 0.00222181f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B2_M1003_g Y 5.53979e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_132 N_B2_c_112_n Y 0.017214f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_133 N_B2_c_113_n Y 0.00222181f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B2_M1003_g N_VPWR_c_613_n 0.00357835f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B2_M1005_g N_VPWR_c_613_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B2_M1021_g N_VPWR_c_613_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B2_M1028_g N_VPWR_c_613_n 0.00357877f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B2_M1003_g N_VPWR_c_607_n 0.00617934f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_139 N_B2_M1005_g N_VPWR_c_607_n 0.00522516f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B2_M1021_g N_VPWR_c_607_n 0.00522516f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B2_M1028_g N_VPWR_c_607_n 0.00525237f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B2_c_108_n N_A_27_47#_c_709_n 0.00630972f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B2_c_109_n N_A_27_47#_c_709_n 5.22228e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B2_c_108_n N_A_27_47#_c_710_n 0.00869873f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B2_c_109_n N_A_27_47#_c_710_n 0.00869873f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B2_c_112_n N_A_27_47#_c_710_n 0.0363039f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_147 N_B2_c_113_n N_A_27_47#_c_710_n 0.00222006f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B2_c_108_n N_A_27_47#_c_711_n 0.00129412f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_149 N_B2_c_112_n N_A_27_47#_c_711_n 0.0279679f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_150 N_B2_c_108_n N_A_27_47#_c_724_n 5.22228e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B2_c_109_n N_A_27_47#_c_724_n 0.00630972f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B2_c_110_n N_A_27_47#_c_724_n 0.00630972f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B2_c_111_n N_A_27_47#_c_724_n 5.22228e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B2_c_110_n N_A_27_47#_c_712_n 0.00865195f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B2_c_111_n N_A_27_47#_c_712_n 0.00869873f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B2_c_112_n N_A_27_47#_c_712_n 0.0363039f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B2_c_113_n N_A_27_47#_c_712_n 0.00222006f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_158 N_B2_c_111_n N_A_27_47#_c_732_n 0.00255288f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B2_c_110_n N_A_27_47#_c_713_n 4.58193e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B2_c_111_n N_A_27_47#_c_713_n 0.00485712f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B2_c_112_n N_A_27_47#_c_713_n 0.00992523f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_162 N_B2_c_109_n N_A_27_47#_c_715_n 0.00113159f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B2_c_110_n N_A_27_47#_c_715_n 0.00113159f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B2_c_112_n N_A_27_47#_c_715_n 0.0266779f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B2_c_113_n N_A_27_47#_c_715_n 0.00230167f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_166 N_B2_c_108_n N_VGND_c_777_n 0.00268723f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B2_c_109_n N_VGND_c_777_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B2_c_110_n N_VGND_c_778_n 0.00146448f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B2_c_111_n N_VGND_c_778_n 0.00268723f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B2_c_108_n N_VGND_c_781_n 0.00423334f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B2_c_109_n N_VGND_c_783_n 0.00423334f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B2_c_110_n N_VGND_c_783_n 0.00423334f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B2_c_111_n N_VGND_c_787_n 0.00421816f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B2_c_108_n N_VGND_c_789_n 0.00667051f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B2_c_109_n N_VGND_c_789_n 0.0057163f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B2_c_110_n N_VGND_c_789_n 0.0057163f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B2_c_111_n N_VGND_c_789_n 0.00575258f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B1_c_193_n N_A1_c_261_n 2.11242e-19 $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B1_c_194_n N_A1_c_261_n 0.0138294f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B1_c_193_n N_A1_c_262_n 0.00655684f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B1_c_194_n N_A1_c_262_n 9.97586e-19 $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_182 N_B1_M1000_g N_A_27_297#_c_414_n 0.00985793f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_M1006_g N_A_27_297#_c_414_n 0.00988743f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_M1024_g N_A_27_297#_c_416_n 0.00988743f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B1_M1029_g N_A_27_297#_c_416_n 0.0121747f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_M1029_g N_A_27_297#_c_397_n 7.27237e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B1_c_193_n N_A_27_297#_c_397_n 0.00406365f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B1_c_194_n N_A_27_297#_c_397_n 0.0440535f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B1_M1000_g N_Y_c_512_n 0.0127518f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B1_c_189_n N_Y_c_535_n 0.00292615f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B1_c_189_n N_Y_c_510_n 0.00275063f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B1_M1000_g N_Y_c_510_n 0.0031628f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B1_c_190_n N_Y_c_510_n 0.00279934f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B1_M1006_g N_Y_c_510_n 0.00306065f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_c_193_n N_Y_c_510_n 0.024791f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B1_c_194_n N_Y_c_510_n 0.0154944f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_197 N_B1_c_190_n N_Y_c_511_n 0.0116354f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B1_c_191_n N_Y_c_511_n 0.0103351f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_c_192_n N_Y_c_511_n 0.0133144f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B1_c_193_n N_Y_c_511_n 0.00854882f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B1_c_194_n N_Y_c_511_n 0.0864193f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_M1006_g N_Y_c_514_n 0.0127578f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B1_M1024_g N_Y_c_514_n 0.0112944f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_204 N_B1_c_193_n N_Y_c_514_n 0.00214321f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B1_c_194_n N_Y_c_514_n 0.0327326f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B1_M1000_g N_Y_c_517_n 0.00180885f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1029_g N_Y_c_518_n 5.90444e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_c_193_n N_Y_c_518_n 0.00222344f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_209 N_B1_c_194_n N_Y_c_518_n 0.0203891f $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B1_M1000_g N_VPWR_c_613_n 0.00357877f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1006_g N_VPWR_c_613_n 0.00357877f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1024_g N_VPWR_c_613_n 0.00357877f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1029_g N_VPWR_c_613_n 0.00357877f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1000_g N_VPWR_c_607_n 0.00525237f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1006_g N_VPWR_c_607_n 0.00522516f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B1_M1024_g N_VPWR_c_607_n 0.00522516f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_217 N_B1_M1029_g N_VPWR_c_607_n 0.00655123f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B1_c_189_n N_A_27_47#_c_714_n 0.0127015f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_190_n N_A_27_47#_c_714_n 0.00892725f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B1_c_191_n N_A_27_47#_c_714_n 0.00892725f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B1_c_192_n N_A_27_47#_c_714_n 0.00892725f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_193_n N_A_27_47#_c_714_n 3.07604e-19 $X=3.495 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B1_c_189_n N_VGND_c_787_n 0.00357877f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B1_c_190_n N_VGND_c_787_n 0.00357877f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B1_c_191_n N_VGND_c_787_n 0.00357877f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B1_c_192_n N_VGND_c_787_n 0.00357877f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_227 N_B1_c_189_n N_VGND_c_789_n 0.00525237f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B1_c_190_n N_VGND_c_789_n 0.00522516f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B1_c_191_n N_VGND_c_789_n 0.00522516f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B1_c_192_n N_VGND_c_789_n 0.00655123f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A1_c_260_n N_A2_c_320_n 0.0151343f $X=5.61 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_232 N_A1_M1030_g N_A2_M1002_g 0.0151343f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_c_261_n N_A2_c_324_n 0.0150082f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A1_c_262_n N_A2_c_324_n 8.87282e-19 $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A1_c_261_n N_A2_c_325_n 2.42383e-19 $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A1_c_262_n N_A2_c_325_n 0.0151343f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A1_M1001_g N_A_27_297#_c_398_n 0.0136219f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A1_M1009_g N_A_27_297#_c_398_n 0.0132714f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A1_c_261_n N_A_27_297#_c_398_n 0.0409754f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A1_c_262_n N_A_27_297#_c_398_n 0.00211509f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A1_M1012_g N_A_27_297#_c_399_n 0.0132714f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A1_M1030_g N_A_27_297#_c_399_n 0.0132641f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A1_c_261_n N_A_27_297#_c_399_n 0.0409754f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A1_c_262_n N_A_27_297#_c_399_n 0.00211509f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A1_c_261_n N_A_27_297#_c_403_n 0.0204549f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A1_c_262_n N_A_27_297#_c_403_n 0.00220041f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A1_c_257_n N_Y_c_511_n 0.0133144f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A1_c_258_n N_Y_c_511_n 0.0103351f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A1_c_259_n N_Y_c_511_n 0.0103351f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A1_c_260_n N_Y_c_511_n 0.00331492f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_261_n N_Y_c_511_n 0.0733505f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A1_c_262_n N_Y_c_511_n 0.00663066f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A1_M1001_g N_VPWR_c_608_n 0.00302074f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A1_M1009_g N_VPWR_c_608_n 0.00157837f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A1_M1009_g N_VPWR_c_609_n 0.00585385f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A1_M1012_g N_VPWR_c_609_n 0.00585385f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A1_M1012_g N_VPWR_c_610_n 0.00157837f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A1_M1030_g N_VPWR_c_610_n 0.00157837f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A1_M1001_g N_VPWR_c_613_n 0.00585385f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A1_M1030_g N_VPWR_c_617_n 0.00585385f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A1_M1001_g N_VPWR_c_607_n 0.0117628f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A1_M1009_g N_VPWR_c_607_n 0.0104367f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A1_M1012_g N_VPWR_c_607_n 0.0104367f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A1_M1030_g N_VPWR_c_607_n 0.010464f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A1_c_257_n N_VGND_c_787_n 0.00357877f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A1_c_258_n N_VGND_c_787_n 0.00357877f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A1_c_259_n N_VGND_c_787_n 0.00357877f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A1_c_260_n N_VGND_c_787_n 0.00357877f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A1_c_257_n N_VGND_c_789_n 0.00655123f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A1_c_258_n N_VGND_c_789_n 0.00522516f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_c_259_n N_VGND_c_789_n 0.00522516f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A1_c_260_n N_VGND_c_789_n 0.00525237f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A1_c_257_n N_A_803_47#_c_883_n 0.00892725f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A1_c_258_n N_A_803_47#_c_883_n 0.00892725f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A1_c_259_n N_A_803_47#_c_883_n 0.00892725f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A1_c_260_n N_A_803_47#_c_883_n 0.0105669f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A1_c_261_n N_A_803_47#_c_883_n 0.00295908f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_278 N_A1_c_260_n N_A_803_47#_c_884_n 6.06509e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A2_M1002_g N_A_27_297#_c_400_n 0.0132641f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_280 N_A2_M1004_g N_A_27_297#_c_400_n 0.0132714f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A2_c_324_n N_A_27_297#_c_400_n 0.041703f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A2_c_325_n N_A_27_297#_c_400_n 0.00211509f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A2_M1007_g N_A_27_297#_c_401_n 0.0132273f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A2_M1025_g N_A_27_297#_c_401_n 0.0134927f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A2_c_324_n N_A_27_297#_c_401_n 0.041703f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A2_c_325_n N_A_27_297#_c_401_n 0.00211509f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A2_c_324_n N_A_27_297#_c_402_n 0.0214236f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A2_c_324_n N_A_27_297#_c_404_n 0.0029993f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A2_c_324_n N_A_27_297#_c_405_n 0.0204549f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A2_c_325_n N_A_27_297#_c_405_n 0.00220041f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A2_M1002_g N_VPWR_c_611_n 0.00157837f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A2_M1004_g N_VPWR_c_611_n 0.00157837f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_293 N_A2_M1007_g N_VPWR_c_612_n 0.00157837f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A2_M1025_g N_VPWR_c_612_n 0.00302074f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A2_M1004_g N_VPWR_c_615_n 0.00585385f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_296 N_A2_M1007_g N_VPWR_c_615_n 0.00585385f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A2_M1002_g N_VPWR_c_617_n 0.00585385f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A2_M1025_g N_VPWR_c_618_n 0.00585385f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A2_M1002_g N_VPWR_c_607_n 0.010464f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A2_M1004_g N_VPWR_c_607_n 0.0104367f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A2_M1007_g N_VPWR_c_607_n 0.0104367f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_302 N_A2_M1025_g N_VPWR_c_607_n 0.0114438f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A2_c_320_n N_VGND_c_779_n 0.00268723f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A2_c_321_n N_VGND_c_779_n 0.00146448f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A2_c_322_n N_VGND_c_780_n 0.00146448f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A2_c_323_n N_VGND_c_780_n 0.00268723f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A2_c_321_n N_VGND_c_785_n 0.00423334f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A2_c_322_n N_VGND_c_785_n 0.00423334f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A2_c_320_n N_VGND_c_787_n 0.00421816f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A2_c_323_n N_VGND_c_788_n 0.00423334f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A2_c_320_n N_VGND_c_789_n 0.00575258f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A2_c_321_n N_VGND_c_789_n 0.0057163f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A2_c_322_n N_VGND_c_789_n 0.0057163f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A2_c_323_n N_VGND_c_789_n 0.00672331f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A2_c_320_n N_A_803_47#_c_895_n 0.00255288f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A2_c_320_n N_A_803_47#_c_884_n 0.00485843f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A2_c_321_n N_A_803_47#_c_884_n 4.58193e-19 $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A2_c_324_n N_A_803_47#_c_884_n 0.0061524f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A2_c_320_n N_A_803_47#_c_885_n 0.00870364f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A2_c_321_n N_A_803_47#_c_885_n 0.00865686f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A2_c_324_n N_A_803_47#_c_885_n 0.0362443f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A2_c_325_n N_A_803_47#_c_885_n 0.00222133f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A2_c_320_n N_A_803_47#_c_903_n 5.22228e-19 $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A2_c_321_n N_A_803_47#_c_903_n 0.00630972f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A2_c_322_n N_A_803_47#_c_903_n 0.00630972f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A2_c_323_n N_A_803_47#_c_903_n 5.22228e-19 $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A2_c_322_n N_A_803_47#_c_886_n 0.00870364f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A2_c_323_n N_A_803_47#_c_886_n 0.00999903f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A2_c_324_n N_A_803_47#_c_886_n 0.0641689f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A2_c_325_n N_A_803_47#_c_886_n 0.00222133f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A2_c_322_n N_A_803_47#_c_887_n 5.22228e-19 $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A2_c_323_n N_A_803_47#_c_887_n 0.00630972f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A2_c_321_n N_A_803_47#_c_888_n 0.00113286f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A2_c_322_n N_A_803_47#_c_888_n 0.00113286f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A2_c_324_n N_A_803_47#_c_888_n 0.0266272f $X=7.14 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A2_c_325_n N_A_803_47#_c_888_n 0.00230339f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_27_297#_c_410_n N_Y_M1003_d 0.00312348f $X=0.975 $Y=2.38 $X2=0 $Y2=0
cc_338 N_A_27_297#_c_412_n N_Y_M1021_d 0.00312348f $X=1.815 $Y=2.38 $X2=0 $Y2=0
cc_339 N_A_27_297#_c_414_n N_Y_M1000_d 0.00312348f $X=2.655 $Y=2.38 $X2=0 $Y2=0
cc_340 N_A_27_297#_c_416_n N_Y_M1024_d 0.00312348f $X=3.495 $Y=2.38 $X2=0 $Y2=0
cc_341 N_A_27_297#_M1028_s N_Y_c_512_n 0.00166124f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_342 N_A_27_297#_c_412_n N_Y_c_512_n 0.00322336f $X=1.815 $Y=2.38 $X2=0 $Y2=0
cc_343 N_A_27_297#_c_449_p N_Y_c_512_n 0.0127256f $X=1.94 $Y=1.96 $X2=0 $Y2=0
cc_344 N_A_27_297#_c_414_n N_Y_c_512_n 0.00257436f $X=2.655 $Y=2.38 $X2=0 $Y2=0
cc_345 N_A_27_297#_c_397_n N_Y_c_511_n 0.00728694f $X=3.88 $Y=1.625 $X2=0 $Y2=0
cc_346 N_A_27_297#_M1006_s N_Y_c_514_n 0.00166124f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_347 N_A_27_297#_c_414_n N_Y_c_514_n 0.00322336f $X=2.655 $Y=2.38 $X2=0 $Y2=0
cc_348 N_A_27_297#_c_454_p N_Y_c_514_n 0.0127256f $X=2.78 $Y=1.96 $X2=0 $Y2=0
cc_349 N_A_27_297#_c_416_n N_Y_c_514_n 0.00322336f $X=3.495 $Y=2.38 $X2=0 $Y2=0
cc_350 N_A_27_297#_M1005_s N_Y_c_515_n 0.00166124f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_351 N_A_27_297#_c_410_n N_Y_c_515_n 0.00322336f $X=0.975 $Y=2.38 $X2=0 $Y2=0
cc_352 N_A_27_297#_c_458_p N_Y_c_515_n 0.0127256f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_353 N_A_27_297#_c_412_n N_Y_c_515_n 0.00322336f $X=1.815 $Y=2.38 $X2=0 $Y2=0
cc_354 N_A_27_297#_c_412_n N_Y_c_516_n 0.0118865f $X=1.815 $Y=2.38 $X2=0 $Y2=0
cc_355 N_A_27_297#_c_414_n N_Y_c_517_n 0.0125836f $X=2.655 $Y=2.38 $X2=0 $Y2=0
cc_356 N_A_27_297#_c_416_n N_Y_c_518_n 0.0118865f $X=3.495 $Y=2.38 $X2=0 $Y2=0
cc_357 N_A_27_297#_c_397_n N_Y_c_518_n 0.00271526f $X=3.88 $Y=1.625 $X2=0 $Y2=0
cc_358 N_A_27_297#_c_396_n Y 0.00777584f $X=0.26 $Y=1.64 $X2=0 $Y2=0
cc_359 N_A_27_297#_c_410_n Y 0.0118865f $X=0.975 $Y=2.38 $X2=0 $Y2=0
cc_360 N_A_27_297#_c_398_n N_VPWR_M1001_d 0.00165831f $X=4.855 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_361 N_A_27_297#_c_399_n N_VPWR_M1012_d 0.00165831f $X=5.695 $Y=1.54 $X2=0
+ $Y2=0
cc_362 N_A_27_297#_c_400_n N_VPWR_M1002_d 0.00165831f $X=6.535 $Y=1.54 $X2=0
+ $Y2=0
cc_363 N_A_27_297#_c_401_n N_VPWR_M1007_d 0.00165831f $X=7.375 $Y=1.54 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_c_398_n N_VPWR_c_608_n 0.0126919f $X=4.855 $Y=1.54 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_c_471_p N_VPWR_c_609_n 0.0142343f $X=4.98 $Y=2.3 $X2=0 $Y2=0
cc_366 N_A_27_297#_c_399_n N_VPWR_c_610_n 0.0126919f $X=5.695 $Y=1.54 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_c_400_n N_VPWR_c_611_n 0.0126919f $X=6.535 $Y=1.54 $X2=0
+ $Y2=0
cc_368 N_A_27_297#_c_401_n N_VPWR_c_612_n 0.0126919f $X=7.375 $Y=1.54 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_395_n N_VPWR_c_613_n 0.0215365f $X=0.257 $Y=2.295 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_410_n N_VPWR_c_613_n 0.0308192f $X=0.975 $Y=2.38 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_412_n N_VPWR_c_613_n 0.0330174f $X=1.815 $Y=2.38 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_414_n N_VPWR_c_613_n 0.0330174f $X=2.655 $Y=2.38 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_416_n N_VPWR_c_613_n 0.0330174f $X=3.495 $Y=2.38 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_c_480_p N_VPWR_c_613_n 0.050872f $X=3.88 $Y=2.295 $X2=0 $Y2=0
cc_375 N_A_27_297#_c_481_p N_VPWR_c_613_n 0.0142933f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_376 N_A_27_297#_c_482_p N_VPWR_c_613_n 0.0142933f $X=1.94 $Y=2.38 $X2=0 $Y2=0
cc_377 N_A_27_297#_c_483_p N_VPWR_c_613_n 0.0142933f $X=2.78 $Y=2.38 $X2=0 $Y2=0
cc_378 N_A_27_297#_c_484_p N_VPWR_c_615_n 0.0142343f $X=6.66 $Y=2.3 $X2=0 $Y2=0
cc_379 N_A_27_297#_c_485_p N_VPWR_c_617_n 0.0142343f $X=5.82 $Y=2.3 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_486_p N_VPWR_c_618_n 0.0158369f $X=7.5 $Y=2.3 $X2=0 $Y2=0
cc_381 N_A_27_297#_M1003_s N_VPWR_c_607_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_M1005_s N_VPWR_c_607_n 0.00215203f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_M1028_s N_VPWR_c_607_n 0.00215203f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_M1006_s N_VPWR_c_607_n 0.00215203f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_385 N_A_27_297#_M1029_s N_VPWR_c_607_n 0.00671229f $X=3.485 $Y=1.485 $X2=0
+ $Y2=0
cc_386 N_A_27_297#_M1009_s N_VPWR_c_607_n 0.00284632f $X=4.845 $Y=1.485 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_M1030_s N_VPWR_c_607_n 0.00284632f $X=5.685 $Y=1.485 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_M1004_s N_VPWR_c_607_n 0.00284632f $X=6.525 $Y=1.485 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_M1025_s N_VPWR_c_607_n 0.00419161f $X=7.365 $Y=1.485 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_c_395_n N_VPWR_c_607_n 0.0126918f $X=0.257 $Y=2.295 $X2=0
+ $Y2=0
cc_391 N_A_27_297#_c_410_n N_VPWR_c_607_n 0.0191798f $X=0.975 $Y=2.38 $X2=0
+ $Y2=0
cc_392 N_A_27_297#_c_412_n N_VPWR_c_607_n 0.0204627f $X=1.815 $Y=2.38 $X2=0
+ $Y2=0
cc_393 N_A_27_297#_c_414_n N_VPWR_c_607_n 0.0204627f $X=2.655 $Y=2.38 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_416_n N_VPWR_c_607_n 0.0204627f $X=3.495 $Y=2.38 $X2=0
+ $Y2=0
cc_395 N_A_27_297#_c_480_p N_VPWR_c_607_n 0.0296541f $X=3.88 $Y=2.295 $X2=0
+ $Y2=0
cc_396 N_A_27_297#_c_471_p N_VPWR_c_607_n 0.00955092f $X=4.98 $Y=2.3 $X2=0 $Y2=0
cc_397 N_A_27_297#_c_485_p N_VPWR_c_607_n 0.00955092f $X=5.82 $Y=2.3 $X2=0 $Y2=0
cc_398 N_A_27_297#_c_484_p N_VPWR_c_607_n 0.00955092f $X=6.66 $Y=2.3 $X2=0 $Y2=0
cc_399 N_A_27_297#_c_486_p N_VPWR_c_607_n 0.00955092f $X=7.5 $Y=2.3 $X2=0 $Y2=0
cc_400 N_A_27_297#_c_481_p N_VPWR_c_607_n 0.00962421f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_482_p N_VPWR_c_607_n 0.00962421f $X=1.94 $Y=2.38 $X2=0
+ $Y2=0
cc_402 N_A_27_297#_c_483_p N_VPWR_c_607_n 0.00962421f $X=2.78 $Y=2.38 $X2=0
+ $Y2=0
cc_403 N_A_27_297#_c_404_n N_A_803_47#_c_884_n 0.00719897f $X=5.82 $Y=1.62 $X2=0
+ $Y2=0
cc_404 N_Y_M1003_d N_VPWR_c_607_n 0.00216833f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_405 N_Y_M1021_d N_VPWR_c_607_n 0.00216833f $X=1.385 $Y=1.485 $X2=0 $Y2=0
cc_406 N_Y_M1000_d N_VPWR_c_607_n 0.00216833f $X=2.225 $Y=1.485 $X2=0 $Y2=0
cc_407 N_Y_M1024_d N_VPWR_c_607_n 0.00216833f $X=3.065 $Y=1.485 $X2=0 $Y2=0
cc_408 N_Y_c_511_n N_A_27_47#_M1022_s 0.00314455f $X=5.4 $Y=0.73 $X2=0 $Y2=0
cc_409 N_Y_c_511_n N_A_27_47#_M1027_s 0.0051435f $X=5.4 $Y=0.73 $X2=0 $Y2=0
cc_410 N_Y_c_512_n N_A_27_47#_c_713_n 0.00495371f $X=2.195 $Y=1.535 $X2=0 $Y2=0
cc_411 N_Y_c_510_n N_A_27_47#_c_713_n 0.00157225f $X=2.32 $Y=1.445 $X2=0 $Y2=0
cc_412 N_Y_M1017_d N_A_27_47#_c_714_n 0.00304656f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_413 N_Y_M1026_d N_A_27_47#_c_714_n 0.00305026f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_414 N_Y_c_535_n N_A_27_47#_c_714_n 0.0143975f $X=2.32 $Y=0.885 $X2=0 $Y2=0
cc_415 N_Y_c_511_n N_A_27_47#_c_714_n 0.0703475f $X=5.4 $Y=0.73 $X2=0 $Y2=0
cc_416 N_Y_c_511_n N_VGND_c_787_n 0.00348529f $X=5.4 $Y=0.73 $X2=0 $Y2=0
cc_417 N_Y_M1017_d N_VGND_c_789_n 0.00216833f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_418 N_Y_M1026_d N_VGND_c_789_n 0.00216833f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_419 N_Y_M1010_d N_VGND_c_789_n 0.00216833f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_420 N_Y_M1018_d N_VGND_c_789_n 0.00216833f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_421 N_Y_c_511_n N_VGND_c_789_n 0.0110378f $X=5.4 $Y=0.73 $X2=0 $Y2=0
cc_422 N_Y_c_511_n N_A_803_47#_M1010_s 0.0069299f $X=5.4 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_423 N_Y_c_511_n N_A_803_47#_M1014_s 0.00314455f $X=5.4 $Y=0.73 $X2=0 $Y2=0
cc_424 N_Y_M1010_d N_A_803_47#_c_883_n 0.00305026f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_425 N_Y_M1018_d N_A_803_47#_c_883_n 0.00305026f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_426 N_Y_c_511_n N_A_803_47#_c_883_n 0.0836052f $X=5.4 $Y=0.73 $X2=0 $Y2=0
cc_427 N_A_27_47#_c_710_n N_VGND_M1013_s 0.00162089f $X=0.935 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_428 N_A_27_47#_c_712_n N_VGND_M1020_s 0.00162089f $X=1.775 $Y=0.815 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_710_n N_VGND_c_777_n 0.0122559f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_712_n N_VGND_c_778_n 0.0122559f $X=1.775 $Y=0.815 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_c_709_n N_VGND_c_781_n 0.0209752f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_710_n N_VGND_c_781_n 0.00198695f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_710_n N_VGND_c_783_n 0.00198695f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_724_n N_VGND_c_783_n 0.0188551f $X=1.1 $Y=0.39 $X2=0 $Y2=0
cc_435 N_A_27_47#_c_712_n N_VGND_c_783_n 0.00198695f $X=1.775 $Y=0.815 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_712_n N_VGND_c_787_n 0.00198695f $X=1.775 $Y=0.815 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_732_n N_VGND_c_787_n 0.0152108f $X=1.9 $Y=0.475 $X2=0 $Y2=0
cc_438 N_A_27_47#_c_714_n N_VGND_c_787_n 0.0991765f $X=3.62 $Y=0.39 $X2=0 $Y2=0
cc_439 N_A_27_47#_M1013_d N_VGND_c_789_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_M1016_d N_VGND_c_789_n 0.00215201f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_M1031_d N_VGND_c_789_n 0.00215206f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_M1022_s N_VGND_c_789_n 0.00215227f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_M1027_s N_VGND_c_789_n 0.00209344f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_709_n N_VGND_c_789_n 0.0124119f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_445 N_A_27_47#_c_710_n N_VGND_c_789_n 0.00835832f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_c_724_n N_VGND_c_789_n 0.0122069f $X=1.1 $Y=0.39 $X2=0 $Y2=0
cc_447 N_A_27_47#_c_712_n N_VGND_c_789_n 0.00835832f $X=1.775 $Y=0.815 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_732_n N_VGND_c_789_n 0.00940698f $X=1.9 $Y=0.475 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_714_n N_VGND_c_789_n 0.0628989f $X=3.62 $Y=0.39 $X2=0 $Y2=0
cc_450 N_A_27_47#_c_714_n N_A_803_47#_c_883_n 0.0188707f $X=3.62 $Y=0.39 $X2=0
+ $Y2=0
cc_451 N_VGND_c_789_n N_A_803_47#_M1010_s 0.00209344f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_452 N_VGND_c_789_n N_A_803_47#_M1014_s 0.00215227f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_c_789_n N_A_803_47#_M1023_s 0.00215206f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_789_n N_A_803_47#_M1011_s 0.00215201f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_455 N_VGND_c_789_n N_A_803_47#_M1019_s 0.00209319f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_456 N_VGND_c_787_n N_A_803_47#_c_883_n 0.0991765f $X=6.155 $Y=0 $X2=0 $Y2=0
cc_457 N_VGND_c_789_n N_A_803_47#_c_883_n 0.0628989f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_787_n N_A_803_47#_c_895_n 0.0152108f $X=6.155 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_789_n N_A_803_47#_c_895_n 0.00940698f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_460 N_VGND_M1008_d N_A_803_47#_c_885_n 0.00162089f $X=6.105 $Y=0.235 $X2=0
+ $Y2=0
cc_461 N_VGND_c_779_n N_A_803_47#_c_885_n 0.0122559f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_462 N_VGND_c_785_n N_A_803_47#_c_885_n 0.00198695f $X=6.995 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_c_787_n N_A_803_47#_c_885_n 0.00198695f $X=6.155 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_789_n N_A_803_47#_c_885_n 0.00835832f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_465 N_VGND_c_785_n N_A_803_47#_c_903_n 0.0188551f $X=6.995 $Y=0 $X2=0 $Y2=0
cc_466 N_VGND_c_789_n N_A_803_47#_c_903_n 0.0122069f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_M1015_d N_A_803_47#_c_886_n 0.00162089f $X=6.945 $Y=0.235 $X2=0
+ $Y2=0
cc_468 N_VGND_c_780_n N_A_803_47#_c_886_n 0.0122559f $X=7.08 $Y=0.39 $X2=0 $Y2=0
cc_469 N_VGND_c_785_n N_A_803_47#_c_886_n 0.00198695f $X=6.995 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_788_n N_A_803_47#_c_886_n 0.00198695f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_789_n N_A_803_47#_c_886_n 0.00835832f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_788_n N_A_803_47#_c_887_n 0.0209752f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_789_n N_A_803_47#_c_887_n 0.0124119f $X=7.59 $Y=0 $X2=0 $Y2=0

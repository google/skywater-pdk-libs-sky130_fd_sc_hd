* File: sky130_fd_sc_hd__sedfxtp_1.pxi.spice
* Created: Tue Sep  1 19:32:08 2020
* 
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%CLK N_CLK_c_275_n N_CLK_c_279_n N_CLK_c_276_n
+ N_CLK_M1040_g N_CLK_c_280_n N_CLK_M1014_g N_CLK_c_281_n CLK
+ PM_SKY130_FD_SC_HD__SEDFXTP_1%CLK
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_27_47# N_A_27_47#_M1040_s N_A_27_47#_M1014_s
+ N_A_27_47#_M1021_g N_A_27_47#_M1000_g N_A_27_47#_M1027_g N_A_27_47#_M1016_g
+ N_A_27_47#_M1025_g N_A_27_47#_c_317_n N_A_27_47#_M1028_g N_A_27_47#_c_577_p
+ N_A_27_47#_c_319_n N_A_27_47#_c_320_n N_A_27_47#_c_332_n N_A_27_47#_c_464_p
+ N_A_27_47#_c_321_n N_A_27_47#_c_322_n N_A_27_47#_c_323_n N_A_27_47#_c_324_n
+ N_A_27_47#_c_335_n N_A_27_47#_c_336_n N_A_27_47#_c_337_n N_A_27_47#_c_338_n
+ N_A_27_47#_c_339_n N_A_27_47#_c_340_n N_A_27_47#_c_341_n N_A_27_47#_c_325_n
+ N_A_27_47#_c_343_n N_A_27_47#_c_326_n N_A_27_47#_c_327_n
+ PM_SKY130_FD_SC_HD__SEDFXTP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%D N_D_M1002_g N_D_M1029_g N_D_c_591_n
+ N_D_c_595_n D N_D_c_593_n PM_SKY130_FD_SC_HD__SEDFXTP_1%D
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_423_343# N_A_423_343#_M1038_s
+ N_A_423_343#_M1011_s N_A_423_343#_c_647_n N_A_423_343#_M1032_g
+ N_A_423_343#_M1022_g N_A_423_343#_c_648_n N_A_423_343#_c_642_n
+ N_A_423_343#_c_643_n N_A_423_343#_c_644_n N_A_423_343#_c_645_n
+ N_A_423_343#_c_646_n PM_SKY130_FD_SC_HD__SEDFXTP_1%A_423_343#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%DE N_DE_M1003_g N_DE_c_730_n N_DE_c_731_n
+ N_DE_M1038_g N_DE_c_733_n N_DE_M1011_g N_DE_c_738_n N_DE_M1015_g N_DE_c_734_n
+ N_DE_c_740_n DE PM_SKY130_FD_SC_HD__SEDFXTP_1%DE
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_791_264# N_A_791_264#_M1031_s
+ N_A_791_264#_M1023_s N_A_791_264#_M1041_g N_A_791_264#_M1036_g
+ N_A_791_264#_M1007_g N_A_791_264#_M1001_g N_A_791_264#_c_827_n
+ N_A_791_264#_c_828_n N_A_791_264#_c_829_n N_A_791_264#_c_816_n
+ N_A_791_264#_c_830_n N_A_791_264#_c_831_n N_A_791_264#_c_832_n
+ N_A_791_264#_c_817_n N_A_791_264#_c_818_n N_A_791_264#_c_819_n
+ N_A_791_264#_c_820_n N_A_791_264#_c_821_n N_A_791_264#_c_822_n
+ PM_SKY130_FD_SC_HD__SEDFXTP_1%A_791_264#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_885_21# N_A_885_21#_M1005_s
+ N_A_885_21#_M1033_s N_A_885_21#_c_1002_n N_A_885_21#_M1034_g
+ N_A_885_21#_c_1003_n N_A_885_21#_c_1004_n N_A_885_21#_c_1005_n
+ N_A_885_21#_M1030_g N_A_885_21#_c_1006_n N_A_885_21#_c_1007_n
+ N_A_885_21#_c_1008_n N_A_885_21#_c_1009_n N_A_885_21#_c_1015_n
+ N_A_885_21#_c_1010_n N_A_885_21#_c_1011_n N_A_885_21#_c_1018_n
+ N_A_885_21#_c_1012_n PM_SKY130_FD_SC_HD__SEDFXTP_1%A_885_21#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%SCD N_SCD_M1024_g N_SCD_M1020_g SCD
+ N_SCD_c_1133_n PM_SKY130_FD_SC_HD__SEDFXTP_1%SCD
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%SCE N_SCE_M1013_g N_SCE_c_1179_n N_SCE_c_1188_n
+ N_SCE_M1033_g N_SCE_M1005_g N_SCE_c_1181_n N_SCE_c_1182_n N_SCE_M1009_g SCE
+ N_SCE_c_1184_n N_SCE_c_1185_n PM_SKY130_FD_SC_HD__SEDFXTP_1%SCE
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_193_47# N_A_193_47#_M1021_d
+ N_A_193_47#_M1000_d N_A_193_47#_M1008_g N_A_193_47#_c_1273_n
+ N_A_193_47#_M1012_g N_A_193_47#_c_1275_n N_A_193_47#_M1026_g
+ N_A_193_47#_M1018_g N_A_193_47#_c_1276_n N_A_193_47#_c_1277_n
+ N_A_193_47#_c_1285_n N_A_193_47#_c_1286_n N_A_193_47#_c_1287_n
+ N_A_193_47#_c_1288_n N_A_193_47#_c_1331_n N_A_193_47#_c_1278_n
+ N_A_193_47#_c_1279_n N_A_193_47#_c_1280_n N_A_193_47#_c_1292_n
+ N_A_193_47#_c_1281_n PM_SKY130_FD_SC_HD__SEDFXTP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_1610_159# N_A_1610_159#_M1004_d
+ N_A_1610_159#_M1017_d N_A_1610_159#_M1006_g N_A_1610_159#_M1019_g
+ N_A_1610_159#_M1037_g N_A_1610_159#_M1039_g N_A_1610_159#_c_1492_n
+ N_A_1610_159#_c_1493_n N_A_1610_159#_c_1494_n N_A_1610_159#_c_1495_n
+ N_A_1610_159#_c_1504_n N_A_1610_159#_c_1496_n N_A_1610_159#_c_1497_n
+ N_A_1610_159#_c_1498_n N_A_1610_159#_c_1499_n
+ PM_SKY130_FD_SC_HD__SEDFXTP_1%A_1610_159#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_1446_413# N_A_1446_413#_M1027_d
+ N_A_1446_413#_M1008_d N_A_1446_413#_c_1607_n N_A_1446_413#_M1017_g
+ N_A_1446_413#_M1004_g N_A_1446_413#_c_1608_n N_A_1446_413#_c_1609_n
+ N_A_1446_413#_c_1610_n N_A_1446_413#_c_1611_n N_A_1446_413#_c_1621_n
+ N_A_1446_413#_c_1627_n N_A_1446_413#_c_1612_n N_A_1446_413#_c_1617_n
+ N_A_1446_413#_c_1613_n PM_SKY130_FD_SC_HD__SEDFXTP_1%A_1446_413#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_2051_413# N_A_2051_413#_M1026_d
+ N_A_2051_413#_M1025_d N_A_2051_413#_M1031_g N_A_2051_413#_M1023_g
+ N_A_2051_413#_c_1714_n N_A_2051_413#_c_1715_n N_A_2051_413#_M1035_g
+ N_A_2051_413#_M1010_g N_A_2051_413#_c_1716_n N_A_2051_413#_c_1717_n
+ N_A_2051_413#_c_1718_n N_A_2051_413#_c_1730_n N_A_2051_413#_c_1733_n
+ N_A_2051_413#_c_1719_n N_A_2051_413#_c_1728_n N_A_2051_413#_c_1720_n
+ N_A_2051_413#_c_1721_n PM_SKY130_FD_SC_HD__SEDFXTP_1%A_2051_413#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%VPWR N_VPWR_M1014_d N_VPWR_M1032_d
+ N_VPWR_M1011_d N_VPWR_M1033_d N_VPWR_M1006_d N_VPWR_M1037_s N_VPWR_M1007_d
+ N_VPWR_M1023_d N_VPWR_c_1824_n N_VPWR_c_1825_n N_VPWR_c_1826_n N_VPWR_c_1827_n
+ N_VPWR_c_1828_n N_VPWR_c_1829_n N_VPWR_c_1830_n N_VPWR_c_1831_n
+ N_VPWR_c_1832_n N_VPWR_c_1833_n N_VPWR_c_1834_n N_VPWR_c_1835_n
+ N_VPWR_c_1836_n N_VPWR_c_1837_n N_VPWR_c_1838_n VPWR N_VPWR_c_1839_n
+ N_VPWR_c_1840_n N_VPWR_c_1841_n N_VPWR_c_1842_n N_VPWR_c_1843_n
+ N_VPWR_c_1823_n N_VPWR_c_1845_n N_VPWR_c_1846_n N_VPWR_c_1847_n
+ N_VPWR_c_1848_n N_VPWR_c_1849_n PM_SKY130_FD_SC_HD__SEDFXTP_1%VPWR
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_299_47# N_A_299_47#_M1002_s
+ N_A_299_47#_M1041_d N_A_299_47#_M1029_s N_A_299_47#_M1036_d
+ N_A_299_47#_c_2016_n N_A_299_47#_c_2009_n N_A_299_47#_c_2018_n
+ N_A_299_47#_c_2010_n N_A_299_47#_c_2011_n N_A_299_47#_c_2012_n
+ N_A_299_47#_c_2040_n N_A_299_47#_c_2013_n N_A_299_47#_c_2014_n
+ N_A_299_47#_c_2015_n PM_SKY130_FD_SC_HD__SEDFXTP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%A_915_47# N_A_915_47#_M1034_d
+ N_A_915_47#_M1009_d N_A_915_47#_M1013_d N_A_915_47#_M1030_d
+ N_A_915_47#_c_2138_n N_A_915_47#_c_2139_n N_A_915_47#_c_2130_n
+ N_A_915_47#_c_2151_n N_A_915_47#_c_2131_n N_A_915_47#_c_2140_n
+ N_A_915_47#_c_2132_n N_A_915_47#_c_2133_n N_A_915_47#_c_2155_n
+ N_A_915_47#_c_2134_n N_A_915_47#_c_2135_n N_A_915_47#_c_2168_n
+ N_A_915_47#_c_2136_n N_A_915_47#_c_2192_n N_A_915_47#_c_2137_n
+ PM_SKY130_FD_SC_HD__SEDFXTP_1%A_915_47#
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%Q N_Q_M1035_d N_Q_M1010_d Q N_Q_c_2269_n
+ PM_SKY130_FD_SC_HD__SEDFXTP_1%Q
x_PM_SKY130_FD_SC_HD__SEDFXTP_1%VGND N_VGND_M1040_d N_VGND_M1003_d
+ N_VGND_M1038_d N_VGND_M1005_d N_VGND_M1019_d N_VGND_M1039_s N_VGND_M1001_d
+ N_VGND_M1031_d N_VGND_c_2286_n N_VGND_c_2287_n N_VGND_c_2288_n N_VGND_c_2289_n
+ N_VGND_c_2290_n N_VGND_c_2291_n N_VGND_c_2292_n N_VGND_c_2293_n
+ N_VGND_c_2294_n N_VGND_c_2295_n N_VGND_c_2296_n N_VGND_c_2297_n
+ N_VGND_c_2298_n N_VGND_c_2299_n N_VGND_c_2300_n N_VGND_c_2301_n
+ N_VGND_c_2302_n N_VGND_c_2303_n VGND N_VGND_c_2304_n N_VGND_c_2305_n
+ N_VGND_c_2306_n N_VGND_c_2307_n N_VGND_c_2308_n N_VGND_c_2309_n
+ N_VGND_c_2310_n N_VGND_c_2311_n PM_SKY130_FD_SC_HD__SEDFXTP_1%VGND
cc_1 VNB N_CLK_c_275_n 0.0573151f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_276_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0185843f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1021_g 0.0373293f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1027_g 0.0216935f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_6 VNB N_A_27_47#_c_317_n 0.0139254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1028_g 0.0461694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_319_n 0.00191938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_320_n 0.00646065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_321_n 0.0024678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_322_n 0.00363529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_323_n 0.0294633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_324_n 0.00457671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_325_n 0.0236749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_326_n 0.00915868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_327_n 0.00210612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_M1002_g 0.0308382f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_18 VNB N_D_c_591_n 0.0161793f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_19 VNB D 0.00399003f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_20 VNB N_D_c_593_n 0.0145063f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_21 VNB N_A_423_343#_M1022_g 0.0217809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_423_343#_c_642_n 0.00769004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_423_343#_c_643_n 0.00185686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_423_343#_c_644_n 0.00333068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_423_343#_c_645_n 0.0291606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_423_343#_c_646_n 0.00198824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_DE_M1003_g 0.0211774f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_28 VNB N_DE_c_730_n 0.0423212f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_29 VNB N_DE_c_731_n 0.032977f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_30 VNB N_DE_M1038_g 0.0242274f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_31 VNB N_DE_c_733_n 0.0180937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_DE_c_734_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB DE 0.0110099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_791_264#_M1041_g 0.0476987f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_35 VNB N_A_791_264#_M1001_g 0.0480681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_791_264#_c_816_n 0.00377528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_791_264#_c_817_n 0.00469958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_791_264#_c_818_n 0.0371933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_791_264#_c_819_n 0.00419717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_791_264#_c_820_n 0.0132319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_791_264#_c_821_n 0.0013422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_791_264#_c_822_n 0.00158979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_885_21#_c_1002_n 0.0185371f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_44 VNB N_A_885_21#_c_1003_n 0.0301762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_885_21#_c_1004_n 0.00817921f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_46 VNB N_A_885_21#_c_1005_n 0.0151729f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_47 VNB N_A_885_21#_c_1006_n 0.00514919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_885_21#_c_1007_n 0.0328426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_885_21#_c_1008_n 0.00206328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_885_21#_c_1009_n 0.00322383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_885_21#_c_1010_n 0.00155169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_885_21#_c_1011_n 0.0108423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_885_21#_c_1012_n 0.00171304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_SCD_M1024_g 0.025414f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_55 VNB SCD 0.00875808f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_56 VNB N_SCD_c_1133_n 0.00758678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_SCE_c_1179_n 0.00191916f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_58 VNB N_SCE_M1005_g 0.0223821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_SCE_c_1181_n 0.054228f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_60 VNB N_SCE_c_1182_n 0.011117f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_61 VNB N_SCE_M1009_g 0.032127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_SCE_c_1184_n 0.00506878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_SCE_c_1185_n 0.0492389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_193_47#_c_1273_n 0.0136524f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_65 VNB N_A_193_47#_M1012_g 0.0429795f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_66 VNB N_A_193_47#_c_1275_n 0.0180286f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_67 VNB N_A_193_47#_c_1276_n 0.00392862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_193_47#_c_1277_n 0.0296727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_193_47#_c_1278_n 0.0032859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_193_47#_c_1279_n 0.017087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_193_47#_c_1280_n 0.00243891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_193_47#_c_1281_n 0.0122334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1610_159#_M1006_g 0.0138674f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_74 VNB N_A_1610_159#_M1019_g 0.0197771f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_75 VNB N_A_1610_159#_M1039_g 0.0283997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1610_159#_c_1492_n 0.0223712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1610_159#_c_1493_n 0.00481399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1610_159#_c_1494_n 0.00932364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1610_159#_c_1495_n 0.00611738f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1610_159#_c_1496_n 0.0048611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1610_159#_c_1497_n 0.0162827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1610_159#_c_1498_n 0.00249997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1610_159#_c_1499_n 0.0317753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1446_413#_c_1607_n 0.0113827f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_85 VNB N_A_1446_413#_c_1608_n 0.0181892f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_86 VNB N_A_1446_413#_c_1609_n 0.0133197f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_87 VNB N_A_1446_413#_c_1610_n 0.00937183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1446_413#_c_1611_n 0.00117523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1446_413#_c_1612_n 0.0117046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1446_413#_c_1613_n 0.00182328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_2051_413#_M1031_g 0.0350674f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_92 VNB N_A_2051_413#_c_1714_n 0.0145702f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_93 VNB N_A_2051_413#_c_1715_n 0.0205457f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_94 VNB N_A_2051_413#_c_1716_n 0.0384709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2051_413#_c_1717_n 0.004935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_2051_413#_c_1718_n 0.0137821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_2051_413#_c_1719_n 0.00719187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_2051_413#_c_1720_n 0.00330077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_2051_413#_c_1721_n 0.002763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VPWR_c_1823_n 0.554392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_299_47#_c_2009_n 0.0139151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_A_299_47#_c_2010_n 0.00281199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_A_299_47#_c_2011_n 0.00489253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_A_299_47#_c_2012_n 0.00419923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_A_299_47#_c_2013_n 0.00440827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_A_299_47#_c_2014_n 0.0029736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_A_299_47#_c_2015_n 0.00400821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_A_915_47#_c_2130_n 2.84745e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_A_915_47#_c_2131_n 0.00181891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_A_915_47#_c_2132_n 0.00904269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_A_915_47#_c_2133_n 0.00845782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_A_915_47#_c_2134_n 0.00538797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_A_915_47#_c_2135_n 5.21438e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_A_915_47#_c_2136_n 0.00569869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_A_915_47#_c_2137_n 0.00349341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_Q_c_2269_n 0.0401252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2286_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2287_n 0.00461568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2288_n 4.14e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2289_n 0.00410737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2290_n 0.00284902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2291_n 0.00256722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2292_n 0.00698438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2293_n 0.00947199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2294_n 0.0365941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2295_n 0.00507461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2296_n 0.0577149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2297_n 0.00332923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2298_n 0.0222458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2299_n 0.00408091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2300_n 0.042635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2301_n 0.0049096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2302_n 0.0189086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2303_n 0.00471252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2304_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2305_n 0.0165213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2306_n 0.0559261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2307_n 0.0230523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2308_n 0.622858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2309_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2310_n 0.00436942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2311_n 0.00597188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_143 VPB N_CLK_c_275_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_144 VPB N_CLK_c_279_n 0.0162092f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_145 VPB N_CLK_c_280_n 0.01861f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_146 VPB N_CLK_c_281_n 0.0230979f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_147 VPB CLK 0.0175757f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_148 VPB N_A_27_47#_M1000_g 0.0377949f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_149 VPB N_A_27_47#_M1016_g 0.0194267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_27_47#_M1025_g 0.033317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_27_47#_c_317_n 0.0198419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_27_47#_c_332_n 0.0018131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_27_47#_c_321_n 0.00333071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_27_47#_c_324_n 0.00290992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_27_47#_c_335_n 0.00357396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_27_47#_c_336_n 0.030972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_27_47#_c_337_n 0.00167507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_27_47#_c_338_n 0.0139626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_27_47#_c_339_n 9.75121e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_27_47#_c_340_n 0.00779662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_27_47#_c_341_n 0.0048201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_27_47#_c_325_n 0.0117983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_27_47#_c_343_n 0.0276115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_27_47#_c_326_n 0.0212228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_27_47#_c_327_n 0.00662783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_D_M1029_g 0.0238916f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_167 VPB N_D_c_595_n 0.0159446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB D 0.00181411f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_169 VPB N_D_c_593_n 0.0165468f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_170 VPB N_A_423_343#_c_647_n 0.0753975f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_171 VPB N_A_423_343#_c_648_n 0.0076426f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_172 VPB N_A_423_343#_c_643_n 0.00615569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_DE_c_733_n 0.0104063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_DE_M1011_g 0.0255037f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_175 VPB N_DE_c_738_n 0.0220855f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_176 VPB N_DE_M1015_g 0.0236724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_DE_c_740_n 0.00456175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB DE 0.00246649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_791_264#_M1041_g 8.35311e-19 $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_180 VPB N_A_791_264#_M1036_g 0.0220687f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_181 VPB N_A_791_264#_M1007_g 0.0241837f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_182 VPB N_A_791_264#_M1001_g 0.0184691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_791_264#_c_827_n 0.011879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_791_264#_c_828_n 0.040689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_791_264#_c_829_n 0.00761748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_791_264#_c_830_n 0.00659101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_791_264#_c_831_n 0.0286821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_791_264#_c_832_n 0.00248001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_791_264#_c_820_n 6.77134e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_791_264#_c_822_n 0.00225466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_885_21#_M1030_g 0.0202861f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_192 VPB N_A_885_21#_c_1009_n 0.00284214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_885_21#_c_1015_n 0.00513925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_885_21#_c_1010_n 0.00161367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_885_21#_c_1011_n 0.0191218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_885_21#_c_1018_n 0.00825295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_SCD_M1020_g 0.0202451f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_198 VPB SCD 0.00341946f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_199 VPB N_SCD_c_1133_n 0.016157f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_SCE_M1013_g 0.0280489f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_201 VPB N_SCE_c_1179_n 0.0191123f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_202 VPB N_SCE_c_1188_n 0.00795493f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_203 VPB N_SCE_M1033_g 0.0311924f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_204 VPB N_SCE_c_1184_n 0.00279238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_SCE_c_1185_n 0.0246671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_193_47#_M1008_g 0.0441742f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_207 VPB N_A_193_47#_c_1273_n 0.0138415f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_208 VPB N_A_193_47#_M1018_g 0.0210318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_193_47#_c_1285_n 0.0413295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_193_47#_c_1286_n 0.00566519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_A_193_47#_c_1287_n 0.0211513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_193_47#_c_1288_n 0.00119312f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_193_47#_c_1278_n 0.00673154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_193_47#_c_1279_n 0.0140385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_A_193_47#_c_1280_n 0.00152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_193_47#_c_1292_n 0.0265183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_193_47#_c_1281_n 0.00945279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_1610_159#_M1006_g 0.0519779f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_219 VPB N_A_1610_159#_M1037_g 0.0564064f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_220 VPB N_A_1610_159#_c_1493_n 0.00955004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1610_159#_c_1494_n 0.00154645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_1610_159#_c_1504_n 0.0154933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1610_159#_c_1496_n 0.00366659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1446_413#_M1017_g 0.0274355f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_225 VPB N_A_1446_413#_c_1610_n 0.018904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1446_413#_c_1611_n 0.0102534f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1446_413#_c_1617_n 0.00394568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1446_413#_c_1613_n 0.00924579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_2051_413#_M1023_g 0.0451789f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_230 VPB N_A_2051_413#_c_1714_n 0.00439136f $X=-0.19 $Y=1.305 $X2=0.33
+ $Y2=1.16
cc_231 VPB N_A_2051_413#_M1010_g 0.0237506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_2051_413#_c_1716_n 0.0157863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_2051_413#_c_1717_n 3.18387e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_2051_413#_c_1718_n 8.89166e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_2051_413#_c_1728_n 0.00704026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_2051_413#_c_1720_n 0.00292829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1824_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1825_n 0.00843162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1826_n 0.00704186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1827_n 0.0029826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1828_n 0.00505269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1829_n 0.0192928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1830_n 0.00629264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1831_n 0.00924361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1832_n 0.010598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1833_n 0.0365367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1834_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1835_n 0.0432692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1836_n 0.00497475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1837_n 0.0224066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1838_n 0.00468329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1839_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1840_n 0.0193581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1841_n 0.0595987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1842_n 0.0622872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1843_n 0.0230248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1823_n 0.0756964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1845_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1846_n 0.00372488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1847_n 0.00550927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1848_n 0.00449095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1849_n 0.00442865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_A_299_47#_c_2016_n 0.00772563f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_A_299_47#_c_2009_n 0.00994696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_A_299_47#_c_2018_n 0.00164603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_A_299_47#_c_2010_n 0.0037017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_A_915_47#_c_2138_n 0.00236345f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_268 VPB N_A_915_47#_c_2139_n 0.00246853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_A_915_47#_c_2140_n 0.00256118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_A_915_47#_c_2132_n 0.00506969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_A_915_47#_c_2134_n 0.00653972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_Q_c_2269_n 0.0436448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 N_CLK_c_275_n N_A_27_47#_M1021_g 0.00520193f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_274 N_CLK_c_276_n N_A_27_47#_M1021_g 0.0200589f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_275 CLK N_A_27_47#_M1021_g 3.12184e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_276 N_CLK_c_279_n N_A_27_47#_M1000_g 0.00541775f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_277 N_CLK_c_281_n N_A_27_47#_M1000_g 0.0276441f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_278 CLK N_A_27_47#_M1000_g 5.77812e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_279 N_CLK_c_275_n N_A_27_47#_c_319_n 0.00775742f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_280 N_CLK_c_276_n N_A_27_47#_c_319_n 0.00684762f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_281 CLK N_A_27_47#_c_319_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_282 N_CLK_c_275_n N_A_27_47#_c_320_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_283 CLK N_A_27_47#_c_320_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_284 N_CLK_c_280_n N_A_27_47#_c_332_n 0.0126874f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_285 N_CLK_c_281_n N_A_27_47#_c_332_n 0.00142281f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_286 CLK N_A_27_47#_c_332_n 0.00766156f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_287 N_CLK_c_275_n N_A_27_47#_c_321_n 0.0046428f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_288 N_CLK_c_279_n N_A_27_47#_c_321_n 7.07325e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_289 N_CLK_c_281_n N_A_27_47#_c_321_n 0.00436768f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_290 CLK N_A_27_47#_c_321_n 0.0511211f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_291 N_CLK_c_275_n N_A_27_47#_c_335_n 2.46885e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_292 N_CLK_c_280_n N_A_27_47#_c_335_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_293 N_CLK_c_281_n N_A_27_47#_c_335_n 0.00343236f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_294 CLK N_A_27_47#_c_335_n 0.0153591f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_295 N_CLK_c_280_n N_A_27_47#_c_337_n 0.00101286f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_296 N_CLK_c_275_n N_A_27_47#_c_325_n 0.0169118f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_297 CLK N_A_27_47#_c_325_n 0.00161603f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_298 N_CLK_c_280_n N_VPWR_c_1824_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_299 N_CLK_c_280_n N_VPWR_c_1839_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_300 N_CLK_c_280_n N_VPWR_c_1823_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_301 N_CLK_c_276_n N_VGND_c_2286_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_302 N_CLK_c_275_n N_VGND_c_2304_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_303 N_CLK_c_276_n N_VGND_c_2304_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_304 N_CLK_c_276_n N_VGND_c_2308_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_336_n N_D_M1029_g 0.00440395f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_306 N_A_27_47#_M1021_g N_D_c_591_n 0.00269191f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_307 N_A_27_47#_M1000_g N_D_c_595_n 0.00269191f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_336_n N_D_c_595_n 0.00153919f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_309 N_A_27_47#_c_336_n D 0.00497736f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_325_n N_D_c_593_n 0.00269191f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_336_n N_A_423_343#_c_647_n 0.0120018f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_336_n N_A_423_343#_c_648_n 0.0221661f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_336_n N_A_423_343#_c_643_n 0.00660521f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_336_n N_DE_M1011_g 0.00347932f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_315 N_A_27_47#_c_336_n N_DE_c_738_n 0.00132678f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_336_n N_DE_M1015_g 0.00575563f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_336_n N_A_791_264#_M1036_g 0.00424046f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_M1028_g N_A_791_264#_M1001_g 0.0443098f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_319 N_A_27_47#_c_336_n N_A_791_264#_c_830_n 0.00923372f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_336_n N_A_791_264#_c_831_n 0.00184708f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_M1028_g N_A_791_264#_c_818_n 0.00644693f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_c_322_n N_A_791_264#_c_818_n 0.0282618f $X=7.45 $Y=0.845 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_323_n N_A_791_264#_c_818_n 0.00156973f $X=7.28 $Y=0.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_326_n N_A_791_264#_c_818_n 8.58822e-19 $X=10.175 $Y=1.32
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_c_327_n N_A_791_264#_c_818_n 0.00521916f $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_326 N_A_27_47#_c_336_n N_A_885_21#_M1030_g 0.00250115f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_336_n N_A_885_21#_c_1009_n 0.00420661f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_336_n N_A_885_21#_c_1015_n 0.037101f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_336_n N_A_885_21#_c_1010_n 0.00530575f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_336_n N_A_885_21#_c_1011_n 3.31125e-19 $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_336_n N_A_885_21#_c_1018_n 0.0213362f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_336_n N_SCD_M1020_g 0.00142656f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_336_n SCD 0.00313621f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_334 N_A_27_47#_c_336_n N_SCD_c_1133_n 0.00198823f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_335 N_A_27_47#_c_336_n N_SCE_M1013_g 0.00338943f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_336 N_A_27_47#_c_336_n N_SCE_c_1179_n 9.29246e-19 $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_337 N_A_27_47#_c_336_n N_SCE_M1033_g 5.07716e-19 $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_338 N_A_27_47#_c_336_n N_SCE_c_1184_n 0.00477001f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_339 N_A_27_47#_c_336_n N_A_193_47#_M1000_d 0.00126326f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_324_n N_A_193_47#_M1008_g 7.3078e-19 $X=7.535 $Y=1.655 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_336_n N_A_193_47#_M1008_g 0.00621666f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_340_n N_A_193_47#_M1008_g 0.00238373f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_343_n N_A_193_47#_M1008_g 0.0270669f $X=7.705 $Y=1.74 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_324_n N_A_193_47#_c_1273_n 0.0120754f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_340_n N_A_193_47#_c_1273_n 0.00149465f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_c_343_n N_A_193_47#_c_1273_n 0.018371f $X=7.705 $Y=1.74 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_M1027_g N_A_193_47#_M1012_g 0.0124733f $X=7.29 $Y=0.415 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_322_n N_A_193_47#_M1012_g 0.00145899f $X=7.45 $Y=0.845 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_323_n N_A_193_47#_M1012_g 0.0168195f $X=7.28 $Y=0.87 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_324_n N_A_193_47#_M1012_g 0.00509325f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_M1028_g N_A_193_47#_c_1275_n 0.0144865f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_M1025_g N_A_193_47#_M1018_g 0.0175064f $X=10.18 $Y=2.275 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_M1028_g N_A_193_47#_c_1276_n 0.00658103f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_326_n N_A_193_47#_c_1276_n 9.61914e-19 $X=10.175 $Y=1.32
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_M1028_g N_A_193_47#_c_1277_n 0.0213226f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_326_n N_A_193_47#_c_1277_n 0.0204217f $X=10.175 $Y=1.32
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_c_327_n N_A_193_47#_c_1277_n 5.64291e-19 $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_c_336_n N_A_193_47#_c_1285_n 0.459939f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_M1000_g N_A_193_47#_c_1286_n 0.00457449f $X=0.89 $Y=2.135
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_c_321_n N_A_193_47#_c_1286_n 0.00673509f $X=0.76 $Y=1.235
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_336_n N_A_193_47#_c_1286_n 0.0262177f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_317_n N_A_193_47#_c_1287_n 0.00218822f $X=10.735 $Y=1.32
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_322_n N_A_193_47#_c_1287_n 0.00220528f $X=7.45 $Y=0.845
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_324_n N_A_193_47#_c_1287_n 0.0122906f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_336_n N_A_193_47#_c_1287_n 0.00995021f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_338_n N_A_193_47#_c_1287_n 0.185323f $X=10.04 $Y=1.87 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_339_n N_A_193_47#_c_1287_n 0.0254049f $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_340_n N_A_193_47#_c_1287_n 0.00659382f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_341_n N_A_193_47#_c_1287_n 0.026031f $X=10.185 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_343_n N_A_193_47#_c_1287_n 0.00183443f $X=7.705 $Y=1.74
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_326_n N_A_193_47#_c_1287_n 0.00372733f $X=10.175 $Y=1.32
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_327_n N_A_193_47#_c_1287_n 0.0147985f $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_322_n N_A_193_47#_c_1288_n 0.00129557f $X=7.45 $Y=0.845
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_324_n N_A_193_47#_c_1288_n 0.00254764f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_336_n N_A_193_47#_c_1288_n 0.0267692f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_327_n N_A_193_47#_c_1331_n 6.47753e-19 $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_M1025_g N_A_193_47#_c_1278_n 0.0020271f $X=10.18 $Y=2.275
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_317_n N_A_193_47#_c_1278_n 0.0169581f $X=10.735 $Y=1.32
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_M1028_g N_A_193_47#_c_1278_n 0.00640774f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_341_n N_A_193_47#_c_1278_n 0.00821717f $X=10.185 $Y=1.87
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_326_n N_A_193_47#_c_1278_n 0.00345899f $X=10.175 $Y=1.32
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_327_n N_A_193_47#_c_1278_n 0.051449f $X=10.175 $Y=1.41 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_322_n N_A_193_47#_c_1279_n 0.00116173f $X=7.45 $Y=0.845
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_323_n N_A_193_47#_c_1279_n 0.0213517f $X=7.28 $Y=0.87 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_324_n N_A_193_47#_c_1279_n 0.00139632f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_336_n N_A_193_47#_c_1279_n 5.87167e-19 $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_322_n N_A_193_47#_c_1280_n 0.0115307f $X=7.45 $Y=0.845 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_323_n N_A_193_47#_c_1280_n 0.00111596f $X=7.28 $Y=0.87 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_324_n N_A_193_47#_c_1280_n 0.0369678f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_336_n N_A_193_47#_c_1280_n 0.00453285f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_340_n N_A_193_47#_c_1280_n 0.00526954f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_343_n N_A_193_47#_c_1280_n 3.45729e-19 $X=7.705 $Y=1.74
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_M1025_g N_A_193_47#_c_1292_n 0.0130792f $X=10.18 $Y=2.275
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_317_n N_A_193_47#_c_1292_n 0.0224153f $X=10.735 $Y=1.32
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_327_n N_A_193_47#_c_1292_n 6.57469e-19 $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_M1021_g N_A_193_47#_c_1281_n 0.0188272f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_319_n N_A_193_47#_c_1281_n 0.0127744f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_464_p N_A_193_47#_c_1281_n 0.00850019f $X=0.73 $Y=1.795
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_321_n N_A_193_47#_c_1281_n 0.0695916f $X=0.76 $Y=1.235 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_336_n N_A_193_47#_c_1281_n 0.0124318f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_337_n N_A_193_47#_c_1281_n 0.00241841f $X=0.865 $Y=1.87
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_M1016_g N_A_1610_159#_M1006_g 0.0243723f $X=7.61 $Y=2.275
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_324_n N_A_1610_159#_M1006_g 0.00146118f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_338_n N_A_1610_159#_M1006_g 0.0013651f $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_340_n N_A_1610_159#_M1006_g 0.00196903f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_343_n N_A_1610_159#_M1006_g 0.0206078f $X=7.705 $Y=1.74
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_M1025_g N_A_1610_159#_M1037_g 0.0428173f $X=10.18 $Y=2.275
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_338_n N_A_1610_159#_M1037_g 0.00780647f $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_341_n N_A_1610_159#_M1037_g 0.00131932f $X=10.185 $Y=1.87
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_327_n N_A_1610_159#_M1037_g 0.00605027f $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_326_n N_A_1610_159#_c_1493_n 0.0189308f $X=10.175 $Y=1.32
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_327_n N_A_1610_159#_c_1493_n 0.00198129f $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_338_n N_A_1610_159#_c_1504_n 0.0261908f $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_326_n N_A_1610_159#_c_1496_n 5.17694e-19 $X=10.175 $Y=1.32
+ $X2=0 $Y2=0
cc_415 N_A_27_47#_c_327_n N_A_1610_159#_c_1496_n 0.00546887f $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_338_n N_A_1446_413#_M1017_g 0.00324412f $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_417 N_A_27_47#_c_338_n N_A_1446_413#_c_1610_n 2.40114e-19 $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_418 N_A_27_47#_M1016_g N_A_1446_413#_c_1621_n 0.00947181f $X=7.61 $Y=2.275
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_c_336_n N_A_1446_413#_c_1621_n 0.00579806f $X=7.45 $Y=1.87
+ $X2=0 $Y2=0
cc_420 N_A_27_47#_c_338_n N_A_1446_413#_c_1621_n 0.0054742f $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_c_339_n N_A_1446_413#_c_1621_n 0.00117338f $X=7.74 $Y=1.87
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_340_n N_A_1446_413#_c_1621_n 0.0279213f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_343_n N_A_1446_413#_c_1621_n 7.4902e-19 $X=7.705 $Y=1.74
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_M1027_g N_A_1446_413#_c_1627_n 0.00529747f $X=7.29 $Y=0.415
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_c_322_n N_A_1446_413#_c_1627_n 0.0197321f $X=7.45 $Y=0.845
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_323_n N_A_1446_413#_c_1627_n 0.00160367f $X=7.28 $Y=0.87
+ $X2=0 $Y2=0
cc_427 N_A_27_47#_c_322_n N_A_1446_413#_c_1612_n 0.0151383f $X=7.45 $Y=0.845
+ $X2=0 $Y2=0
cc_428 N_A_27_47#_c_324_n N_A_1446_413#_c_1612_n 0.024597f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_M1016_g N_A_1446_413#_c_1617_n 0.00104479f $X=7.61 $Y=2.275
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_324_n N_A_1446_413#_c_1617_n 0.00207816f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_338_n N_A_1446_413#_c_1617_n 0.0129147f $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_339_n N_A_1446_413#_c_1617_n 4.13019e-19 $X=7.74 $Y=1.87
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_340_n N_A_1446_413#_c_1617_n 0.0255803f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_c_343_n N_A_1446_413#_c_1617_n 6.18409e-19 $X=7.705 $Y=1.74
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_324_n N_A_1446_413#_c_1613_n 0.0144717f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_338_n N_A_1446_413#_c_1613_n 0.00326146f $X=10.04 $Y=1.87
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_340_n N_A_1446_413#_c_1613_n 0.00725124f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_343_n N_A_1446_413#_c_1613_n 5.89706e-19 $X=7.705 $Y=1.74
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_M1025_g N_A_2051_413#_c_1730_n 0.00428769f $X=10.18 $Y=2.275
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_341_n N_A_2051_413#_c_1730_n 0.0021332f $X=10.185 $Y=1.87
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_327_n N_A_2051_413#_c_1730_n 0.00225822f $X=10.175 $Y=1.41
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_M1028_g N_A_2051_413#_c_1733_n 0.0121553f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_M1028_g N_A_2051_413#_c_1719_n 0.00499822f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_317_n N_A_2051_413#_c_1728_n 6.71564e-19 $X=10.735 $Y=1.32
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_M1028_g N_A_2051_413#_c_1721_n 0.00301916f $X=10.81 $Y=0.415
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_464_p N_VPWR_M1014_d 6.67509e-19 $X=0.73 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_447 N_A_27_47#_c_337_n N_VPWR_M1014_d 0.00178771f $X=0.865 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_448 N_A_27_47#_c_336_n N_VPWR_M1011_d 0.00132004f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_338_n N_VPWR_M1006_d 0.00515584f $X=10.04 $Y=1.87 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_M1000_g N_VPWR_c_1824_n 0.00944765f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_332_n N_VPWR_c_1824_n 0.00346278f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_464_p N_VPWR_c_1824_n 0.013292f $X=0.73 $Y=1.795 $X2=0 $Y2=0
cc_453 N_A_27_47#_c_335_n N_VPWR_c_1824_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_454 N_A_27_47#_c_337_n N_VPWR_c_1824_n 0.003216f $X=0.865 $Y=1.87 $X2=0 $Y2=0
cc_455 N_A_27_47#_c_336_n N_VPWR_c_1825_n 0.0177398f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_456 N_A_27_47#_c_336_n N_VPWR_c_1826_n 0.0144415f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_457 N_A_27_47#_c_336_n N_VPWR_c_1827_n 0.00158709f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_338_n N_VPWR_c_1828_n 0.0124077f $X=10.04 $Y=1.87 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_M1025_g N_VPWR_c_1830_n 0.00239883f $X=10.18 $Y=2.275 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_338_n N_VPWR_c_1830_n 0.010979f $X=10.04 $Y=1.87 $X2=0 $Y2=0
cc_461 N_A_27_47#_M1000_g N_VPWR_c_1833_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_M1025_g N_VPWR_c_1835_n 0.00429356f $X=10.18 $Y=2.275 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_327_n N_VPWR_c_1835_n 0.00157744f $X=10.175 $Y=1.41 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_332_n N_VPWR_c_1839_n 0.0018545f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_335_n N_VPWR_c_1839_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_466 N_A_27_47#_M1016_g N_VPWR_c_1842_n 0.00375986f $X=7.61 $Y=2.275 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_M1000_g N_VPWR_c_1823_n 0.00534571f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_M1016_g N_VPWR_c_1823_n 0.00556927f $X=7.61 $Y=2.275 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_M1025_g N_VPWR_c_1823_n 0.00573395f $X=10.18 $Y=2.275 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_332_n N_VPWR_c_1823_n 0.00404038f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_335_n N_VPWR_c_1823_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_336_n N_VPWR_c_1823_n 0.311577f $X=7.45 $Y=1.87 $X2=0 $Y2=0
cc_473 N_A_27_47#_c_337_n N_VPWR_c_1823_n 0.0145601f $X=0.865 $Y=1.87 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_338_n N_VPWR_c_1823_n 0.11007f $X=10.04 $Y=1.87 $X2=0 $Y2=0
cc_475 N_A_27_47#_c_339_n N_VPWR_c_1823_n 0.0144472f $X=7.74 $Y=1.87 $X2=0 $Y2=0
cc_476 N_A_27_47#_c_341_n N_VPWR_c_1823_n 0.0159851f $X=10.185 $Y=1.87 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_327_n N_VPWR_c_1823_n 0.00101559f $X=10.175 $Y=1.41 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_336_n N_A_299_47#_c_2016_n 0.020151f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_336_n N_A_299_47#_c_2009_n 0.00810658f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_c_336_n N_A_299_47#_c_2018_n 0.0217319f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_336_n N_A_299_47#_c_2010_n 0.00317487f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_M1021_g N_A_299_47#_c_2015_n 0.00143698f $X=0.89 $Y=0.445
+ $X2=0 $Y2=0
cc_483 N_A_27_47#_c_336_n A_381_369# 0.00298073f $X=7.45 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_484 N_A_27_47#_c_336_n A_729_369# 0.00510983f $X=7.45 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_485 N_A_27_47#_c_336_n N_A_915_47#_M1013_d 6.61893e-19 $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_336_n N_A_915_47#_M1030_d 0.00115845f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_336_n N_A_915_47#_c_2138_n 0.0107002f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_336_n N_A_915_47#_c_2139_n 0.00859404f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_M1027_g N_A_915_47#_c_2130_n 0.00568611f $X=7.29 $Y=0.415
+ $X2=0 $Y2=0
cc_490 N_A_27_47#_c_322_n N_A_915_47#_c_2130_n 0.0143216f $X=7.45 $Y=0.845 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_c_323_n N_A_915_47#_c_2130_n 0.00163085f $X=7.28 $Y=0.87 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_324_n N_A_915_47#_c_2130_n 0.00612681f $X=7.535 $Y=1.655
+ $X2=0 $Y2=0
cc_493 N_A_27_47#_c_336_n N_A_915_47#_c_2151_n 0.0129167f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_339_n N_A_915_47#_c_2151_n 3.14279e-19 $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_340_n N_A_915_47#_c_2151_n 0.00378437f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_496 N_A_27_47#_c_336_n N_A_915_47#_c_2140_n 0.0014312f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_336_n N_A_915_47#_c_2155_n 0.00255293f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_c_336_n N_A_915_47#_c_2134_n 0.00590396f $X=7.45 $Y=1.87 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_339_n N_A_915_47#_c_2134_n 2.89444e-19 $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_340_n N_A_915_47#_c_2134_n 0.00358872f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_501 N_A_27_47#_M1027_g N_A_915_47#_c_2137_n 0.00683036f $X=7.29 $Y=0.415
+ $X2=0 $Y2=0
cc_502 N_A_27_47#_c_322_n N_A_915_47#_c_2137_n 0.00131254f $X=7.45 $Y=0.845
+ $X2=0 $Y2=0
cc_503 N_A_27_47#_c_323_n N_A_915_47#_c_2137_n 4.36817e-19 $X=7.28 $Y=0.87 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_c_319_n N_VGND_M1040_d 0.00164502f $X=0.615 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_505 N_A_27_47#_M1021_g N_VGND_c_2286_n 0.0090859f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_c_319_n N_VGND_c_2286_n 0.0172929f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_325_n N_VGND_c_2286_n 5.70216e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_M1028_g N_VGND_c_2292_n 0.00155843f $X=10.81 $Y=0.415 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_M1021_g N_VGND_c_2294_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_M1028_g N_VGND_c_2300_n 0.00373071f $X=10.81 $Y=0.415 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_c_577_p N_VGND_c_2304_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_512 N_A_27_47#_c_319_n N_VGND_c_2304_n 0.00243651f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_M1027_g N_VGND_c_2306_n 0.00406674f $X=7.29 $Y=0.415 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_322_n N_VGND_c_2306_n 0.00226614f $X=7.45 $Y=0.845 $X2=0
+ $Y2=0
cc_515 N_A_27_47#_c_323_n N_VGND_c_2306_n 0.00108996f $X=7.28 $Y=0.87 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_M1040_s N_VGND_c_2308_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_M1021_g N_VGND_c_2308_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_518 N_A_27_47#_M1027_g N_VGND_c_2308_n 0.00693963f $X=7.29 $Y=0.415 $X2=0
+ $Y2=0
cc_519 N_A_27_47#_M1028_g N_VGND_c_2308_n 0.00568812f $X=10.81 $Y=0.415 $X2=0
+ $Y2=0
cc_520 N_A_27_47#_c_577_p N_VGND_c_2308_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_c_319_n N_VGND_c_2308_n 0.00580457f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_322_n N_VGND_c_2308_n 0.00188658f $X=7.45 $Y=0.845 $X2=0
+ $Y2=0
cc_523 N_A_27_47#_c_323_n N_VGND_c_2308_n 0.0011282f $X=7.28 $Y=0.87 $X2=0 $Y2=0
cc_524 N_D_M1029_g N_A_423_343#_c_647_n 0.059369f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_525 N_D_c_595_n N_A_423_343#_c_647_n 0.00202148f $X=1.765 $Y=1.65 $X2=0 $Y2=0
cc_526 D N_A_423_343#_c_647_n 0.00175679f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_527 N_D_c_593_n N_A_423_343#_c_647_n 0.00564261f $X=1.78 $Y=1.145 $X2=0 $Y2=0
cc_528 D N_A_423_343#_c_643_n 0.00775821f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_529 N_D_c_593_n N_A_423_343#_c_643_n 0.00112085f $X=1.78 $Y=1.145 $X2=0 $Y2=0
cc_530 N_D_M1002_g N_DE_M1003_g 0.0501357f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_531 D N_DE_M1003_g 3.59802e-19 $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_532 N_D_M1002_g N_DE_c_731_n 0.00609422f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_533 N_D_c_591_n N_DE_c_731_n 0.0121267f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_534 D N_DE_c_731_n 5.46011e-19 $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_535 N_D_M1002_g DE 7.68806e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_536 N_D_c_591_n DE 0.00538864f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_537 D DE 0.0433254f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_538 N_D_c_595_n N_A_193_47#_c_1285_n 0.00238342f $X=1.765 $Y=1.65 $X2=0 $Y2=0
cc_539 D N_A_193_47#_c_1285_n 0.0215563f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_540 N_D_c_593_n N_A_193_47#_c_1285_n 0.00384385f $X=1.78 $Y=1.145 $X2=0 $Y2=0
cc_541 N_D_M1029_g N_VPWR_c_1825_n 0.00282543f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_542 N_D_M1029_g N_VPWR_c_1833_n 0.00541359f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_543 N_D_M1029_g N_VPWR_c_1823_n 0.00735355f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_544 N_D_M1029_g N_A_299_47#_c_2016_n 0.00949347f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_545 N_D_c_595_n N_A_299_47#_c_2016_n 0.00320688f $X=1.765 $Y=1.65 $X2=0 $Y2=0
cc_546 D N_A_299_47#_c_2016_n 0.00525464f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_547 N_D_M1002_g N_A_299_47#_c_2009_n 0.00738489f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_548 N_D_M1029_g N_A_299_47#_c_2009_n 0.00462667f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_549 N_D_c_591_n N_A_299_47#_c_2009_n 0.00752867f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_550 D N_A_299_47#_c_2009_n 0.0697065f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_551 N_D_M1002_g N_A_299_47#_c_2012_n 7.51093e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_552 N_D_M1002_g N_A_299_47#_c_2013_n 0.00320603f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_553 N_D_c_591_n N_A_299_47#_c_2013_n 0.00203556f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_554 D N_A_299_47#_c_2013_n 0.00827304f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_555 N_D_M1002_g N_A_299_47#_c_2015_n 0.00424642f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_556 N_D_c_591_n N_A_299_47#_c_2015_n 0.00228287f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_557 D N_A_299_47#_c_2015_n 0.00347931f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_558 N_D_M1002_g N_VGND_c_2287_n 0.00200661f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_559 N_D_M1002_g N_VGND_c_2294_n 0.00539883f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_560 N_D_M1002_g N_VGND_c_2308_n 0.00608889f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_561 N_A_423_343#_c_642_n N_DE_M1003_g 0.00526826f $X=2.92 $Y=0.51 $X2=0 $Y2=0
cc_562 N_A_423_343#_c_647_n N_DE_c_730_n 0.0080968f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_563 N_A_423_343#_c_643_n N_DE_c_730_n 0.005738f $X=2.932 $Y=1.355 $X2=0 $Y2=0
cc_564 N_A_423_343#_c_646_n N_DE_c_730_n 0.0178991f $X=2.932 $Y=1.01 $X2=0 $Y2=0
cc_565 N_A_423_343#_c_647_n N_DE_c_731_n 0.00919986f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_566 N_A_423_343#_c_646_n N_DE_c_731_n 6.99116e-19 $X=2.932 $Y=1.01 $X2=0
+ $Y2=0
cc_567 N_A_423_343#_M1022_g N_DE_M1038_g 0.0148047f $X=3.57 $Y=0.445 $X2=0 $Y2=0
cc_568 N_A_423_343#_c_642_n N_DE_M1038_g 0.00862574f $X=2.92 $Y=0.51 $X2=0 $Y2=0
cc_569 N_A_423_343#_c_644_n N_DE_M1038_g 0.00220234f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_570 N_A_423_343#_c_645_n N_DE_M1038_g 0.0213224f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_571 N_A_423_343#_c_646_n N_DE_M1038_g 5.67233e-19 $X=2.932 $Y=1.01 $X2=0
+ $Y2=0
cc_572 N_A_423_343#_c_647_n N_DE_c_733_n 0.0152313f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_573 N_A_423_343#_c_643_n N_DE_c_733_n 0.0179184f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_574 N_A_423_343#_c_644_n N_DE_c_733_n 0.00575309f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_575 N_A_423_343#_c_646_n N_DE_c_733_n 0.00317696f $X=2.932 $Y=1.01 $X2=0
+ $Y2=0
cc_576 N_A_423_343#_c_648_n N_DE_M1011_g 0.0105135f $X=2.92 $Y=1.99 $X2=0 $Y2=0
cc_577 N_A_423_343#_c_643_n N_DE_M1011_g 0.00362978f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_578 N_A_423_343#_c_644_n N_DE_c_738_n 0.00580736f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_579 N_A_423_343#_c_645_n N_DE_c_738_n 0.0122629f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_580 N_A_423_343#_c_648_n N_DE_M1015_g 8.04992e-19 $X=2.92 $Y=1.99 $X2=0 $Y2=0
cc_581 N_A_423_343#_c_643_n N_DE_M1015_g 5.26012e-19 $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_582 N_A_423_343#_c_644_n N_DE_c_734_n 0.00305763f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_583 N_A_423_343#_c_646_n N_DE_c_734_n 4.2374e-19 $X=2.932 $Y=1.01 $X2=0 $Y2=0
cc_584 N_A_423_343#_c_643_n N_DE_c_740_n 0.00610053f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_585 N_A_423_343#_c_647_n DE 0.00845936f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_586 N_A_423_343#_c_642_n DE 0.00561932f $X=2.92 $Y=0.51 $X2=0 $Y2=0
cc_587 N_A_423_343#_c_643_n DE 0.0143622f $X=2.932 $Y=1.355 $X2=0 $Y2=0
cc_588 N_A_423_343#_c_646_n DE 0.0240519f $X=2.932 $Y=1.01 $X2=0 $Y2=0
cc_589 N_A_423_343#_M1022_g N_A_791_264#_M1041_g 0.0251313f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_590 N_A_423_343#_c_645_n N_A_791_264#_M1041_g 0.0108934f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_591 N_A_423_343#_M1022_g N_A_791_264#_c_819_n 0.0021118f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_592 N_A_423_343#_c_644_n N_A_791_264#_c_819_n 0.00406567f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_593 N_A_423_343#_c_645_n N_A_791_264#_c_819_n 0.00242559f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_594 N_A_423_343#_M1022_g N_A_791_264#_c_820_n 0.00307938f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_595 N_A_423_343#_c_644_n N_A_791_264#_c_820_n 0.0248957f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_596 N_A_423_343#_c_645_n N_A_791_264#_c_820_n 0.00233652f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_597 N_A_423_343#_c_647_n N_A_193_47#_c_1285_n 0.00463103f $X=2.19 $Y=1.77
+ $X2=0 $Y2=0
cc_598 N_A_423_343#_c_648_n N_A_193_47#_c_1285_n 3.18139e-19 $X=2.92 $Y=1.99
+ $X2=0 $Y2=0
cc_599 N_A_423_343#_c_643_n N_A_193_47#_c_1285_n 0.0327297f $X=2.932 $Y=1.355
+ $X2=0 $Y2=0
cc_600 N_A_423_343#_c_644_n N_A_193_47#_c_1285_n 0.0177671f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_601 N_A_423_343#_c_645_n N_A_193_47#_c_1285_n 0.00228465f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_602 N_A_423_343#_c_647_n N_VPWR_c_1825_n 0.0251559f $X=2.19 $Y=1.77 $X2=0
+ $Y2=0
cc_603 N_A_423_343#_c_648_n N_VPWR_c_1825_n 0.0405714f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_604 N_A_423_343#_c_643_n N_VPWR_c_1825_n 0.00458578f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_605 N_A_423_343#_c_648_n N_VPWR_c_1826_n 0.0418939f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_606 N_A_423_343#_c_644_n N_VPWR_c_1826_n 0.00271398f $X=3.55 $Y=1.01 $X2=0
+ $Y2=0
cc_607 N_A_423_343#_c_647_n N_VPWR_c_1833_n 0.0046653f $X=2.19 $Y=1.77 $X2=0
+ $Y2=0
cc_608 N_A_423_343#_c_648_n N_VPWR_c_1840_n 0.0167964f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_609 N_A_423_343#_M1011_s N_VPWR_c_1823_n 0.00173907f $X=2.795 $Y=1.845 $X2=0
+ $Y2=0
cc_610 N_A_423_343#_c_647_n N_VPWR_c_1823_n 0.00430483f $X=2.19 $Y=1.77 $X2=0
+ $Y2=0
cc_611 N_A_423_343#_c_648_n N_VPWR_c_1823_n 0.00581267f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_612 N_A_423_343#_c_647_n N_A_299_47#_c_2016_n 0.00159809f $X=2.19 $Y=1.77
+ $X2=0 $Y2=0
cc_613 N_A_423_343#_M1022_g N_A_299_47#_c_2040_n 2.04373e-19 $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_614 N_A_423_343#_M1038_s N_A_299_47#_c_2013_n 6.77802e-19 $X=2.795 $Y=0.235
+ $X2=0 $Y2=0
cc_615 N_A_423_343#_M1022_g N_A_299_47#_c_2013_n 0.00414801f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_616 N_A_423_343#_c_642_n N_A_299_47#_c_2013_n 0.0183276f $X=2.92 $Y=0.51
+ $X2=0 $Y2=0
cc_617 N_A_423_343#_c_644_n N_A_299_47#_c_2013_n 0.0107001f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_618 N_A_423_343#_c_645_n N_A_299_47#_c_2013_n 9.48498e-19 $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_619 N_A_423_343#_c_646_n N_A_299_47#_c_2013_n 0.00351536f $X=2.932 $Y=1.01
+ $X2=0 $Y2=0
cc_620 N_A_423_343#_M1022_g N_A_299_47#_c_2014_n 0.00155158f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_621 N_A_423_343#_c_642_n N_VGND_c_2287_n 0.0164318f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_622 N_A_423_343#_M1022_g N_VGND_c_2288_n 0.0113899f $X=3.57 $Y=0.445 $X2=0
+ $Y2=0
cc_623 N_A_423_343#_c_642_n N_VGND_c_2288_n 0.0148662f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_624 N_A_423_343#_c_644_n N_VGND_c_2288_n 0.0151977f $X=3.55 $Y=1.01 $X2=0
+ $Y2=0
cc_625 N_A_423_343#_c_645_n N_VGND_c_2288_n 0.00159308f $X=3.55 $Y=1.01 $X2=0
+ $Y2=0
cc_626 N_A_423_343#_M1022_g N_VGND_c_2296_n 0.00505556f $X=3.57 $Y=0.445 $X2=0
+ $Y2=0
cc_627 N_A_423_343#_c_642_n N_VGND_c_2305_n 0.0154917f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_628 N_A_423_343#_M1038_s N_VGND_c_2308_n 0.00120778f $X=2.795 $Y=0.235 $X2=0
+ $Y2=0
cc_629 N_A_423_343#_M1022_g N_VGND_c_2308_n 0.00379888f $X=3.57 $Y=0.445 $X2=0
+ $Y2=0
cc_630 N_A_423_343#_c_642_n N_VGND_c_2308_n 0.00215984f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_631 N_DE_M1015_g N_A_791_264#_M1036_g 0.033024f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_632 N_DE_c_733_n N_A_791_264#_c_830_n 0.00334239f $X=3.13 $Y=1.46 $X2=0 $Y2=0
cc_633 N_DE_c_738_n N_A_791_264#_c_830_n 0.00386505f $X=3.495 $Y=1.535 $X2=0
+ $Y2=0
cc_634 N_DE_c_738_n N_A_791_264#_c_831_n 0.00786818f $X=3.495 $Y=1.535 $X2=0
+ $Y2=0
cc_635 N_DE_c_733_n N_A_791_264#_c_820_n 0.00317814f $X=3.13 $Y=1.46 $X2=0 $Y2=0
cc_636 N_DE_c_738_n N_A_193_47#_c_1285_n 0.0079741f $X=3.495 $Y=1.535 $X2=0
+ $Y2=0
cc_637 N_DE_c_740_n N_A_193_47#_c_1285_n 0.00255711f $X=3.13 $Y=1.535 $X2=0
+ $Y2=0
cc_638 DE N_A_193_47#_c_1285_n 0.0181093f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_639 N_DE_M1011_g N_VPWR_c_1825_n 0.00292738f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_640 DE N_VPWR_c_1825_n 0.00131185f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_641 N_DE_M1011_g N_VPWR_c_1826_n 0.00567389f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_642 N_DE_c_738_n N_VPWR_c_1826_n 0.00241702f $X=3.495 $Y=1.535 $X2=0 $Y2=0
cc_643 N_DE_M1015_g N_VPWR_c_1826_n 0.00345066f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_644 N_DE_M1011_g N_VPWR_c_1840_n 0.00542953f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_645 N_DE_M1015_g N_VPWR_c_1841_n 0.00585385f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_646 N_DE_M1011_g N_VPWR_c_1823_n 0.00739796f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_647 N_DE_M1015_g N_VPWR_c_1823_n 0.00652437f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_648 N_DE_M1015_g N_A_299_47#_c_2018_n 0.00208296f $X=3.57 $Y=2.165 $X2=0
+ $Y2=0
cc_649 N_DE_M1003_g N_A_299_47#_c_2013_n 0.00328866f $X=2.19 $Y=0.445 $X2=0
+ $Y2=0
cc_650 N_DE_c_730_n N_A_299_47#_c_2013_n 0.00449574f $X=3.055 $Y=0.925 $X2=0
+ $Y2=0
cc_651 N_DE_M1038_g N_A_299_47#_c_2013_n 0.00212954f $X=3.13 $Y=0.445 $X2=0
+ $Y2=0
cc_652 DE N_A_299_47#_c_2013_n 0.014806f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_653 N_DE_M1003_g N_A_299_47#_c_2015_n 7.72933e-19 $X=2.19 $Y=0.445 $X2=0
+ $Y2=0
cc_654 N_DE_M1003_g N_VGND_c_2287_n 0.0103332f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_655 N_DE_c_730_n N_VGND_c_2287_n 5.49262e-19 $X=3.055 $Y=0.925 $X2=0 $Y2=0
cc_656 N_DE_c_731_n N_VGND_c_2287_n 9.86308e-19 $X=2.455 $Y=0.925 $X2=0 $Y2=0
cc_657 N_DE_M1038_g N_VGND_c_2287_n 0.00200593f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_658 DE N_VGND_c_2287_n 0.0147118f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_659 N_DE_M1038_g N_VGND_c_2288_n 0.00765346f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_660 N_DE_M1003_g N_VGND_c_2294_n 0.0046653f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_661 N_DE_M1038_g N_VGND_c_2305_n 0.00505556f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_662 N_DE_M1003_g N_VGND_c_2308_n 0.00313929f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_663 N_DE_M1038_g N_VGND_c_2308_n 0.00491778f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_664 N_A_791_264#_M1041_g N_A_885_21#_c_1002_n 0.0204071f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_665 N_A_791_264#_c_818_n N_A_885_21#_c_1003_n 0.00530549f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_666 N_A_791_264#_c_818_n N_A_885_21#_c_1004_n 0.00376476f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_667 N_A_791_264#_c_818_n N_A_885_21#_c_1006_n 0.00179302f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_668 N_A_791_264#_c_818_n N_A_885_21#_c_1010_n 0.0032108f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_669 N_A_791_264#_c_818_n N_A_885_21#_c_1012_n 0.0218496f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_670 N_A_791_264#_c_818_n N_SCD_M1024_g 0.00331392f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_671 N_A_791_264#_c_818_n SCD 0.00963209f $X=11.94 $Y=0.85 $X2=0 $Y2=0
cc_672 N_A_791_264#_M1036_g N_SCE_M1013_g 0.0130813f $X=4.08 $Y=2.165 $X2=0
+ $Y2=0
cc_673 N_A_791_264#_c_830_n N_SCE_c_1188_n 2.77563e-19 $X=4.09 $Y=1.485 $X2=0
+ $Y2=0
cc_674 N_A_791_264#_c_831_n N_SCE_c_1188_n 0.0124712f $X=4.09 $Y=1.485 $X2=0
+ $Y2=0
cc_675 N_A_791_264#_c_818_n N_SCE_c_1188_n 0.00151081f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_676 N_A_791_264#_c_818_n N_SCE_M1005_g 0.00275998f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_677 N_A_791_264#_c_818_n N_SCE_M1009_g 0.00395652f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_678 N_A_791_264#_c_818_n N_SCE_c_1184_n 0.00399796f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_679 N_A_791_264#_c_818_n N_SCE_c_1185_n 5.58043e-19 $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_680 N_A_791_264#_c_818_n N_A_193_47#_c_1273_n 4.65473e-19 $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_681 N_A_791_264#_c_818_n N_A_193_47#_M1012_g 0.00493455f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_682 N_A_791_264#_c_828_n N_A_193_47#_M1018_g 0.0199779f $X=11.365 $Y=1.74
+ $X2=0 $Y2=0
cc_683 N_A_791_264#_M1001_g N_A_193_47#_c_1276_n 3.66194e-19 $X=11.285 $Y=0.445
+ $X2=0 $Y2=0
cc_684 N_A_791_264#_c_818_n N_A_193_47#_c_1276_n 0.0311489f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_685 N_A_791_264#_c_818_n N_A_193_47#_c_1277_n 0.00343724f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_686 N_A_791_264#_c_830_n N_A_193_47#_c_1285_n 0.0212f $X=4.09 $Y=1.485 $X2=0
+ $Y2=0
cc_687 N_A_791_264#_c_831_n N_A_193_47#_c_1285_n 0.00126879f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_688 N_A_791_264#_c_818_n N_A_193_47#_c_1285_n 0.128587f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_689 N_A_791_264#_c_819_n N_A_193_47#_c_1285_n 0.013239f $X=4.035 $Y=0.85
+ $X2=0 $Y2=0
cc_690 N_A_791_264#_c_820_n N_A_193_47#_c_1285_n 3.15466e-19 $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_691 N_A_791_264#_c_818_n N_A_193_47#_c_1287_n 0.132905f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_692 N_A_791_264#_c_818_n N_A_193_47#_c_1288_n 0.0130915f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_693 N_A_791_264#_c_818_n N_A_193_47#_c_1331_n 0.012252f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_694 N_A_791_264#_c_828_n N_A_193_47#_c_1278_n 7.03497e-19 $X=11.365 $Y=1.74
+ $X2=0 $Y2=0
cc_695 N_A_791_264#_c_818_n N_A_193_47#_c_1279_n 0.00127009f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_696 N_A_791_264#_c_818_n N_A_193_47#_c_1280_n 0.00111342f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_697 N_A_791_264#_c_828_n N_A_193_47#_c_1292_n 0.0137111f $X=11.365 $Y=1.74
+ $X2=0 $Y2=0
cc_698 N_A_791_264#_c_818_n N_A_1610_159#_M1039_g 0.00577171f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_699 N_A_791_264#_c_818_n N_A_1610_159#_c_1492_n 0.00619242f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_700 N_A_791_264#_c_818_n N_A_1610_159#_c_1494_n 0.0564626f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_701 N_A_791_264#_c_818_n N_A_1610_159#_c_1496_n 0.012477f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_702 N_A_791_264#_c_818_n N_A_1610_159#_c_1498_n 0.0112362f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_703 N_A_791_264#_c_818_n N_A_1610_159#_c_1499_n 0.00300444f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_704 N_A_791_264#_c_818_n N_A_1446_413#_c_1627_n 0.00659708f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_705 N_A_791_264#_c_818_n N_A_1446_413#_c_1612_n 0.0152331f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_706 N_A_791_264#_c_818_n N_A_1446_413#_c_1613_n 0.00619733f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_707 N_A_791_264#_c_816_n N_A_2051_413#_M1031_g 0.00561498f $X=12.015 $Y=0.385
+ $X2=0 $Y2=0
cc_708 N_A_791_264#_c_817_n N_A_2051_413#_M1031_g 0.00477121f $X=12.015 $Y=0.825
+ $X2=0 $Y2=0
cc_709 N_A_791_264#_c_821_n N_A_2051_413#_M1031_g 0.00517962f $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_710 N_A_791_264#_c_822_n N_A_2051_413#_M1031_g 0.0052888f $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_711 N_A_791_264#_c_828_n N_A_2051_413#_M1023_g 0.00345271f $X=11.365 $Y=1.74
+ $X2=0 $Y2=0
cc_712 N_A_791_264#_c_829_n N_A_2051_413#_M1023_g 0.00613006f $X=12.005 $Y=1.99
+ $X2=0 $Y2=0
cc_713 N_A_791_264#_c_832_n N_A_2051_413#_M1023_g 0.0104703f $X=12.01 $Y=1.717
+ $X2=0 $Y2=0
cc_714 N_A_791_264#_c_822_n N_A_2051_413#_M1023_g 0.00721223f $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_715 N_A_791_264#_c_816_n N_A_2051_413#_c_1715_n 5.51494e-19 $X=12.015
+ $Y=0.385 $X2=0 $Y2=0
cc_716 N_A_791_264#_c_821_n N_A_2051_413#_c_1715_n 3.16115e-19 $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_717 N_A_791_264#_c_822_n N_A_2051_413#_M1010_g 4.45214e-19 $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_718 N_A_791_264#_M1001_g N_A_2051_413#_c_1716_n 0.0191523f $X=11.285 $Y=0.445
+ $X2=0 $Y2=0
cc_719 N_A_791_264#_c_827_n N_A_2051_413#_c_1716_n 0.00609226f $X=11.84 $Y=1.717
+ $X2=0 $Y2=0
cc_720 N_A_791_264#_c_832_n N_A_2051_413#_c_1716_n 0.00641947f $X=12.01 $Y=1.717
+ $X2=0 $Y2=0
cc_721 N_A_791_264#_c_817_n N_A_2051_413#_c_1716_n 0.00500691f $X=12.015
+ $Y=0.825 $X2=0 $Y2=0
cc_722 N_A_791_264#_c_818_n N_A_2051_413#_c_1716_n 0.00892528f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_723 N_A_791_264#_c_821_n N_A_2051_413#_c_1716_n 0.00143362f $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_724 N_A_791_264#_c_822_n N_A_2051_413#_c_1716_n 0.0170494f $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_725 N_A_791_264#_c_822_n N_A_2051_413#_c_1717_n 0.00983534f $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_726 N_A_791_264#_M1007_g N_A_2051_413#_c_1730_n 0.00510852f $X=11.17 $Y=2.275
+ $X2=0 $Y2=0
cc_727 N_A_791_264#_M1001_g N_A_2051_413#_c_1733_n 0.00188481f $X=11.285
+ $Y=0.445 $X2=0 $Y2=0
cc_728 N_A_791_264#_c_818_n N_A_2051_413#_c_1733_n 0.00605628f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_729 N_A_791_264#_M1001_g N_A_2051_413#_c_1719_n 0.0088172f $X=11.285 $Y=0.445
+ $X2=0 $Y2=0
cc_730 N_A_791_264#_c_818_n N_A_2051_413#_c_1719_n 0.0223085f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_731 N_A_791_264#_M1007_g N_A_2051_413#_c_1728_n 0.0120201f $X=11.17 $Y=2.275
+ $X2=0 $Y2=0
cc_732 N_A_791_264#_M1001_g N_A_2051_413#_c_1728_n 0.00751613f $X=11.285
+ $Y=0.445 $X2=0 $Y2=0
cc_733 N_A_791_264#_c_827_n N_A_2051_413#_c_1728_n 0.0282373f $X=11.84 $Y=1.717
+ $X2=0 $Y2=0
cc_734 N_A_791_264#_c_828_n N_A_2051_413#_c_1728_n 0.0079118f $X=11.365 $Y=1.74
+ $X2=0 $Y2=0
cc_735 N_A_791_264#_M1001_g N_A_2051_413#_c_1720_n 0.0183255f $X=11.285 $Y=0.445
+ $X2=0 $Y2=0
cc_736 N_A_791_264#_c_827_n N_A_2051_413#_c_1720_n 0.0359416f $X=11.84 $Y=1.717
+ $X2=0 $Y2=0
cc_737 N_A_791_264#_c_828_n N_A_2051_413#_c_1720_n 0.00495398f $X=11.365 $Y=1.74
+ $X2=0 $Y2=0
cc_738 N_A_791_264#_c_818_n N_A_2051_413#_c_1720_n 0.0291683f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_739 N_A_791_264#_c_822_n N_A_2051_413#_c_1720_n 0.0240437f $X=12.085 $Y=0.85
+ $X2=0 $Y2=0
cc_740 N_A_791_264#_M1007_g N_VPWR_c_1831_n 0.00462747f $X=11.17 $Y=2.275 $X2=0
+ $Y2=0
cc_741 N_A_791_264#_c_827_n N_VPWR_c_1831_n 0.0155824f $X=11.84 $Y=1.717 $X2=0
+ $Y2=0
cc_742 N_A_791_264#_c_828_n N_VPWR_c_1831_n 0.00514677f $X=11.365 $Y=1.74 $X2=0
+ $Y2=0
cc_743 N_A_791_264#_c_829_n N_VPWR_c_1831_n 0.0182471f $X=12.005 $Y=1.99 $X2=0
+ $Y2=0
cc_744 N_A_791_264#_c_832_n N_VPWR_c_1832_n 0.0283369f $X=12.01 $Y=1.717 $X2=0
+ $Y2=0
cc_745 N_A_791_264#_c_822_n N_VPWR_c_1832_n 0.00515656f $X=12.085 $Y=0.85 $X2=0
+ $Y2=0
cc_746 N_A_791_264#_M1007_g N_VPWR_c_1835_n 0.00564808f $X=11.17 $Y=2.275 $X2=0
+ $Y2=0
cc_747 N_A_791_264#_c_829_n N_VPWR_c_1837_n 0.0217414f $X=12.005 $Y=1.99 $X2=0
+ $Y2=0
cc_748 N_A_791_264#_M1036_g N_VPWR_c_1841_n 0.00541359f $X=4.08 $Y=2.165 $X2=0
+ $Y2=0
cc_749 N_A_791_264#_M1023_s N_VPWR_c_1823_n 0.00217517f $X=11.88 $Y=1.845 $X2=0
+ $Y2=0
cc_750 N_A_791_264#_M1036_g N_VPWR_c_1823_n 0.00652616f $X=4.08 $Y=2.165 $X2=0
+ $Y2=0
cc_751 N_A_791_264#_M1007_g N_VPWR_c_1823_n 0.0117199f $X=11.17 $Y=2.275 $X2=0
+ $Y2=0
cc_752 N_A_791_264#_c_827_n N_VPWR_c_1823_n 0.0122998f $X=11.84 $Y=1.717 $X2=0
+ $Y2=0
cc_753 N_A_791_264#_c_828_n N_VPWR_c_1823_n 8.92751e-19 $X=11.365 $Y=1.74 $X2=0
+ $Y2=0
cc_754 N_A_791_264#_c_829_n N_VPWR_c_1823_n 0.0128119f $X=12.005 $Y=1.99 $X2=0
+ $Y2=0
cc_755 N_A_791_264#_M1036_g N_A_299_47#_c_2018_n 0.0132707f $X=4.08 $Y=2.165
+ $X2=0 $Y2=0
cc_756 N_A_791_264#_c_830_n N_A_299_47#_c_2018_n 0.00318555f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_757 N_A_791_264#_c_831_n N_A_299_47#_c_2018_n 0.00178853f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_758 N_A_791_264#_M1041_g N_A_299_47#_c_2010_n 0.00247582f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_759 N_A_791_264#_M1036_g N_A_299_47#_c_2010_n 0.00245488f $X=4.08 $Y=2.165
+ $X2=0 $Y2=0
cc_760 N_A_791_264#_c_830_n N_A_299_47#_c_2010_n 0.0238925f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_761 N_A_791_264#_c_831_n N_A_299_47#_c_2010_n 0.00361751f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_762 N_A_791_264#_c_820_n N_A_299_47#_c_2010_n 0.00525839f $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_763 N_A_791_264#_M1041_g N_A_299_47#_c_2011_n 0.00526337f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_764 N_A_791_264#_c_830_n N_A_299_47#_c_2011_n 0.00212358f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_765 N_A_791_264#_c_831_n N_A_299_47#_c_2011_n 0.00197416f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_766 N_A_791_264#_c_818_n N_A_299_47#_c_2011_n 0.00430154f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_767 N_A_791_264#_M1041_g N_A_299_47#_c_2040_n 0.00100352f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_768 N_A_791_264#_c_818_n N_A_299_47#_c_2040_n 0.0250725f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_769 N_A_791_264#_M1041_g N_A_299_47#_c_2013_n 0.00367101f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_770 N_A_791_264#_c_818_n N_A_299_47#_c_2013_n 0.00735691f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_771 N_A_791_264#_c_819_n N_A_299_47#_c_2013_n 0.0273168f $X=4.035 $Y=0.85
+ $X2=0 $Y2=0
cc_772 N_A_791_264#_c_820_n N_A_299_47#_c_2013_n 0.00264974f $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_773 N_A_791_264#_M1041_g N_A_299_47#_c_2014_n 0.0129918f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_774 N_A_791_264#_c_818_n N_A_299_47#_c_2014_n 0.0173013f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_775 N_A_791_264#_c_819_n N_A_299_47#_c_2014_n 0.00238395f $X=4.035 $Y=0.85
+ $X2=0 $Y2=0
cc_776 N_A_791_264#_c_820_n N_A_299_47#_c_2014_n 0.0329237f $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_777 N_A_791_264#_c_818_n N_A_915_47#_M1009_d 0.00214089f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_778 N_A_791_264#_c_818_n N_A_915_47#_c_2130_n 0.027265f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_779 N_A_791_264#_c_818_n N_A_915_47#_c_2131_n 0.00714473f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_780 N_A_791_264#_M1041_g N_A_915_47#_c_2132_n 0.00169341f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_781 N_A_791_264#_c_818_n N_A_915_47#_c_2132_n 0.00947367f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_782 N_A_791_264#_c_818_n N_A_915_47#_c_2135_n 0.0252919f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_783 N_A_791_264#_c_818_n N_A_915_47#_c_2168_n 0.0249712f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_784 N_A_791_264#_c_818_n N_A_915_47#_c_2136_n 0.130603f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_785 N_A_791_264#_c_818_n N_A_915_47#_c_2137_n 0.00623535f $X=11.94 $Y=0.85
+ $X2=0 $Y2=0
cc_786 N_A_791_264#_c_821_n N_Q_c_2269_n 0.00151602f $X=12.085 $Y=0.85 $X2=0
+ $Y2=0
cc_787 N_A_791_264#_c_822_n N_Q_c_2269_n 0.0137869f $X=12.085 $Y=0.85 $X2=0
+ $Y2=0
cc_788 N_A_791_264#_c_818_n N_VGND_M1005_d 0.00270061f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_789 N_A_791_264#_M1041_g N_VGND_c_2288_n 0.00210691f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_790 N_A_791_264#_c_818_n N_VGND_c_2289_n 0.0117651f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_791 N_A_791_264#_c_818_n N_VGND_c_2290_n 0.00209284f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_792 N_A_791_264#_c_818_n N_VGND_c_2291_n 0.00448688f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_793 N_A_791_264#_M1001_g N_VGND_c_2292_n 0.010757f $X=11.285 $Y=0.445 $X2=0
+ $Y2=0
cc_794 N_A_791_264#_c_816_n N_VGND_c_2292_n 0.0246268f $X=12.015 $Y=0.385 $X2=0
+ $Y2=0
cc_795 N_A_791_264#_c_818_n N_VGND_c_2292_n 0.00490532f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_796 N_A_791_264#_c_816_n N_VGND_c_2293_n 0.0299916f $X=12.015 $Y=0.385 $X2=0
+ $Y2=0
cc_797 N_A_791_264#_c_821_n N_VGND_c_2293_n 0.00495351f $X=12.085 $Y=0.85 $X2=0
+ $Y2=0
cc_798 N_A_791_264#_M1041_g N_VGND_c_2296_n 0.00571722f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_799 N_A_791_264#_c_820_n N_VGND_c_2296_n 0.00260398f $X=3.89 $Y=0.85 $X2=0
+ $Y2=0
cc_800 N_A_791_264#_M1001_g N_VGND_c_2300_n 0.00544582f $X=11.285 $Y=0.445 $X2=0
+ $Y2=0
cc_801 N_A_791_264#_c_816_n N_VGND_c_2302_n 0.016199f $X=12.015 $Y=0.385 $X2=0
+ $Y2=0
cc_802 N_A_791_264#_M1031_s N_VGND_c_2308_n 0.00169299f $X=11.89 $Y=0.235 $X2=0
+ $Y2=0
cc_803 N_A_791_264#_M1041_g N_VGND_c_2308_n 0.00552168f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_804 N_A_791_264#_M1001_g N_VGND_c_2308_n 0.00524744f $X=11.285 $Y=0.445 $X2=0
+ $Y2=0
cc_805 N_A_791_264#_c_816_n N_VGND_c_2308_n 0.00555624f $X=12.015 $Y=0.385 $X2=0
+ $Y2=0
cc_806 N_A_791_264#_c_818_n N_VGND_c_2308_n 0.252627f $X=11.94 $Y=0.85 $X2=0
+ $Y2=0
cc_807 N_A_791_264#_c_821_n N_VGND_c_2308_n 0.0146996f $X=12.085 $Y=0.85 $X2=0
+ $Y2=0
cc_808 N_A_791_264#_c_818_n A_1226_119# 0.00414878f $X=11.94 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_809 N_A_885_21#_c_1008_n N_SCD_M1024_g 2.23202e-19 $X=5.425 $Y=0.75 $X2=0
+ $Y2=0
cc_810 N_A_885_21#_c_1009_n N_SCD_M1024_g 2.06692e-19 $X=5.505 $Y=1.835 $X2=0
+ $Y2=0
cc_811 N_A_885_21#_c_1012_n N_SCD_M1024_g 9.76068e-19 $X=5.425 $Y=0.935 $X2=0
+ $Y2=0
cc_812 N_A_885_21#_M1030_g N_SCD_M1020_g 0.0341463f $X=6.56 $Y=2.165 $X2=0 $Y2=0
cc_813 N_A_885_21#_c_1009_n N_SCD_M1020_g 9.31983e-19 $X=5.505 $Y=1.835 $X2=0
+ $Y2=0
cc_814 N_A_885_21#_c_1015_n N_SCD_M1020_g 0.0119239f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_815 N_A_885_21#_c_1010_n N_SCD_M1020_g 0.00285156f $X=6.5 $Y=1.52 $X2=0 $Y2=0
cc_816 N_A_885_21#_c_1018_n N_SCD_M1020_g 9.97145e-19 $X=5.32 $Y=2 $X2=0 $Y2=0
cc_817 N_A_885_21#_c_1009_n SCD 0.0422189f $X=5.505 $Y=1.835 $X2=0 $Y2=0
cc_818 N_A_885_21#_c_1015_n SCD 0.031117f $X=6.385 $Y=1.92 $X2=0 $Y2=0
cc_819 N_A_885_21#_c_1010_n SCD 0.0229756f $X=6.5 $Y=1.52 $X2=0 $Y2=0
cc_820 N_A_885_21#_c_1011_n SCD 0.00162041f $X=6.5 $Y=1.52 $X2=0 $Y2=0
cc_821 N_A_885_21#_c_1009_n N_SCD_c_1133_n 4.99203e-19 $X=5.505 $Y=1.835 $X2=0
+ $Y2=0
cc_822 N_A_885_21#_c_1015_n N_SCD_c_1133_n 0.00279837f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_823 N_A_885_21#_c_1010_n N_SCD_c_1133_n 5.39908e-19 $X=6.5 $Y=1.52 $X2=0
+ $Y2=0
cc_824 N_A_885_21#_c_1011_n N_SCD_c_1133_n 0.0212159f $X=6.5 $Y=1.52 $X2=0 $Y2=0
cc_825 N_A_885_21#_c_1003_n N_SCE_c_1179_n 0.00553839f $X=4.995 $Y=0.84 $X2=0
+ $Y2=0
cc_826 N_A_885_21#_c_1004_n N_SCE_c_1188_n 0.00553839f $X=4.575 $Y=0.84 $X2=0
+ $Y2=0
cc_827 N_A_885_21#_c_1009_n N_SCE_M1033_g 0.0102925f $X=5.505 $Y=1.835 $X2=0
+ $Y2=0
cc_828 N_A_885_21#_c_1015_n N_SCE_M1033_g 0.00378294f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_829 N_A_885_21#_c_1018_n N_SCE_M1033_g 0.0115767f $X=5.32 $Y=2 $X2=0 $Y2=0
cc_830 N_A_885_21#_c_1005_n N_SCE_M1005_g 0.00660962f $X=5.07 $Y=0.765 $X2=0
+ $Y2=0
cc_831 N_A_885_21#_c_1006_n N_SCE_M1005_g 0.0055978f $X=5.26 $Y=0.385 $X2=0
+ $Y2=0
cc_832 N_A_885_21#_c_1008_n N_SCE_M1005_g 0.00346462f $X=5.425 $Y=0.75 $X2=0
+ $Y2=0
cc_833 N_A_885_21#_c_1009_n N_SCE_M1005_g 0.00553447f $X=5.505 $Y=1.835 $X2=0
+ $Y2=0
cc_834 N_A_885_21#_c_1012_n N_SCE_M1005_g 0.00160804f $X=5.425 $Y=0.935 $X2=0
+ $Y2=0
cc_835 N_A_885_21#_c_1006_n N_SCE_c_1182_n 2.57001e-19 $X=5.26 $Y=0.385 $X2=0
+ $Y2=0
cc_836 N_A_885_21#_c_1007_n N_SCE_c_1182_n 0.0145162f $X=5.13 $Y=0.34 $X2=0
+ $Y2=0
cc_837 N_A_885_21#_c_1015_n N_SCE_M1009_g 5.19778e-19 $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_838 N_A_885_21#_c_1010_n N_SCE_M1009_g 7.94182e-19 $X=6.5 $Y=1.52 $X2=0 $Y2=0
cc_839 N_A_885_21#_c_1011_n N_SCE_M1009_g 0.00852721f $X=6.5 $Y=1.52 $X2=0 $Y2=0
cc_840 N_A_885_21#_c_1003_n N_SCE_c_1184_n 0.0014425f $X=4.995 $Y=0.84 $X2=0
+ $Y2=0
cc_841 N_A_885_21#_c_1006_n N_SCE_c_1184_n 0.00321461f $X=5.26 $Y=0.385 $X2=0
+ $Y2=0
cc_842 N_A_885_21#_c_1007_n N_SCE_c_1184_n 6.16455e-19 $X=5.13 $Y=0.34 $X2=0
+ $Y2=0
cc_843 N_A_885_21#_c_1009_n N_SCE_c_1184_n 0.0365192f $X=5.505 $Y=1.835 $X2=0
+ $Y2=0
cc_844 N_A_885_21#_c_1018_n N_SCE_c_1184_n 0.00528494f $X=5.32 $Y=2 $X2=0 $Y2=0
cc_845 N_A_885_21#_c_1003_n N_SCE_c_1185_n 0.00637023f $X=4.995 $Y=0.84 $X2=0
+ $Y2=0
cc_846 N_A_885_21#_c_1009_n N_SCE_c_1185_n 0.0190301f $X=5.505 $Y=1.835 $X2=0
+ $Y2=0
cc_847 N_A_885_21#_c_1015_n N_SCE_c_1185_n 0.00218618f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_848 N_A_885_21#_c_1018_n N_SCE_c_1185_n 0.00370055f $X=5.32 $Y=2 $X2=0 $Y2=0
cc_849 N_A_885_21#_c_1012_n N_SCE_c_1185_n 0.0057535f $X=5.425 $Y=0.935 $X2=0
+ $Y2=0
cc_850 N_A_885_21#_c_1011_n N_A_193_47#_M1008_g 0.0249846f $X=6.5 $Y=1.52 $X2=0
+ $Y2=0
cc_851 N_A_885_21#_c_1004_n N_A_193_47#_c_1285_n 4.56595e-19 $X=4.575 $Y=0.84
+ $X2=0 $Y2=0
cc_852 N_A_885_21#_c_1009_n N_A_193_47#_c_1285_n 0.0126257f $X=5.505 $Y=1.835
+ $X2=0 $Y2=0
cc_853 N_A_885_21#_c_1015_n N_A_193_47#_c_1285_n 0.00300896f $X=6.385 $Y=1.92
+ $X2=0 $Y2=0
cc_854 N_A_885_21#_c_1010_n N_A_193_47#_c_1285_n 0.0123204f $X=6.5 $Y=1.52 $X2=0
+ $Y2=0
cc_855 N_A_885_21#_c_1011_n N_A_193_47#_c_1285_n 0.00302472f $X=6.5 $Y=1.52
+ $X2=0 $Y2=0
cc_856 N_A_885_21#_c_1018_n N_A_193_47#_c_1285_n 0.00120533f $X=5.32 $Y=2 $X2=0
+ $Y2=0
cc_857 N_A_885_21#_c_1012_n N_A_193_47#_c_1285_n 0.00398102f $X=5.425 $Y=0.935
+ $X2=0 $Y2=0
cc_858 N_A_885_21#_c_1011_n N_A_193_47#_c_1279_n 0.0035473f $X=6.5 $Y=1.52 $X2=0
+ $Y2=0
cc_859 N_A_885_21#_c_1015_n N_VPWR_M1033_d 0.00321876f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_860 N_A_885_21#_M1030_g N_VPWR_c_1827_n 0.00188336f $X=6.56 $Y=2.165 $X2=0
+ $Y2=0
cc_861 N_A_885_21#_c_1015_n N_VPWR_c_1827_n 0.0201793f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_862 N_A_885_21#_c_1015_n N_VPWR_c_1841_n 6.97462e-19 $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_863 N_A_885_21#_c_1018_n N_VPWR_c_1841_n 0.0230574f $X=5.32 $Y=2 $X2=0 $Y2=0
cc_864 N_A_885_21#_M1030_g N_VPWR_c_1842_n 0.00486028f $X=6.56 $Y=2.165 $X2=0
+ $Y2=0
cc_865 N_A_885_21#_c_1015_n N_VPWR_c_1842_n 0.00763017f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_866 N_A_885_21#_M1033_s N_VPWR_c_1823_n 0.00175811f $X=5.195 $Y=1.845 $X2=0
+ $Y2=0
cc_867 N_A_885_21#_M1030_g N_VPWR_c_1823_n 0.00653909f $X=6.56 $Y=2.165 $X2=0
+ $Y2=0
cc_868 N_A_885_21#_c_1015_n N_VPWR_c_1823_n 0.00792805f $X=6.385 $Y=1.92 $X2=0
+ $Y2=0
cc_869 N_A_885_21#_c_1018_n N_VPWR_c_1823_n 0.00708842f $X=5.32 $Y=2 $X2=0 $Y2=0
cc_870 N_A_885_21#_c_1004_n N_A_299_47#_c_2011_n 0.00354861f $X=4.575 $Y=0.84
+ $X2=0 $Y2=0
cc_871 N_A_885_21#_c_1002_n N_A_299_47#_c_2014_n 0.00261058f $X=4.5 $Y=0.765
+ $X2=0 $Y2=0
cc_872 N_A_885_21#_c_1018_n N_A_915_47#_c_2138_n 0.01209f $X=5.32 $Y=2 $X2=0
+ $Y2=0
cc_873 N_A_885_21#_c_1018_n N_A_915_47#_c_2139_n 0.0352313f $X=5.32 $Y=2 $X2=0
+ $Y2=0
cc_874 N_A_885_21#_M1030_g N_A_915_47#_c_2151_n 0.00426855f $X=6.56 $Y=2.165
+ $X2=0 $Y2=0
cc_875 N_A_885_21#_c_1003_n N_A_915_47#_c_2131_n 0.00828733f $X=4.995 $Y=0.84
+ $X2=0 $Y2=0
cc_876 N_A_885_21#_c_1005_n N_A_915_47#_c_2131_n 0.00126502f $X=5.07 $Y=0.765
+ $X2=0 $Y2=0
cc_877 N_A_885_21#_c_1008_n N_A_915_47#_c_2131_n 0.00512039f $X=5.425 $Y=0.75
+ $X2=0 $Y2=0
cc_878 N_A_885_21#_c_1003_n N_A_915_47#_c_2132_n 0.00645336f $X=4.995 $Y=0.84
+ $X2=0 $Y2=0
cc_879 N_A_885_21#_c_1009_n N_A_915_47#_c_2132_n 0.00942669f $X=5.505 $Y=1.835
+ $X2=0 $Y2=0
cc_880 N_A_885_21#_c_1012_n N_A_915_47#_c_2132_n 0.00512039f $X=5.425 $Y=0.935
+ $X2=0 $Y2=0
cc_881 N_A_885_21#_c_1010_n N_A_915_47#_c_2133_n 0.00529702f $X=6.5 $Y=1.52
+ $X2=0 $Y2=0
cc_882 N_A_885_21#_c_1011_n N_A_915_47#_c_2133_n 0.00295115f $X=6.5 $Y=1.52
+ $X2=0 $Y2=0
cc_883 N_A_885_21#_c_1015_n N_A_915_47#_c_2134_n 0.0123117f $X=6.385 $Y=1.92
+ $X2=0 $Y2=0
cc_884 N_A_885_21#_c_1010_n N_A_915_47#_c_2134_n 0.0336064f $X=6.5 $Y=1.52 $X2=0
+ $Y2=0
cc_885 N_A_885_21#_c_1011_n N_A_915_47#_c_2134_n 0.00426855f $X=6.5 $Y=1.52
+ $X2=0 $Y2=0
cc_886 N_A_885_21#_c_1002_n N_A_915_47#_c_2135_n 9.60356e-19 $X=4.5 $Y=0.765
+ $X2=0 $Y2=0
cc_887 N_A_885_21#_c_1005_n N_A_915_47#_c_2135_n 7.37078e-19 $X=5.07 $Y=0.765
+ $X2=0 $Y2=0
cc_888 N_A_885_21#_c_1008_n N_A_915_47#_c_2135_n 0.00115128f $X=5.425 $Y=0.75
+ $X2=0 $Y2=0
cc_889 N_A_885_21#_c_1003_n N_A_915_47#_c_2136_n 6.24142e-19 $X=4.995 $Y=0.84
+ $X2=0 $Y2=0
cc_890 N_A_885_21#_c_1005_n N_A_915_47#_c_2136_n 0.00237108f $X=5.07 $Y=0.765
+ $X2=0 $Y2=0
cc_891 N_A_885_21#_c_1006_n N_A_915_47#_c_2136_n 0.0202599f $X=5.26 $Y=0.385
+ $X2=0 $Y2=0
cc_892 N_A_885_21#_c_1008_n N_A_915_47#_c_2136_n 0.00951737f $X=5.425 $Y=0.75
+ $X2=0 $Y2=0
cc_893 N_A_885_21#_c_1002_n N_A_915_47#_c_2192_n 0.0014936f $X=4.5 $Y=0.765
+ $X2=0 $Y2=0
cc_894 N_A_885_21#_c_1005_n N_A_915_47#_c_2192_n 0.00107169f $X=5.07 $Y=0.765
+ $X2=0 $Y2=0
cc_895 N_A_885_21#_c_1006_n N_A_915_47#_c_2192_n 0.0201338f $X=5.26 $Y=0.385
+ $X2=0 $Y2=0
cc_896 N_A_885_21#_c_1007_n N_A_915_47#_c_2192_n 8.02625e-19 $X=5.13 $Y=0.34
+ $X2=0 $Y2=0
cc_897 N_A_885_21#_c_1008_n N_A_915_47#_c_2192_n 0.00329508f $X=5.425 $Y=0.75
+ $X2=0 $Y2=0
cc_898 N_A_885_21#_c_1015_n A_1231_369# 0.00410624f $X=6.385 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_899 N_A_885_21#_c_1006_n N_VGND_c_2289_n 0.0196608f $X=5.26 $Y=0.385 $X2=0
+ $Y2=0
cc_900 N_A_885_21#_c_1007_n N_VGND_c_2289_n 4.91263e-19 $X=5.13 $Y=0.34 $X2=0
+ $Y2=0
cc_901 N_A_885_21#_c_1008_n N_VGND_c_2289_n 0.0187439f $X=5.425 $Y=0.75 $X2=0
+ $Y2=0
cc_902 N_A_885_21#_c_1002_n N_VGND_c_2296_n 0.00585385f $X=4.5 $Y=0.765 $X2=0
+ $Y2=0
cc_903 N_A_885_21#_c_1003_n N_VGND_c_2296_n 0.00127181f $X=4.995 $Y=0.84 $X2=0
+ $Y2=0
cc_904 N_A_885_21#_c_1006_n N_VGND_c_2296_n 0.0422697f $X=5.26 $Y=0.385 $X2=0
+ $Y2=0
cc_905 N_A_885_21#_c_1007_n N_VGND_c_2296_n 0.00544529f $X=5.13 $Y=0.34 $X2=0
+ $Y2=0
cc_906 N_A_885_21#_c_1002_n N_VGND_c_2308_n 0.00720023f $X=4.5 $Y=0.765 $X2=0
+ $Y2=0
cc_907 N_A_885_21#_c_1006_n N_VGND_c_2308_n 0.00545326f $X=5.26 $Y=0.385 $X2=0
+ $Y2=0
cc_908 N_A_885_21#_c_1007_n N_VGND_c_2308_n 0.00670392f $X=5.13 $Y=0.34 $X2=0
+ $Y2=0
cc_909 N_SCD_M1020_g N_SCE_M1033_g 0.022868f $X=6.08 $Y=2.165 $X2=0 $Y2=0
cc_910 N_SCD_M1024_g N_SCE_M1005_g 0.0200438f $X=6.055 $Y=0.805 $X2=0 $Y2=0
cc_911 N_SCD_M1024_g N_SCE_c_1181_n 0.0100965f $X=6.055 $Y=0.805 $X2=0 $Y2=0
cc_912 N_SCD_M1024_g N_SCE_M1009_g 0.0428375f $X=6.055 $Y=0.805 $X2=0 $Y2=0
cc_913 SCD N_SCE_M1009_g 3.13488e-19 $X=5.895 $Y=1.105 $X2=0 $Y2=0
cc_914 N_SCD_M1024_g N_SCE_c_1185_n 0.00342493f $X=6.055 $Y=0.805 $X2=0 $Y2=0
cc_915 SCD N_SCE_c_1185_n 0.00397767f $X=5.895 $Y=1.105 $X2=0 $Y2=0
cc_916 N_SCD_c_1133_n N_SCE_c_1185_n 0.0154611f $X=6.02 $Y=1.52 $X2=0 $Y2=0
cc_917 SCD N_A_193_47#_c_1285_n 0.024323f $X=5.895 $Y=1.105 $X2=0 $Y2=0
cc_918 N_SCD_M1020_g N_VPWR_c_1827_n 0.0142327f $X=6.08 $Y=2.165 $X2=0 $Y2=0
cc_919 N_SCD_M1020_g N_VPWR_c_1842_n 0.00421152f $X=6.08 $Y=2.165 $X2=0 $Y2=0
cc_920 N_SCD_M1020_g N_VPWR_c_1823_n 0.00471179f $X=6.08 $Y=2.165 $X2=0 $Y2=0
cc_921 N_SCD_M1024_g N_A_915_47#_c_2133_n 2.50449e-19 $X=6.055 $Y=0.805 $X2=0
+ $Y2=0
cc_922 SCD N_A_915_47#_c_2133_n 0.00467347f $X=5.895 $Y=1.105 $X2=0 $Y2=0
cc_923 N_SCD_M1024_g N_A_915_47#_c_2134_n 7.86841e-19 $X=6.055 $Y=0.805 $X2=0
+ $Y2=0
cc_924 SCD N_A_915_47#_c_2134_n 0.00619056f $X=5.895 $Y=1.105 $X2=0 $Y2=0
cc_925 N_SCD_M1024_g N_A_915_47#_c_2168_n 2.02646e-19 $X=6.055 $Y=0.805 $X2=0
+ $Y2=0
cc_926 N_SCD_M1024_g N_A_915_47#_c_2136_n 0.00162107f $X=6.055 $Y=0.805 $X2=0
+ $Y2=0
cc_927 N_SCD_M1024_g N_VGND_c_2289_n 0.00812902f $X=6.055 $Y=0.805 $X2=0 $Y2=0
cc_928 SCD N_VGND_c_2289_n 0.0141356f $X=5.895 $Y=1.105 $X2=0 $Y2=0
cc_929 N_SCD_c_1133_n N_VGND_c_2289_n 3.1502e-19 $X=6.02 $Y=1.52 $X2=0 $Y2=0
cc_930 N_SCE_M1013_g N_A_193_47#_c_1285_n 0.00139967f $X=4.54 $Y=2.165 $X2=0
+ $Y2=0
cc_931 N_SCE_c_1179_n N_A_193_47#_c_1285_n 0.00230653f $X=4.955 $Y=1.5 $X2=0
+ $Y2=0
cc_932 N_SCE_c_1188_n N_A_193_47#_c_1285_n 8.85046e-19 $X=4.615 $Y=1.5 $X2=0
+ $Y2=0
cc_933 N_SCE_M1033_g N_A_193_47#_c_1285_n 2.76439e-19 $X=5.535 $Y=2.165 $X2=0
+ $Y2=0
cc_934 N_SCE_M1009_g N_A_193_47#_c_1285_n 5.39536e-19 $X=6.415 $Y=0.805 $X2=0
+ $Y2=0
cc_935 N_SCE_c_1184_n N_A_193_47#_c_1285_n 0.0130697f $X=5.12 $Y=1.44 $X2=0
+ $Y2=0
cc_936 N_SCE_c_1185_n N_A_193_47#_c_1285_n 0.00676958f $X=5.535 $Y=1.332 $X2=0
+ $Y2=0
cc_937 N_SCE_M1033_g N_VPWR_c_1827_n 0.00304048f $X=5.535 $Y=2.165 $X2=0 $Y2=0
cc_938 N_SCE_M1013_g N_VPWR_c_1841_n 0.00536022f $X=4.54 $Y=2.165 $X2=0 $Y2=0
cc_939 N_SCE_M1033_g N_VPWR_c_1841_n 0.00419527f $X=5.535 $Y=2.165 $X2=0 $Y2=0
cc_940 N_SCE_M1013_g N_VPWR_c_1823_n 0.00755353f $X=4.54 $Y=2.165 $X2=0 $Y2=0
cc_941 N_SCE_M1033_g N_VPWR_c_1823_n 0.0070231f $X=5.535 $Y=2.165 $X2=0 $Y2=0
cc_942 N_SCE_M1013_g N_A_299_47#_c_2018_n 0.00348858f $X=4.54 $Y=2.165 $X2=0
+ $Y2=0
cc_943 N_SCE_M1013_g N_A_299_47#_c_2010_n 0.00476513f $X=4.54 $Y=2.165 $X2=0
+ $Y2=0
cc_944 N_SCE_c_1188_n N_A_299_47#_c_2010_n 0.00370037f $X=4.615 $Y=1.5 $X2=0
+ $Y2=0
cc_945 N_SCE_c_1179_n N_A_915_47#_c_2138_n 0.00385829f $X=4.955 $Y=1.5 $X2=0
+ $Y2=0
cc_946 N_SCE_M1033_g N_A_915_47#_c_2138_n 0.00153514f $X=5.535 $Y=2.165 $X2=0
+ $Y2=0
cc_947 N_SCE_M1009_g N_A_915_47#_c_2130_n 0.00701148f $X=6.415 $Y=0.805 $X2=0
+ $Y2=0
cc_948 N_SCE_c_1188_n N_A_915_47#_c_2131_n 7.51487e-19 $X=4.615 $Y=1.5 $X2=0
+ $Y2=0
cc_949 N_SCE_M1013_g N_A_915_47#_c_2132_n 0.00680013f $X=4.54 $Y=2.165 $X2=0
+ $Y2=0
cc_950 N_SCE_c_1179_n N_A_915_47#_c_2132_n 0.0116261f $X=4.955 $Y=1.5 $X2=0
+ $Y2=0
cc_951 N_SCE_M1033_g N_A_915_47#_c_2132_n 8.62346e-19 $X=5.535 $Y=2.165 $X2=0
+ $Y2=0
cc_952 N_SCE_c_1184_n N_A_915_47#_c_2132_n 0.0369704f $X=5.12 $Y=1.44 $X2=0
+ $Y2=0
cc_953 N_SCE_c_1185_n N_A_915_47#_c_2132_n 0.00363922f $X=5.535 $Y=1.332 $X2=0
+ $Y2=0
cc_954 N_SCE_M1009_g N_A_915_47#_c_2168_n 0.00354275f $X=6.415 $Y=0.805 $X2=0
+ $Y2=0
cc_955 N_SCE_M1005_g N_A_915_47#_c_2136_n 0.00345261f $X=5.635 $Y=0.805 $X2=0
+ $Y2=0
cc_956 N_SCE_c_1181_n N_A_915_47#_c_2136_n 0.0018451f $X=6.34 $Y=0.18 $X2=0
+ $Y2=0
cc_957 N_SCE_M1009_g N_A_915_47#_c_2136_n 0.00407187f $X=6.415 $Y=0.805 $X2=0
+ $Y2=0
cc_958 N_SCE_M1009_g N_A_915_47#_c_2137_n 0.00841094f $X=6.415 $Y=0.805 $X2=0
+ $Y2=0
cc_959 N_SCE_M1005_g N_VGND_c_2289_n 0.00321091f $X=5.635 $Y=0.805 $X2=0 $Y2=0
cc_960 N_SCE_c_1181_n N_VGND_c_2289_n 0.0192645f $X=6.34 $Y=0.18 $X2=0 $Y2=0
cc_961 N_SCE_M1009_g N_VGND_c_2289_n 0.00320475f $X=6.415 $Y=0.805 $X2=0 $Y2=0
cc_962 N_SCE_c_1182_n N_VGND_c_2296_n 0.00731067f $X=5.71 $Y=0.18 $X2=0 $Y2=0
cc_963 N_SCE_c_1181_n N_VGND_c_2306_n 0.0177988f $X=6.34 $Y=0.18 $X2=0 $Y2=0
cc_964 N_SCE_c_1181_n N_VGND_c_2308_n 0.0135574f $X=6.34 $Y=0.18 $X2=0 $Y2=0
cc_965 N_SCE_c_1182_n N_VGND_c_2308_n 0.00505206f $X=5.71 $Y=0.18 $X2=0 $Y2=0
cc_966 N_A_193_47#_c_1273_n N_A_1610_159#_M1006_g 0.0138337f $X=7.655 $Y=1.29
+ $X2=0 $Y2=0
cc_967 N_A_193_47#_c_1287_n N_A_1610_159#_M1006_g 0.00185536f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_968 N_A_193_47#_c_1279_n N_A_1610_159#_M1006_g 0.00119103f $X=7.18 $Y=1.29
+ $X2=0 $Y2=0
cc_969 N_A_193_47#_M1012_g N_A_1610_159#_M1019_g 0.0189994f $X=7.73 $Y=0.415
+ $X2=0 $Y2=0
cc_970 N_A_193_47#_c_1287_n N_A_1610_159#_M1037_g 0.00722181f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_971 N_A_193_47#_c_1275_n N_A_1610_159#_M1039_g 0.0181756f $X=10.28 $Y=0.705
+ $X2=0 $Y2=0
cc_972 N_A_193_47#_c_1276_n N_A_1610_159#_M1039_g 0.00208129f $X=10.39 $Y=0.87
+ $X2=0 $Y2=0
cc_973 N_A_193_47#_c_1277_n N_A_1610_159#_c_1492_n 0.0181756f $X=10.39 $Y=0.87
+ $X2=0 $Y2=0
cc_974 N_A_193_47#_c_1287_n N_A_1610_159#_c_1492_n 0.00123775f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_975 N_A_193_47#_c_1278_n N_A_1610_159#_c_1492_n 2.51226e-19 $X=10.605 $Y=1.53
+ $X2=0 $Y2=0
cc_976 N_A_193_47#_c_1287_n N_A_1610_159#_c_1493_n 0.00252648f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_977 N_A_193_47#_c_1287_n N_A_1610_159#_c_1494_n 0.00787458f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_978 N_A_193_47#_c_1287_n N_A_1610_159#_c_1504_n 0.0260184f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_979 N_A_193_47#_c_1287_n N_A_1610_159#_c_1496_n 0.0182403f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_980 N_A_193_47#_c_1278_n N_A_1610_159#_c_1497_n 0.00478379f $X=10.605 $Y=1.53
+ $X2=0 $Y2=0
cc_981 N_A_193_47#_c_1287_n N_A_1610_159#_c_1498_n 7.49207e-19 $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_982 N_A_193_47#_M1012_g N_A_1610_159#_c_1499_n 0.0138337f $X=7.73 $Y=0.415
+ $X2=0 $Y2=0
cc_983 N_A_193_47#_c_1287_n N_A_1446_413#_M1017_g 0.00174404f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_984 N_A_193_47#_c_1287_n N_A_1446_413#_c_1610_n 8.02119e-19 $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_985 N_A_193_47#_c_1287_n N_A_1446_413#_c_1611_n 0.00120348f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_986 N_A_193_47#_M1008_g N_A_1446_413#_c_1621_n 0.00259696f $X=7.155 $Y=2.275
+ $X2=0 $Y2=0
cc_987 N_A_193_47#_c_1279_n N_A_1446_413#_c_1621_n 9.99101e-19 $X=7.18 $Y=1.29
+ $X2=0 $Y2=0
cc_988 N_A_193_47#_c_1280_n N_A_1446_413#_c_1621_n 7.25987e-19 $X=7.18 $Y=1.35
+ $X2=0 $Y2=0
cc_989 N_A_193_47#_c_1273_n N_A_1446_413#_c_1627_n 4.77975e-19 $X=7.655 $Y=1.29
+ $X2=0 $Y2=0
cc_990 N_A_193_47#_M1012_g N_A_1446_413#_c_1627_n 0.0112915f $X=7.73 $Y=0.415
+ $X2=0 $Y2=0
cc_991 N_A_193_47#_M1012_g N_A_1446_413#_c_1612_n 0.00847049f $X=7.73 $Y=0.415
+ $X2=0 $Y2=0
cc_992 N_A_193_47#_c_1287_n N_A_1446_413#_c_1617_n 0.0041331f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_993 N_A_193_47#_c_1273_n N_A_1446_413#_c_1613_n 5.3564e-19 $X=7.655 $Y=1.29
+ $X2=0 $Y2=0
cc_994 N_A_193_47#_c_1287_n N_A_1446_413#_c_1613_n 0.0376331f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_995 N_A_193_47#_M1018_g N_A_2051_413#_c_1730_n 0.00963552f $X=10.6 $Y=2.275
+ $X2=0 $Y2=0
cc_996 N_A_193_47#_c_1287_n N_A_2051_413#_c_1730_n 0.00391921f $X=10.46 $Y=1.53
+ $X2=0 $Y2=0
cc_997 N_A_193_47#_c_1331_n N_A_2051_413#_c_1730_n 0.00103138f $X=10.605 $Y=1.53
+ $X2=0 $Y2=0
cc_998 N_A_193_47#_c_1278_n N_A_2051_413#_c_1730_n 0.0198599f $X=10.605 $Y=1.53
+ $X2=0 $Y2=0
cc_999 N_A_193_47#_c_1292_n N_A_2051_413#_c_1730_n 0.00303787f $X=10.685 $Y=1.74
+ $X2=0 $Y2=0
cc_1000 N_A_193_47#_c_1275_n N_A_2051_413#_c_1733_n 0.00459251f $X=10.28
+ $Y=0.705 $X2=0 $Y2=0
cc_1001 N_A_193_47#_c_1276_n N_A_2051_413#_c_1733_n 0.0278532f $X=10.39 $Y=0.87
+ $X2=0 $Y2=0
cc_1002 N_A_193_47#_c_1277_n N_A_2051_413#_c_1733_n 0.00108492f $X=10.39 $Y=0.87
+ $X2=0 $Y2=0
cc_1003 N_A_193_47#_c_1276_n N_A_2051_413#_c_1719_n 0.0210561f $X=10.39 $Y=0.87
+ $X2=0 $Y2=0
cc_1004 N_A_193_47#_M1018_g N_A_2051_413#_c_1728_n 0.00365921f $X=10.6 $Y=2.275
+ $X2=0 $Y2=0
cc_1005 N_A_193_47#_c_1331_n N_A_2051_413#_c_1728_n 0.00161073f $X=10.605
+ $Y=1.53 $X2=0 $Y2=0
cc_1006 N_A_193_47#_c_1278_n N_A_2051_413#_c_1728_n 0.0495718f $X=10.605 $Y=1.53
+ $X2=0 $Y2=0
cc_1007 N_A_193_47#_c_1292_n N_A_2051_413#_c_1728_n 0.00182086f $X=10.685
+ $Y=1.74 $X2=0 $Y2=0
cc_1008 N_A_193_47#_c_1276_n N_A_2051_413#_c_1721_n 0.0277807f $X=10.39 $Y=0.87
+ $X2=0 $Y2=0
cc_1009 N_A_193_47#_c_1281_n N_VPWR_c_1824_n 0.012721f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_1010 N_A_193_47#_c_1285_n N_VPWR_c_1825_n 0.00138291f $X=7.04 $Y=1.53 $X2=0
+ $Y2=0
cc_1011 N_A_193_47#_c_1285_n N_VPWR_c_1826_n 7.40558e-19 $X=7.04 $Y=1.53 $X2=0
+ $Y2=0
cc_1012 N_A_193_47#_c_1287_n N_VPWR_c_1828_n 8.15834e-19 $X=10.46 $Y=1.53 $X2=0
+ $Y2=0
cc_1013 N_A_193_47#_c_1281_n N_VPWR_c_1833_n 0.0120448f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_1014 N_A_193_47#_M1018_g N_VPWR_c_1835_n 0.0037981f $X=10.6 $Y=2.275 $X2=0
+ $Y2=0
cc_1015 N_A_193_47#_M1008_g N_VPWR_c_1842_n 0.00564445f $X=7.155 $Y=2.275 $X2=0
+ $Y2=0
cc_1016 N_A_193_47#_M1008_g N_VPWR_c_1823_n 0.00684774f $X=7.155 $Y=2.275 $X2=0
+ $Y2=0
cc_1017 N_A_193_47#_M1018_g N_VPWR_c_1823_n 0.0057367f $X=10.6 $Y=2.275 $X2=0
+ $Y2=0
cc_1018 N_A_193_47#_c_1281_n N_VPWR_c_1823_n 0.00308197f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_1019 N_A_193_47#_c_1285_n N_A_299_47#_c_2016_n 0.0010389f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1020 N_A_193_47#_c_1285_n N_A_299_47#_c_2009_n 0.0170784f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1021 N_A_193_47#_c_1286_n N_A_299_47#_c_2009_n 0.00275409f $X=1.245 $Y=1.53
+ $X2=0 $Y2=0
cc_1022 N_A_193_47#_c_1281_n N_A_299_47#_c_2009_n 0.145237f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_1023 N_A_193_47#_c_1285_n N_A_299_47#_c_2018_n 8.15261e-19 $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1024 N_A_193_47#_c_1285_n N_A_299_47#_c_2010_n 0.0126011f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1025 N_A_193_47#_c_1285_n N_A_299_47#_c_2011_n 0.00275532f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1026 N_A_193_47#_c_1281_n N_A_299_47#_c_2012_n 0.00796831f $X=1.1 $Y=0.51
+ $X2=0 $Y2=0
cc_1027 N_A_193_47#_c_1281_n N_A_299_47#_c_2015_n 0.0117897f $X=1.1 $Y=0.51
+ $X2=0 $Y2=0
cc_1028 N_A_193_47#_c_1285_n N_A_915_47#_c_2138_n 0.00360434f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1029 N_A_193_47#_M1008_g N_A_915_47#_c_2151_n 0.0107721f $X=7.155 $Y=2.275
+ $X2=0 $Y2=0
cc_1030 N_A_193_47#_c_1285_n N_A_915_47#_c_2151_n 4.75993e-19 $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1031 N_A_193_47#_c_1285_n N_A_915_47#_c_2132_n 0.0125927f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1032 N_A_193_47#_c_1285_n N_A_915_47#_c_2133_n 0.00592292f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1033 N_A_193_47#_c_1280_n N_A_915_47#_c_2133_n 0.0419872f $X=7.18 $Y=1.35
+ $X2=0 $Y2=0
cc_1034 N_A_193_47#_M1008_g N_A_915_47#_c_2134_n 0.00298978f $X=7.155 $Y=2.275
+ $X2=0 $Y2=0
cc_1035 N_A_193_47#_c_1285_n N_A_915_47#_c_2134_n 0.0128597f $X=7.04 $Y=1.53
+ $X2=0 $Y2=0
cc_1036 N_A_193_47#_c_1288_n N_A_915_47#_c_2134_n 0.00256294f $X=7.33 $Y=1.53
+ $X2=0 $Y2=0
cc_1037 N_A_193_47#_c_1279_n N_A_915_47#_c_2134_n 0.00514864f $X=7.18 $Y=1.29
+ $X2=0 $Y2=0
cc_1038 N_A_193_47#_c_1279_n N_A_915_47#_c_2137_n 0.00207603f $X=7.18 $Y=1.29
+ $X2=0 $Y2=0
cc_1039 N_A_193_47#_c_1280_n N_A_915_47#_c_2137_n 2.86271e-19 $X=7.18 $Y=1.35
+ $X2=0 $Y2=0
cc_1040 N_A_193_47#_c_1285_n N_VGND_c_2289_n 2.10897e-19 $X=7.04 $Y=1.53 $X2=0
+ $Y2=0
cc_1041 N_A_193_47#_M1012_g N_VGND_c_2290_n 0.00140802f $X=7.73 $Y=0.415 $X2=0
+ $Y2=0
cc_1042 N_A_193_47#_c_1275_n N_VGND_c_2291_n 0.00237285f $X=10.28 $Y=0.705 $X2=0
+ $Y2=0
cc_1043 N_A_193_47#_c_1281_n N_VGND_c_2294_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_1044 N_A_193_47#_c_1275_n N_VGND_c_2300_n 0.00523869f $X=10.28 $Y=0.705 $X2=0
+ $Y2=0
cc_1045 N_A_193_47#_c_1276_n N_VGND_c_2300_n 2.78187e-19 $X=10.39 $Y=0.87 $X2=0
+ $Y2=0
cc_1046 N_A_193_47#_M1012_g N_VGND_c_2306_n 0.00357877f $X=7.73 $Y=0.415 $X2=0
+ $Y2=0
cc_1047 N_A_193_47#_M1021_d N_VGND_c_2308_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_1048 N_A_193_47#_M1012_g N_VGND_c_2308_n 0.00553273f $X=7.73 $Y=0.415 $X2=0
+ $Y2=0
cc_1049 N_A_193_47#_c_1275_n N_VGND_c_2308_n 0.00656556f $X=10.28 $Y=0.705 $X2=0
+ $Y2=0
cc_1050 N_A_193_47#_c_1276_n N_VGND_c_2308_n 0.00106975f $X=10.39 $Y=0.87 $X2=0
+ $Y2=0
cc_1051 N_A_193_47#_c_1281_n N_VGND_c_2308_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_1052 N_A_1610_159#_c_1494_n N_A_1446_413#_c_1607_n 0.00661847f $X=8.83
+ $Y=0.915 $X2=0 $Y2=0
cc_1053 N_A_1610_159#_c_1496_n N_A_1446_413#_c_1607_n 2.83663e-19 $X=9.66
+ $Y=1.21 $X2=0 $Y2=0
cc_1054 N_A_1610_159#_c_1497_n N_A_1446_413#_c_1607_n 0.00149495f $X=9.66
+ $Y=1.21 $X2=0 $Y2=0
cc_1055 N_A_1610_159#_M1006_g N_A_1446_413#_M1017_g 0.0142214f $X=8.125 $Y=2.275
+ $X2=0 $Y2=0
cc_1056 N_A_1610_159#_c_1504_n N_A_1446_413#_M1017_g 0.0168148f $X=8.995 $Y=1.88
+ $X2=0 $Y2=0
cc_1057 N_A_1610_159#_M1019_g N_A_1446_413#_c_1608_n 0.0121471f $X=8.26 $Y=0.445
+ $X2=0 $Y2=0
cc_1058 N_A_1610_159#_c_1492_n N_A_1446_413#_c_1608_n 0.00145117f $X=9.697
+ $Y=1.045 $X2=0 $Y2=0
cc_1059 N_A_1610_159#_c_1494_n N_A_1446_413#_c_1608_n 0.00790103f $X=8.83
+ $Y=0.915 $X2=0 $Y2=0
cc_1060 N_A_1610_159#_c_1495_n N_A_1446_413#_c_1608_n 0.0110908f $X=9.065
+ $Y=0.39 $X2=0 $Y2=0
cc_1061 N_A_1610_159#_c_1499_n N_A_1446_413#_c_1608_n 0.00500472f $X=8.26
+ $Y=0.93 $X2=0 $Y2=0
cc_1062 N_A_1610_159#_M1006_g N_A_1446_413#_c_1609_n 0.00465771f $X=8.125
+ $Y=2.275 $X2=0 $Y2=0
cc_1063 N_A_1610_159#_c_1494_n N_A_1446_413#_c_1609_n 0.0132603f $X=8.83
+ $Y=0.915 $X2=0 $Y2=0
cc_1064 N_A_1610_159#_c_1497_n N_A_1446_413#_c_1609_n 0.00145117f $X=9.66
+ $Y=1.21 $X2=0 $Y2=0
cc_1065 N_A_1610_159#_c_1498_n N_A_1446_413#_c_1609_n 2.46982e-19 $X=8.37
+ $Y=0.93 $X2=0 $Y2=0
cc_1066 N_A_1610_159#_c_1499_n N_A_1446_413#_c_1609_n 0.0049948f $X=8.26 $Y=0.93
+ $X2=0 $Y2=0
cc_1067 N_A_1610_159#_M1006_g N_A_1446_413#_c_1610_n 0.0173823f $X=8.125
+ $Y=2.275 $X2=0 $Y2=0
cc_1068 N_A_1610_159#_c_1494_n N_A_1446_413#_c_1610_n 0.00455719f $X=8.83
+ $Y=0.915 $X2=0 $Y2=0
cc_1069 N_A_1610_159#_c_1499_n N_A_1446_413#_c_1610_n 5.95332e-19 $X=8.26
+ $Y=0.93 $X2=0 $Y2=0
cc_1070 N_A_1610_159#_c_1493_n N_A_1446_413#_c_1611_n 0.00149495f $X=9.662
+ $Y=1.375 $X2=0 $Y2=0
cc_1071 N_A_1610_159#_c_1494_n N_A_1446_413#_c_1611_n 0.00339078f $X=8.83
+ $Y=0.915 $X2=0 $Y2=0
cc_1072 N_A_1610_159#_c_1504_n N_A_1446_413#_c_1611_n 0.0056425f $X=8.995
+ $Y=1.88 $X2=0 $Y2=0
cc_1073 N_A_1610_159#_M1006_g N_A_1446_413#_c_1621_n 0.00989606f $X=8.125
+ $Y=2.275 $X2=0 $Y2=0
cc_1074 N_A_1610_159#_M1019_g N_A_1446_413#_c_1627_n 0.00266694f $X=8.26
+ $Y=0.445 $X2=0 $Y2=0
cc_1075 N_A_1610_159#_M1019_g N_A_1446_413#_c_1612_n 0.00424924f $X=8.26
+ $Y=0.445 $X2=0 $Y2=0
cc_1076 N_A_1610_159#_c_1498_n N_A_1446_413#_c_1612_n 0.0222086f $X=8.37 $Y=0.93
+ $X2=0 $Y2=0
cc_1077 N_A_1610_159#_c_1499_n N_A_1446_413#_c_1612_n 0.00620582f $X=8.26
+ $Y=0.93 $X2=0 $Y2=0
cc_1078 N_A_1610_159#_M1006_g N_A_1446_413#_c_1617_n 0.0163963f $X=8.125
+ $Y=2.275 $X2=0 $Y2=0
cc_1079 N_A_1610_159#_c_1504_n N_A_1446_413#_c_1617_n 0.00686804f $X=8.995
+ $Y=1.88 $X2=0 $Y2=0
cc_1080 N_A_1610_159#_M1006_g N_A_1446_413#_c_1613_n 0.0131936f $X=8.125
+ $Y=2.275 $X2=0 $Y2=0
cc_1081 N_A_1610_159#_c_1494_n N_A_1446_413#_c_1613_n 0.0417632f $X=8.83
+ $Y=0.915 $X2=0 $Y2=0
cc_1082 N_A_1610_159#_c_1498_n N_A_1446_413#_c_1613_n 0.0114411f $X=8.37 $Y=0.93
+ $X2=0 $Y2=0
cc_1083 N_A_1610_159#_c_1499_n N_A_1446_413#_c_1613_n 0.00198791f $X=8.26
+ $Y=0.93 $X2=0 $Y2=0
cc_1084 N_A_1610_159#_M1037_g N_A_2051_413#_c_1730_n 5.6946e-19 $X=9.725
+ $Y=2.275 $X2=0 $Y2=0
cc_1085 N_A_1610_159#_M1039_g N_A_2051_413#_c_1733_n 6.23163e-19 $X=9.795
+ $Y=0.445 $X2=0 $Y2=0
cc_1086 N_A_1610_159#_M1006_g N_VPWR_c_1828_n 0.00644429f $X=8.125 $Y=2.275
+ $X2=0 $Y2=0
cc_1087 N_A_1610_159#_c_1504_n N_VPWR_c_1828_n 0.0249957f $X=8.995 $Y=1.88 $X2=0
+ $Y2=0
cc_1088 N_A_1610_159#_c_1504_n N_VPWR_c_1829_n 0.0210382f $X=8.995 $Y=1.88 $X2=0
+ $Y2=0
cc_1089 N_A_1610_159#_M1037_g N_VPWR_c_1830_n 0.0123787f $X=9.725 $Y=2.275 $X2=0
+ $Y2=0
cc_1090 N_A_1610_159#_c_1504_n N_VPWR_c_1830_n 0.0256005f $X=8.995 $Y=1.88 $X2=0
+ $Y2=0
cc_1091 N_A_1610_159#_M1037_g N_VPWR_c_1835_n 0.00544582f $X=9.725 $Y=2.275
+ $X2=0 $Y2=0
cc_1092 N_A_1610_159#_M1006_g N_VPWR_c_1842_n 0.00375838f $X=8.125 $Y=2.275
+ $X2=0 $Y2=0
cc_1093 N_A_1610_159#_M1017_d N_VPWR_c_1823_n 0.00172424f $X=8.86 $Y=1.735 $X2=0
+ $Y2=0
cc_1094 N_A_1610_159#_M1006_g N_VPWR_c_1823_n 0.0060313f $X=8.125 $Y=2.275 $X2=0
+ $Y2=0
cc_1095 N_A_1610_159#_M1037_g N_VPWR_c_1823_n 0.0052001f $X=9.725 $Y=2.275 $X2=0
+ $Y2=0
cc_1096 N_A_1610_159#_c_1504_n N_VPWR_c_1823_n 0.00592003f $X=8.995 $Y=1.88
+ $X2=0 $Y2=0
cc_1097 N_A_1610_159#_c_1494_n N_VGND_M1019_d 0.00294965f $X=8.83 $Y=0.915 $X2=0
+ $Y2=0
cc_1098 N_A_1610_159#_M1019_g N_VGND_c_2290_n 0.013797f $X=8.26 $Y=0.445 $X2=0
+ $Y2=0
cc_1099 N_A_1610_159#_c_1495_n N_VGND_c_2290_n 0.02237f $X=9.065 $Y=0.39 $X2=0
+ $Y2=0
cc_1100 N_A_1610_159#_c_1498_n N_VGND_c_2290_n 0.0221165f $X=8.37 $Y=0.93 $X2=0
+ $Y2=0
cc_1101 N_A_1610_159#_c_1499_n N_VGND_c_2290_n 4.43315e-19 $X=8.26 $Y=0.93 $X2=0
+ $Y2=0
cc_1102 N_A_1610_159#_M1039_g N_VGND_c_2291_n 0.0133742f $X=9.795 $Y=0.445 $X2=0
+ $Y2=0
cc_1103 N_A_1610_159#_c_1492_n N_VGND_c_2291_n 0.00332209f $X=9.697 $Y=1.045
+ $X2=0 $Y2=0
cc_1104 N_A_1610_159#_c_1495_n N_VGND_c_2291_n 0.0237563f $X=9.065 $Y=0.39 $X2=0
+ $Y2=0
cc_1105 N_A_1610_159#_c_1496_n N_VGND_c_2291_n 0.00471991f $X=9.66 $Y=1.21 $X2=0
+ $Y2=0
cc_1106 N_A_1610_159#_c_1495_n N_VGND_c_2298_n 0.0261692f $X=9.065 $Y=0.39 $X2=0
+ $Y2=0
cc_1107 N_A_1610_159#_M1039_g N_VGND_c_2300_n 0.00505556f $X=9.795 $Y=0.445
+ $X2=0 $Y2=0
cc_1108 N_A_1610_159#_M1019_g N_VGND_c_2306_n 0.00232377f $X=8.26 $Y=0.445 $X2=0
+ $Y2=0
cc_1109 N_A_1610_159#_M1004_d N_VGND_c_2308_n 0.00172424f $X=8.93 $Y=0.235 $X2=0
+ $Y2=0
cc_1110 N_A_1610_159#_M1019_g N_VGND_c_2308_n 0.00261449f $X=8.26 $Y=0.445 $X2=0
+ $Y2=0
cc_1111 N_A_1610_159#_M1039_g N_VGND_c_2308_n 0.00494779f $X=9.795 $Y=0.445
+ $X2=0 $Y2=0
cc_1112 N_A_1610_159#_c_1494_n N_VGND_c_2308_n 0.00432725f $X=8.83 $Y=0.915
+ $X2=0 $Y2=0
cc_1113 N_A_1610_159#_c_1495_n N_VGND_c_2308_n 0.00714477f $X=9.065 $Y=0.39
+ $X2=0 $Y2=0
cc_1114 N_A_1610_159#_c_1498_n N_VGND_c_2308_n 0.00255175f $X=8.37 $Y=0.93 $X2=0
+ $Y2=0
cc_1115 N_A_1610_159#_c_1499_n N_VGND_c_2308_n 7.19298e-19 $X=8.26 $Y=0.93 $X2=0
+ $Y2=0
cc_1116 N_A_1446_413#_M1017_g N_VPWR_c_1828_n 0.0032365f $X=8.785 $Y=2.11 $X2=0
+ $Y2=0
cc_1117 N_A_1446_413#_c_1610_n N_VPWR_c_1828_n 0.00132475f $X=8.71 $Y=1.41 $X2=0
+ $Y2=0
cc_1118 N_A_1446_413#_c_1617_n N_VPWR_c_1828_n 0.0209688f $X=8.17 $Y=2.175 $X2=0
+ $Y2=0
cc_1119 N_A_1446_413#_c_1613_n N_VPWR_c_1828_n 0.0108482f $X=8.17 $Y=1.41 $X2=0
+ $Y2=0
cc_1120 N_A_1446_413#_M1017_g N_VPWR_c_1829_n 0.00541359f $X=8.785 $Y=2.11 $X2=0
+ $Y2=0
cc_1121 N_A_1446_413#_M1017_g N_VPWR_c_1830_n 0.00292103f $X=8.785 $Y=2.11 $X2=0
+ $Y2=0
cc_1122 N_A_1446_413#_c_1621_n N_VPWR_c_1842_n 0.0372444f $X=8.085 $Y=2.275
+ $X2=0 $Y2=0
cc_1123 N_A_1446_413#_M1008_d N_VPWR_c_1823_n 0.00206096f $X=7.23 $Y=2.065 $X2=0
+ $Y2=0
cc_1124 N_A_1446_413#_M1017_g N_VPWR_c_1823_n 0.00782689f $X=8.785 $Y=2.11 $X2=0
+ $Y2=0
cc_1125 N_A_1446_413#_c_1621_n N_VPWR_c_1823_n 0.0160193f $X=8.085 $Y=2.275
+ $X2=0 $Y2=0
cc_1126 N_A_1446_413#_c_1621_n N_A_915_47#_c_2155_n 0.0138511f $X=8.085 $Y=2.275
+ $X2=0 $Y2=0
cc_1127 N_A_1446_413#_c_1627_n N_A_915_47#_c_2168_n 5.93115e-19 $X=7.81 $Y=0.41
+ $X2=0 $Y2=0
cc_1128 N_A_1446_413#_c_1627_n N_A_915_47#_c_2137_n 0.0263002f $X=7.81 $Y=0.41
+ $X2=0 $Y2=0
cc_1129 N_A_1446_413#_c_1621_n A_1537_413# 0.00553919f $X=8.085 $Y=2.275
+ $X2=-0.19 $Y2=-0.24
cc_1130 N_A_1446_413#_c_1608_n N_VGND_c_2290_n 0.00570804f $X=8.82 $Y=0.95 $X2=0
+ $Y2=0
cc_1131 N_A_1446_413#_c_1627_n N_VGND_c_2290_n 0.0181194f $X=7.81 $Y=0.41 $X2=0
+ $Y2=0
cc_1132 N_A_1446_413#_c_1608_n N_VGND_c_2291_n 0.00214573f $X=8.82 $Y=0.95 $X2=0
+ $Y2=0
cc_1133 N_A_1446_413#_c_1608_n N_VGND_c_2298_n 0.00435091f $X=8.82 $Y=0.95 $X2=0
+ $Y2=0
cc_1134 N_A_1446_413#_c_1627_n N_VGND_c_2306_n 0.0393557f $X=7.81 $Y=0.41 $X2=0
+ $Y2=0
cc_1135 N_A_1446_413#_M1027_d N_VGND_c_2308_n 0.00190253f $X=7.365 $Y=0.235
+ $X2=0 $Y2=0
cc_1136 N_A_1446_413#_c_1608_n N_VGND_c_2308_n 0.00708984f $X=8.82 $Y=0.95 $X2=0
+ $Y2=0
cc_1137 N_A_1446_413#_c_1627_n N_VGND_c_2308_n 0.0114791f $X=7.81 $Y=0.41 $X2=0
+ $Y2=0
cc_1138 N_A_1446_413#_c_1627_n A_1561_47# 0.00436463f $X=7.81 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1139 N_A_1446_413#_c_1612_n A_1561_47# 0.00105811f $X=7.895 $Y=1.315
+ $X2=-0.19 $Y2=-0.24
cc_1140 N_A_2051_413#_c_1730_n N_VPWR_c_1830_n 0.00551479f $X=10.94 $Y=2.26
+ $X2=0 $Y2=0
cc_1141 N_A_2051_413#_M1023_g N_VPWR_c_1831_n 0.00188178f $X=12.225 $Y=2.165
+ $X2=0 $Y2=0
cc_1142 N_A_2051_413#_M1023_g N_VPWR_c_1832_n 0.00910498f $X=12.225 $Y=2.165
+ $X2=0 $Y2=0
cc_1143 N_A_2051_413#_c_1714_n N_VPWR_c_1832_n 0.00466622f $X=12.635 $Y=1.16
+ $X2=0 $Y2=0
cc_1144 N_A_2051_413#_M1010_g N_VPWR_c_1832_n 0.00310362f $X=12.71 $Y=1.985
+ $X2=0 $Y2=0
cc_1145 N_A_2051_413#_c_1730_n N_VPWR_c_1835_n 0.0295685f $X=10.94 $Y=2.26 $X2=0
+ $Y2=0
cc_1146 N_A_2051_413#_M1023_g N_VPWR_c_1837_n 0.00541359f $X=12.225 $Y=2.165
+ $X2=0 $Y2=0
cc_1147 N_A_2051_413#_M1010_g N_VPWR_c_1843_n 0.00557712f $X=12.71 $Y=1.985
+ $X2=0 $Y2=0
cc_1148 N_A_2051_413#_M1025_d N_VPWR_c_1823_n 0.00215743f $X=10.255 $Y=2.065
+ $X2=0 $Y2=0
cc_1149 N_A_2051_413#_M1023_g N_VPWR_c_1823_n 0.0110723f $X=12.225 $Y=2.165
+ $X2=0 $Y2=0
cc_1150 N_A_2051_413#_M1010_g N_VPWR_c_1823_n 0.0110874f $X=12.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1151 N_A_2051_413#_c_1730_n N_VPWR_c_1823_n 0.0280716f $X=10.94 $Y=2.26 $X2=0
+ $Y2=0
cc_1152 N_A_2051_413#_c_1730_n A_2135_413# 0.00905112f $X=10.94 $Y=2.26
+ $X2=-0.19 $Y2=-0.24
cc_1153 N_A_2051_413#_c_1728_n A_2135_413# 0.00123507f $X=11.025 $Y=2.165
+ $X2=-0.19 $Y2=-0.24
cc_1154 N_A_2051_413#_M1031_g N_Q_c_2269_n 4.27936e-19 $X=12.225 $Y=0.445 $X2=0
+ $Y2=0
cc_1155 N_A_2051_413#_M1023_g N_Q_c_2269_n 6.50973e-19 $X=12.225 $Y=2.165 $X2=0
+ $Y2=0
cc_1156 N_A_2051_413#_c_1715_n N_Q_c_2269_n 0.00994181f $X=12.71 $Y=0.995 $X2=0
+ $Y2=0
cc_1157 N_A_2051_413#_M1010_g N_Q_c_2269_n 0.0153574f $X=12.71 $Y=1.985 $X2=0
+ $Y2=0
cc_1158 N_A_2051_413#_c_1718_n N_Q_c_2269_n 0.0164431f $X=12.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1159 N_A_2051_413#_c_1733_n N_VGND_c_2291_n 0.00574753f $X=10.94 $Y=0.432
+ $X2=0 $Y2=0
cc_1160 N_A_2051_413#_M1031_g N_VGND_c_2292_n 0.00357154f $X=12.225 $Y=0.445
+ $X2=0 $Y2=0
cc_1161 N_A_2051_413#_c_1716_n N_VGND_c_2292_n 0.00151274f $X=12.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1162 N_A_2051_413#_c_1733_n N_VGND_c_2292_n 0.0129405f $X=10.94 $Y=0.432
+ $X2=0 $Y2=0
cc_1163 N_A_2051_413#_c_1719_n N_VGND_c_2292_n 0.00448678f $X=11.025 $Y=0.995
+ $X2=0 $Y2=0
cc_1164 N_A_2051_413#_c_1720_n N_VGND_c_2292_n 0.00691913f $X=11.725 $Y=1.16
+ $X2=0 $Y2=0
cc_1165 N_A_2051_413#_M1031_g N_VGND_c_2293_n 0.0069333f $X=12.225 $Y=0.445
+ $X2=0 $Y2=0
cc_1166 N_A_2051_413#_c_1714_n N_VGND_c_2293_n 0.00495621f $X=12.635 $Y=1.16
+ $X2=0 $Y2=0
cc_1167 N_A_2051_413#_c_1715_n N_VGND_c_2293_n 0.00306265f $X=12.71 $Y=0.995
+ $X2=0 $Y2=0
cc_1168 N_A_2051_413#_c_1733_n N_VGND_c_2300_n 0.0312214f $X=10.94 $Y=0.432
+ $X2=0 $Y2=0
cc_1169 N_A_2051_413#_M1031_g N_VGND_c_2302_n 0.00543148f $X=12.225 $Y=0.445
+ $X2=0 $Y2=0
cc_1170 N_A_2051_413#_c_1715_n N_VGND_c_2307_n 0.00557839f $X=12.71 $Y=0.995
+ $X2=0 $Y2=0
cc_1171 N_A_2051_413#_M1026_d N_VGND_c_2308_n 0.00256476f $X=10.355 $Y=0.235
+ $X2=0 $Y2=0
cc_1172 N_A_2051_413#_M1031_g N_VGND_c_2308_n 0.00952759f $X=12.225 $Y=0.445
+ $X2=0 $Y2=0
cc_1173 N_A_2051_413#_c_1715_n N_VGND_c_2308_n 0.0110878f $X=12.71 $Y=0.995
+ $X2=0 $Y2=0
cc_1174 N_A_2051_413#_c_1733_n N_VGND_c_2308_n 0.0125713f $X=10.94 $Y=0.432
+ $X2=0 $Y2=0
cc_1175 N_A_2051_413#_c_1733_n A_2177_47# 0.00443949f $X=10.94 $Y=0.432
+ $X2=-0.19 $Y2=-0.24
cc_1176 N_A_2051_413#_c_1719_n A_2177_47# 0.00147825f $X=11.025 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_1177 N_VPWR_c_1823_n N_A_299_47#_M1029_s 0.00172424f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1178 N_VPWR_c_1823_n N_A_299_47#_M1036_d 0.00205179f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1179 N_VPWR_c_1825_n N_A_299_47#_c_2016_n 0.0192069f $X=2.4 $Y=2 $X2=0 $Y2=0
cc_1180 N_VPWR_c_1833_n N_A_299_47#_c_2016_n 0.0280365f $X=2.235 $Y=2.72 $X2=0
+ $Y2=0
cc_1181 N_VPWR_c_1823_n N_A_299_47#_c_2016_n 0.00771147f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1182 N_VPWR_c_1826_n N_A_299_47#_c_2018_n 0.00729213f $X=3.35 $Y=1.99 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1841_n N_A_299_47#_c_2018_n 0.0201764f $X=5.665 $Y=2.72 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1823_n N_A_299_47#_c_2018_n 0.00655199f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1823_n A_381_369# 0.00302076f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1186 N_VPWR_c_1823_n A_729_369# 0.00517845f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1187 N_VPWR_c_1823_n N_A_915_47#_M1013_d 0.0022185f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1823_n N_A_915_47#_M1030_d 0.00384946f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1841_n N_A_915_47#_c_2140_n 0.0218032f $X=5.665 $Y=2.72 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1823_n N_A_915_47#_c_2140_n 0.0059727f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1842_n N_A_915_47#_c_2155_n 0.0222204f $X=8.425 $Y=2.72 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1823_n N_A_915_47#_c_2155_n 0.00594985f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1823_n A_1231_369# 0.00309589f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1194 N_VPWR_c_1823_n A_1537_413# 0.00247765f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1195 N_VPWR_c_1823_n A_1960_413# 0.0042834f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1196 N_VPWR_c_1823_n A_2135_413# 0.00357865f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1197 N_VPWR_c_1823_n N_Q_M1010_d 0.00228626f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1198 N_VPWR_c_1832_n N_Q_c_2269_n 0.0365895f $X=12.5 $Y=1.63 $X2=0 $Y2=0
cc_1199 N_VPWR_c_1843_n N_Q_c_2269_n 0.0163462f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1200 N_VPWR_c_1823_n N_Q_c_2269_n 0.0121893f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1201 N_VPWR_c_1832_n N_VGND_c_2293_n 0.00976036f $X=12.5 $Y=1.63 $X2=0 $Y2=0
cc_1202 N_A_299_47#_c_2010_n N_A_915_47#_c_2138_n 0.025473f $X=4.32 $Y=1.82
+ $X2=0 $Y2=0
cc_1203 N_A_299_47#_c_2018_n N_A_915_47#_c_2139_n 0.025473f $X=4.29 $Y=2 $X2=0
+ $Y2=0
cc_1204 N_A_299_47#_c_2011_n N_A_915_47#_c_2132_n 0.025473f $X=4.33 $Y=1.15
+ $X2=0 $Y2=0
cc_1205 N_A_299_47#_c_2014_n N_A_915_47#_c_2132_n 0.0073483f $X=4.29 $Y=0.445
+ $X2=0 $Y2=0
cc_1206 N_A_299_47#_c_2040_n N_A_915_47#_c_2135_n 0.0258206f $X=4.27 $Y=0.51
+ $X2=0 $Y2=0
cc_1207 N_A_299_47#_c_2014_n N_A_915_47#_c_2135_n 8.1654e-19 $X=4.29 $Y=0.445
+ $X2=0 $Y2=0
cc_1208 N_A_299_47#_c_2040_n N_A_915_47#_c_2192_n 8.32699e-19 $X=4.27 $Y=0.51
+ $X2=0 $Y2=0
cc_1209 N_A_299_47#_c_2014_n N_A_915_47#_c_2192_n 0.0200497f $X=4.29 $Y=0.445
+ $X2=0 $Y2=0
cc_1210 N_A_299_47#_c_2013_n N_VGND_M1003_d 0.00213973f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_1211 N_A_299_47#_c_2015_n N_VGND_c_2286_n 0.00316681f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_1212 N_A_299_47#_c_2013_n N_VGND_c_2287_n 0.0145222f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_1213 N_A_299_47#_c_2015_n N_VGND_c_2287_n 0.0070895f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_1214 N_A_299_47#_c_2040_n N_VGND_c_2288_n 5.24197e-19 $X=4.27 $Y=0.51 $X2=0
+ $Y2=0
cc_1215 N_A_299_47#_c_2013_n N_VGND_c_2288_n 0.0213503f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_1216 N_A_299_47#_c_2014_n N_VGND_c_2288_n 0.0056261f $X=4.29 $Y=0.445 $X2=0
+ $Y2=0
cc_1217 N_A_299_47#_c_2012_n N_VGND_c_2294_n 6.17783e-19 $X=1.585 $Y=0.51 $X2=0
+ $Y2=0
cc_1218 N_A_299_47#_c_2013_n N_VGND_c_2294_n 0.00229575f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_1219 N_A_299_47#_c_2015_n N_VGND_c_2294_n 0.0264163f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_1220 N_A_299_47#_c_2013_n N_VGND_c_2296_n 0.00288773f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_1221 N_A_299_47#_c_2014_n N_VGND_c_2296_n 0.0152055f $X=4.29 $Y=0.445 $X2=0
+ $Y2=0
cc_1222 N_A_299_47#_c_2013_n N_VGND_c_2305_n 0.00219701f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_1223 N_A_299_47#_M1002_s N_VGND_c_2308_n 0.00110044f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_1224 N_A_299_47#_M1041_d N_VGND_c_2308_n 0.00123074f $X=4.155 $Y=0.235 $X2=0
+ $Y2=0
cc_1225 N_A_299_47#_c_2012_n N_VGND_c_2308_n 0.305313f $X=1.585 $Y=0.51 $X2=0
+ $Y2=0
cc_1226 N_A_299_47#_c_2014_n N_VGND_c_2308_n 0.00257571f $X=4.29 $Y=0.445 $X2=0
+ $Y2=0
cc_1227 N_A_299_47#_c_2015_n N_VGND_c_2308_n 0.00373095f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_1228 N_A_299_47#_c_2013_n A_381_47# 0.00879585f $X=4.125 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_1229 N_A_299_47#_c_2013_n A_729_47# 0.00632255f $X=4.125 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_1230 N_A_915_47#_c_2130_n N_VGND_c_2289_n 0.00495078f $X=6.72 $Y=0.98 $X2=0
+ $Y2=0
cc_1231 N_A_915_47#_c_2168_n N_VGND_c_2289_n 8.90737e-19 $X=6.615 $Y=0.51 $X2=0
+ $Y2=0
cc_1232 N_A_915_47#_c_2136_n N_VGND_c_2289_n 0.0181298f $X=6.47 $Y=0.51 $X2=0
+ $Y2=0
cc_1233 N_A_915_47#_c_2137_n N_VGND_c_2289_n 0.00906279f $X=6.97 $Y=0.41 $X2=0
+ $Y2=0
cc_1234 N_A_915_47#_c_2131_n N_VGND_c_2296_n 9.76595e-19 $X=4.725 $Y=0.825 $X2=0
+ $Y2=0
cc_1235 N_A_915_47#_c_2135_n N_VGND_c_2296_n 0.0011212f $X=4.845 $Y=0.51 $X2=0
+ $Y2=0
cc_1236 N_A_915_47#_c_2136_n N_VGND_c_2296_n 0.00128268f $X=6.47 $Y=0.51 $X2=0
+ $Y2=0
cc_1237 N_A_915_47#_c_2192_n N_VGND_c_2296_n 0.0126216f $X=4.71 $Y=0.445 $X2=0
+ $Y2=0
cc_1238 N_A_915_47#_c_2136_n N_VGND_c_2306_n 0.00262344f $X=6.47 $Y=0.51 $X2=0
+ $Y2=0
cc_1239 N_A_915_47#_c_2137_n N_VGND_c_2306_n 0.0410021f $X=6.97 $Y=0.41 $X2=0
+ $Y2=0
cc_1240 N_A_915_47#_M1034_d N_VGND_c_2308_n 0.00123805f $X=4.575 $Y=0.235 $X2=0
+ $Y2=0
cc_1241 N_A_915_47#_M1009_d N_VGND_c_2308_n 0.00411937f $X=6.49 $Y=0.595 $X2=0
+ $Y2=0
cc_1242 N_A_915_47#_c_2135_n N_VGND_c_2308_n 0.215868f $X=4.845 $Y=0.51 $X2=0
+ $Y2=0
cc_1243 N_A_915_47#_c_2192_n N_VGND_c_2308_n 0.00190201f $X=4.71 $Y=0.445 $X2=0
+ $Y2=0
cc_1244 N_A_915_47#_c_2137_n N_VGND_c_2308_n 0.00878695f $X=6.97 $Y=0.41 $X2=0
+ $Y2=0
cc_1245 N_Q_c_2269_n N_VGND_c_2293_n 0.022497f $X=12.93 $Y=0.395 $X2=0 $Y2=0
cc_1246 N_Q_c_2269_n N_VGND_c_2307_n 0.0159484f $X=12.93 $Y=0.395 $X2=0 $Y2=0
cc_1247 N_Q_M1035_d N_VGND_c_2308_n 0.00229159f $X=12.785 $Y=0.235 $X2=0 $Y2=0
cc_1248 N_Q_c_2269_n N_VGND_c_2308_n 0.0121559f $X=12.93 $Y=0.395 $X2=0 $Y2=0
cc_1249 N_VGND_c_2308_n A_381_47# 0.00172536f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1250 N_VGND_c_2308_n A_729_47# 0.0025277f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1251 N_VGND_c_2308_n A_1561_47# 0.00379452f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1252 N_VGND_c_2308_n A_1974_47# 0.00481883f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1253 N_VGND_c_2308_n A_2177_47# 0.00296047f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__dlymetal6s6s_1.pex.spice
* Created: Tue Sep  1 19:07:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A 3 7 9 10 15 17
c31 17 0 1.57226e-19 $X=0.65 $Y=1.16
r32 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.425 $Y=1.16
+ $X2=0.65 $Y2=1.16
r33 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.425
+ $Y=1.16 $X2=0.425 $Y2=1.16
r34 9 10 8.29932 $w=4.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.33 $Y=1.19 $X2=0.33
+ $Y2=1.53
r35 9 15 0.732293 $w=4.88e-07 $l=3e-08 $layer=LI1_cond $X=0.33 $Y=1.19 $X2=0.33
+ $Y2=1.16
r36 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.325
+ $X2=0.65 $Y2=1.16
r37 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.65 $Y=1.325 $X2=0.65
+ $Y2=2.275
r38 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=0.995
+ $X2=0.65 $Y2=1.16
r39 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.65 $Y=0.995 $X2=0.65
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_63_47# 1 2 9 12 14 16 21 23 27 33
+ 34 35 38
c60 33 0 1.1704e-19 $X=1.07 $Y=1.16
c61 16 0 1.57226e-19 $X=0.745 $Y=1.955
r62 34 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.16
+ $X2=1.07 $Y2=1.325
r63 34 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.16
+ $X2=1.07 $Y2=0.995
r64 33 36 5.05753 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=1.325
r65 33 35 5.05753 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=0.995
r66 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.16 $X2=1.07 $Y2=1.16
r67 27 30 8.3814 $w=4.38e-07 $l=3.2e-07 $layer=LI1_cond $X=0.305 $Y=1.955
+ $X2=0.305 $Y2=2.275
r68 23 25 7.72661 $w=4.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.305 $Y=0.445
+ $X2=0.305 $Y2=0.74
r69 21 36 18.7487 $w=3.33e-07 $l=5.45e-07 $layer=LI1_cond $X=0.912 $Y=1.87
+ $X2=0.912 $Y2=1.325
r70 18 35 5.84822 $w=3.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.912 $Y=0.825
+ $X2=0.912 $Y2=0.995
r71 17 27 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=1.955
+ $X2=0.305 $Y2=1.955
r72 16 21 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=0.745 $Y=1.955
+ $X2=0.912 $Y2=1.87
r73 16 17 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.745 $Y=1.955
+ $X2=0.525 $Y2=1.955
r74 15 25 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=0.74
+ $X2=0.305 $Y2=0.74
r75 14 18 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=0.745 $Y=0.74
+ $X2=0.912 $Y2=0.825
r76 14 15 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.745 $Y=0.74
+ $X2=0.525 $Y2=0.74
r77 12 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.125 $Y=1.985
+ $X2=1.125 $Y2=1.325
r78 9 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.125 $Y=0.56
+ $X2=1.125 $Y2=0.995
r79 2 30 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=2.065 $X2=0.44 $Y2=2.275
r80 1 23 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.315
+ $Y=0.235 $X2=0.44 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_240_47# 1 2 9 13 17 19 21 24 25 31
r55 28 31 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=2.065 $Y2=1.16
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.84
+ $Y=1.16 $X2=1.84 $Y2=1.16
r57 24 27 9.80533 $w=6.69e-07 $l=2.59711e-07 $layer=LI1_cond $X=1.422 $Y=0.995
+ $X2=1.612 $Y2=1.16
r58 24 25 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=1.422 $Y=0.995
+ $X2=1.422 $Y2=0.825
r59 19 27 13.8675 $w=6.69e-07 $l=6.18167e-07 $layer=LI1_cond $X=1.385 $Y=1.675
+ $X2=1.612 $Y2=1.16
r60 19 21 12.1647 $w=2.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.385 $Y=1.675
+ $X2=1.385 $Y2=1.96
r61 15 25 6.67067 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.385 $Y=0.69
+ $X2=1.385 $Y2=0.825
r62 15 17 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.385 $Y=0.69
+ $X2=1.385 $Y2=0.44
r63 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.325
+ $X2=2.065 $Y2=1.16
r64 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.065 $Y=1.325
+ $X2=2.065 $Y2=2.275
r65 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=0.995
+ $X2=2.065 $Y2=1.16
r66 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.065 $Y=0.995
+ $X2=2.065 $Y2=0.445
r67 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.2
+ $Y=1.485 $X2=1.335 $Y2=1.96
r68 1 17 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.235 $X2=1.335 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_346_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c69 26 0 1.27733e-19 $X=2.32 $Y=1.325
r70 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.16
+ $X2=2.485 $Y2=1.325
r71 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.16
+ $X2=2.485 $Y2=0.995
r72 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.16 $X2=2.485 $Y2=1.16
r73 28 30 13.2746 $w=3.86e-07 $l=4.2e-07 $layer=LI1_cond $X=2.357 $Y=0.74
+ $X2=2.357 $Y2=1.16
r74 26 30 5.34605 $w=3.86e-07 $l=1.82565e-07 $layer=LI1_cond $X=2.32 $Y=1.325
+ $X2=2.357 $Y2=1.16
r75 26 27 17.122 $w=3.48e-07 $l=5.2e-07 $layer=LI1_cond $X=2.32 $Y=1.325
+ $X2=2.32 $Y2=1.845
r76 24 27 7.55928 $w=1.95e-07 $l=2.18174e-07 $layer=LI1_cond $X=2.145 $Y=1.942
+ $X2=2.32 $Y2=1.845
r77 24 25 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=2.145 $Y=1.942
+ $X2=1.94 $Y2=1.942
r78 22 28 5.5624 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.145 $Y=0.74
+ $X2=2.357 $Y2=0.74
r79 22 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.145 $Y=0.74
+ $X2=1.94 $Y2=0.74
r80 18 25 6.9528 $w=1.95e-07 $l=1.66958e-07 $layer=LI1_cond $X=1.815 $Y=2.04
+ $X2=1.94 $Y2=1.942
r81 18 20 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=1.815 $Y=2.04
+ $X2=1.815 $Y2=2.275
r82 14 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.815 $Y=0.655
+ $X2=1.94 $Y2=0.74
r83 14 16 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.815 $Y=0.655
+ $X2=1.815 $Y2=0.44
r84 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.54 $Y=1.985
+ $X2=2.54 $Y2=1.325
r85 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.54 $Y=0.56 $X2=2.54
+ $Y2=0.995
r86 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=2.065 $X2=1.855 $Y2=2.275
r87 1 16 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.73
+ $Y=0.235 $X2=1.855 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_523_47# 1 2 9 13 17 19 21 24 25 31
r55 28 31 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.255 $Y=1.16
+ $X2=3.48 $Y2=1.16
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.255
+ $Y=1.16 $X2=3.255 $Y2=1.16
r57 24 27 10.6023 $w=6.69e-07 $l=2.70185e-07 $layer=LI1_cond $X=2.827 $Y=0.995
+ $X2=3.027 $Y2=1.16
r58 24 25 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=2.827 $Y=0.995
+ $X2=2.827 $Y2=0.825
r59 19 27 14.4032 $w=6.69e-07 $l=6.22318e-07 $layer=LI1_cond $X=2.79 $Y=1.675
+ $X2=3.027 $Y2=1.16
r60 19 21 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=2.79 $Y=1.675
+ $X2=2.79 $Y2=1.96
r61 15 25 6.81244 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.79 $Y=0.7
+ $X2=2.79 $Y2=0.825
r62 15 17 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.79 $Y=0.7 $X2=2.79
+ $Y2=0.44
r63 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.325
+ $X2=3.48 $Y2=1.16
r64 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.48 $Y=1.325
+ $X2=3.48 $Y2=2.275
r65 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=0.995
+ $X2=3.48 $Y2=1.16
r66 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.48 $Y=0.995 $X2=3.48
+ $Y2=0.445
r67 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.615
+ $Y=1.485 $X2=2.75 $Y2=1.96
r68 1 17 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.235 $X2=2.75 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_629_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c66 26 0 1.27733e-19 $X=3.735 $Y=1.325
r67 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.16 $X2=3.9
+ $Y2=1.325
r68 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.16 $X2=3.9
+ $Y2=0.995
r69 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9
+ $Y=1.16 $X2=3.9 $Y2=1.16
r70 28 30 13.2746 $w=3.86e-07 $l=4.2e-07 $layer=LI1_cond $X=3.772 $Y=0.74
+ $X2=3.772 $Y2=1.16
r71 26 30 5.34605 $w=3.86e-07 $l=1.82565e-07 $layer=LI1_cond $X=3.735 $Y=1.325
+ $X2=3.772 $Y2=1.16
r72 26 27 17.122 $w=3.48e-07 $l=5.2e-07 $layer=LI1_cond $X=3.735 $Y=1.325
+ $X2=3.735 $Y2=1.845
r73 24 27 7.55928 $w=1.95e-07 $l=2.18174e-07 $layer=LI1_cond $X=3.56 $Y=1.942
+ $X2=3.735 $Y2=1.845
r74 24 25 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.56 $Y=1.942
+ $X2=3.355 $Y2=1.942
r75 22 28 5.5624 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.56 $Y=0.74
+ $X2=3.772 $Y2=0.74
r76 22 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.56 $Y=0.74
+ $X2=3.355 $Y2=0.74
r77 18 25 7.04969 $w=1.95e-07 $l=1.77356e-07 $layer=LI1_cond $X=3.22 $Y=2.04
+ $X2=3.355 $Y2=1.942
r78 18 20 10.0305 $w=2.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.22 $Y=2.04
+ $X2=3.22 $Y2=2.275
r79 14 23 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.22 $Y=0.655
+ $X2=3.355 $Y2=0.74
r80 14 16 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.22 $Y=0.655
+ $X2=3.22 $Y2=0.44
r81 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.955 $Y=1.985
+ $X2=3.955 $Y2=1.325
r82 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.955 $Y=0.56
+ $X2=3.955 $Y2=0.995
r83 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=2.065 $X2=3.27 $Y2=2.275
r84 1 16 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.27 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%VPWR 1 2 3 12 16 20 23 24 26 27 29 30
+ 31 50 51 56
r63 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r64 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r65 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 44 47 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 42 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r71 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r72 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r73 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 35 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 35 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 31 56 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 29 47 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.525 $Y=2.72
+ $X2=3.45 $Y2=2.72
r79 29 30 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.525 $Y=2.72
+ $X2=3.717 $Y2=2.72
r80 28 50 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r81 28 30 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=3.717 $Y2=2.72
r82 26 41 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.11 $Y=2.72 $X2=2.07
+ $Y2=2.72
r83 26 27 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.11 $Y=2.72
+ $X2=2.302 $Y2=2.72
r84 25 44 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.495 $Y=2.72
+ $X2=2.53 $Y2=2.72
r85 25 27 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.495 $Y=2.72
+ $X2=2.302 $Y2=2.72
r86 23 34 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=0.69 $Y2=2.72
r87 23 24 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.695 $Y=2.72
+ $X2=0.887 $Y2=2.72
r88 22 38 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.08 $Y=2.72 $X2=1.15
+ $Y2=2.72
r89 22 24 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.08 $Y=2.72
+ $X2=0.887 $Y2=2.72
r90 18 30 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.717 $Y=2.635
+ $X2=3.717 $Y2=2.72
r91 18 20 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.717 $Y=2.635
+ $X2=3.717 $Y2=2.36
r92 14 27 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.302 $Y=2.635
+ $X2=2.302 $Y2=2.72
r93 14 16 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=2.302 $Y=2.635
+ $X2=2.302 $Y2=2.36
r94 10 24 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.887 $Y=2.635
+ $X2=0.887 $Y2=2.72
r95 10 12 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=0.887 $Y=2.635
+ $X2=0.887 $Y2=2.36
r96 3 20 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=2.065 $X2=3.72 $Y2=2.36
r97 2 16 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=2.065 $X2=2.305 $Y2=2.36
r98 1 12 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=0.725
+ $Y=2.065 $X2=0.89 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%X 1 2 7 8 9 10 11 12 24 38 45
r16 45 46 1.30392 $w=4.33e-07 $l=3.5e-08 $layer=LI1_cond $X=4.297 $Y=1.53
+ $X2=4.297 $Y2=1.495
r17 24 43 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=4.335 $Y=0.85
+ $X2=4.335 $Y2=0.825
r18 12 33 6.62324 $w=4.33e-07 $l=2.5e-07 $layer=LI1_cond $X=4.297 $Y=2.21
+ $X2=4.297 $Y2=1.96
r19 11 33 2.38436 $w=4.33e-07 $l=9e-08 $layer=LI1_cond $X=4.297 $Y=1.87
+ $X2=4.297 $Y2=1.96
r20 11 29 4.18588 $w=4.33e-07 $l=1.58e-07 $layer=LI1_cond $X=4.297 $Y=1.87
+ $X2=4.297 $Y2=1.712
r21 10 29 4.15939 $w=4.33e-07 $l=1.57e-07 $layer=LI1_cond $X=4.297 $Y=1.555
+ $X2=4.297 $Y2=1.712
r22 10 45 0.662324 $w=4.33e-07 $l=2.5e-08 $layer=LI1_cond $X=4.297 $Y=1.555
+ $X2=4.297 $Y2=1.53
r23 10 46 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=4.335 $Y=1.47
+ $X2=4.335 $Y2=1.495
r24 9 10 8.96345 $w=3.58e-07 $l=2.8e-07 $layer=LI1_cond $X=4.335 $Y=1.19
+ $X2=4.335 $Y2=1.47
r25 8 43 1.17145 $w=4.33e-07 $l=3e-08 $layer=LI1_cond $X=4.297 $Y=0.795
+ $X2=4.297 $Y2=0.825
r26 8 9 9.92381 $w=3.58e-07 $l=3.1e-07 $layer=LI1_cond $X=4.335 $Y=0.88
+ $X2=4.335 $Y2=1.19
r27 8 24 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=4.335 $Y=0.88
+ $X2=4.335 $Y2=0.85
r28 7 8 7.55049 $w=4.33e-07 $l=2.85e-07 $layer=LI1_cond $X=4.297 $Y=0.51
+ $X2=4.297 $Y2=0.795
r29 7 38 1.85451 $w=4.33e-07 $l=7e-08 $layer=LI1_cond $X=4.297 $Y=0.51 $X2=4.297
+ $Y2=0.44
r30 2 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.03
+ $Y=1.485 $X2=4.165 $Y2=1.96
r31 1 38 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.235 $X2=4.165 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%VGND 1 2 3 12 16 20 23 24 26 27 29 30
+ 31 50 51 56
r66 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r67 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r68 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r69 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r70 44 47 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r71 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r72 42 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r73 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r74 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r75 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r76 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r77 35 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r78 35 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r79 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r80 31 56 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=0 $X2=0.23
+ $Y2=0
r81 29 47 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.45
+ $Y2=0
r82 29 30 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.717
+ $Y2=0
r83 28 50 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r84 28 30 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=3.717
+ $Y2=0
r85 26 41 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.07
+ $Y2=0
r86 26 27 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.302
+ $Y2=0
r87 25 44 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.53
+ $Y2=0
r88 25 27 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.302
+ $Y2=0
r89 23 34 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.695 $Y=0 $X2=0.69
+ $Y2=0
r90 23 24 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.695 $Y=0 $X2=0.887
+ $Y2=0
r91 22 38 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.08 $Y=0 $X2=1.15
+ $Y2=0
r92 22 24 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.887
+ $Y2=0
r93 18 30 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.717 $Y=0.085
+ $X2=3.717 $Y2=0
r94 18 20 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=3.717 $Y=0.085
+ $X2=3.717 $Y2=0.38
r95 14 27 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.302 $Y=0.085
+ $X2=2.302 $Y2=0
r96 14 16 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=2.302 $Y=0.085
+ $X2=2.302 $Y2=0.38
r97 10 24 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.887 $Y=0.085
+ $X2=0.887 $Y2=0
r98 10 12 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.887 $Y=0.085
+ $X2=0.887 $Y2=0.38
r99 3 20 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.235 $X2=3.715 $Y2=0.38
r100 2 16 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.235 $X2=2.3 $Y2=0.38
r101 1 12 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.725
+ $Y=0.235 $X2=0.885 $Y2=0.38
.ends


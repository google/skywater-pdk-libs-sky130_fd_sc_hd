* File: sky130_fd_sc_hd__o2111a_2.pex.spice
* Created: Tue Sep  1 19:19:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2111A_2%A_80_21# 1 2 3 10 12 15 17 19 22 27 28 29
+ 30 31 33 37 39 41 48
c84 31 0 1.37404e-19 $X=1.64 $Y=0.715
r85 51 53 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.16
+ $X2=0.905 $Y2=1.16
r86 39 50 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=3.03 $Y=2.025
+ $X2=3.03 $Y2=1.905
r87 39 41 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.03 $Y=2.025
+ $X2=3.03 $Y2=2.34
r88 38 48 5.86152 $w=2.4e-07 $l=1.4e-07 $layer=LI1_cond $X=2.14 $Y=1.905 $X2=2
+ $Y2=1.905
r89 37 50 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=1.905
+ $X2=3.03 $Y2=1.905
r90 37 38 34.8134 $w=2.38e-07 $l=7.25e-07 $layer=LI1_cond $X=2.865 $Y=1.905
+ $X2=2.14 $Y2=1.905
r91 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.64 $Y=0.715
+ $X2=1.64 $Y2=0.4
r92 29 48 5.86152 $w=2.4e-07 $l=1.4e-07 $layer=LI1_cond $X=1.86 $Y=1.905 $X2=2
+ $Y2=1.905
r93 29 30 26.6502 $w=2.38e-07 $l=5.55e-07 $layer=LI1_cond $X=1.86 $Y=1.905
+ $X2=1.305 $Y2=1.905
r94 28 53 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.115 $Y=1.16
+ $X2=0.905 $Y2=1.16
r95 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.16 $X2=1.115 $Y2=1.16
r96 25 30 6.85752 $w=2.4e-07 $l=1.8869e-07 $layer=LI1_cond $X=1.167 $Y=1.785
+ $X2=1.305 $Y2=1.905
r97 25 27 26.1919 $w=2.73e-07 $l=6.25e-07 $layer=LI1_cond $X=1.167 $Y=1.785
+ $X2=1.167 $Y2=1.16
r98 24 31 30.8588 $w=1.68e-07 $l=4.73e-07 $layer=LI1_cond $X=1.167 $Y=0.8
+ $X2=1.64 $Y2=0.8
r99 24 27 11.5244 $w=2.73e-07 $l=2.75e-07 $layer=LI1_cond $X=1.167 $Y=0.885
+ $X2=1.167 $Y2=1.16
r100 20 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r101 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r102 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r103 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r104 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.16
r105 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.985
r106 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r107 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r108 3 50 600 $w=1.7e-07 $l=4.89898e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.485 $X2=3.03 $Y2=1.885
r109 3 41 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.485 $X2=3.03 $Y2=2.34
r110 2 48 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.485 $X2=2 $Y2=1.885
r111 1 33 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.235 $X2=1.64 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%D1 3 5 7 8 9 17
r33 16 17 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.785 $Y=1.16
+ $X2=1.855 $Y2=1.16
r34 13 16 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=1.67 $Y=1.16
+ $X2=1.785 $Y2=1.16
r35 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.67 $Y=1.16 $X2=1.67
+ $Y2=1.53
r36 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r37 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=1.16
r38 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=0.56
r39 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.16
r40 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.785 $Y=1.325
+ $X2=1.785 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%C1 3 7 9 10 11 12 18
c40 3 0 1.37404e-19 $X=2.215 $Y=0.56
r41 18 21 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.305 $Y=1.16
+ $X2=2.305 $Y2=1.295
r42 18 20 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.305 $Y=1.16
+ $X2=2.305 $Y2=1.025
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=1.16 $X2=2.305 $Y2=1.16
r44 11 12 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.197 $Y=1.19
+ $X2=2.197 $Y2=1.53
r45 11 19 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=2.197 $Y=1.19
+ $X2=2.197 $Y2=1.16
r46 10 19 9.27941 $w=3.83e-07 $l=3.1e-07 $layer=LI1_cond $X=2.197 $Y=0.85
+ $X2=2.197 $Y2=1.16
r47 9 10 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.197 $Y=0.51
+ $X2=2.197 $Y2=0.85
r48 7 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.215 $Y=1.985
+ $X2=2.215 $Y2=1.295
r49 3 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.215 $Y=0.56
+ $X2=2.215 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%B1 3 7 9 10 14 15
c34 7 0 2.30545e-20 $X=2.755 $Y=1.985
c35 3 0 1.45039e-19 $X=2.755 $Y=0.56
r36 14 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.845 $Y=1.16
+ $X2=2.845 $Y2=1.295
r37 14 16 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.845 $Y=1.16
+ $X2=2.845 $Y2=1.025
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.16 $X2=2.845 $Y2=1.16
r39 9 10 9.3293 $w=4.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.89 $Y=1.19 $X2=2.89
+ $Y2=1.53
r40 9 15 0.823174 $w=4.18e-07 $l=3e-08 $layer=LI1_cond $X=2.89 $Y=1.19 $X2=2.89
+ $Y2=1.16
r41 7 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.755 $Y=1.985
+ $X2=2.755 $Y2=1.295
r42 3 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.755 $Y=0.56
+ $X2=2.755 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%A2 3 7 9 10 14 15
c35 15 0 3.18111e-19 $X=3.385 $Y=1.16
c36 7 0 1.38914e-20 $X=3.295 $Y=1.985
c37 3 0 1.38914e-20 $X=3.295 $Y=0.56
r38 14 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.385 $Y=1.16
+ $X2=3.385 $Y2=1.295
r39 14 16 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.385 $Y=1.16
+ $X2=3.385 $Y2=1.025
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.16 $X2=3.385 $Y2=1.16
r41 10 26 35.1694 $w=2.88e-07 $l=8.85e-07 $layer=LI1_cond $X=3.515 $Y=2.21
+ $X2=3.515 $Y2=1.325
r42 9 26 4.79093 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=3.48 $Y=1.19
+ $X2=3.48 $Y2=1.325
r43 9 15 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=3.48 $Y=1.19 $X2=3.48
+ $Y2=1.16
r44 7 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.295 $Y=1.985
+ $X2=3.295 $Y2=1.295
r45 3 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.295 $Y=0.56
+ $X2=3.295 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%A1 3 7 9 10 11 12 13 23 32
c32 10 0 2.77828e-20 $X=4.395 $Y=1.19
r33 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.16 $X2=4.05 $Y2=1.16
r34 20 23 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=3.835 $Y=1.16
+ $X2=4.05 $Y2=1.16
r35 12 13 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=4.412 $Y=1.87
+ $X2=4.412 $Y2=2.21
r36 11 12 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=4.412 $Y=1.53
+ $X2=4.412 $Y2=1.87
r37 11 32 11.6319 $w=2.03e-07 $l=2.15e-07 $layer=LI1_cond $X=4.412 $Y=1.53
+ $X2=4.412 $Y2=1.315
r38 10 32 4.33736 $w=2.05e-07 $l=1.55e-07 $layer=LI1_cond $X=4.412 $Y=1.16
+ $X2=4.412 $Y2=1.315
r39 10 24 7.97574 $w=4.78e-07 $l=2.6e-07 $layer=LI1_cond $X=4.31 $Y=1.16
+ $X2=4.05 $Y2=1.16
r40 9 24 4.27519 $w=3.08e-07 $l=1.15e-07 $layer=LI1_cond $X=3.935 $Y=1.16
+ $X2=4.05 $Y2=1.16
r41 5 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.835 $Y=1.295
+ $X2=3.835 $Y2=1.16
r42 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.835 $Y=1.295
+ $X2=3.835 $Y2=1.985
r43 1 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.835 $Y=1.025
+ $X2=3.835 $Y2=1.16
r44 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.835 $Y=1.025
+ $X2=3.835 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%VPWR 1 2 3 4 13 15 21 25 29 36 41 48 49 57
+ 60 62 65
r68 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 59 60 8.65265 $w=6.08e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.5
+ $X2=1.655 $Y2=2.5
r71 55 59 8.23529 $w=6.08e-07 $l=4.2e-07 $layer=LI1_cond $X=1.15 $Y=2.5 $X2=1.57
+ $Y2=2.5
r72 55 57 9.24088 $w=6.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.15 $Y=2.5
+ $X2=1.035 $Y2=2.5
r73 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 49 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r76 46 65 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.14 $Y=2.72
+ $X2=4.012 $Y2=2.72
r77 46 48 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.14 $Y=2.72
+ $X2=4.37 $Y2=2.72
r78 45 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 45 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 42 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.49 $Y2=2.72
r82 42 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 41 65 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.012 $Y2=2.72
r84 41 44 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=2.99 $Y2=2.72
r85 40 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r86 40 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 39 60 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=1.655 $Y2=2.72
r88 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r89 36 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.49 $Y2=2.72
r90 36 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.07 $Y2=2.72
r91 35 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r92 34 57 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.035 $Y2=2.72
r93 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 32 52 3.66972 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r95 32 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r97 29 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r98 25 28 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=4.012 $Y=1.66
+ $X2=4.012 $Y2=2.34
r99 23 65 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.012 $Y=2.635
+ $X2=4.012 $Y2=2.72
r100 23 28 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=4.012 $Y=2.635
+ $X2=4.012 $Y2=2.34
r101 19 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=2.635
+ $X2=2.49 $Y2=2.72
r102 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.49 $Y=2.635
+ $X2=2.49 $Y2=2.34
r103 15 18 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=1.66
+ $X2=0.24 $Y2=2.34
r104 13 52 3.24547 $w=2.1e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.172 $Y2=2.72
r105 13 18 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.34
r106 4 28 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.485 $X2=4.05 $Y2=2.34
r107 4 25 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.485 $X2=4.05 $Y2=1.66
r108 3 21 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.485 $X2=2.49 $Y2=2.34
r109 2 59 300 $w=1.7e-07 $l=1.1322e-06 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.57 $Y2=2.36
r110 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r111 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%X 1 2 7 8 12
r13 8 21 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.685 $Y=2.21
+ $X2=0.685 $Y2=2.34
r14 8 17 18.6425 $w=3.38e-07 $l=5.5e-07 $layer=LI1_cond $X=0.685 $Y=2.21
+ $X2=0.685 $Y2=1.66
r15 7 17 38.9797 $w=3.38e-07 $l=1.15e-06 $layer=LI1_cond $X=0.685 $Y=0.51
+ $X2=0.685 $Y2=1.66
r16 7 12 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=0.685 $Y=0.51 $X2=0.685
+ $Y2=0.42
r17 2 21 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=2.34
r18 2 17 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.66
r19 1 12 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r57 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r58 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r59 37 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r60 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r61 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.55
+ $Y2=0
r62 34 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=4.37
+ $Y2=0
r63 33 47 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.45
+ $Y2=0
r64 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r65 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r66 30 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.16
+ $Y2=0
r67 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.61
+ $Y2=0
r68 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.55
+ $Y2=0
r69 29 32 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=1.61 $Y2=0
r70 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r71 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 25 40 3.66972 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r73 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r74 24 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.16
+ $Y2=0
r75 24 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r76 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r77 22 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r78 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r79 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.37
r80 14 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0
r81 14 16 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0.38
r82 10 40 3.24547 $w=2.1e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.172 $Y2=0
r83 10 12 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r84 3 20 182 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.235 $X2=3.55 $Y2=0.37
r85 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.38
r86 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O2111A_2%A_566_47# 1 2 7 9 11 15
r23 13 15 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=4.05 $Y=0.625
+ $X2=4.05 $Y2=0.4
r24 12 18 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=0.725
+ $X2=3.03 $Y2=0.725
r25 11 13 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=3.885 $Y=0.725
+ $X2=4.05 $Y2=0.625
r26 11 12 38.2636 $w=1.98e-07 $l=6.9e-07 $layer=LI1_cond $X=3.885 $Y=0.725
+ $X2=3.195 $Y2=0.725
r27 7 18 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=3.03 $Y=0.625 $X2=3.03
+ $Y2=0.725
r28 7 9 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.03 $Y=0.625
+ $X2=3.03 $Y2=0.4
r29 2 15 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=3.91
+ $Y=0.235 $X2=4.05 $Y2=0.4
r30 1 18 182 $w=1.7e-07 $l=5.96678e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.235 $X2=3.03 $Y2=0.74
r31 1 9 182 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.235 $X2=3.03 $Y2=0.4
.ends


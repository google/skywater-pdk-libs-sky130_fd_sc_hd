* File: sky130_fd_sc_hd__ha_1.spice
* Created: Thu Aug 27 14:21:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__ha_1.spice.pex"
.subckt sky130_fd_sc_hd__ha_1  VNB VPB B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_79_21#_M1012_g N_SUM_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_297_47#_M1003_d N_A_250_199#_M1003_g N_A_79_21#_M1003_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_A_297_47#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_297_47#_M1008_d N_A_M1008_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 A_674_47# N_B_M1004_g N_A_250_199#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g A_674_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.0441 PD=0.765421 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1010 N_COUT_M1010_d N_A_250_199#_M1010_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_A_79_21#_M1011_g N_SUM_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.332465 AS=0.26 PD=2.48592 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1005 N_A_79_21#_M1005_d N_A_250_199#_M1005_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.139635 PD=0.69 PS=1.04408 NRD=0 NRS=133.665 M=1 R=2.8
+ SA=75001.1 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1001 A_376_413# N_B_M1001_g N_A_79_21#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.084 AS=0.0567 PD=0.82 PS=0.69 NRD=68.0044 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_376_413# VPB PHIGHVT L=0.15 W=0.42 AD=0.1491
+ AS=0.084 PD=1.13 PS=0.82 NRD=21.0987 NRS=68.0044 M=1 R=2.8 SA=75002.1 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_250_199#_M1009_d N_B_M1009_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0609 AS=0.1491 PD=0.71 PS=1.13 NRD=2.3443 NRS=21.0987 M=1 R=2.8
+ SA=75002.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_250_199#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0832606 AS=0.0609 PD=0.783803 PS=0.71 NRD=23.443 NRS=2.3443 M=1 R=2.8
+ SA=75003.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_COUT_M1013_d N_A_250_199#_M1013_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.198239 PD=2.52 PS=1.8662 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__ha_1.spice.SKY130_FD_SC_HD__HA_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_inputiso0n_1.pex.spice
* Created: Tue Sep  1 19:12:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%A 3 7 9 10 11 19 21
r34 17 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.455 $Y=1.2 $X2=0.365
+ $Y2=1.2
r35 16 19 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.455 $Y=1.16
+ $X2=0.65 $Y2=1.16
r36 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.455
+ $Y=1.16 $X2=0.455 $Y2=1.16
r37 11 17 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=1.2
+ $X2=0.455 $Y2=1.2
r38 10 21 8.91512 $w=2.63e-07 $l=2.05e-07 $layer=LI1_cond $X=0.232 $Y=1.53
+ $X2=0.232 $Y2=1.325
r39 9 21 3.30621 $w=2.65e-07 $l=1.25e-07 $layer=LI1_cond $X=0.232 $Y=1.2
+ $X2=0.232 $Y2=1.325
r40 9 24 3.51781 $w=2.5e-07 $l=1.33e-07 $layer=LI1_cond $X=0.232 $Y=1.2
+ $X2=0.365 $Y2=1.2
r41 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.325
+ $X2=0.65 $Y2=1.16
r42 5 7 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.65 $Y=1.325 $X2=0.65
+ $Y2=2.065
r43 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=0.995
+ $X2=0.65 $Y2=1.16
r44 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.65 $Y=0.995 $X2=0.65
+ $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%SLEEP_B 3 7 9 12
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=1.16 $Y2=1.325
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=1.16 $Y2=0.995
r38 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.16 $X2=1.16 $Y2=1.16
r39 7 15 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.07 $Y=2.065
+ $X2=1.07 $Y2=1.325
r40 3 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.07 $Y=0.585
+ $X2=1.07 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%A_59_75# 1 2 9 12 16 18 19 22 24
+ 25 26 27 31 33
r76 31 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.16 $X2=1.7
+ $Y2=1.325
r77 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.16 $X2=1.7
+ $Y2=0.995
r78 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.16 $X2=1.7 $Y2=1.16
r79 28 30 18.2479 $w=2.34e-07 $l=3.5e-07 $layer=LI1_cond $X=1.65 $Y=0.81
+ $X2=1.65 $Y2=1.16
r80 26 30 9.53671 $w=2.34e-07 $l=1.92678e-07 $layer=LI1_cond $X=1.59 $Y=1.325
+ $X2=1.65 $Y2=1.16
r81 26 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.59 $Y=1.325
+ $X2=1.59 $Y2=1.575
r82 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=1.66
+ $X2=1.59 $Y2=1.575
r83 24 25 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.505 $Y=1.66
+ $X2=1.035 $Y2=1.66
r84 20 25 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.885 $Y=1.745
+ $X2=1.035 $Y2=1.66
r85 20 22 14.7897 $w=2.98e-07 $l=3.85e-07 $layer=LI1_cond $X=0.885 $Y=1.745
+ $X2=0.885 $Y2=2.13
r86 18 28 1.95941 $w=1.9e-07 $l=1.45e-07 $layer=LI1_cond $X=1.505 $Y=0.81
+ $X2=1.65 $Y2=0.81
r87 18 19 51.9522 $w=1.88e-07 $l=8.9e-07 $layer=LI1_cond $X=1.505 $Y=0.81
+ $X2=0.615 $Y2=0.81
r88 14 19 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.45 $Y=0.715
+ $X2=0.615 $Y2=0.81
r89 14 16 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.45 $Y=0.715
+ $X2=0.45 $Y2=0.52
r90 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.61 $Y=1.985
+ $X2=1.61 $Y2=1.325
r91 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.61 $Y=0.56 $X2=1.61
+ $Y2=0.995
r92 2 22 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.725
+ $Y=1.855 $X2=0.86 $Y2=2.13
r93 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.295
+ $Y=0.375 $X2=0.44 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%VPWR 1 2 9 13 16 17 19 20 21 30
+ 31
r31 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r33 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r34 21 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 21 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r36 19 27 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.4 $Y2=2.72
r38 18 30 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=1.4 $Y2=2.72
r40 16 24 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.285 $Y=2.72
+ $X2=0.23 $Y2=2.72
r41 16 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.285 $Y=2.72
+ $X2=0.425 $Y2=2.72
r42 15 27 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=1.15 $Y2=2.72
r43 15 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.425 $Y2=2.72
r44 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=2.635 $X2=1.4
+ $Y2=2.72
r45 11 13 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.4 $Y=2.635
+ $X2=1.4 $Y2=2
r46 7 17 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.425 $Y=2.635
+ $X2=0.425 $Y2=2.72
r47 7 9 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=0.425 $Y=2.635
+ $X2=0.425 $Y2=2.13
r48 2 13 300 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=1.855 $X2=1.4 $Y2=2
r49 1 9 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.295
+ $Y=1.855 $X2=0.44 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%X 1 2 7 11 12 13 14 15 16 25 36
r25 36 40 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=2.09 $Y=1.87 $X2=2.09
+ $Y2=1.915
r26 16 42 5.46036 $w=4.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.985 $Y=2.21
+ $X2=1.985 $Y2=2
r27 15 42 1.69011 $w=4.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.985 $Y=1.935
+ $X2=1.985 $Y2=2
r28 15 40 2.99563 $w=4.58e-07 $l=2e-08 $layer=LI1_cond $X=1.985 $Y=1.935
+ $X2=1.985 $Y2=1.915
r29 15 36 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=2.09 $Y=1.85 $X2=2.09
+ $Y2=1.87
r30 14 15 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.09 $Y=1.53
+ $X2=2.09 $Y2=1.85
r31 13 14 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.09 $Y=1.19
+ $X2=2.09 $Y2=1.53
r32 12 13 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.09 $Y=0.85
+ $X2=2.09 $Y2=1.19
r33 11 25 3.6869 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=2.09 $Y=0.4 $X2=2.09
+ $Y2=0.545
r34 11 12 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.09 $Y=0.57
+ $X2=2.09 $Y2=0.85
r35 11 25 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.09 $Y=0.57
+ $X2=2.09 $Y2=0.545
r36 7 11 3.17836 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=1.965 $Y=0.4 $X2=2.09
+ $Y2=0.4
r37 7 9 5.76222 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.965 $Y=0.4 $X2=1.82
+ $Y2=0.4
r38 2 42 300 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=1.485 $X2=1.92 $Y2=2
r39 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.235 $X2=1.82 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%VGND 1 6 9 10 11 21 22
r27 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r28 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r29 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r30 14 18 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r31 11 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r32 11 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r33 9 18 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.15
+ $Y2=0
r34 9 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.36
+ $Y2=0
r35 8 21 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=2.07
+ $Y2=0
r36 8 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.36
+ $Y2=0
r37 4 10 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0
r38 4 6 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0.38
r39 1 6 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.375 $X2=1.4 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a21boi_2.pex.spice
* Created: Thu Aug 27 14:00:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21BOI_2%B1_N 3 5 7 11 14 15 18
c33 15 0 1.55253e-19 $X=0.23 $Y=0.85
r34 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.34
+ $Y=0.93 $X2=0.34 $Y2=0.93
r35 15 19 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=0.272 $Y=0.85 $X2=0.272
+ $Y2=0.93
r36 13 18 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=0.362 $Y=1.248
+ $X2=0.362 $Y2=0.93
r37 13 14 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.362 $Y=1.248
+ $X2=0.362 $Y2=1.435
r38 9 18 7.41538 $w=3.75e-07 $l=5e-08 $layer=POLY_cond $X=0.362 $Y=0.88
+ $X2=0.362 $Y2=0.93
r39 9 11 163.06 $w=1.5e-07 $l=3.18e-07 $layer=POLY_cond $X=0.362 $Y=0.805
+ $X2=0.68 $Y2=0.805
r40 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.68 $Y=0.73 $X2=0.68
+ $Y2=0.805
r41 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.68 $Y=0.73 $X2=0.68
+ $Y2=0.445
r42 3 14 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=0.475 $Y=2.1
+ $X2=0.475 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_2%A_61_47# 1 2 9 13 17 21 23 25 27 32 35 39
+ 42
c69 23 0 1.55253e-19 $X=1.345 $Y=1.16
c70 13 0 6.77984e-20 $X=1.42 $Y=1.985
r71 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.16 $X2=1.16 $Y2=1.16
r72 37 42 1.58651 $w=2.15e-07 $l=1.3e-07 $layer=LI1_cond $X=0.855 $Y=1.177
+ $X2=0.725 $Y2=1.177
r73 37 39 16.3486 $w=2.13e-07 $l=3.05e-07 $layer=LI1_cond $X=0.855 $Y=1.177
+ $X2=1.16 $Y2=1.177
r74 33 42 4.8823 $w=2.3e-07 $l=1.08e-07 $layer=LI1_cond $X=0.725 $Y=1.285
+ $X2=0.725 $Y2=1.177
r75 33 35 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=0.725 $Y=1.285
+ $X2=0.725 $Y2=2.1
r76 32 42 4.8823 $w=2.3e-07 $l=1.21074e-07 $layer=LI1_cond $X=0.695 $Y=1.07
+ $X2=0.725 $Y2=1.177
r77 31 32 29.9455 $w=1.98e-07 $l=5.4e-07 $layer=LI1_cond $X=0.695 $Y=0.53
+ $X2=0.695 $Y2=1.07
r78 27 31 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.595 $Y=0.445
+ $X2=0.695 $Y2=0.53
r79 27 29 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=0.445
+ $X2=0.43 $Y2=0.445
r80 24 25 86.8776 $w=2.9e-07 $l=4.2e-07 $layer=POLY_cond $X=1.42 $Y=1.16
+ $X2=1.84 $Y2=1.16
r81 23 40 38.2675 $w=2.9e-07 $l=1.85e-07 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.16 $Y2=1.16
r82 23 24 15.5139 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.42 $Y2=1.16
r83 19 25 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.84 $Y=1.305
+ $X2=1.84 $Y2=1.16
r84 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.84 $Y=1.305
+ $X2=1.84 $Y2=1.985
r85 15 25 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.84 $Y=1.015
+ $X2=1.84 $Y2=1.16
r86 15 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.84 $Y=1.015
+ $X2=1.84 $Y2=0.56
r87 11 24 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.42 $Y=1.305
+ $X2=1.42 $Y2=1.16
r88 11 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.42 $Y=1.305
+ $X2=1.42 $Y2=1.985
r89 7 24 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.42 $Y=1.015
+ $X2=1.42 $Y2=1.16
r90 7 9 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.42 $Y=1.015
+ $X2=1.42 $Y2=0.56
r91 2 35 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.89 $X2=0.69 $Y2=2.1
r92 1 29 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.305
+ $Y=0.235 $X2=0.43 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_2%A2 3 7 10 14 17 18 19 21 22 27 28 31 35 39
c82 31 0 1.68189e-19 $X=3.475 $Y=1.53
c83 22 0 2.65731e-19 $X=2.26 $Y=1.16
c84 17 0 2.22276e-19 $X=2.262 $Y=1.495
r85 31 39 2.80098 $w=2.9e-07 $l=9e-08 $layer=LI1_cond $X=3.53 $Y=1.585 $X2=3.53
+ $Y2=1.495
r86 31 39 0.993485 $w=2.88e-07 $l=2.5e-08 $layer=LI1_cond $X=3.53 $Y=1.47
+ $X2=3.53 $Y2=1.495
r87 30 31 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=3.53 $Y=1.295
+ $X2=3.53 $Y2=1.47
r88 28 38 42.7143 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.63 $Y=1.16
+ $X2=3.63 $Y2=1.305
r89 28 37 42.7143 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.63 $Y=1.16
+ $X2=3.63 $Y2=1.015
r90 27 30 4.79698 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=3.59 $Y=1.16
+ $X2=3.59 $Y2=1.295
r91 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.63
+ $Y=1.16 $X2=3.63 $Y2=1.16
r92 22 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.26 $Y2=0.995
r93 21 24 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=1.16
+ $X2=2.26 $Y2=1.245
r94 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r95 18 31 4.5127 $w=1.8e-07 $l=1.45e-07 $layer=LI1_cond $X=3.385 $Y=1.585
+ $X2=3.53 $Y2=1.585
r96 18 19 59.1515 $w=1.78e-07 $l=9.6e-07 $layer=LI1_cond $X=3.385 $Y=1.585
+ $X2=2.425 $Y2=1.585
r97 17 19 7.57412 $w=1.8e-07 $l=2.03074e-07 $layer=LI1_cond $X=2.262 $Y=1.495
+ $X2=2.425 $Y2=1.585
r98 17 24 8.86495 $w=3.23e-07 $l=2.5e-07 $layer=LI1_cond $X=2.262 $Y=1.495
+ $X2=2.262 $Y2=1.245
r99 14 38 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.54 $Y=1.985
+ $X2=3.54 $Y2=1.305
r100 10 37 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.54 $Y=0.56
+ $X2=3.54 $Y2=1.015
r101 7 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.32 $Y=0.56
+ $X2=2.32 $Y2=0.995
r102 1 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.325
+ $X2=2.26 $Y2=1.16
r103 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.26 $Y=1.325
+ $X2=2.26 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_2%A1 1 3 6 8 10 13 15 22
r48 20 22 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.08 $Y=1.16 $X2=3.11
+ $Y2=1.16
r49 17 20 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=2.68 $Y=1.16 $X2=3.08
+ $Y2=1.16
r50 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.08
+ $Y=1.16 $X2=3.08 $Y2=1.16
r51 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r52 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.985
r53 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=1.16
r54 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=0.56
r55 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.325
+ $X2=2.68 $Y2=1.16
r56 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.68 $Y=1.325 $X2=2.68
+ $Y2=1.985
r57 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=0.995
+ $X2=2.68 $Y2=1.16
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.68 $Y=0.995 $X2=2.68
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_2%VPWR 1 2 3 10 12 16 20 23 24 26 27 28 41 42
c64 3 0 1.13712e-19 $X=3.185 $Y=1.485
c65 2 0 1.13651e-19 $X=2.335 $Y=1.485
r66 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r71 33 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r72 32 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r73 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r74 30 45 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r75 30 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 28 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 28 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 26 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.16 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=2.72
+ $X2=3.325 $Y2=2.72
r80 25 41 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.49 $Y=2.72
+ $X2=3.91 $Y2=2.72
r81 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.49 $Y=2.72
+ $X2=3.325 $Y2=2.72
r82 23 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.07 $Y2=2.72
r83 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.47 $Y2=2.72
r84 22 38 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.99 $Y2=2.72
r85 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.47 $Y2=2.72
r86 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.635
+ $X2=3.325 $Y2=2.72
r87 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.325 $Y=2.635
+ $X2=3.325 $Y2=2.36
r88 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=2.635
+ $X2=2.47 $Y2=2.72
r89 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.47 $Y=2.635
+ $X2=2.47 $Y2=2.36
r90 10 45 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r91 10 12 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.165
r92 3 20 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.485 $X2=3.325 $Y2=2.36
r93 2 16 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.47 $Y2=2.36
r94 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.89 $X2=0.26 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_2%A_217_297# 1 2 3 4 15 17 18 19 20 21 25 27
+ 29 31 36
c61 21 0 1.30898e-19 $X=2.81 $Y=1.94
c62 19 0 1.34834e-19 $X=2.05 $Y=2.025
c63 18 0 6.77984e-20 $X=1.35 $Y=2.375
c64 2 0 1.08624e-19 $X=1.915 $Y=1.485
r65 29 38 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=3.79 $Y=2.105
+ $X2=3.79 $Y2=1.98
r66 29 31 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=3.79 $Y=2.105
+ $X2=3.79 $Y2=2.3
r67 28 36 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=1.98 $X2=2.895
+ $Y2=1.98
r68 27 38 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=3.66 $Y=1.98 $X2=3.79
+ $Y2=1.98
r69 27 28 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.66 $Y=1.98
+ $X2=2.98 $Y2=1.98
r70 23 36 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.895 $Y=2.105
+ $X2=2.895 $Y2=1.98
r71 23 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.895 $Y=2.105
+ $X2=2.895 $Y2=2.3
r72 22 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=1.94
+ $X2=2.05 $Y2=1.94
r73 21 36 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.81 $Y=1.94
+ $X2=2.895 $Y2=1.98
r74 21 22 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.81 $Y=1.94
+ $X2=2.215 $Y2=1.94
r75 19 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.025 $X2=2.05
+ $Y2=1.94
r76 19 20 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.05 $Y=2.025
+ $X2=2.05 $Y2=2.285
r77 17 20 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.885 $Y=2.375
+ $X2=2.05 $Y2=2.285
r78 17 18 32.9646 $w=1.78e-07 $l=5.35e-07 $layer=LI1_cond $X=1.885 $Y=2.375
+ $X2=1.35 $Y2=2.375
r79 13 18 7.42255 $w=1.8e-07 $l=1.92819e-07 $layer=LI1_cond $X=1.197 $Y=2.285
+ $X2=1.35 $Y2=2.375
r80 13 15 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=1.197 $Y=2.285
+ $X2=1.197 $Y2=1.96
r81 4 38 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=1.485 $X2=3.755 $Y2=1.96
r82 4 31 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=1.485 $X2=3.755 $Y2=2.3
r83 3 36 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.485 $X2=2.895 $Y2=1.94
r84 3 25 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.485 $X2=2.895 $Y2=2.3
r85 2 34 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.915
+ $Y=1.485 $X2=2.05 $Y2=2.02
r86 1 15 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.485 $X2=1.21 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_2%Y 1 2 3 12 14 18 23 26
r41 23 26 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=1.62 $Y=0.51 $X2=1.62
+ $Y2=0.42
r42 20 23 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=1.62 $Y=0.615
+ $X2=1.62 $Y2=0.51
r43 20 22 4.55203 $w=1.97e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.615
+ $X2=1.62 $Y2=0.7
r44 16 18 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=0.615
+ $X2=2.895 $Y2=0.36
r45 15 22 1.88765 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.72 $Y=0.7 $X2=1.62
+ $Y2=0.7
r46 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.73 $Y=0.7
+ $X2=2.895 $Y2=0.615
r47 14 15 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.73 $Y=0.7
+ $X2=1.72 $Y2=0.7
r48 10 22 4.55203 $w=1.97e-07 $l=8.6487e-08 $layer=LI1_cond $X=1.617 $Y=0.785
+ $X2=1.62 $Y2=0.7
r49 10 12 46.9231 $w=1.93e-07 $l=8.25e-07 $layer=LI1_cond $X=1.617 $Y=0.785
+ $X2=1.617 $Y2=1.61
r50 3 12 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.485 $X2=1.63 $Y2=1.61
r51 2 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.235 $X2=2.895 $Y2=0.36
r52 1 26 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.63 $Y2=0.42
r53 1 22 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.63 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_2%VGND 1 2 3 12 16 18 20 23 24 25 31 35 44 48
+ 50
r55 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r56 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r57 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r58 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r59 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r60 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r61 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r62 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r63 36 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.105
+ $Y2=0
r64 36 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.53
+ $Y2=0
r65 35 47 4.2632 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.887
+ $Y2=0
r66 35 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.45
+ $Y2=0
r67 34 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r68 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r69 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.105
+ $Y2=0
r70 31 33 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.61
+ $Y2=0
r71 29 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r72 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r73 25 29 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r74 25 50 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r75 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.69
+ $Y2=0
r76 23 24 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.105
+ $Y2=0
r77 22 33 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.61
+ $Y2=0
r78 22 24 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.105
+ $Y2=0
r79 18 47 3.21432 $w=2.95e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.782 $Y=0.085
+ $X2=3.887 $Y2=0
r80 18 20 10.7431 $w=2.93e-07 $l=2.75e-07 $layer=LI1_cond $X=3.782 $Y=0.085
+ $X2=3.782 $Y2=0.36
r81 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r82 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.36
r83 10 24 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=0.085
+ $X2=1.105 $Y2=0
r84 10 12 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=1.105 $Y=0.085
+ $X2=1.105 $Y2=0.38
r85 3 20 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.615
+ $Y=0.235 $X2=3.755 $Y2=0.36
r86 2 16 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.235 $X2=2.105 $Y2=0.36
r87 1 12 91 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_NDIFF $count=2 $X=0.755
+ $Y=0.235 $X2=1.105 $Y2=0.38
.ends


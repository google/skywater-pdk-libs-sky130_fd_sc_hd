* File: sky130_fd_sc_hd__o2bb2ai_2.spice.SKY130_FD_SC_HD__O2BB2AI_2.pxi
* Created: Thu Aug 27 14:38:42 2020
* 
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%A1_N N_A1_N_M1010_g N_A1_N_M1002_g
+ N_A1_N_M1011_g N_A1_N_M1013_g N_A1_N_c_98_n N_A1_N_c_99_n N_A1_N_c_91_n A1_N
+ N_A1_N_c_92_n N_A1_N_c_93_n N_A1_N_c_94_n N_A1_N_c_95_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_2%A1_N
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%A2_N N_A2_N_c_168_n N_A2_N_M1004_g
+ N_A2_N_M1014_g N_A2_N_c_169_n N_A2_N_M1005_g N_A2_N_M1017_g A2_N
+ N_A2_N_c_171_n PM_SKY130_FD_SC_HD__O2BB2AI_2%A2_N
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%A_113_297# N_A_113_297#_M1004_s
+ N_A_113_297#_M1002_d N_A_113_297#_M1017_d N_A_113_297#_c_213_n
+ N_A_113_297#_M1012_g N_A_113_297#_M1016_g N_A_113_297#_c_214_n
+ N_A_113_297#_M1015_g N_A_113_297#_M1019_g N_A_113_297#_c_227_n
+ N_A_113_297#_c_215_n N_A_113_297#_c_232_n N_A_113_297#_c_216_n
+ N_A_113_297#_c_222_n N_A_113_297#_c_241_n N_A_113_297#_c_217_n
+ N_A_113_297#_c_243_n N_A_113_297#_c_218_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_2%A_113_297#
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%B1 N_B1_c_317_n N_B1_M1006_g N_B1_M1000_g
+ N_B1_M1007_g N_B1_M1018_g N_B1_c_318_n N_B1_c_319_n N_B1_c_327_n B1
+ N_B1_c_321_n N_B1_c_322_n N_B1_c_330_n PM_SKY130_FD_SC_HD__O2BB2AI_2%B1
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%B2 N_B2_c_400_n N_B2_M1001_g N_B2_M1003_g
+ N_B2_c_401_n N_B2_M1009_g N_B2_M1008_g B2 N_B2_c_403_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_2%B2
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%VPWR N_VPWR_M1002_s N_VPWR_M1014_s
+ N_VPWR_M1013_s N_VPWR_M1019_d N_VPWR_M1018_d N_VPWR_c_449_n N_VPWR_c_450_n
+ N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n
+ VPWR N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n N_VPWR_c_448_n
+ N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n N_VPWR_c_463_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%Y N_Y_M1012_d N_Y_M1016_s N_Y_M1003_s
+ N_Y_c_533_n N_Y_c_537_n N_Y_c_550_n N_Y_c_531_n N_Y_c_540_n N_Y_c_556_n Y
+ PM_SKY130_FD_SC_HD__O2BB2AI_2%Y
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%A_730_297# N_A_730_297#_M1000_s
+ N_A_730_297#_M1008_d N_A_730_297#_c_582_n N_A_730_297#_c_581_n
+ N_A_730_297#_c_588_n PM_SKY130_FD_SC_HD__O2BB2AI_2%A_730_297#
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%VGND N_VGND_M1010_d N_VGND_M1011_d
+ N_VGND_M1006_d N_VGND_M1009_s N_VGND_c_595_n N_VGND_c_596_n N_VGND_c_597_n
+ N_VGND_c_598_n N_VGND_c_599_n N_VGND_c_600_n N_VGND_c_601_n N_VGND_c_602_n
+ N_VGND_c_603_n N_VGND_c_604_n N_VGND_c_605_n VGND N_VGND_c_606_n
+ N_VGND_c_607_n PM_SKY130_FD_SC_HD__O2BB2AI_2%VGND
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%A_113_47# N_A_113_47#_M1010_s
+ N_A_113_47#_M1005_d N_A_113_47#_c_677_n N_A_113_47#_c_676_n
+ N_A_113_47#_c_682_n PM_SKY130_FD_SC_HD__O2BB2AI_2%A_113_47#
x_PM_SKY130_FD_SC_HD__O2BB2AI_2%A_471_47# N_A_471_47#_M1012_s
+ N_A_471_47#_M1015_s N_A_471_47#_M1001_d N_A_471_47#_M1007_s
+ N_A_471_47#_c_704_n N_A_471_47#_c_709_n N_A_471_47#_c_710_n
+ N_A_471_47#_c_698_n N_A_471_47#_c_699_n N_A_471_47#_c_718_n
+ N_A_471_47#_c_700_n N_A_471_47#_c_701_n N_A_471_47#_c_702_n
+ N_A_471_47#_c_703_n PM_SKY130_FD_SC_HD__O2BB2AI_2%A_471_47#
cc_1 VNB N_A1_N_c_91_n 0.027272f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_2 VNB N_A1_N_c_92_n 0.0322882f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_3 VNB N_A1_N_c_93_n 0.0143983f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_4 VNB N_A1_N_c_94_n 0.0218917f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=0.995
cc_5 VNB N_A1_N_c_95_n 0.0196176f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=0.995
cc_6 VNB N_A2_N_c_168_n 0.0161504f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_7 VNB N_A2_N_c_169_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_8 VNB A2_N 0.00221934f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.53
cc_9 VNB N_A2_N_c_171_n 0.0299959f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_10 VNB N_A_113_297#_c_213_n 0.0191083f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_11 VNB N_A_113_297#_c_214_n 0.0160918f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.445
cc_12 VNB N_A_113_297#_c_215_n 0.0106771f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.325
cc_13 VNB N_A_113_297#_c_216_n 0.014236f $X=-0.19 $Y=-0.24 $X2=0.357 $Y2=1.16
cc_14 VNB N_A_113_297#_c_217_n 0.00219468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_113_297#_c_218_n 0.0493388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_c_317_n 0.0165399f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_17 VNB N_B1_c_318_n 0.00366635f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.445
cc_18 VNB N_B1_c_319_n 0.0195026f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_19 VNB B1 0.0239041f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_B1_c_321_n 0.0267828f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_21 VNB N_B1_c_322_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.325
cc_22 VNB N_B2_c_400_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_23 VNB N_B2_c_401_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_24 VNB B2 0.0015795f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.53
cc_25 VNB N_B2_c_403_n 0.0308136f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_26 VNB N_VPWR_c_448_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_531_n 0.00181832f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_28 VNB N_VGND_c_595_n 0.0116911f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.985
cc_29 VNB N_VGND_c_596_n 0.00651208f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.53
cc_30 VNB N_VGND_c_597_n 0.00469239f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_31 VNB N_VGND_c_598_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_599_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=0.995
cc_33 VNB N_VGND_c_600_n 0.0373934f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=0.995
cc_34 VNB N_VGND_c_601_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.325
cc_35 VNB N_VGND_c_602_n 0.0393939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_603_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0.357 $Y2=1.19
cc_37 VNB N_VGND_c_604_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0.357 $Y2=1.53
cc_38 VNB N_VGND_c_605_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_606_n 0.0240673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_607_n 0.29083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_113_47#_c_676_n 0.00290328f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_42 VNB N_A_471_47#_c_698_n 0.00332606f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_43 VNB N_A_471_47#_c_699_n 0.00748893f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_44 VNB N_A_471_47#_c_700_n 0.0138471f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_45 VNB N_A_471_47#_c_701_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_46 VNB N_A_471_47#_c_702_n 0.00341654f $X=-0.19 $Y=-0.24 $X2=0.357 $Y2=1.19
cc_47 VNB N_A_471_47#_c_703_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VPB N_A1_N_M1002_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_49 VPB N_A1_N_M1013_g 0.0223541f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_50 VPB N_A1_N_c_98_n 0.00888011f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.53
cc_51 VPB N_A1_N_c_99_n 0.00220702f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_52 VPB N_A1_N_c_91_n 0.00655093f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_53 VPB N_A1_N_c_92_n 0.00672428f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_54 VPB N_A1_N_c_93_n 0.0158086f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_55 VPB N_A2_N_M1014_g 0.0183602f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_56 VPB N_A2_N_M1017_g 0.0183587f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_57 VPB N_A2_N_c_171_n 0.00400475f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_58 VPB N_A_113_297#_M1016_g 0.0218037f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.53
cc_59 VPB N_A_113_297#_M1019_g 0.0176027f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_60 VPB N_A_113_297#_c_216_n 0.0109534f $X=-0.19 $Y=1.305 $X2=0.357 $Y2=1.16
cc_61 VPB N_A_113_297#_c_222_n 0.00263893f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_113_297#_c_218_n 0.014681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_B1_M1000_g 0.0176435f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_64 VPB N_B1_M1018_g 0.0223957f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_65 VPB N_B1_c_318_n 0.00235779f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.445
cc_66 VPB N_B1_c_319_n 0.00444401f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_67 VPB N_B1_c_327_n 2.61886e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB B1 0.0264276f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_69 VPB N_B1_c_321_n 0.00483422f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_70 VPB N_B1_c_330_n 0.00841978f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.325
cc_71 VPB N_B2_M1003_g 0.0183389f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_72 VPB N_B2_M1008_g 0.0183442f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_73 VPB N_B2_c_403_n 0.00405367f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_74 VPB N_VPWR_c_449_n 0.0117686f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.53
cc_75 VPB N_VPWR_c_450_n 0.00456855f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_76 VPB N_VPWR_c_451_n 0.00393511f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_77 VPB N_VPWR_c_452_n 0.00478931f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_78 VPB N_VPWR_c_453_n 0.00492724f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=0.995
cc_79 VPB N_VPWR_c_454_n 0.0363617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_455_n 0.00391723f $X=-0.19 $Y=1.305 $X2=0.357 $Y2=1.19
cc_81 VPB N_VPWR_c_456_n 0.0159336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_457_n 0.017149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_458_n 0.013281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_448_n 0.0545127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_460_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_461_n 0.0163086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_462_n 0.0208855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_463_n 0.00545601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB Y 0.00116797f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_90 N_A1_N_c_94_n N_A2_N_c_168_n 0.012379f $X=0.46 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A1_N_M1002_g N_A2_N_M1014_g 0.0277995f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A1_N_c_98_n N_A2_N_M1014_g 0.00985724f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_93 N_A1_N_c_93_n N_A2_N_M1014_g 0.00311269f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A1_N_c_95_n N_A2_N_c_169_n 0.0269138f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A1_N_M1013_g N_A2_N_M1017_g 0.0420013f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A1_N_c_98_n N_A2_N_M1017_g 0.01034f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_97 N_A1_N_c_99_n N_A2_N_M1017_g 0.00265828f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A1_N_c_98_n A2_N 0.0428438f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_99 N_A1_N_c_99_n A2_N 0.0129639f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A1_N_c_91_n A2_N 6.836e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A1_N_c_92_n A2_N 0.00119077f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A1_N_c_93_n A2_N 0.0171095f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A1_N_c_98_n N_A2_N_c_171_n 0.00214031f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_104 N_A1_N_c_99_n N_A2_N_c_171_n 0.00115736f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A1_N_c_91_n N_A2_N_c_171_n 0.0224479f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A1_N_c_92_n N_A2_N_c_171_n 0.0222728f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A1_N_c_93_n N_A2_N_c_171_n 6.05453e-19 $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A1_N_c_98_n N_A_113_297#_M1002_d 0.00193053f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_109 N_A1_N_c_93_n N_A_113_297#_M1002_d 3.15855e-19 $X=0.46 $Y=1.16 $X2=0
+ $Y2=0
cc_110 N_A1_N_c_98_n N_A_113_297#_M1017_d 0.00161579f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_111 N_A1_N_c_98_n N_A_113_297#_c_227_n 0.0317352f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_112 N_A1_N_c_98_n N_A_113_297#_c_215_n 0.00724488f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_113 N_A1_N_c_99_n N_A_113_297#_c_215_n 0.0252775f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A1_N_c_91_n N_A_113_297#_c_215_n 0.00447326f $X=1.78 $Y=1.16 $X2=0
+ $Y2=0
cc_115 N_A1_N_c_95_n N_A_113_297#_c_215_n 0.0140641f $X=1.78 $Y=0.995 $X2=0
+ $Y2=0
cc_116 N_A1_N_M1013_g N_A_113_297#_c_232_n 0.0123658f $X=1.75 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A1_N_c_98_n N_A_113_297#_c_232_n 0.0162711f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_118 N_A1_N_c_91_n N_A_113_297#_c_232_n 3.71138e-19 $X=1.78 $Y=1.16 $X2=0
+ $Y2=0
cc_119 N_A1_N_c_99_n N_A_113_297#_c_216_n 0.0204179f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A1_N_c_91_n N_A_113_297#_c_216_n 0.00416282f $X=1.78 $Y=1.16 $X2=0
+ $Y2=0
cc_121 N_A1_N_c_95_n N_A_113_297#_c_216_n 0.00270192f $X=1.78 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_A1_N_M1013_g N_A_113_297#_c_222_n 0.00664027f $X=1.75 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A1_N_c_98_n N_A_113_297#_c_222_n 0.0139547f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_124 N_A1_N_c_99_n N_A_113_297#_c_222_n 0.00943421f $X=1.78 $Y=1.16 $X2=0
+ $Y2=0
cc_125 N_A1_N_c_98_n N_A_113_297#_c_241_n 0.0124479f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_126 N_A1_N_c_95_n N_A_113_297#_c_217_n 3.91234e-19 $X=1.78 $Y=0.995 $X2=0
+ $Y2=0
cc_127 N_A1_N_c_98_n N_A_113_297#_c_243_n 0.0119948f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_128 N_A1_N_c_99_n N_A_113_297#_c_218_n 2.28984e-19 $X=1.78 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A1_N_c_91_n N_A_113_297#_c_218_n 0.00929877f $X=1.78 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A1_N_c_93_n N_VPWR_M1002_s 0.00364133f $X=0.46 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A1_N_c_98_n N_VPWR_M1014_s 0.00166235f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_132 N_A1_N_c_98_n N_VPWR_M1013_s 0.00202599f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_133 N_A1_N_M1002_g N_VPWR_c_450_n 0.00335371f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A1_N_c_92_n N_VPWR_c_450_n 3.6579e-19 $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A1_N_c_93_n N_VPWR_c_450_n 0.0175772f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A1_N_M1002_g N_VPWR_c_456_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A1_N_M1002_g N_VPWR_c_448_n 0.0114494f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A1_N_M1013_g N_VPWR_c_448_n 0.00725698f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_N_M1013_g N_VPWR_c_461_n 0.00441875f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A1_N_M1013_g N_VPWR_c_462_n 0.00353572f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A1_N_c_92_n N_VGND_c_596_n 0.00176179f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A1_N_c_93_n N_VGND_c_596_n 0.0145468f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A1_N_c_94_n N_VGND_c_596_n 0.00460417f $X=0.46 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_N_c_95_n N_VGND_c_597_n 0.00438629f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A1_N_c_94_n N_VGND_c_600_n 0.00541892f $X=0.46 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A1_N_c_95_n N_VGND_c_600_n 0.00423906f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A1_N_c_94_n N_VGND_c_607_n 0.0104687f $X=0.46 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A1_N_c_95_n N_VGND_c_607_n 0.0070828f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A1_N_c_94_n N_A_113_47#_c_677_n 0.00217882f $X=0.46 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A1_N_c_98_n N_A_113_47#_c_676_n 0.00586387f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_151 N_A1_N_c_92_n N_A_113_47#_c_676_n 0.0015436f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A1_N_c_93_n N_A_113_47#_c_676_n 0.00717578f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A1_N_c_94_n N_A_113_47#_c_676_n 0.00511542f $X=0.46 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_A1_N_c_95_n N_A_113_47#_c_682_n 0.00265651f $X=1.78 $Y=0.995 $X2=0
+ $Y2=0
cc_155 N_A2_N_M1014_g N_A_113_297#_c_227_n 0.0104429f $X=0.91 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A2_N_M1017_g N_A_113_297#_c_227_n 0.0103881f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A2_N_c_169_n N_A_113_297#_c_215_n 0.00768885f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_158 N_A2_N_c_168_n N_A_113_297#_c_217_n 0.00381649f $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A2_N_c_169_n N_A_113_297#_c_217_n 0.00298551f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_160 A2_N N_A_113_297#_c_217_n 0.0323718f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A2_N_c_171_n N_A_113_297#_c_217_n 0.00224214f $X=1.33 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A2_N_M1014_g N_VPWR_c_451_n 0.00158508f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_N_M1017_g N_VPWR_c_451_n 0.00157702f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A2_N_M1014_g N_VPWR_c_456_n 0.00441875f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A2_N_M1014_g N_VPWR_c_448_n 0.00588739f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A2_N_M1017_g N_VPWR_c_448_n 0.00593338f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A2_N_M1017_g N_VPWR_c_461_n 0.00441875f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A2_N_c_168_n N_VGND_c_600_n 0.00368123f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A2_N_c_169_n N_VGND_c_600_n 0.00368123f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A2_N_c_168_n N_VGND_c_607_n 0.00527354f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A2_N_c_169_n N_VGND_c_607_n 0.00527354f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_N_c_168_n N_A_113_47#_c_682_n 0.00957565f $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A2_N_c_169_n N_A_113_47#_c_682_n 0.00826183f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_174 A2_N N_A_113_47#_c_682_n 0.00353291f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_175 N_A_113_297#_c_214_n N_B1_c_317_n 0.0103783f $X=3.12 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_113_297#_M1019_g N_B1_M1000_g 0.0370974f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_113_297#_c_218_n N_B1_c_318_n 0.00126243f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_113_297#_c_218_n N_B1_c_319_n 0.0184166f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_113_297#_M1019_g N_B1_c_327_n 6.89304e-19 $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_113_297#_c_227_n N_VPWR_M1014_s 0.00317395f $X=1.415 $Y=1.875 $X2=0
+ $Y2=0
cc_181 N_A_113_297#_c_232_n N_VPWR_M1013_s 0.016629f $X=2.115 $Y=1.875 $X2=0
+ $Y2=0
cc_182 N_A_113_297#_c_222_n N_VPWR_M1013_s 0.0100007f $X=2.2 $Y=1.785 $X2=0
+ $Y2=0
cc_183 N_A_113_297#_c_227_n N_VPWR_c_451_n 0.0123469f $X=1.415 $Y=1.875 $X2=0
+ $Y2=0
cc_184 N_A_113_297#_M1019_g N_VPWR_c_452_n 0.00170597f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_113_297#_c_227_n N_VPWR_c_456_n 0.0020229f $X=1.415 $Y=1.875 $X2=0
+ $Y2=0
cc_186 N_A_113_297#_c_241_n N_VPWR_c_456_n 0.0141298f $X=0.7 $Y=1.96 $X2=0 $Y2=0
cc_187 N_A_113_297#_M1016_g N_VPWR_c_457_n 0.00541359f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_113_297#_M1019_g N_VPWR_c_457_n 0.00585385f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_113_297#_M1002_d N_VPWR_c_448_n 0.00253991f $X=0.565 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A_113_297#_M1017_d N_VPWR_c_448_n 0.00302071f $X=1.405 $Y=1.485 $X2=0
+ $Y2=0
cc_191 N_A_113_297#_M1016_g N_VPWR_c_448_n 0.0108251f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_113_297#_M1019_g N_VPWR_c_448_n 0.00599344f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_113_297#_c_227_n N_VPWR_c_448_n 0.00806641f $X=1.415 $Y=1.875 $X2=0
+ $Y2=0
cc_194 N_A_113_297#_c_232_n N_VPWR_c_448_n 0.00530436f $X=2.115 $Y=1.875 $X2=0
+ $Y2=0
cc_195 N_A_113_297#_c_241_n N_VPWR_c_448_n 0.00953524f $X=0.7 $Y=1.96 $X2=0
+ $Y2=0
cc_196 N_A_113_297#_c_243_n N_VPWR_c_448_n 0.00745459f $X=1.54 $Y=1.875 $X2=0
+ $Y2=0
cc_197 N_A_113_297#_c_227_n N_VPWR_c_461_n 0.0020229f $X=1.415 $Y=1.875 $X2=0
+ $Y2=0
cc_198 N_A_113_297#_c_232_n N_VPWR_c_461_n 0.0020229f $X=2.115 $Y=1.875 $X2=0
+ $Y2=0
cc_199 N_A_113_297#_c_243_n N_VPWR_c_461_n 0.00414246f $X=1.54 $Y=1.875 $X2=0
+ $Y2=0
cc_200 N_A_113_297#_M1016_g N_VPWR_c_462_n 0.00331225f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_113_297#_c_232_n N_VPWR_c_462_n 0.0329633f $X=2.115 $Y=1.875 $X2=0
+ $Y2=0
cc_202 N_A_113_297#_c_213_n N_Y_c_533_n 0.0100687f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_113_297#_c_214_n N_Y_c_533_n 0.00607626f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_113_297#_c_216_n N_Y_c_533_n 0.0364002f $X=2.2 $Y=1.325 $X2=0 $Y2=0
cc_205 N_A_113_297#_c_218_n N_Y_c_533_n 0.00665189f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_113_297#_M1016_g N_Y_c_537_n 0.011388f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_113_297#_c_232_n N_Y_c_537_n 3.59749e-19 $X=2.115 $Y=1.875 $X2=0
+ $Y2=0
cc_208 N_A_113_297#_c_218_n N_Y_c_531_n 0.0174032f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_113_297#_M1016_g N_Y_c_540_n 0.00310918f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_113_297#_M1019_g N_Y_c_540_n 0.00831614f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_113_297#_c_232_n N_Y_c_540_n 0.00679272f $X=2.115 $Y=1.875 $X2=0
+ $Y2=0
cc_212 N_A_113_297#_M1016_g Y 0.0101677f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_113_297#_M1019_g Y 0.0101353f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_113_297#_c_222_n Y 0.0162945f $X=2.2 $Y=1.785 $X2=0 $Y2=0
cc_215 N_A_113_297#_c_218_n Y 0.00304388f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_113_297#_c_215_n N_VGND_M1011_d 0.00315681f $X=2.115 $Y=0.815 $X2=0
+ $Y2=0
cc_217 N_A_113_297#_c_213_n N_VGND_c_597_n 0.00192498f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_113_297#_c_215_n N_VGND_c_597_n 0.0127273f $X=2.115 $Y=0.815 $X2=0
+ $Y2=0
cc_219 N_A_113_297#_c_215_n N_VGND_c_600_n 0.00199263f $X=2.115 $Y=0.815 $X2=0
+ $Y2=0
cc_220 N_A_113_297#_c_213_n N_VGND_c_602_n 0.00357877f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_113_297#_c_214_n N_VGND_c_602_n 0.00357877f $X=3.12 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_113_297#_c_215_n N_VGND_c_602_n 0.00102539f $X=2.115 $Y=0.815 $X2=0
+ $Y2=0
cc_223 N_A_113_297#_c_216_n N_VGND_c_602_n 0.00289403f $X=2.2 $Y=1.325 $X2=0
+ $Y2=0
cc_224 N_A_113_297#_M1004_s N_VGND_c_607_n 0.00220248f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_225 N_A_113_297#_c_213_n N_VGND_c_607_n 0.00655123f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_113_297#_c_214_n N_VGND_c_607_n 0.00533624f $X=3.12 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_113_297#_c_215_n N_VGND_c_607_n 0.00733587f $X=2.115 $Y=0.815 $X2=0
+ $Y2=0
cc_228 N_A_113_297#_c_216_n N_VGND_c_607_n 0.00478629f $X=2.2 $Y=1.325 $X2=0
+ $Y2=0
cc_229 N_A_113_297#_c_215_n N_A_113_47#_M1005_d 0.00191752f $X=2.115 $Y=0.815
+ $X2=0 $Y2=0
cc_230 N_A_113_297#_c_217_n N_A_113_47#_c_676_n 0.0105027f $X=1.285 $Y=0.775
+ $X2=0 $Y2=0
cc_231 N_A_113_297#_M1004_s N_A_113_47#_c_682_n 0.00318958f $X=0.985 $Y=0.235
+ $X2=0 $Y2=0
cc_232 N_A_113_297#_c_215_n N_A_113_47#_c_682_n 0.014624f $X=2.115 $Y=0.815
+ $X2=0 $Y2=0
cc_233 N_A_113_297#_c_217_n N_A_113_47#_c_682_n 0.015032f $X=1.285 $Y=0.775
+ $X2=0 $Y2=0
cc_234 N_A_113_297#_c_213_n N_A_471_47#_c_704_n 0.0127333f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_113_297#_c_214_n N_A_471_47#_c_704_n 0.010549f $X=3.12 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_113_297#_c_218_n N_A_471_47#_c_704_n 3.07604e-19 $X=3.12 $Y=1.16
+ $X2=0 $Y2=0
cc_237 N_A_113_297#_c_216_n N_A_471_47#_c_702_n 0.00917889f $X=2.2 $Y=1.325
+ $X2=0 $Y2=0
cc_238 N_A_113_297#_c_218_n N_A_471_47#_c_702_n 0.00150181f $X=3.12 $Y=1.16
+ $X2=0 $Y2=0
cc_239 N_B1_c_317_n N_B2_c_400_n 0.0258191f $X=3.575 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_240 N_B1_M1000_g N_B2_M1003_g 0.0440009f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_241 N_B1_c_330_n N_B2_M1003_g 0.0108086f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_242 N_B1_c_322_n N_B2_c_401_n 0.0234969f $X=4.895 $Y=0.995 $X2=0 $Y2=0
cc_243 N_B1_M1018_g N_B2_M1008_g 0.0234969f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_244 N_B1_c_330_n N_B2_M1008_g 0.0149047f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_245 N_B1_c_318_n B2 0.0134455f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_246 N_B1_c_319_n B2 2.20976e-19 $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_247 B1 B2 0.0147638f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_248 N_B1_c_321_n B2 7.56849e-19 $X=4.895 $Y=1.16 $X2=0 $Y2=0
cc_249 N_B1_c_330_n B2 0.0381541f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_250 N_B1_c_318_n N_B2_c_403_n 0.00527477f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_251 N_B1_c_319_n N_B2_c_403_n 0.022397f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_252 B1 N_B2_c_403_n 0.00517996f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_253 N_B1_c_321_n N_B2_c_403_n 0.0234969f $X=4.895 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_c_330_n N_B2_c_403_n 0.00214031f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_255 N_B1_c_327_n N_VPWR_M1019_d 0.00156637f $X=3.74 $Y=1.53 $X2=0 $Y2=0
cc_256 B1 N_VPWR_M1018_d 0.00405314f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_257 N_B1_M1000_g N_VPWR_c_452_n 0.0031196f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B1_M1018_g N_VPWR_c_453_n 0.00439972f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_259 B1 N_VPWR_c_453_n 0.0170768f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_260 N_B1_c_321_n N_VPWR_c_453_n 2.70076e-19 $X=4.895 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B1_M1000_g N_VPWR_c_454_n 0.00585385f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_262 N_B1_M1018_g N_VPWR_c_454_n 0.00585385f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_263 N_B1_M1000_g N_VPWR_c_448_n 0.00602311f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_264 N_B1_M1018_g N_VPWR_c_448_n 0.0116831f $X=4.835 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B1_c_330_n N_Y_M1003_s 0.00165831f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_266 N_B1_c_317_n N_Y_c_533_n 5.12048e-19 $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B1_c_319_n N_Y_c_533_n 4.20265e-19 $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B1_M1000_g N_Y_c_550_n 0.0117106f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B1_c_319_n N_Y_c_550_n 3.01349e-19 $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B1_c_327_n N_Y_c_550_n 0.0164816f $X=3.74 $Y=1.53 $X2=0 $Y2=0
cc_271 N_B1_c_330_n N_Y_c_550_n 0.0190307f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_272 N_B1_c_318_n N_Y_c_531_n 0.0286572f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B1_c_319_n N_Y_c_531_n 8.75389e-19 $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B1_c_330_n N_Y_c_556_n 0.0120079f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_275 N_B1_M1000_g Y 6.03153e-19 $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B1_c_327_n Y 0.00852039f $X=3.74 $Y=1.53 $X2=0 $Y2=0
cc_277 N_B1_c_327_n N_A_730_297#_M1000_s 3.52503e-19 $X=3.74 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_278 N_B1_c_330_n N_A_730_297#_M1000_s 0.00130005f $X=4.73 $Y=1.345 $X2=-0.19
+ $Y2=-0.24
cc_279 N_B1_c_330_n N_A_730_297#_M1008_d 0.00165831f $X=4.73 $Y=1.345 $X2=0
+ $Y2=0
cc_280 N_B1_c_330_n N_A_730_297#_c_581_n 0.0126919f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_281 N_B1_c_317_n N_VGND_c_598_n 0.00268723f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B1_c_322_n N_VGND_c_599_n 0.00268723f $X=4.895 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B1_c_317_n N_VGND_c_602_n 0.00422898f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B1_c_322_n N_VGND_c_606_n 0.00423334f $X=4.895 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B1_c_317_n N_VGND_c_607_n 0.00588342f $X=3.575 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B1_c_322_n N_VGND_c_607_n 0.00684971f $X=4.895 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B1_c_317_n N_A_471_47#_c_709_n 0.00255288f $X=3.575 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_B1_c_317_n N_A_471_47#_c_710_n 0.00393886f $X=3.575 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_B1_c_317_n N_A_471_47#_c_698_n 0.00845282f $X=3.575 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_B1_c_318_n N_A_471_47#_c_698_n 0.0160434f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_291 N_B1_c_319_n N_A_471_47#_c_698_n 0.001478f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B1_c_330_n N_A_471_47#_c_698_n 0.0071189f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_293 N_B1_c_317_n N_A_471_47#_c_699_n 0.00109291f $X=3.575 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_B1_c_318_n N_A_471_47#_c_699_n 0.010391f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_295 N_B1_c_319_n N_A_471_47#_c_699_n 0.00153445f $X=3.575 $Y=1.16 $X2=0 $Y2=0
cc_296 N_B1_c_317_n N_A_471_47#_c_718_n 5.22228e-19 $X=3.575 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_B1_c_322_n N_A_471_47#_c_718_n 5.22228e-19 $X=4.895 $Y=0.995 $X2=0
+ $Y2=0
cc_298 B1 N_A_471_47#_c_700_n 0.0407659f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_299 N_B1_c_321_n N_A_471_47#_c_700_n 0.00307118f $X=4.895 $Y=1.16 $X2=0 $Y2=0
cc_300 N_B1_c_322_n N_A_471_47#_c_700_n 0.00995225f $X=4.895 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_B1_c_330_n N_A_471_47#_c_700_n 0.00779194f $X=4.73 $Y=1.345 $X2=0 $Y2=0
cc_302 N_B1_c_322_n N_A_471_47#_c_701_n 0.00630972f $X=4.895 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_B2_M1003_g N_VPWR_c_454_n 0.00357877f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_304 N_B2_M1008_g N_VPWR_c_454_n 0.00357877f $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_305 N_B2_M1003_g N_VPWR_c_448_n 0.00525237f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_306 N_B2_M1008_g N_VPWR_c_448_n 0.00525237f $X=4.415 $Y=1.985 $X2=0 $Y2=0
cc_307 N_B2_M1003_g N_Y_c_550_n 0.00924026f $X=3.995 $Y=1.985 $X2=0 $Y2=0
cc_308 N_B2_M1003_g N_A_730_297#_c_582_n 0.00851673f $X=3.995 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_B2_M1008_g N_A_730_297#_c_582_n 0.0121306f $X=4.415 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_B2_c_400_n N_VGND_c_598_n 0.00146448f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_311 N_B2_c_401_n N_VGND_c_599_n 0.00146448f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_312 N_B2_c_400_n N_VGND_c_604_n 0.00424416f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B2_c_401_n N_VGND_c_604_n 0.00423334f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B2_c_400_n N_VGND_c_607_n 0.00576327f $X=3.995 $Y=0.995 $X2=0 $Y2=0
cc_315 N_B2_c_401_n N_VGND_c_607_n 0.0057435f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B2_c_400_n N_A_471_47#_c_710_n 4.87042e-19 $X=3.995 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_B2_c_400_n N_A_471_47#_c_698_n 0.00894278f $X=3.995 $Y=0.995 $X2=0
+ $Y2=0
cc_318 B2 N_A_471_47#_c_698_n 0.00545718f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_319 N_B2_c_400_n N_A_471_47#_c_718_n 0.00630972f $X=3.995 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_B2_c_401_n N_A_471_47#_c_718_n 0.00630972f $X=4.415 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_B2_c_401_n N_A_471_47#_c_700_n 0.00865686f $X=4.415 $Y=0.995 $X2=0
+ $Y2=0
cc_322 B2 N_A_471_47#_c_700_n 0.00900407f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_323 N_B2_c_401_n N_A_471_47#_c_701_n 5.22228e-19 $X=4.415 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_B2_c_400_n N_A_471_47#_c_703_n 0.00128009f $X=3.995 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_B2_c_401_n N_A_471_47#_c_703_n 0.00113286f $X=4.415 $Y=0.995 $X2=0
+ $Y2=0
cc_326 B2 N_A_471_47#_c_703_n 0.0265405f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_327 N_B2_c_403_n N_A_471_47#_c_703_n 0.00230339f $X=4.415 $Y=1.16 $X2=0 $Y2=0
cc_328 N_VPWR_c_448_n N_Y_M1016_s 0.00219397f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_329 N_VPWR_c_448_n N_Y_M1003_s 0.0021603f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_330 N_VPWR_c_457_n N_Y_c_537_n 0.0165691f $X=3.205 $Y=2.72 $X2=0 $Y2=0
cc_331 N_VPWR_c_448_n N_Y_c_537_n 0.0108863f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_332 N_VPWR_M1019_d N_Y_c_550_n 0.0083378f $X=3.195 $Y=1.485 $X2=0 $Y2=0
cc_333 N_VPWR_c_452_n N_Y_c_550_n 0.0150965f $X=3.33 $Y=2.3 $X2=0 $Y2=0
cc_334 N_VPWR_c_448_n N_Y_c_550_n 0.00691349f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_335 N_VPWR_c_448_n N_Y_c_540_n 0.00587149f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_336 N_VPWR_c_448_n N_A_730_297#_M1000_s 0.00219968f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_337 N_VPWR_c_448_n N_A_730_297#_M1008_d 0.00246446f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_454_n N_A_730_297#_c_582_n 0.0473226f $X=4.965 $Y=2.72 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_448_n N_A_730_297#_c_582_n 0.0300947f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_454_n N_A_730_297#_c_588_n 0.0137033f $X=4.965 $Y=2.72 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_448_n N_A_730_297#_c_588_n 0.00938745f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_342 N_Y_c_550_n N_A_730_297#_M1000_s 0.00325521f $X=4.08 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_343 N_Y_M1003_s N_A_730_297#_c_582_n 0.00312348f $X=4.07 $Y=1.485 $X2=0 $Y2=0
cc_344 N_Y_c_550_n N_A_730_297#_c_582_n 0.00506389f $X=4.08 $Y=1.87 $X2=0 $Y2=0
cc_345 N_Y_c_556_n N_A_730_297#_c_582_n 0.0112811f $X=4.205 $Y=1.87 $X2=0 $Y2=0
cc_346 N_Y_c_550_n N_A_730_297#_c_588_n 0.0116461f $X=4.08 $Y=1.87 $X2=0 $Y2=0
cc_347 N_Y_M1012_d N_VGND_c_607_n 0.00216833f $X=2.775 $Y=0.235 $X2=0 $Y2=0
cc_348 N_Y_M1012_d N_A_471_47#_c_704_n 0.00304656f $X=2.775 $Y=0.235 $X2=0 $Y2=0
cc_349 N_Y_c_533_n N_A_471_47#_c_704_n 0.0164158f $X=2.91 $Y=0.73 $X2=0 $Y2=0
cc_350 N_Y_c_531_n N_A_471_47#_c_704_n 0.00362427f $X=2.98 $Y=1.31 $X2=0 $Y2=0
cc_351 N_Y_c_533_n N_A_471_47#_c_699_n 0.00729487f $X=2.91 $Y=0.73 $X2=0 $Y2=0
cc_352 N_VGND_c_607_n N_A_113_47#_M1010_s 0.00218529f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_353 N_VGND_c_607_n N_A_113_47#_M1005_d 0.00218617f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_600_n N_A_113_47#_c_677_n 0.0114667f $X=1.875 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_607_n N_A_113_47#_c_677_n 0.00913547f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_596_n N_A_113_47#_c_676_n 0.0154056f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_357 N_VGND_c_600_n N_A_113_47#_c_682_n 0.0378883f $X=1.875 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_607_n N_A_113_47#_c_682_n 0.031469f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_359 N_VGND_c_607_n N_A_471_47#_M1012_s 0.00217543f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_360 N_VGND_c_607_n N_A_471_47#_M1015_s 0.0024331f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_607_n N_A_471_47#_M1001_d 0.00215201f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_607_n N_A_471_47#_M1007_s 0.00209319f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_602_n N_A_471_47#_c_709_n 0.0176639f $X=3.7 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_607_n N_A_471_47#_c_709_n 0.0107533f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_M1006_d N_A_471_47#_c_698_n 0.00165819f $X=3.65 $Y=0.235 $X2=0
+ $Y2=0
cc_366 N_VGND_c_598_n N_A_471_47#_c_698_n 0.0116528f $X=3.785 $Y=0.39 $X2=0
+ $Y2=0
cc_367 N_VGND_c_602_n N_A_471_47#_c_698_n 0.00193763f $X=3.7 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_604_n N_A_471_47#_c_698_n 0.00193763f $X=4.54 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_607_n N_A_471_47#_c_698_n 0.00827287f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_604_n N_A_471_47#_c_718_n 0.0188551f $X=4.54 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_607_n N_A_471_47#_c_718_n 0.0122069f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_M1009_s N_A_471_47#_c_700_n 0.00162089f $X=4.49 $Y=0.235 $X2=0
+ $Y2=0
cc_373 N_VGND_c_599_n N_A_471_47#_c_700_n 0.0122559f $X=4.625 $Y=0.39 $X2=0
+ $Y2=0
cc_374 N_VGND_c_604_n N_A_471_47#_c_700_n 0.00198695f $X=4.54 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_606_n N_A_471_47#_c_700_n 0.00198695f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_c_607_n N_A_471_47#_c_700_n 0.00835832f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_377 N_VGND_c_606_n N_A_471_47#_c_701_n 0.0209752f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_607_n N_A_471_47#_c_701_n 0.0124119f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_597_n N_A_471_47#_c_702_n 0.0169665f $X=1.96 $Y=0.39 $X2=0 $Y2=0
cc_380 N_VGND_c_602_n N_A_471_47#_c_702_n 0.0526207f $X=3.7 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_c_607_n N_A_471_47#_c_702_n 0.0330071f $X=5.29 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a32oi_1.pxi.spice
* Created: Tue Sep  1 18:55:53 2020
* 
x_PM_SKY130_FD_SC_HD__A32OI_1%B2 N_B2_c_54_n N_B2_M1008_g N_B2_M1006_g B2
+ N_B2_c_56_n PM_SKY130_FD_SC_HD__A32OI_1%B2
x_PM_SKY130_FD_SC_HD__A32OI_1%B1 N_B1_M1000_g N_B1_M1001_g N_B1_c_80_n
+ N_B1_c_81_n B1 N_B1_c_82_n PM_SKY130_FD_SC_HD__A32OI_1%B1
x_PM_SKY130_FD_SC_HD__A32OI_1%A1 N_A1_M1003_g N_A1_M1007_g N_A1_c_124_n
+ N_A1_c_125_n N_A1_c_126_n A1 N_A1_c_127_n PM_SKY130_FD_SC_HD__A32OI_1%A1
x_PM_SKY130_FD_SC_HD__A32OI_1%A2 N_A2_M1004_g N_A2_M1005_g N_A2_c_169_n
+ N_A2_c_170_n N_A2_c_171_n A2 A2 A2 N_A2_c_174_n PM_SKY130_FD_SC_HD__A32OI_1%A2
x_PM_SKY130_FD_SC_HD__A32OI_1%A3 N_A3_M1009_g N_A3_M1002_g A3 N_A3_c_209_n
+ N_A3_c_210_n N_A3_c_213_n A3 PM_SKY130_FD_SC_HD__A32OI_1%A3
x_PM_SKY130_FD_SC_HD__A32OI_1%A_27_297# N_A_27_297#_M1006_s N_A_27_297#_M1001_d
+ N_A_27_297#_M1005_d N_A_27_297#_c_232_n N_A_27_297#_c_233_n
+ N_A_27_297#_c_236_n N_A_27_297#_c_240_n N_A_27_297#_c_242_n
+ N_A_27_297#_c_245_n N_A_27_297#_c_249_n PM_SKY130_FD_SC_HD__A32OI_1%A_27_297#
x_PM_SKY130_FD_SC_HD__A32OI_1%Y N_Y_M1000_d N_Y_M1006_d N_Y_c_278_n N_Y_c_272_n
+ N_Y_c_273_n Y PM_SKY130_FD_SC_HD__A32OI_1%Y
x_PM_SKY130_FD_SC_HD__A32OI_1%VPWR N_VPWR_M1007_d N_VPWR_M1002_d N_VPWR_c_309_n
+ N_VPWR_c_310_n VPWR N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n
+ N_VPWR_c_308_n N_VPWR_c_315_n N_VPWR_c_316_n PM_SKY130_FD_SC_HD__A32OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A32OI_1%VGND N_VGND_M1008_s N_VGND_M1009_d N_VGND_c_349_n
+ N_VGND_c_350_n N_VGND_c_351_n VGND N_VGND_c_352_n N_VGND_c_353_n
+ N_VGND_c_354_n N_VGND_c_355_n PM_SKY130_FD_SC_HD__A32OI_1%VGND
cc_1 VNB N_B2_c_54_n 0.0202658f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB B2 0.0153414f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_B2_c_56_n 0.0349095f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B1_c_80_n 9.56732e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_5 VNB N_B1_c_81_n 0.0253422f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_6 VNB N_B1_c_82_n 0.0176733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A1_c_124_n 0.00147725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_c_125_n 0.0055817f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_9 VNB N_A1_c_126_n 0.0222373f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_10 VNB N_A1_c_127_n 0.0169271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_169_n 0.0121906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_170_n 0.0146127f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_13 VNB N_A2_c_171_n 0.00166423f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_14 VNB A2 0.00195631f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_15 VNB A2 0.00226642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_174_n 0.00984986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A3_c_209_n 0.0401975f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_18 VNB N_A3_c_210_n 0.0188436f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_19 VNB A3 0.0132445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB Y 0.0028102f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_21 VNB N_VPWR_c_308_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_349_n 0.010303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_350_n 0.0120801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_351_n 0.025126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_352_n 0.0515977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_353_n 0.0188498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_354_n 0.197873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_355_n 0.00523789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_B2_M1006_g 0.0253571f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_30 VPB B2 0.00454807f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_31 VPB N_B2_c_56_n 0.0111443f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_32 VPB N_B1_M1001_g 0.0197495f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB N_B1_c_80_n 0.00130595f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_34 VPB N_B1_c_81_n 0.00610571f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_35 VPB B1 0.00525172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A1_M1007_g 0.0205227f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A1_c_126_n 0.00478553f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_38 VPB N_A2_c_171_n 0.0246285f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_39 VPB A2 0.0018642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A3_c_209_n 0.0186734f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_41 VPB N_A3_c_213_n 0.0184936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB A3 0.00288317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_297#_c_232_n 0.00929745f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_44 VPB N_A_27_297#_c_233_n 0.0165453f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_45 VPB Y 0.00105516f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_46 VPB N_VPWR_c_309_n 0.00449567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_310_n 0.041319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_311_n 0.0395083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_312_n 0.0148112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_313_n 0.0188498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_308_n 0.0611355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_315_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_316_n 0.005212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 N_B2_M1006_g N_B1_M1001_g 0.0407931f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_55 N_B2_c_56_n N_B1_c_80_n 3.66234e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_56 N_B2_c_56_n N_B1_c_81_n 0.0203794f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_57 N_B2_c_54_n N_B1_c_82_n 0.0492854f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_58 B2 N_A_27_297#_c_233_n 0.0090825f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_59 N_B2_c_56_n N_A_27_297#_c_233_n 0.0015323f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_60 N_B2_M1006_g N_A_27_297#_c_236_n 0.0123483f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_61 N_B2_c_54_n N_Y_c_272_n 0.0103957f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_62 N_B2_c_54_n N_Y_c_273_n 0.00128602f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_63 N_B2_c_54_n Y 0.00877717f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_64 N_B2_M1006_g Y 0.0275786f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_65 B2 Y 0.023122f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B2_c_56_n Y 0.00719527f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B2_M1006_g N_VPWR_c_311_n 0.00357877f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_68 N_B2_M1006_g N_VPWR_c_308_n 0.00620762f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 N_B2_c_54_n N_VGND_c_350_n 0.0113548f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_70 B2 N_VGND_c_350_n 0.00830991f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_71 N_B2_c_56_n N_VGND_c_350_n 0.00148403f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B2_c_54_n N_VGND_c_352_n 0.00434443f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_73 N_B2_c_54_n N_VGND_c_354_n 0.00690194f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_74 N_B1_M1001_g N_A1_M1007_g 0.0220324f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_75 N_B1_c_80_n N_A1_M1007_g 0.00173558f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_76 B1 N_A1_M1007_g 0.00507615f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_77 N_B1_c_80_n N_A1_c_124_n 0.0028638f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B1_c_81_n N_A1_c_124_n 2.39197e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B1_c_82_n N_A1_c_124_n 0.0010221f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B1_c_80_n N_A1_c_125_n 0.0118357f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B1_c_81_n N_A1_c_125_n 0.00113072f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_82 B1 N_A1_c_125_n 0.0019068f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_83 N_B1_c_80_n N_A1_c_126_n 9.10793e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B1_c_81_n N_A1_c_126_n 0.0208367f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_85 N_B1_c_82_n N_A1_c_127_n 0.0160279f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_86 B1 N_A_27_297#_M1001_d 0.00554787f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_87 N_B1_M1001_g N_A_27_297#_c_236_n 0.0131406f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_88 B1 N_A_27_297#_c_236_n 0.00430008f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_89 N_B1_M1001_g N_A_27_297#_c_240_n 0.00165031f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_90 B1 N_A_27_297#_c_240_n 0.0131155f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_91 N_B1_M1001_g N_A_27_297#_c_242_n 0.00537132f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B1_c_80_n N_Y_c_278_n 0.00989733f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B1_c_81_n N_Y_c_278_n 0.00201029f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_94 B1 N_Y_c_278_n 0.00447179f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_95 N_B1_c_82_n N_Y_c_278_n 0.0126382f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B1_c_82_n N_Y_c_273_n 0.00594627f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B1_M1001_g Y 0.0123247f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B1_c_80_n Y 0.0307182f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B1_c_81_n Y 0.00317882f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_100 B1 Y 0.0149198f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_101 N_B1_c_82_n Y 0.00419585f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_M1001_g N_VPWR_c_311_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_M1001_g N_VPWR_c_308_n 0.00567715f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B1_c_82_n N_VGND_c_350_n 0.00188123f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B1_c_82_n N_VGND_c_352_n 0.00422612f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B1_c_82_n N_VGND_c_354_n 0.00620852f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A1_c_125_n N_A2_c_169_n 0.00108368f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A1_c_126_n N_A2_c_169_n 0.0205778f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A1_c_124_n N_A2_c_170_n 0.00158817f $X=1.5 $Y=1.075 $X2=0 $Y2=0
cc_110 A1 N_A2_c_170_n 0.0036992f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_111 N_A1_c_127_n N_A2_c_170_n 0.0511901f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A1_M1007_g N_A2_c_171_n 0.0457588f $X=1.47 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A1_c_124_n A2 0.00474205f $X=1.5 $Y=1.075 $X2=0 $Y2=0
cc_114 N_A1_c_124_n A2 0.00516426f $X=1.5 $Y=1.075 $X2=0 $Y2=0
cc_115 N_A1_c_125_n A2 0.0122656f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_c_126_n A2 7.22727e-19 $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A1_c_125_n N_A_27_297#_c_240_n 0.00292515f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A1_c_126_n N_A_27_297#_c_240_n 0.00115446f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A1_M1007_g N_A_27_297#_c_245_n 0.0113304f $X=1.47 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A1_c_125_n N_A_27_297#_c_245_n 0.00551178f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_121 A1 N_Y_c_278_n 0.0105542f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_122 N_A1_c_127_n N_Y_c_278_n 0.00141321f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_123 A1 N_Y_c_273_n 0.0167625f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_124 N_A1_c_127_n N_Y_c_273_n 0.0033207f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A1_M1007_g N_VPWR_c_309_n 0.00302074f $X=1.47 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A1_M1007_g N_VPWR_c_311_n 0.00585385f $X=1.47 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A1_M1007_g N_VPWR_c_308_n 0.00628264f $X=1.47 $Y=1.985 $X2=0 $Y2=0
cc_128 A1 N_VGND_c_351_n 0.00186073f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_129 A1 N_VGND_c_352_n 0.011626f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_130 N_A1_c_127_n N_VGND_c_352_n 0.00391163f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_131 A1 N_VGND_c_354_n 0.0102069f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_132 N_A1_c_127_n N_VGND_c_354_n 0.00607465f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_133 A1 A_309_47# 0.00996883f $X=1.535 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_134 N_A2_c_169_n N_A3_c_209_n 0.0293426f $X=1.9 $Y=1.095 $X2=0 $Y2=0
cc_135 A2 N_A3_c_209_n 0.00271019f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A2_c_170_n N_A3_c_210_n 0.027053f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_137 A2 N_A3_c_210_n 0.00760279f $X=1.995 $Y=0.425 $X2=0 $Y2=0
cc_138 N_A2_c_171_n N_A3_c_213_n 0.0208129f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A2_c_169_n A3 2.59282e-19 $X=1.9 $Y=1.095 $X2=0 $Y2=0
cc_140 A2 A3 0.0251977f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A2_c_171_n N_A_27_297#_c_245_n 0.0110474f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_142 A2 N_A_27_297#_c_245_n 0.00576625f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A2_c_171_n N_A_27_297#_c_249_n 4.30096e-19 $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_144 A2 N_A_27_297#_c_249_n 0.0065805f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A2_c_171_n N_VPWR_c_309_n 0.00152357f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_171_n N_VPWR_c_310_n 0.00182011f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A2_c_171_n N_VPWR_c_312_n 0.00585385f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A2_c_171_n N_VPWR_c_308_n 0.00596375f $X=1.9 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A2_c_170_n N_VGND_c_351_n 0.00185475f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_150 A2 N_VGND_c_351_n 0.026809f $X=1.995 $Y=0.425 $X2=0 $Y2=0
cc_151 N_A2_c_170_n N_VGND_c_352_n 0.00585385f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_152 A2 N_VGND_c_352_n 0.00662354f $X=1.995 $Y=0.425 $X2=0 $Y2=0
cc_153 N_A2_c_170_n N_VGND_c_354_n 0.0108797f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_154 A2 N_VGND_c_354_n 0.00691408f $X=1.995 $Y=0.425 $X2=0 $Y2=0
cc_155 A2 A_383_47# 0.0106711f $X=1.995 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_156 N_A3_c_209_n N_VPWR_c_310_n 0.00775775f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A3_c_213_n N_VPWR_c_310_n 0.0189473f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_158 A3 N_VPWR_c_310_n 0.0251877f $X=2.57 $Y=1.19 $X2=0 $Y2=0
cc_159 N_A3_c_213_n N_VPWR_c_312_n 0.00427505f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A3_c_213_n N_VPWR_c_308_n 0.00732923f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A3_c_209_n N_VGND_c_351_n 0.00729453f $X=2.51 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A3_c_210_n N_VGND_c_351_n 0.0150941f $X=2.465 $Y=0.96 $X2=0 $Y2=0
cc_163 A3 N_VGND_c_351_n 0.021388f $X=2.57 $Y=1.19 $X2=0 $Y2=0
cc_164 N_A3_c_210_n N_VGND_c_352_n 0.00427505f $X=2.465 $Y=0.96 $X2=0 $Y2=0
cc_165 N_A3_c_210_n N_VGND_c_354_n 0.00752764f $X=2.465 $Y=0.96 $X2=0 $Y2=0
cc_166 N_A_27_297#_c_236_n N_Y_M1006_d 0.00314797f $X=1.095 $Y=2.36 $X2=0 $Y2=0
cc_167 N_A_27_297#_c_236_n Y 0.0167443f $X=1.095 $Y=2.36 $X2=0 $Y2=0
cc_168 N_A_27_297#_c_240_n Y 0.0111439f $X=1.22 $Y=1.955 $X2=0 $Y2=0
cc_169 N_A_27_297#_c_242_n Y 0.00780437f $X=1.22 $Y=2.255 $X2=0 $Y2=0
cc_170 N_A_27_297#_c_245_n N_VPWR_M1007_d 0.00761626f $X=2.015 $Y=1.87 $X2=-0.19
+ $Y2=1.305
cc_171 N_A_27_297#_c_245_n N_VPWR_c_309_n 0.0117423f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_c_249_n N_VPWR_c_310_n 0.054752f $X=2.1 $Y=1.91 $X2=0 $Y2=0
cc_173 N_A_27_297#_c_232_n N_VPWR_c_311_n 0.0179721f $X=0.215 $Y=2.255 $X2=0
+ $Y2=0
cc_174 N_A_27_297#_c_236_n N_VPWR_c_311_n 0.0411774f $X=1.095 $Y=2.36 $X2=0
+ $Y2=0
cc_175 N_A_27_297#_c_242_n N_VPWR_c_311_n 0.0173363f $X=1.22 $Y=2.255 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_c_249_n N_VPWR_c_312_n 0.0116529f $X=2.1 $Y=1.91 $X2=0 $Y2=0
cc_177 N_A_27_297#_M1006_s N_VPWR_c_308_n 0.00209324f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_M1001_d N_VPWR_c_308_n 0.0037296f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_179 N_A_27_297#_M1005_d N_VPWR_c_308_n 0.0045801f $X=1.965 $Y=1.485 $X2=0
+ $Y2=0
cc_180 N_A_27_297#_c_232_n N_VPWR_c_308_n 0.00998795f $X=0.215 $Y=2.255 $X2=0
+ $Y2=0
cc_181 N_A_27_297#_c_236_n N_VPWR_c_308_n 0.0266165f $X=1.095 $Y=2.36 $X2=0
+ $Y2=0
cc_182 N_A_27_297#_c_242_n N_VPWR_c_308_n 0.00962794f $X=1.22 $Y=2.255 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_c_245_n N_VPWR_c_308_n 0.0138845f $X=2.015 $Y=1.87 $X2=0
+ $Y2=0
cc_184 N_A_27_297#_c_249_n N_VPWR_c_308_n 0.00647979f $X=2.1 $Y=1.91 $X2=0 $Y2=0
cc_185 N_Y_M1006_d N_VPWR_c_308_n 0.00216833f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_186 N_Y_c_273_n N_VGND_c_350_n 0.00527345f $X=1.08 $Y=0.53 $X2=0 $Y2=0
cc_187 N_Y_c_278_n N_VGND_c_352_n 0.00341195f $X=0.915 $Y=0.72 $X2=0 $Y2=0
cc_188 N_Y_c_272_n N_VGND_c_352_n 0.002702f $X=0.685 $Y=0.72 $X2=0 $Y2=0
cc_189 N_Y_c_273_n N_VGND_c_352_n 0.0120832f $X=1.08 $Y=0.53 $X2=0 $Y2=0
cc_190 N_Y_M1000_d N_VGND_c_354_n 0.0118326f $X=0.925 $Y=0.235 $X2=0 $Y2=0
cc_191 N_Y_c_278_n N_VGND_c_354_n 0.005807f $X=0.915 $Y=0.72 $X2=0 $Y2=0
cc_192 N_Y_c_272_n N_VGND_c_354_n 0.00496107f $X=0.685 $Y=0.72 $X2=0 $Y2=0
cc_193 N_Y_c_273_n N_VGND_c_354_n 0.00924136f $X=1.08 $Y=0.53 $X2=0 $Y2=0
cc_194 N_Y_c_278_n A_109_47# 0.00177909f $X=0.915 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_195 N_Y_c_272_n A_109_47# 0.00151733f $X=0.685 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_196 Y A_109_47# 8.77739e-19 $X=0.595 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_197 N_VGND_c_354_n A_109_47# 0.00268395f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_198 N_VGND_c_354_n A_309_47# 0.00393634f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_199 N_VGND_c_354_n A_383_47# 0.00740685f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__nand4bb_4.spice
* Created: Thu Aug 27 14:31:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand4bb_4.pex.spice"
.subckt sky130_fd_sc_hd__nand4bb_4  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_A_N_M1031_g N_A_27_47#_M1031_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1015 N_A_193_47#_M1015_d N_B_N_M1015_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.65
+ AD=0.32175 AS=0.08775 PD=2.29 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1014_d N_A_27_47#_M1014_g N_A_432_47#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1014_d N_A_27_47#_M1019_g N_A_432_47#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1021 N_Y_M1021_d N_A_27_47#_M1021_g N_A_432_47#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1027 N_Y_M1021_d N_A_27_47#_M1027_g N_A_432_47#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1017 N_A_432_47#_M1027_s N_A_193_47#_M1017_g N_A_850_47#_M1017_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1025 N_A_432_47#_M1025_d N_A_193_47#_M1025_g N_A_850_47#_M1017_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1028 N_A_432_47#_M1025_d N_A_193_47#_M1028_g N_A_850_47#_M1028_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1034 N_A_432_47#_M1034_d N_A_193_47#_M1034_g N_A_850_47#_M1028_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_1266_47#_M1003_d N_C_M1003_g N_A_850_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1885 AS=0.08775 PD=1.88 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1022 N_A_1266_47#_M1022_d N_C_M1022_g N_A_850_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1032 N_A_1266_47#_M1022_d N_C_M1032_g N_A_850_47#_M1032_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1033 N_A_1266_47#_M1033_d N_C_M1033_g N_A_850_47#_M1032_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1002 N_A_1266_47#_M1033_d N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1005 N_A_1266_47#_M1005_d N_D_M1005_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1008 N_A_1266_47#_M1005_d N_D_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1029 N_A_1266_47#_M1029_d N_D_M1029_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.08775 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1023 N_VPWR_M1023_d N_A_N_M1023_g N_A_27_47#_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1006 N_A_193_47#_M1006_d N_B_N_M1006_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=1
+ AD=0.495 AS=0.135 PD=2.99 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.4 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_27_47#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75007.3 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_47#_M1010_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75006.9 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1010_d N_A_27_47#_M1018_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75006.5 A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_A_27_47#_M1024_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75006.1 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1024_d N_A_193_47#_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75005.7 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_193_47#_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1001_d N_A_193_47#_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1030 N_VPWR_M1030_d N_A_193_47#_M1030_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.555 AS=0.135 PD=2.11 PS=1.27 NRD=8.8453 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1030_d N_C_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.555
+ AS=0.135 PD=2.11 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75004.4 SB=75003.1
+ A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_C_M1016_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.8 SB=75002.7
+ A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1016_d N_C_M1020_g N_Y_M1020_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.2 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1026 N_VPWR_M1026_d N_C_M1026_g N_Y_M1020_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.6 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.1 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1009 N_Y_M1004_d N_D_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.5 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1013 N_Y_M1013_d N_D_M1013_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.9 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1035 N_Y_M1013_d N_D_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.3 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX36_noxref VNB VPB NWDIODE A=16.8525 P=24.21
c_75 VNB 0 2.7311e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__nand4bb_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__einvp_4.pex.spice
* Created: Tue Sep  1 19:08:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVP_4%TE 1 3 6 8 9 10 12 13 15 17 18 20 22 23 25
+ 27 28 29 30 31 32
c82 30 0 9.62962e-20 $X=1.75 $Y=1.035
c83 29 0 9.62962e-20 $X=1.33 $Y=1.035
c84 23 0 4.50788e-20 $X=2.095 $Y=1.035
c85 18 0 1.96823e-19 $X=1.675 $Y=1.035
r86 36 38 31.8035 $w=3.41e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.142
+ $X2=0.47 $Y2=1.142
r87 31 32 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r88 31 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r89 25 27 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.17 $Y=0.96 $X2=2.17
+ $Y2=0.56
r90 24 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.035
+ $X2=1.75 $Y2=1.035
r91 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.095 $Y=1.035
+ $X2=2.17 $Y2=0.96
r92 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.095 $Y=1.035
+ $X2=1.825 $Y2=1.035
r93 20 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=0.96
+ $X2=1.75 $Y2=1.035
r94 20 22 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.75 $Y=0.96 $X2=1.75
+ $Y2=0.56
r95 19 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.405 $Y=1.035
+ $X2=1.33 $Y2=1.035
r96 18 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.035
+ $X2=1.75 $Y2=1.035
r97 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.675 $Y=1.035
+ $X2=1.405 $Y2=1.035
r98 15 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.33 $Y=0.96
+ $X2=1.33 $Y2=1.035
r99 15 17 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.33 $Y=0.96 $X2=1.33
+ $Y2=0.56
r100 14 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.965 $Y=1.035
+ $X2=0.89 $Y2=1.035
r101 13 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.255 $Y=1.035
+ $X2=1.33 $Y2=1.035
r102 13 14 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.255 $Y=1.035
+ $X2=0.965 $Y2=1.035
r103 10 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=0.96
+ $X2=0.89 $Y2=1.035
r104 10 12 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.89 $Y=0.96 $X2=0.89
+ $Y2=0.56
r105 9 38 25.9675 $w=3.41e-07 $l=1.39549e-07 $layer=POLY_cond $X=0.545 $Y=1.035
+ $X2=0.47 $Y2=1.142
r106 8 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.815 $Y=1.035
+ $X2=0.89 $Y2=1.035
r107 8 9 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.815 $Y=1.035
+ $X2=0.545 $Y2=1.035
r108 4 38 22.0049 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.142
r109 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r110 1 38 22.0049 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.47 $Y=0.96
+ $X2=0.47 $Y2=1.142
r111 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.47 $Y=0.96 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_4%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 23 27 31 35 37 38 40 43 44 54
c105 54 0 1.9418e-19 $X=0.687 $Y=1.16
c106 23 0 1.50055e-19 $X=1.83 $Y=1.395
c107 20 0 2.43799e-19 $X=2.67 $Y=1.47
c108 15 0 7.37964e-20 $X=2.175 $Y=1.395
c109 11 0 1.86371e-19 $X=1.485 $Y=1.395
c110 10 0 7.37964e-20 $X=1.755 $Y=1.395
r111 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.16 $X2=2.61 $Y2=1.16
r112 41 54 0.820356 $w=3.3e-07 $l=1.88e-07 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=0.687 $Y2=1.16
r113 41 43 60.5906 $w=3.28e-07 $l=1.735e-06 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=2.61 $Y2=1.16
r114 39 54 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=0.687 $Y=1.325
+ $X2=0.687 $Y2=1.16
r115 39 40 14.1366 $w=3.73e-07 $l=4.6e-07 $layer=LI1_cond $X=0.687 $Y=1.325
+ $X2=0.687 $Y2=1.785
r116 38 54 5.82594 $w=2.85e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.597 $Y=0.995
+ $X2=0.687 $Y2=1.16
r117 37 38 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.597 $Y=0.825
+ $X2=0.597 $Y2=0.995
r118 33 40 30.7936 $w=1.68e-07 $l=4.72e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.687 $Y2=1.87
r119 33 35 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=1.955
+ $X2=0.215 $Y2=2.165
r120 29 37 24.9219 $w=1.68e-07 $l=3.82e-07 $layer=LI1_cond $X=0.215 $Y=0.74
+ $X2=0.597 $Y2=0.74
r121 29 31 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r122 26 44 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=2.61 $Y=1.32
+ $X2=2.61 $Y2=1.16
r123 26 27 30.766 $w=1.5e-07 $l=6e-08 $layer=POLY_cond $X=2.61 $Y=1.395 $X2=2.67
+ $Y2=1.395
r124 24 26 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.25 $Y=1.395
+ $X2=2.61 $Y2=1.395
r125 20 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=1.47
+ $X2=2.67 $Y2=1.395
r126 20 22 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.67 $Y=1.47
+ $X2=2.67 $Y2=2.015
r127 17 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=1.47
+ $X2=2.25 $Y2=1.395
r128 17 19 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.25 $Y=1.47
+ $X2=2.25 $Y2=2.015
r129 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.395
+ $X2=1.83 $Y2=1.395
r130 15 24 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.175 $Y=1.395
+ $X2=2.25 $Y2=1.395
r131 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.175 $Y=1.395
+ $X2=1.905 $Y2=1.395
r132 12 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.47
+ $X2=1.83 $Y2=1.395
r133 12 14 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.83 $Y=1.47
+ $X2=1.83 $Y2=2.015
r134 10 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=1.395
+ $X2=1.83 $Y2=1.395
r135 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.755 $Y=1.395
+ $X2=1.485 $Y2=1.395
r136 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.47
+ $X2=1.485 $Y2=1.395
r137 7 9 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.41 $Y=1.47
+ $X2=1.41 $Y2=2.015
r138 2 35 600 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.165
r139 1 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_4%A 1 3 6 8 10 13 17 21 23 25 29 31 32 33
r75 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.585
+ $Y=1.16 $X2=4.585 $Y2=1.16
r76 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.245
+ $Y=1.16 $X2=4.245 $Y2=1.16
r77 38 40 55.5525 $w=2.95e-07 $l=3.4e-07 $layer=POLY_cond $X=3.565 $Y=1.16
+ $X2=3.905 $Y2=1.16
r78 37 38 68.6237 $w=2.95e-07 $l=4.2e-07 $layer=POLY_cond $X=3.145 $Y=1.16
+ $X2=3.565 $Y2=1.16
r79 33 49 12.2023 $w=2.53e-07 $l=2.7e-07 $layer=LI1_cond $X=4.855 $Y=1.147
+ $X2=4.585 $Y2=1.147
r80 32 49 8.58683 $w=2.53e-07 $l=1.9e-07 $layer=LI1_cond $X=4.395 $Y=1.147
+ $X2=4.585 $Y2=1.147
r81 32 45 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=4.395 $Y=1.147
+ $X2=4.245 $Y2=1.147
r82 31 45 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=3.905 $Y=1.147
+ $X2=4.245 $Y2=1.147
r83 31 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.905
+ $Y=1.16 $X2=3.905 $Y2=1.16
r84 23 48 29.4102 $w=2.95e-07 $l=1.8e-07 $layer=POLY_cond $X=4.405 $Y=1.16
+ $X2=4.585 $Y2=1.16
r85 23 44 26.1424 $w=2.95e-07 $l=1.6e-07 $layer=POLY_cond $X=4.405 $Y=1.16
+ $X2=4.245 $Y2=1.16
r86 23 29 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.405 $Y=1.305
+ $X2=4.405 $Y2=1.985
r87 23 25 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.405 $Y=1.015
+ $X2=4.405 $Y2=0.56
r88 15 44 42.4814 $w=2.95e-07 $l=2.6e-07 $layer=POLY_cond $X=3.985 $Y=1.16
+ $X2=4.245 $Y2=1.16
r89 15 40 13.0712 $w=2.95e-07 $l=8e-08 $layer=POLY_cond $X=3.985 $Y=1.16
+ $X2=3.905 $Y2=1.16
r90 15 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.985 $Y=1.295
+ $X2=3.985 $Y2=1.985
r91 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.985 $Y=1.025
+ $X2=3.985 $Y2=0.56
r92 11 38 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=1.16
r93 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=1.985
r94 8 38 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=1.16
r95 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=0.56
r96 4 37 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.325
+ $X2=3.145 $Y2=1.16
r97 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.145 $Y=1.325
+ $X2=3.145 $Y2=1.985
r98 1 37 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=1.16
r99 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_4%VPWR 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
r71 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r74 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r75 42 45 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r76 42 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 41 44 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r78 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 39 54 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.475 $Y2=2.72
r80 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.655 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r82 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r83 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r84 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r85 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r86 34 54 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.475 $Y2=2.72
r87 34 37 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r89 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r91 30 48 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.695 $Y2=2.72
r92 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r93 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r94 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r95 24 48 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.695 $Y2=2.72
r96 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r98 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r99 18 54 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=2.635
+ $X2=2.475 $Y2=2.72
r100 18 20 19.6876 $w=3.58e-07 $l=6.15e-07 $layer=LI1_cond $X=2.475 $Y=2.635
+ $X2=2.475 $Y2=2.02
r101 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r102 14 16 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.02
r103 10 48 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r104 10 12 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.34
r105 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=1.545 $X2=2.46 $Y2=2.02
r106 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.545 $X2=1.62 $Y2=2.02
r107 1 12 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_4%A_215_309# 1 2 3 4 5 18 20 21 24 26 31 32 33
+ 36 38 40 43 44
c64 26 0 4.50788e-20 $X=2.825 $Y=1.64
c65 20 0 3.89415e-19 $X=1.955 $Y=1.64
r66 40 42 9.18427 $w=4.45e-07 $l=3.35e-07 $layer=LI1_cond $X=4.752 $Y=2.295
+ $X2=4.752 $Y2=1.96
r67 39 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=2.38
+ $X2=3.775 $Y2=2.38
r68 38 40 8.76165 $w=1.7e-07 $l=2.61063e-07 $layer=LI1_cond $X=4.53 $Y=2.38
+ $X2=4.752 $Y2=2.295
r69 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.53 $Y=2.38
+ $X2=3.86 $Y2=2.38
r70 34 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=2.295
+ $X2=3.775 $Y2=2.38
r71 34 36 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.775 $Y=2.295
+ $X2=3.775 $Y2=1.96
r72 32 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.38
+ $X2=3.775 $Y2=2.38
r73 32 33 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.69 $Y=2.38
+ $X2=2.995 $Y2=2.38
r74 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.91 $Y=2.295
+ $X2=2.995 $Y2=2.38
r75 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.91 $Y=2.295
+ $X2=2.91 $Y2=1.96
r76 28 31 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.91 $Y=1.725
+ $X2=2.91 $Y2=1.96
r77 27 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=1.64
+ $X2=2.04 $Y2=1.64
r78 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.825 $Y=1.64
+ $X2=2.91 $Y2=1.725
r79 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.825 $Y=1.64
+ $X2=2.125 $Y2=1.64
r80 22 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=1.725
+ $X2=2.04 $Y2=1.64
r81 22 24 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.04 $Y=1.725
+ $X2=2.04 $Y2=1.96
r82 20 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.64
+ $X2=2.04 $Y2=1.64
r83 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=1.64
+ $X2=1.285 $Y2=1.64
r84 16 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.18 $Y=1.725
+ $X2=1.285 $Y2=1.64
r85 16 18 27.1991 $w=2.08e-07 $l=5.15e-07 $layer=LI1_cond $X=1.18 $Y=1.725
+ $X2=1.18 $Y2=2.24
r86 5 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.48
+ $Y=1.485 $X2=4.615 $Y2=1.96
r87 4 36 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.64
+ $Y=1.485 $X2=3.775 $Y2=1.96
r88 3 31 300 $w=1.7e-07 $l=4.90612e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.545 $X2=2.91 $Y2=1.96
r89 2 24 300 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.545 $X2=2.04 $Y2=1.96
r90 1 18 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.545 $X2=1.2 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_4%Z 1 2 3 4 15 19 21 22 23 24 25 47
c55 47 0 1.99481e-19 $X=3.455 $Y=1.87
c56 24 0 4.43179e-20 $X=3.475 $Y=1.53
r57 44 47 2.34525 $w=5.08e-07 $l=1e-07 $layer=LI1_cond $X=3.355 $Y=1.87
+ $X2=3.455 $Y2=1.87
r58 44 45 3.28461 $w=3.3e-07 $l=2.55e-07 $layer=LI1_cond $X=3.355 $Y=1.87
+ $X2=3.355 $Y2=1.615
r59 25 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.935 $Y=1.53
+ $X2=3.57 $Y2=1.53
r60 24 41 4.08752 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.38 $Y=1.53 $X2=3.57
+ $Y2=1.53
r61 24 45 2.70057 $w=3.55e-07 $l=9.66954e-08 $layer=LI1_cond $X=3.38 $Y=1.53
+ $X2=3.355 $Y2=1.615
r62 24 47 9.00371 $w=1.3e-07 $l=2.55e-07 $layer=LI1_cond $X=3.455 $Y=1.615
+ $X2=3.455 $Y2=1.87
r63 23 24 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.38 $Y=1.19
+ $X2=3.38 $Y2=1.445
r64 22 23 9.03758 $w=3.78e-07 $l=2.98e-07 $layer=LI1_cond $X=3.38 $Y=0.892
+ $X2=3.38 $Y2=1.19
r65 19 25 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.03 $Y=1.53
+ $X2=3.935 $Y2=1.53
r66 19 21 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=1.53
+ $X2=4.195 $Y2=1.53
r67 13 22 4.79554 $w=2.15e-07 $l=1.9e-07 $layer=LI1_cond $X=3.57 $Y=0.742
+ $X2=3.38 $Y2=0.742
r68 13 15 33.5013 $w=2.13e-07 $l=6.25e-07 $layer=LI1_cond $X=3.57 $Y=0.742
+ $X2=4.195 $Y2=0.742
r69 4 21 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=4.06
+ $Y=1.485 $X2=4.195 $Y2=1.61
r70 3 24 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.485 $X2=3.355 $Y2=1.61
r71 2 15 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.195 $Y2=0.76
r72 1 22 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.235 $X2=3.355 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_4%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r77 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r78 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r79 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r80 42 52 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.83 $Y=0 $X2=2.53
+ $Y2=0
r81 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r82 39 51 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.555 $Y=0 $X2=2.385
+ $Y2=0
r83 39 41 148.422 $w=1.68e-07 $l=2.275e-06 $layer=LI1_cond $X=2.555 $Y=0
+ $X2=4.83 $Y2=0
r84 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r85 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r86 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r87 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.54
+ $Y2=0
r88 35 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=2.07
+ $Y2=0
r89 34 51 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.385
+ $Y2=0
r90 34 37 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.07
+ $Y2=0
r91 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r92 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r93 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r94 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r95 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r96 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.54
+ $Y2=0
r97 29 32 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.15
+ $Y2=0
r98 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r99 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r100 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r101 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r102 18 51 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0
r103 18 20 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0.36
r104 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0
r105 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0.36
r106 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r107 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r108 3 20 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.36
r109 2 16 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.36
r110 1 12 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_4%A_193_47# 1 2 3 4 5 18 20 21 24 26 31 32 36
+ 38
c57 38 0 1.50055e-19 $X=1.96 $Y=0.74
c58 26 0 7.37964e-20 $X=2.735 $Y=0.74
c59 20 0 2.60168e-19 $X=1.875 $Y=0.74
r60 34 36 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=3.775 $Y=0.36
+ $X2=4.615 $Y2=0.36
r61 32 34 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=3.02 $Y=0.36
+ $X2=3.775 $Y2=0.36
r62 29 31 4.85239 $w=2.83e-07 $l=1.2e-07 $layer=LI1_cond $X=2.877 $Y=0.655
+ $X2=2.877 $Y2=0.535
r63 28 32 7.02201 $w=2.1e-07 $l=1.88319e-07 $layer=LI1_cond $X=2.877 $Y=0.465
+ $X2=3.02 $Y2=0.36
r64 28 31 2.83056 $w=2.83e-07 $l=7e-08 $layer=LI1_cond $X=2.877 $Y=0.465
+ $X2=2.877 $Y2=0.535
r65 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.74
+ $X2=1.96 $Y2=0.74
r66 26 29 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.735 $Y=0.74
+ $X2=2.877 $Y2=0.655
r67 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.735 $Y=0.74
+ $X2=2.045 $Y2=0.74
r68 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.655
+ $X2=1.96 $Y2=0.74
r69 22 24 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.96 $Y=0.655
+ $X2=1.96 $Y2=0.535
r70 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.96 $Y2=0.74
r71 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.205 $Y2=0.74
r72 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.655
+ $X2=1.205 $Y2=0.74
r73 16 18 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.12 $Y=0.655
+ $X2=1.12 $Y2=0.535
r74 5 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.235 $X2=4.615 $Y2=0.36
r75 4 34 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.235 $X2=3.775 $Y2=0.36
r76 3 31 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.235 $X2=2.935 $Y2=0.535
r77 2 24 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.535
r78 1 18 182 $w=1.7e-07 $l=3.69459e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.12 $Y2=0.535
.ends


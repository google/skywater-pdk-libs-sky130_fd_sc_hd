* File: sky130_fd_sc_hd__decap_3.spice
* Created: Thu Aug 27 14:13:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__decap_3.spice.pex"
.subckt sky130_fd_sc_hd__decap_3  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_VPWR_M1001_g N_VGND_M1001_s VNB NSHORT L=0.59 W=0.55
+ AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 M=1 R=0.932203 SA=295000
+ SB=295000 A=0.3245 P=2.28 MULT=1
MM1000 N_VPWR_M1000_s N_VGND_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.59 W=0.87
+ AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 M=1 R=1.47458 SA=295000
+ SB=295000 A=0.5133 P=2.92 MULT=1
DX2_noxref VNB VPB NWDIODE A=2.8248 P=6.73
*
.include "sky130_fd_sc_hd__decap_3.spice.SKY130_FD_SC_HD__DECAP_3.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__o31ai_4.spice.pex
* Created: Thu Aug 27 14:40:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O31AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 54
r91 52 54 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.615 $Y=1.16
+ $X2=1.75 $Y2=1.16
r92 50 52 63.3195 $w=2.7e-07 $l=2.85e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.615 $Y2=1.16
r93 48 50 12.2196 $w=2.7e-07 $l=5.5e-08 $layer=POLY_cond $X=1.275 $Y=1.16
+ $X2=1.33 $Y2=1.16
r94 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.275
+ $Y=1.16 $X2=1.275 $Y2=1.16
r95 46 48 81.0934 $w=2.7e-07 $l=3.65e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.275 $Y2=1.16
r96 44 46 69.9847 $w=2.7e-07 $l=3.15e-07 $layer=POLY_cond $X=0.595 $Y=1.16
+ $X2=0.91 $Y2=1.16
r97 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r98 41 44 23.3282 $w=2.7e-07 $l=1.05e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.595 $Y2=1.16
r99 36 49 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.615 $Y=1.24
+ $X2=1.275 $Y2=1.24
r100 36 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.615
+ $Y=1.16 $X2=1.615 $Y2=1.16
r101 35 49 3.73765 $w=3.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.155 $Y=1.24
+ $X2=1.275 $Y2=1.24
r102 34 35 14.3277 $w=3.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.24
+ $X2=1.155 $Y2=1.24
r103 34 45 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=0.695 $Y=1.24
+ $X2=0.595 $Y2=1.24
r104 33 45 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.235 $Y=1.24
+ $X2=0.595 $Y2=1.24
r105 29 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.75 $Y=1.295
+ $X2=1.75 $Y2=1.16
r106 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.75 $Y=1.295
+ $X2=1.75 $Y2=1.985
r107 25 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.75 $Y=1.025
+ $X2=1.75 $Y2=1.16
r108 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.75 $Y=1.025
+ $X2=1.75 $Y2=0.56
r109 21 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.33 $Y=1.295
+ $X2=1.33 $Y2=1.16
r110 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.33 $Y=1.295
+ $X2=1.33 $Y2=1.985
r111 17 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.33 $Y=1.025
+ $X2=1.33 $Y2=1.16
r112 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.33 $Y=1.025
+ $X2=1.33 $Y2=0.56
r113 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.91 $Y=1.295
+ $X2=0.91 $Y2=1.16
r114 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.91 $Y=1.295
+ $X2=0.91 $Y2=1.985
r115 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.91 $Y=1.025
+ $X2=0.91 $Y2=1.16
r116 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.91 $Y=1.025
+ $X2=0.91 $Y2=0.56
r117 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.49 $Y=1.295
+ $X2=0.49 $Y2=1.16
r118 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.49 $Y=1.295
+ $X2=0.49 $Y2=1.985
r119 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.49 $Y=1.025
+ $X2=0.49 $Y2=1.16
r120 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.49 $Y=1.025
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%A2 3 7 11 15 19 23 27 31 33 34 35 36 54
r92 52 54 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.28 $Y=1.16
+ $X2=3.43 $Y2=1.16
r93 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.28
+ $Y=1.16 $X2=3.28 $Y2=1.16
r94 50 52 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=3.28 $Y2=1.16
r95 48 50 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=2.94 $Y=1.16 $X2=3.01
+ $Y2=1.16
r96 46 48 77.7608 $w=2.7e-07 $l=3.5e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.94 $Y2=1.16
r97 44 46 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.59 $Y2=1.16
r98 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r99 41 44 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.17 $Y=1.16 $X2=2.26
+ $Y2=1.16
r100 36 53 5.45074 $w=3.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.455 $Y=1.24
+ $X2=3.28 $Y2=1.24
r101 35 53 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.94 $Y=1.24 $X2=3.28
+ $Y2=1.24
r102 35 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.94
+ $Y=1.16 $X2=2.94 $Y2=1.16
r103 34 35 12.6146 $w=3.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.535 $Y=1.24
+ $X2=2.94 $Y2=1.24
r104 34 45 8.56545 $w=3.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.535 $Y=1.24
+ $X2=2.26 $Y2=1.24
r105 33 45 5.76222 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.075 $Y=1.24
+ $X2=2.26 $Y2=1.24
r106 29 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.43 $Y=1.295
+ $X2=3.43 $Y2=1.16
r107 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.43 $Y=1.295
+ $X2=3.43 $Y2=1.985
r108 25 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.43 $Y=1.025
+ $X2=3.43 $Y2=1.16
r109 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.43 $Y=1.025
+ $X2=3.43 $Y2=0.56
r110 21 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.01 $Y=1.295
+ $X2=3.01 $Y2=1.16
r111 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.01 $Y=1.295
+ $X2=3.01 $Y2=1.985
r112 17 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.01 $Y=1.025
+ $X2=3.01 $Y2=1.16
r113 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.01 $Y=1.025
+ $X2=3.01 $Y2=0.56
r114 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.59 $Y=1.295
+ $X2=2.59 $Y2=1.16
r115 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.59 $Y=1.295
+ $X2=2.59 $Y2=1.985
r116 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.59 $Y=1.025
+ $X2=2.59 $Y2=1.16
r117 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.59 $Y=1.025
+ $X2=2.59 $Y2=0.56
r118 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.17 $Y=1.295
+ $X2=2.17 $Y2=1.16
r119 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.17 $Y=1.295
+ $X2=2.17 $Y2=1.985
r120 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.17 $Y=1.025
+ $X2=2.17 $Y2=1.16
r121 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.17 $Y=1.025
+ $X2=2.17 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 37 38
+ 44 56
c76 27 0 1.07318e-19 $X=5.645 $Y=0.56
r77 54 56 76.6499 $w=2.7e-07 $l=3.45e-07 $layer=POLY_cond $X=5.3 $Y=1.16
+ $X2=5.645 $Y2=1.16
r78 52 54 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.225 $Y=1.16 $X2=5.3
+ $Y2=1.16
r79 51 52 26.6608 $w=2.7e-07 $l=1.2e-07 $layer=POLY_cond $X=5.105 $Y=1.16
+ $X2=5.225 $Y2=1.16
r80 50 51 66.6521 $w=2.7e-07 $l=3e-07 $layer=POLY_cond $X=4.805 $Y=1.16
+ $X2=5.105 $Y2=1.16
r81 49 50 26.6608 $w=2.7e-07 $l=1.2e-07 $layer=POLY_cond $X=4.685 $Y=1.16
+ $X2=4.805 $Y2=1.16
r82 48 49 66.6521 $w=2.7e-07 $l=3e-07 $layer=POLY_cond $X=4.385 $Y=1.16
+ $X2=4.685 $Y2=1.16
r83 44 48 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.31 $Y=1.16
+ $X2=4.385 $Y2=1.16
r84 44 46 82.2043 $w=2.7e-07 $l=3.7e-07 $layer=POLY_cond $X=4.31 $Y=1.16
+ $X2=3.94 $Y2=1.16
r85 37 38 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=5.29 $Y=1.165
+ $X2=5.75 $Y2=1.165
r86 37 54 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.3
+ $Y=1.16 $X2=5.3 $Y2=1.16
r87 36 37 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=4.83 $Y=1.165
+ $X2=5.29 $Y2=1.165
r88 35 36 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=4.37 $Y=1.165
+ $X2=4.83 $Y2=1.165
r89 34 35 23.8346 $w=2.18e-07 $l=4.55e-07 $layer=LI1_cond $X=3.915 $Y=1.165
+ $X2=4.37 $Y2=1.165
r90 34 46 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.94
+ $Y=1.16 $X2=3.94 $Y2=1.16
r91 33 46 3.33261 $w=2.7e-07 $l=1.5e-08 $layer=POLY_cond $X=3.925 $Y=1.16
+ $X2=3.94 $Y2=1.16
r92 29 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.645 $Y=1.295
+ $X2=5.645 $Y2=1.16
r93 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.645 $Y=1.295
+ $X2=5.645 $Y2=1.985
r94 25 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.645 $Y=1.025
+ $X2=5.645 $Y2=1.16
r95 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.645 $Y=1.025
+ $X2=5.645 $Y2=0.56
r96 21 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.225 $Y=1.295
+ $X2=5.225 $Y2=1.16
r97 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.225 $Y=1.295
+ $X2=5.225 $Y2=1.985
r98 17 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.105 $Y=1.025
+ $X2=5.105 $Y2=1.16
r99 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.105 $Y=1.025
+ $X2=5.105 $Y2=0.56
r100 13 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.805 $Y=1.295
+ $X2=4.805 $Y2=1.16
r101 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.805 $Y=1.295
+ $X2=4.805 $Y2=1.985
r102 9 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.685 $Y=1.025
+ $X2=4.685 $Y2=1.16
r103 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.685 $Y=1.025
+ $X2=4.685 $Y2=0.56
r104 5 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.385 $Y=1.295
+ $X2=4.385 $Y2=1.16
r105 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.385 $Y=1.295
+ $X2=4.385 $Y2=1.985
r106 1 33 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.85 $Y=1.025
+ $X2=3.925 $Y2=1.16
r107 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.85 $Y=1.025
+ $X2=3.85 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%B1 3 7 11 15 19 23 27 31 33 34 35 49
r74 47 49 3.33261 $w=2.7e-07 $l=1.5e-08 $layer=POLY_cond $X=7.31 $Y=1.16
+ $X2=7.325 $Y2=1.16
r75 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.16 $X2=7.31 $Y2=1.16
r76 45 47 89.9803 $w=2.7e-07 $l=4.05e-07 $layer=POLY_cond $X=6.905 $Y=1.16
+ $X2=7.31 $Y2=1.16
r77 43 45 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=6.63 $Y=1.16
+ $X2=6.905 $Y2=1.16
r78 41 43 32.2152 $w=2.7e-07 $l=1.45e-07 $layer=POLY_cond $X=6.485 $Y=1.16
+ $X2=6.63 $Y2=1.16
r79 39 41 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.065 $Y=1.16
+ $X2=6.485 $Y2=1.16
r80 35 48 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=7.59 $Y=1.165
+ $X2=7.31 $Y2=1.165
r81 34 48 9.42908 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=7.13 $Y=1.165
+ $X2=7.31 $Y2=1.165
r82 33 34 26.1919 $w=2.18e-07 $l=5e-07 $layer=LI1_cond $X=6.63 $Y=1.165 $X2=7.13
+ $Y2=1.165
r83 33 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.63
+ $Y=1.16 $X2=6.63 $Y2=1.16
r84 29 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.325 $Y=1.295
+ $X2=7.325 $Y2=1.16
r85 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.325 $Y=1.295
+ $X2=7.325 $Y2=1.985
r86 25 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.325 $Y=1.025
+ $X2=7.325 $Y2=1.16
r87 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.325 $Y=1.025
+ $X2=7.325 $Y2=0.56
r88 21 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.905 $Y=1.295
+ $X2=6.905 $Y2=1.16
r89 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.905 $Y=1.295
+ $X2=6.905 $Y2=1.985
r90 17 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.905 $Y=1.025
+ $X2=6.905 $Y2=1.16
r91 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.905 $Y=1.025
+ $X2=6.905 $Y2=0.56
r92 13 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.485 $Y=1.295
+ $X2=6.485 $Y2=1.16
r93 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.485 $Y=1.295
+ $X2=6.485 $Y2=1.985
r94 9 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.485 $Y=1.025
+ $X2=6.485 $Y2=1.16
r95 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.485 $Y=1.025
+ $X2=6.485 $Y2=0.56
r96 5 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.065 $Y=1.295
+ $X2=6.065 $Y2=1.16
r97 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.065 $Y=1.295
+ $X2=6.065 $Y2=1.985
r98 1 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.065 $Y=1.025
+ $X2=6.065 $Y2=1.16
r99 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.065 $Y=1.025
+ $X2=6.065 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 34 39 45
r73 45 47 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.8 $Y=2.02 $X2=2.8
+ $Y2=2.335
r74 32 47 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=2.335
+ $X2=2.8 $Y2=2.335
r75 32 34 29.9192 $w=2.58e-07 $l=6.75e-07 $layer=LI1_cond $X=2.965 $Y=2.335
+ $X2=3.64 $Y2=2.335
r76 31 43 3.88283 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=2.335
+ $X2=1.96 $Y2=2.335
r77 30 47 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=2.335
+ $X2=2.8 $Y2=2.335
r78 30 31 22.6056 $w=2.58e-07 $l=5.1e-07 $layer=LI1_cond $X=2.635 $Y=2.335
+ $X2=2.125 $Y2=2.335
r79 29 43 3.0592 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=1.96 $Y=2.205 $X2=1.96
+ $Y2=2.335
r80 28 41 3.25553 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.96 $Y=1.895
+ $X2=1.96 $Y2=1.745
r81 28 29 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.96 $Y=1.895
+ $X2=1.96 $Y2=2.205
r82 27 39 5.58832 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=1.745
+ $X2=1.12 $Y2=1.745
r83 26 41 3.58108 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=1.745
+ $X2=1.96 $Y2=1.745
r84 26 27 19.5915 $w=2.98e-07 $l=5.1e-07 $layer=LI1_cond $X=1.795 $Y=1.745
+ $X2=1.285 $Y2=1.745
r85 22 39 1.0017 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.12 $Y=1.895 $X2=1.12
+ $Y2=1.745
r86 22 24 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.12 $Y=1.895
+ $X2=1.12 $Y2=2.36
r87 21 37 3.73322 $w=3e-07 $l=1.78e-07 $layer=LI1_cond $X=0.445 $Y=1.745
+ $X2=0.267 $Y2=1.745
r88 20 39 5.58832 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=1.745
+ $X2=1.12 $Y2=1.745
r89 20 21 19.5915 $w=2.98e-07 $l=5.1e-07 $layer=LI1_cond $X=0.955 $Y=1.745
+ $X2=0.445 $Y2=1.745
r90 16 37 3.14597 $w=3.55e-07 $l=1.5e-07 $layer=LI1_cond $X=0.267 $Y=1.895
+ $X2=0.267 $Y2=1.745
r91 16 18 15.0954 $w=3.53e-07 $l=4.65e-07 $layer=LI1_cond $X=0.267 $Y=1.895
+ $X2=0.267 $Y2=2.36
r92 5 34 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=2.36
r93 4 45 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=2.02
r94 3 43 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.36
r95 3 41 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.68
r96 2 39 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.68
r97 2 24 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.36
r98 1 37 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.68
r99 1 18 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%VPWR 1 2 3 4 17 21 25 29 31 33 38 43 50 51
+ 54 57 60 63
r104 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r105 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r106 57 58 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r108 51 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r109 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r110 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.28 $Y=2.72
+ $X2=7.115 $Y2=2.72
r111 48 50 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.28 $Y=2.72
+ $X2=7.59 $Y2=2.72
r112 47 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r113 47 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r115 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.44 $Y=2.72
+ $X2=6.275 $Y2=2.72
r116 44 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.44 $Y=2.72
+ $X2=6.67 $Y2=2.72
r117 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=2.72
+ $X2=7.115 $Y2=2.72
r118 43 46 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.95 $Y=2.72
+ $X2=6.67 $Y2=2.72
r119 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r120 42 58 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=1.61 $Y2=2.72
r121 41 42 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r122 39 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.54 $Y2=2.72
r123 39 41 269.118 $w=1.68e-07 $l=4.125e-06 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=5.75 $Y2=2.72
r124 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.11 $Y=2.72
+ $X2=6.275 $Y2=2.72
r125 38 41 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.11 $Y=2.72
+ $X2=5.75 $Y2=2.72
r126 37 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r127 37 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r128 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r129 34 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=2.72
+ $X2=0.7 $Y2=2.72
r130 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 33 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.54 $Y2=2.72
r132 33 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r133 31 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r134 27 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.115 $Y=2.635
+ $X2=7.115 $Y2=2.72
r135 27 29 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=7.115 $Y=2.635
+ $X2=7.115 $Y2=2.02
r136 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.275 $Y=2.635
+ $X2=6.275 $Y2=2.72
r137 23 25 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=6.275 $Y=2.635
+ $X2=6.275 $Y2=2.02
r138 19 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2.72
r139 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2.34
r140 15 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2.72
r141 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.34
r142 4 29 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.98
+ $Y=1.485 $X2=7.115 $Y2=2.02
r143 3 25 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.14
+ $Y=1.485 $X2=6.275 $Y2=2.02
r144 2 21 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=2.34
r145 1 17 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%A_449_297# 1 2 3 4 17 19 23 27 28 31
r40 30 31 17.1332 $w=5.98e-07 $l=5.15e-07 $layer=LI1_cond $X=4.595 $Y=2.165
+ $X2=4.08 $Y2=2.165
r41 28 31 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=1.95
+ $X2=4.08 $Y2=1.95
r42 26 28 14.5975 $w=4.38e-07 $l=3.85e-07 $layer=LI1_cond $X=3.22 $Y=1.815
+ $X2=3.605 $Y2=1.815
r43 26 27 6.73996 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=1.815
+ $X2=3.135 $Y2=1.815
r44 17 30 1.69444 $w=5.98e-07 $l=8.5e-08 $layer=LI1_cond $X=4.68 $Y=2.165
+ $X2=4.595 $Y2=2.165
r45 17 19 15.0507 $w=5.98e-07 $l=7.55e-07 $layer=LI1_cond $X=4.68 $Y=2.165
+ $X2=5.435 $Y2=2.165
r46 14 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.68
+ $X2=2.38 $Y2=1.68
r47 14 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.465 $Y=1.68
+ $X2=3.135 $Y2=1.68
r48 4 19 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.3
+ $Y=1.485 $X2=5.435 $Y2=1.95
r49 3 30 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.46
+ $Y=1.485 $X2=4.595 $Y2=1.95
r50 2 26 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.76
r51 1 23 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.76
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%Y 1 2 3 4 5 6 7 24 28 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 62 78 79 85 89 93 101
c75 79 0 1.07318e-19 $X=6.202 $Y=0.885
r76 62 78 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=5.77 $Y=1.57 $X2=5.75
+ $Y2=1.57
r77 41 42 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=7.592 $Y=1.87
+ $X2=7.592 $Y2=2.21
r78 41 93 7.0764 $w=2.83e-07 $l=1.75e-07 $layer=LI1_cond $X=7.592 $Y=1.87
+ $X2=7.592 $Y2=1.695
r79 40 93 3.20904 $w=2.85e-07 $l=1.25e-07 $layer=LI1_cond $X=7.592 $Y=1.57
+ $X2=7.592 $Y2=1.695
r80 40 89 3.64547 $w=2.5e-07 $l=1.42e-07 $layer=LI1_cond $X=7.592 $Y=1.57
+ $X2=7.45 $Y2=1.57
r81 39 89 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=7.13 $Y=1.57
+ $X2=7.45 $Y2=1.57
r82 39 90 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=7.13 $Y=1.57
+ $X2=6.78 $Y2=1.57
r83 38 85 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.695 $Y=1.57
+ $X2=6.61 $Y2=1.57
r84 38 90 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.695 $Y=1.57
+ $X2=6.78 $Y2=1.57
r85 38 85 0.59927 $w=2.48e-07 $l=1.3e-08 $layer=LI1_cond $X=6.597 $Y=1.57
+ $X2=6.61 $Y2=1.57
r86 37 106 0.368782 $w=2.48e-07 $l=8e-09 $layer=LI1_cond $X=6.21 $Y=1.57
+ $X2=6.202 $Y2=1.57
r87 37 106 2.52673 $w=1.85e-07 $l=1.25e-07 $layer=LI1_cond $X=6.202 $Y=1.445
+ $X2=6.202 $Y2=1.57
r88 37 38 10.1596 $w=4.18e-07 $l=3.02e-07 $layer=LI1_cond $X=6.295 $Y=1.57
+ $X2=6.597 $Y2=1.57
r89 36 37 10.9095 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=6.202 $Y=1.19
+ $X2=6.202 $Y2=1.445
r90 35 79 3.92452 $w=1.85e-07 $l=1.2e-07 $layer=LI1_cond $X=6.202 $Y=0.765
+ $X2=6.202 $Y2=0.885
r91 35 101 27.5336 $w=3.58e-07 $l=8.2e-07 $layer=LI1_cond $X=6.295 $Y=0.765
+ $X2=7.115 $Y2=0.765
r92 35 36 16.7862 $w=1.83e-07 $l=2.8e-07 $layer=LI1_cond $X=6.202 $Y=0.91
+ $X2=6.202 $Y2=1.19
r93 35 79 1.49877 $w=1.83e-07 $l=2.5e-08 $layer=LI1_cond $X=6.202 $Y=0.91
+ $X2=6.202 $Y2=0.885
r94 34 106 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=5.802 $Y=1.57
+ $X2=6.202 $Y2=1.57
r95 34 62 1.47513 $w=2.48e-07 $l=3.2e-08 $layer=LI1_cond $X=5.802 $Y=1.57
+ $X2=5.77 $Y2=1.57
r96 34 78 1.52122 $w=2.48e-07 $l=3.3e-08 $layer=LI1_cond $X=5.717 $Y=1.57
+ $X2=5.75 $Y2=1.57
r97 33 34 19.6837 $w=2.48e-07 $l=4.27e-07 $layer=LI1_cond $X=5.29 $Y=1.57
+ $X2=5.717 $Y2=1.57
r98 33 73 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.29 $Y=1.57
+ $X2=5.015 $Y2=1.57
r99 32 73 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=4.83 $Y=1.57
+ $X2=5.015 $Y2=1.57
r100 31 32 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.37 $Y=1.57
+ $X2=4.83 $Y2=1.57
r101 31 67 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=4.37 $Y=1.57
+ $X2=4.175 $Y2=1.57
r102 30 67 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=3.915 $Y=1.57
+ $X2=4.175 $Y2=1.57
r103 26 38 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.695 $Y=1.695
+ $X2=6.695 $Y2=1.57
r104 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.695 $Y=1.695
+ $X2=6.695 $Y2=1.95
r105 22 34 2.99516 $w=1.7e-07 $l=1.49164e-07 $layer=LI1_cond $X=5.855 $Y=1.695
+ $X2=5.802 $Y2=1.57
r106 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.855 $Y=1.695
+ $X2=5.855 $Y2=1.95
r107 7 40 300 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=2 $X=7.4
+ $Y=1.485 $X2=7.535 $Y2=1.69
r108 6 38 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=6.56
+ $Y=1.485 $X2=6.695 $Y2=1.61
r109 6 28 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=6.56
+ $Y=1.485 $X2=6.695 $Y2=1.95
r110 5 34 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.485 $X2=5.855 $Y2=1.61
r111 5 24 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.72
+ $Y=1.485 $X2=5.855 $Y2=1.95
r112 4 73 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.485 $X2=5.015 $Y2=1.61
r113 3 67 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.485 $X2=4.175 $Y2=1.61
r114 2 101 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=6.98
+ $Y=0.235 $X2=7.115 $Y2=0.76
r115 1 35 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=6.14
+ $Y=0.235 $X2=6.275 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%A_31_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 48 50 54 56 60 62 68 69 72 74 76 77 78 79 80
r141 72 82 3.04002 $w=2.85e-07 $l=1.1e-07 $layer=LI1_cond $X=7.592 $Y=0.475
+ $X2=7.592 $Y2=0.365
r142 72 74 9.90697 $w=2.83e-07 $l=2.45e-07 $layer=LI1_cond $X=7.592 $Y=0.475
+ $X2=7.592 $Y2=0.72
r143 69 71 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=5.94 $Y=0.365
+ $X2=6.695 $Y2=0.365
r144 68 82 3.92439 $w=2.2e-07 $l=1.42e-07 $layer=LI1_cond $X=7.45 $Y=0.365
+ $X2=7.592 $Y2=0.365
r145 68 71 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=7.45 $Y=0.365
+ $X2=6.695 $Y2=0.365
r146 65 67 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.855 $Y=0.715
+ $X2=5.855 $Y2=0.56
r147 64 69 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.855 $Y=0.475
+ $X2=5.94 $Y2=0.365
r148 64 67 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.855 $Y=0.475
+ $X2=5.855 $Y2=0.56
r149 63 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.8
+ $X2=4.895 $Y2=0.8
r150 62 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.77 $Y=0.8
+ $X2=5.855 $Y2=0.715
r151 62 63 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.77 $Y=0.8
+ $X2=4.98 $Y2=0.8
r152 58 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0.715
+ $X2=4.895 $Y2=0.8
r153 58 60 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.895 $Y=0.715
+ $X2=4.895 $Y2=0.56
r154 57 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=0.8
+ $X2=3.64 $Y2=0.8
r155 56 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=0.8
+ $X2=4.895 $Y2=0.8
r156 56 57 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.81 $Y=0.8
+ $X2=3.805 $Y2=0.8
r157 52 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.715
+ $X2=3.64 $Y2=0.8
r158 52 54 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.64 $Y=0.715
+ $X2=3.64 $Y2=0.36
r159 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.8
+ $X2=2.8 $Y2=0.8
r160 50 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=0.8
+ $X2=3.64 $Y2=0.8
r161 50 51 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.475 $Y=0.8
+ $X2=2.965 $Y2=0.8
r162 46 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.715 $X2=2.8
+ $Y2=0.8
r163 46 48 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.8 $Y=0.715
+ $X2=2.8 $Y2=0.36
r164 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0.8
+ $X2=1.96 $Y2=0.8
r165 44 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=0.8
+ $X2=2.8 $Y2=0.8
r166 44 45 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.635 $Y=0.8
+ $X2=2.125 $Y2=0.8
r167 40 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.715
+ $X2=1.96 $Y2=0.8
r168 40 42 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.96 $Y=0.715
+ $X2=1.96 $Y2=0.36
r169 39 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0.8
+ $X2=1.12 $Y2=0.8
r170 38 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0.8
+ $X2=1.96 $Y2=0.8
r171 38 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.795 $Y=0.8
+ $X2=1.285 $Y2=0.8
r172 34 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.715
+ $X2=1.12 $Y2=0.8
r173 34 36 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.12 $Y=0.715
+ $X2=1.12 $Y2=0.36
r174 32 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0.8
+ $X2=1.12 $Y2=0.8
r175 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.955 $Y=0.8
+ $X2=0.445 $Y2=0.8
r176 28 33 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.445 $Y2=0.8
r177 28 30 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.267 $Y2=0.38
r178 9 82 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.4
+ $Y=0.235 $X2=7.535 $Y2=0.38
r179 9 74 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=7.4
+ $Y=0.235 $X2=7.535 $Y2=0.72
r180 8 71 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.56
+ $Y=0.235 $X2=6.695 $Y2=0.36
r181 7 67 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=5.72
+ $Y=0.235 $X2=5.855 $Y2=0.56
r182 6 60 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.76
+ $Y=0.235 $X2=4.895 $Y2=0.56
r183 5 54 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.36
r184 4 48 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.36
r185 3 42 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.36
r186 2 36 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.36
r187 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_4%VGND 1 2 3 4 5 6 23 27 31 35 39 42 43 45 46
+ 48 49 50 66 76 77 80 85 88 90
r125 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r126 87 88 10.3517 $w=6.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0.23
+ $X2=4.64 $Y2=0.23
r127 83 87 1.99346 $w=6.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.37 $Y=0.23
+ $X2=4.475 $Y2=0.23
r128 83 85 14.3386 $w=6.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.37 $Y=0.23
+ $X2=3.995 $Y2=0.23
r129 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r130 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r131 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r132 74 77 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=7.59 $Y2=0
r133 74 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r134 73 76 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=7.59
+ $Y2=0
r135 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r136 71 90 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=5.6 $Y=0 $X2=5.375
+ $Y2=0
r137 71 73 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.6 $Y=0 $X2=5.75
+ $Y2=0
r138 70 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r139 70 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r140 69 88 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.64
+ $Y2=0
r141 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r142 66 90 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.375
+ $Y2=0
r143 66 69 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=4.83
+ $Y2=0
r144 65 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r145 64 85 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=0 $X2=3.995
+ $Y2=0
r146 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r147 61 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r148 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r149 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r150 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r151 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r152 55 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r153 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r154 52 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.7
+ $Y2=0
r155 52 54 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=0
+ $X2=1.15 $Y2=0
r156 50 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r157 48 60 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.135 $Y=0
+ $X2=2.99 $Y2=0
r158 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.22
+ $Y2=0
r159 47 64 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.305 $Y=0
+ $X2=3.91 $Y2=0
r160 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.22
+ $Y2=0
r161 45 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=0
+ $X2=2.07 $Y2=0
r162 45 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.38
+ $Y2=0
r163 44 60 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=2.99 $Y2=0
r164 44 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.38
+ $Y2=0
r165 42 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r166 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.54
+ $Y2=0
r167 41 57 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.625 $Y=0
+ $X2=2.07 $Y2=0
r168 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.54
+ $Y2=0
r169 37 90 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0
r170 37 39 7.30937 $w=4.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0.36
r171 33 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0
r172 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0.38
r173 29 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=0.085
+ $X2=2.38 $Y2=0
r174 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.38 $Y=0.085
+ $X2=2.38 $Y2=0.38
r175 25 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0
r176 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0.38
r177 21 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r178 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.38
r179 6 39 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.235 $X2=5.375 $Y2=0.36
r180 5 87 91 $w=1.7e-07 $l=6.09303e-07 $layer=licon1_NDIFF $count=2 $X=3.925
+ $Y=0.235 $X2=4.475 $Y2=0.36
r181 4 35 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.38
r182 3 31 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.38
r183 2 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.38
r184 1 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__or3b_1.spice
* Created: Tue Sep  1 19:28:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or3b_1.pex.spice"
.subckt sky130_fd_sc_hd__or3b_1  VNB VPB C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1009 N_A_109_93#_M1009_d N_C_N_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_109_93#_M1005_g N_A_215_53#_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_215_53#_M1004_d N_B_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_215_53#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.0567 PD=0.773271 PS=0.69 NRD=11.424 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_215_53#_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.121799 PD=1.85 PS=1.19673 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75001 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_109_93#_M1007_d N_C_N_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_297_297# N_A_109_93#_M1000_g N_A_215_53#_M1000_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 A_369_297# N_B_M1002_g A_297_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.06825
+ AS=0.0441 PD=0.745 PS=0.63 NRD=50.4123 NRS=23.443 M=1 R=2.8 SA=75000.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_369_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0876972 AS=0.06825 PD=0.792676 PS=0.745 NRD=72.1217 NRS=50.4123 M=1 R=2.8
+ SA=75001 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_215_53#_M1003_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.208803 PD=2.55 PS=1.88732 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_70 VPB 0 2.34755e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__or3b_1.pxi.spice"
*
.ends
*
*

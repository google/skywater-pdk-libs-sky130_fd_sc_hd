# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__clkdlybuf4s50_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.480000 1.285000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.390500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.185000 0.270000 3.625000 0.640000 ;
        RECT 3.185000 1.530000 3.625000 2.465000 ;
        RECT 3.345000 0.640000 3.625000 1.530000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.140000 0.085000 ;
        RECT 0.585000  0.085000 0.915000 0.565000 ;
        RECT 2.685000  0.085000 3.015000 0.565000 ;
        RECT 3.795000  0.085000 4.055000 0.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.140000 2.805000 ;
        RECT 0.600000 1.800000 0.930000 2.635000 ;
        RECT 2.685000 1.800000 3.015000 2.635000 ;
        RECT 3.795000 1.800000 4.055000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.270000 0.415000 0.735000 ;
      RECT 0.085000 0.735000 1.270000 0.905000 ;
      RECT 0.085000 1.455000 1.270000 1.630000 ;
      RECT 0.085000 1.630000 0.430000 2.465000 ;
      RECT 0.765000 1.075000 1.435000 1.245000 ;
      RECT 0.850000 0.905000 1.270000 1.075000 ;
      RECT 0.850000 1.245000 1.270000 1.455000 ;
      RECT 1.390000 1.785000 1.795000 2.465000 ;
      RECT 1.440000 0.270000 1.795000 0.900000 ;
      RECT 1.625000 0.900000 1.795000 1.075000 ;
      RECT 1.625000 1.075000 2.305000 1.245000 ;
      RECT 1.625000 1.245000 1.795000 1.785000 ;
      RECT 1.985000 0.270000 2.235000 0.735000 ;
      RECT 1.985000 0.735000 2.645000 0.905000 ;
      RECT 1.985000 1.460000 2.645000 1.630000 ;
      RECT 1.985000 1.630000 2.235000 2.465000 ;
      RECT 2.475000 0.905000 2.645000 0.995000 ;
      RECT 2.475000 0.995000 3.175000 1.325000 ;
      RECT 2.475000 1.325000 2.645000 1.460000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_2
END LIBRARY

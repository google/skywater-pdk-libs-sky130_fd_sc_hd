* NGSPICE file created from sky130_fd_sc_hd__einvp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
M1000 a_215_309# a_27_47# VPWR VPB phighvt w=940000u l=150000u
+  ad=1.3487e+12p pd=1.253e+07u as=7.676e+11p ps=7.36e+06u
M1001 VPWR a_27_47# a_215_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_215_309# a_27_47# VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND TE a_193_47# VNB nshort w=650000u l=150000u
+  ad=5.33e+11p pd=5.54e+06u as=8.905e+11p ps=9.24e+06u
M1004 Z A a_215_309# VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1005 a_215_309# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_47# a_215_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_193_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_215_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_193_47# TE VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND TE a_193_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR TE a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1012 a_215_309# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z A a_193_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=0p ps=0u
M1014 a_193_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND TE a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1016 Z A a_193_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_193_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__lpflow_inputiso1n_1.pex.spice
* Created: Thu Aug 27 14:25:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1%SLEEP_B 3 7 9 15 18
r26 12 15 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r27 9 18 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.2 $X2=0.23
+ $Y2=1.2
r28 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r29 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r30 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r31 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r32 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1%A_27_53# 1 2 9 13 17 19 20 23 27
+ 30 37
r48 36 37 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.37 $Y=1.16 $X2=1.43
+ $Y2=1.16
r49 28 36 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.22 $Y=1.16
+ $X2=1.37 $Y2=1.16
r50 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.16 $X2=1.22 $Y2=1.16
r51 25 33 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.16
+ $X2=0.72 $Y2=1.325
r52 25 30 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.72 $Y=1.16
+ $X2=0.72 $Y2=0.82
r53 25 27 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.845 $Y=1.16
+ $X2=1.22 $Y2=1.16
r54 23 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=1.62
+ $X2=0.68 $Y2=1.325
r55 19 30 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.72 $Y2=0.82
r56 19 20 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.42 $Y2=0.82
r57 15 20 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.42 $Y2=0.82
r58 15 17 10.7809 $w=3.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.265 $Y2=0.445
r59 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.43 $Y2=1.16
r60 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.43 $Y2=1.695
r61 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=0.995
+ $X2=1.37 $Y2=1.16
r62 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.37 $Y=0.995 $X2=1.37
+ $Y2=0.475
r63 2 23 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.62
r64 1 17 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1%A 1 5 8 9 15
r36 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=2.28
+ $X2=1.175 $Y2=2.28
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=2.28 $X2=1.01 $Y2=2.28
r38 9 13 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.155 $Y=2.25
+ $X2=1.01 $Y2=2.25
r39 5 8 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=1.79 $Y=0.475
+ $X2=1.79 $Y2=1.695
r40 3 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.79 $Y=2.265 $X2=1.79
+ $Y2=1.695
r41 1 3 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.715 $Y=2.34
+ $X2=1.79 $Y2=2.265
r42 1 15 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.715 $Y=2.34
+ $X2=1.175 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1%A_219_297# 1 2 9 12 14 18 20 21
+ 25 26 32 33 34 37
c58 25 0 1.06604e-19 $X=2.15 $Y=1.495
r59 33 38 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.16
+ $X2=2.215 $Y2=1.325
r60 33 37 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.16
+ $X2=2.215 $Y2=0.995
r61 32 35 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=1.16
+ $X2=2.18 $Y2=1.325
r62 32 34 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=1.16
+ $X2=2.18 $Y2=0.995
r63 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.16 $X2=2.21 $Y2=1.16
r64 26 29 2.88111 $w=4.18e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.58 $X2=1.2
+ $Y2=1.685
r65 25 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.15 $Y=1.495
+ $X2=2.15 $Y2=1.325
r66 22 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.15 $Y=0.825
+ $X2=2.15 $Y2=0.995
r67 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=0.74
+ $X2=2.15 $Y2=0.825
r68 20 21 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.065 $Y=0.74
+ $X2=1.665 $Y2=0.74
r69 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=0.655
+ $X2=1.665 $Y2=0.74
r70 16 18 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.58 $Y=0.655
+ $X2=1.58 $Y2=0.47
r71 15 26 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.41 $Y=1.58 $X2=1.2
+ $Y2=1.58
r72 14 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=1.58
+ $X2=2.15 $Y2=1.495
r73 14 15 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.065 $Y=1.58
+ $X2=1.41 $Y2=1.58
r74 12 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.28 $Y=1.985
+ $X2=2.28 $Y2=1.325
r75 9 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.28 $Y=0.56 $X2=2.28
+ $Y2=0.995
r76 2 29 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.485 $X2=1.22 $Y2=1.685
r77 1 18 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.265 $X2=1.58 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1%VPWR 1 2 7 9 13 15 17 27 28 34
c32 2 0 1.06604e-19 $X=1.865 $Y=1.485
r33 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r35 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 25 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.055 $Y2=2.72
r37 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 21 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r41 20 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 18 31 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r44 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 17 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.055 $Y2=2.72
r46 17 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.61 $Y2=2.72
r47 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 11 34 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2.72
r50 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2
r51 7 31 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r52 7 9 44.064 $w=2.53e-07 $l=9.75e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=1.66
r53 2 13 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.485 $X2=2.065 $Y2=2
r54 1 9 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1%X 1 2 12 14 15 16
r16 14 16 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.54 $Y=1.63
+ $X2=2.54 $Y2=1.845
r17 14 15 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.54 $Y=1.63
+ $X2=2.54 $Y2=1.495
r18 10 12 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=2.49 $Y=0.587 $X2=2.59
+ $Y2=0.587
r19 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.59 $Y=0.76 $X2=2.59
+ $Y2=0.587
r20 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.59 $Y=0.76
+ $X2=2.59 $Y2=1.495
r21 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=1.485 $X2=2.49 $Y2=1.845
r22 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.49 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1N_1%VGND 1 2 9 11 18 25 26 31 37 39
r41 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r42 36 37 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=0.24
+ $X2=1.325 $Y2=0.24
r43 33 36 0.184012 $w=6.48e-07 $l=1e-08 $layer=LI1_cond $X=1.15 $Y=0.24 $X2=1.16
+ $Y2=0.24
r44 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r45 30 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r46 29 33 8.46455 $w=6.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.24
+ $X2=1.15 $Y2=0.24
r47 29 31 9.28585 $w=6.48e-07 $l=1e-07 $layer=LI1_cond $X=0.69 $Y=0.24 $X2=0.59
+ $Y2=0.24
r48 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r49 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r50 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r51 23 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.025
+ $Y2=0
r52 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.53
+ $Y2=0
r53 22 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r54 22 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r55 21 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.325
+ $Y2=0
r56 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r57 18 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.025
+ $Y2=0
r58 18 21 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.61
+ $Y2=0
r59 15 31 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.59
+ $Y2=0
r60 11 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r61 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r62 7 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r63 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.4
r64 2 9 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.265 $X2=2.05 $Y2=0.4
r65 1 36 91 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.265 $X2=1.16 $Y2=0.4
.ends


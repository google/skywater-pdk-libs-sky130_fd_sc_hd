* File: sky130_fd_sc_hd__o32ai_2.pex.spice
* Created: Thu Aug 27 14:41:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O32AI_2%B2 1 3 6 8 10 13 15 16 24
c38 16 0 1.81089e-19 $X=0.695 $Y=1.19
r39 22 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.68 $Y=1.16
+ $X2=0.89 $Y2=1.16
r40 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.68 $Y2=1.16
r41 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=1.16 $X2=0.68 $Y2=1.16
r42 15 16 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.235 $Y=1.2
+ $X2=0.68 $Y2=1.2
r43 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r44 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r45 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r46 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r47 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r49 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%B1 1 3 6 8 10 13 15 16 24
c48 24 0 1.81089e-19 $X=1.73 $Y=1.16
c49 16 0 1.25815e-19 $X=1.615 $Y=1.19
r50 22 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.73 $Y2=1.16
r51 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r52 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r53 16 23 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.2
+ $X2=1.52 $Y2=1.2
r54 15 23 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.2
+ $X2=1.52 $Y2=1.2
r55 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r56 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r57 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r58 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r59 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r60 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r61 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%A3 3 6 9 11 13 16 18 21 24 26
c54 26 0 8.05404e-21 $X=3.15 $Y=1.16
c55 6 0 1.02109e-19 $X=2.225 $Y=1.19
c56 3 0 1.25815e-19 $X=2.15 $Y=0.56
r57 25 26 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.09 $Y=1.16 $X2=3.15
+ $Y2=1.16
r58 23 25 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.9 $Y=1.16 $X2=3.09
+ $Y2=1.16
r59 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.9
+ $Y=1.16 $X2=2.9 $Y2=1.16
r60 20 23 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.73 $Y=1.16 $X2=2.9
+ $Y2=1.16
r61 20 21 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.73 $Y=1.16
+ $X2=2.655 $Y2=1.16
r62 18 24 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.535 $Y=1.2
+ $X2=2.9 $Y2=1.2
r63 14 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.16
r64 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.985
r65 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=1.16
r66 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=0.56
r67 7 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.16
r68 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.73 $Y=1.325 $X2=2.73
+ $Y2=1.985
r69 6 21 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.225 $Y=1.19
+ $X2=2.655 $Y2=1.19
r70 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.15 $Y=1.115
+ $X2=2.225 $Y2=1.19
r71 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.15 $Y=1.115
+ $X2=2.15 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%A2 1 3 6 8 10 13 15 16 26
r46 25 26 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.93 $Y=1.16 $X2=3.99
+ $Y2=1.16
r47 23 25 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.74 $Y=1.16
+ $X2=3.93 $Y2=1.16
r48 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.16 $X2=3.74 $Y2=1.16
r49 21 23 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=3.57 $Y=1.16
+ $X2=3.74 $Y2=1.16
r50 19 21 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.51 $Y=1.16 $X2=3.57
+ $Y2=1.16
r51 16 24 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.375 $Y=1.2
+ $X2=3.74 $Y2=1.2
r52 15 24 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=3.455 $Y=1.2
+ $X2=3.74 $Y2=1.2
r53 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.16
r54 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.985
r55 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.16
r56 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=0.56
r57 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=1.16
r58 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.57 $Y=1.325 $X2=3.57
+ $Y2=1.985
r59 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.16
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995 $X2=3.51
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%A1 1 3 6 8 10 13 15 16 17 28
r39 27 28 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.29 $Y=1.16 $X2=5.37
+ $Y2=1.16
r40 25 27 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=5.09 $Y=1.16 $X2=5.29
+ $Y2=1.16
r41 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.09
+ $Y=1.16 $X2=5.09 $Y2=1.16
r42 23 25 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.95 $Y=1.16
+ $X2=5.09 $Y2=1.16
r43 21 23 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=4.87 $Y=1.16 $X2=4.95
+ $Y2=1.16
r44 16 17 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=5.295 $Y=1.2
+ $X2=5.755 $Y2=1.2
r45 16 26 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=5.295 $Y=1.2
+ $X2=5.09 $Y2=1.2
r46 15 26 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.835 $Y=1.2
+ $X2=5.09 $Y2=1.2
r47 11 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.37 $Y=1.325
+ $X2=5.37 $Y2=1.16
r48 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.37 $Y=1.325
+ $X2=5.37 $Y2=1.985
r49 8 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.29 $Y=0.995
+ $X2=5.29 $Y2=1.16
r50 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.29 $Y=0.995
+ $X2=5.29 $Y2=0.56
r51 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.95 $Y=1.325
+ $X2=4.95 $Y2=1.16
r52 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.95 $Y=1.325 $X2=4.95
+ $Y2=1.985
r53 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.87 $Y=0.995
+ $X2=4.87 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.87 $Y=0.995 $X2=4.87
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%A_27_297# 1 2 3 10 12 14 16 17 18 27
c40 27 0 1.02109e-19 $X=1.94 $Y=2
c41 3 0 1.4598e-19 $X=1.805 $Y=1.485
r42 19 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=1.92
+ $X2=1.14 $Y2=1.92
r43 18 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=1.92
+ $X2=1.94 $Y2=1.92
r44 18 19 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=1.92
+ $X2=1.265 $Y2=1.92
r45 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.005
+ $X2=1.14 $Y2=1.92
r46 16 17 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.14 $Y=2.005
+ $X2=1.14 $Y2=2.295
r47 15 23 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=2.38
+ $X2=0.217 $Y2=2.38
r48 14 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.015 $Y=2.38
+ $X2=1.14 $Y2=2.295
r49 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=2.38
+ $X2=0.345 $Y2=2.38
r50 10 23 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=2.295
+ $X2=0.217 $Y2=2.38
r51 10 12 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.217 $Y=2.295
+ $X2=0.217 $Y2=1.66
r52 3 27 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r53 2 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r54 1 23 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r55 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%Y 1 2 3 4 13 21 23 28 31 32 33 48
c71 32 0 1.54034e-19 $X=1.99 $Y=1.105
r72 39 48 2.42208 $w=2.93e-07 $l=6.2e-08 $layer=LI1_cond $X=2.022 $Y=1.252
+ $X2=2.022 $Y2=1.19
r73 33 40 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.022 $Y=1.58
+ $X2=2.022 $Y2=1.495
r74 33 40 0.976647 $w=2.93e-07 $l=2.5e-08 $layer=LI1_cond $X=2.022 $Y=1.47
+ $X2=2.022 $Y2=1.495
r75 32 48 0.46879 $w=2.93e-07 $l=1.2e-08 $layer=LI1_cond $X=2.022 $Y=1.178
+ $X2=2.022 $Y2=1.19
r76 32 33 8.08663 $w=2.93e-07 $l=2.07e-07 $layer=LI1_cond $X=2.022 $Y=1.263
+ $X2=2.022 $Y2=1.47
r77 32 39 0.429725 $w=2.93e-07 $l=1.1e-08 $layer=LI1_cond $X=2.022 $Y=1.263
+ $X2=2.022 $Y2=1.252
r78 29 32 10.9595 $w=2.23e-07 $l=2e-07 $layer=LI1_cond $X=1.96 $Y=0.905 $X2=1.96
+ $Y2=1.105
r79 24 33 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.17 $Y=1.58
+ $X2=2.022 $Y2=1.58
r80 23 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.94 $Y2=1.58
r81 23 24 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.17 $Y2=1.58
r82 22 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.58
+ $X2=0.68 $Y2=1.58
r83 21 33 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.875 $Y=1.58
+ $X2=2.022 $Y2=1.58
r84 21 22 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=1.875 $Y=1.58
+ $X2=0.845 $Y2=1.58
r85 15 18 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=0.68 $Y=0.78
+ $X2=1.52 $Y2=0.78
r86 13 29 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.875 $Y=0.78
+ $X2=1.96 $Y2=0.905
r87 13 18 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=1.875 $Y=0.78
+ $X2=1.52 $Y2=0.78
r88 4 31 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=2.94 $Y2=1.66
r89 3 28 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r90 2 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.74
r91 1 15 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%VPWR 1 2 3 12 16 18 20 25 26 28 29 30 45 51
r75 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r76 48 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r77 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r78 45 50 3.67125 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.737 $Y2=2.72
r79 45 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.29 $Y2=2.72
r80 44 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r81 43 44 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r82 41 44 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=4.37 $Y2=2.72
r83 40 43 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=4.37 $Y2=2.72
r84 40 41 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r85 38 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r86 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 33 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 30 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 30 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r90 28 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.37 $Y2=2.72
r91 28 29 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.722 $Y2=2.72
r92 27 47 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=5.29 $Y2=2.72
r93 27 29 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.722 $Y2=2.72
r94 25 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r95 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.52 $Y2=2.72
r96 24 40 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.61 $Y2=2.72
r97 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.52 $Y2=2.72
r98 20 23 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=5.605 $Y=1.66
+ $X2=5.605 $Y2=2.34
r99 18 50 3.29199 $w=2.2e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.605 $Y=2.635
+ $X2=5.737 $Y2=2.72
r100 18 23 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=5.605 $Y=2.635
+ $X2=5.605 $Y2=2.34
r101 14 29 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.722 $Y=2.635
+ $X2=4.722 $Y2=2.72
r102 14 16 34.3548 $w=2.03e-07 $l=6.35e-07 $layer=LI1_cond $X=4.722 $Y=2.635
+ $X2=4.722 $Y2=2
r103 10 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r104 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.34
r105 3 23 400 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=1.485 $X2=5.6 $Y2=2.34
r106 3 20 400 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=1.485 $X2=5.6 $Y2=1.66
r107 2 16 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=4.615
+ $Y=1.485 $X2=4.74 $Y2=2
r108 1 12 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%A_475_297# 1 2 3 10 12 14 18 20 22 24 29
r40 22 31 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.26 $Y=2.255
+ $X2=4.26 $Y2=2.35
r41 22 24 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.26 $Y=2.255
+ $X2=4.26 $Y2=2
r42 21 29 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=2.35
+ $X2=3.36 $Y2=2.35
r43 20 31 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.135 $Y=2.35
+ $X2=4.26 $Y2=2.35
r44 20 21 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=4.135 $Y=2.35
+ $X2=3.445 $Y2=2.35
r45 16 29 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.36 $Y=2.255
+ $X2=3.36 $Y2=2.35
r46 16 18 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.36 $Y=2.255
+ $X2=3.36 $Y2=1.66
r47 15 27 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=2.585 $Y=2.35
+ $X2=2.46 $Y2=2.35
r48 14 29 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=2.35
+ $X2=3.36 $Y2=2.35
r49 14 15 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=3.275 $Y=2.35
+ $X2=2.585 $Y2=2.35
r50 10 27 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=2.46 $Y=2.255
+ $X2=2.46 $Y2=2.35
r51 10 12 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.46 $Y=2.255
+ $X2=2.46 $Y2=2
r52 3 31 600 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.485 $X2=4.22 $Y2=2.34
r53 3 24 600 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.485 $X2=4.22 $Y2=2
r54 2 29 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=2.34
r55 2 18 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=1.66
r56 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.485 $X2=2.5 $Y2=2.34
r57 1 12 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.485 $X2=2.5 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%A_729_297# 1 2 9 11 13 16
r29 11 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=1.665 $X2=5.16
+ $Y2=1.58
r30 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.16 $Y=1.665
+ $X2=5.16 $Y2=2.34
r31 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=1.58
+ $X2=3.78 $Y2=1.58
r32 9 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=1.58
+ $X2=5.16 $Y2=1.58
r33 9 10 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=4.995 $Y=1.58
+ $X2=3.945 $Y2=1.58
r34 2 18 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.025
+ $Y=1.485 $X2=5.16 $Y2=1.66
r35 2 13 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.025
+ $Y=1.485 $X2=5.16 $Y2=2.34
r36 1 16 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=3.645
+ $Y=1.485 $X2=3.78 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%A_27_47# 1 2 3 4 5 6 19 21 23 30 31 32 35 39
+ 43 47 50 51
r92 49 51 9.67895 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.56 $Y=0.58
+ $X2=4.725 $Y2=0.58
r93 49 50 15.9354 $w=6.48e-07 $l=5.05e-07 $layer=LI1_cond $X=4.56 $Y=0.58
+ $X2=4.055 $Y2=0.58
r94 41 43 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.59 $Y=0.715
+ $X2=5.59 $Y2=0.38
r95 39 41 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=5.425 $Y=0.81
+ $X2=5.59 $Y2=0.715
r96 39 51 40.8612 $w=1.88e-07 $l=7e-07 $layer=LI1_cond $X=5.425 $Y=0.81
+ $X2=4.725 $Y2=0.81
r97 38 47 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=0.81
+ $X2=3.3 $Y2=0.81
r98 38 50 34.4402 $w=1.88e-07 $l=5.9e-07 $layer=LI1_cond $X=3.465 $Y=0.81
+ $X2=4.055 $Y2=0.81
r99 33 47 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.3 $Y=0.715 $X2=3.3
+ $Y2=0.81
r100 33 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.3 $Y=0.715
+ $X2=3.3 $Y2=0.38
r101 31 47 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0.81
+ $X2=3.3 $Y2=0.81
r102 31 32 42.6124 $w=1.88e-07 $l=7.3e-07 $layer=LI1_cond $X=3.135 $Y=0.81
+ $X2=2.405 $Y2=0.81
r103 30 32 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.32 $Y=0.715
+ $X2=2.405 $Y2=0.81
r104 29 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.32 $Y=0.485
+ $X2=2.32 $Y2=0.715
r105 26 28 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=0.37
+ $X2=1.94 $Y2=0.37
r106 24 46 3.603 $w=2.3e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.37
+ $X2=0.217 $Y2=0.37
r107 24 26 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.345 $Y=0.37
+ $X2=1.1 $Y2=0.37
r108 23 29 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.235 $Y=0.37
+ $X2=2.32 $Y2=0.485
r109 23 28 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.235 $Y=0.37
+ $X2=1.94 $Y2=0.37
r110 19 46 3.23707 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=0.217 $Y=0.485
+ $X2=0.217 $Y2=0.37
r111 19 21 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.217 $Y=0.485
+ $X2=0.217 $Y2=0.74
r112 6 43 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=5.365
+ $Y=0.235 $X2=5.59 $Y2=0.38
r113 5 49 45.5 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_NDIFF $count=4 $X=4.005
+ $Y=0.235 $X2=4.56 $Y2=0.38
r114 4 35 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.38
r115 3 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r116 2 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r117 1 46 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r118 1 21 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__O32AI_2%VGND 1 2 3 12 16 20 23 24 26 27 29 30 31 50
+ 51
r78 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r79 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r80 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r81 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r82 44 47 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r83 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r84 42 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r85 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r86 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r87 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r88 34 38 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r89 31 39 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r90 31 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r91 29 47 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.905 $Y=0 $X2=4.83
+ $Y2=0
r92 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=0 $X2=5.07
+ $Y2=0
r93 28 50 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.75
+ $Y2=0
r94 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.07
+ $Y2=0
r95 26 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.45
+ $Y2=0
r96 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.72
+ $Y2=0
r97 25 44 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.91
+ $Y2=0
r98 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.72
+ $Y2=0
r99 23 38 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.62 $Y=0 $X2=2.53
+ $Y2=0
r100 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=0 $X2=2.785
+ $Y2=0
r101 22 41 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.95 $Y=0 $X2=3.45
+ $Y2=0
r102 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=0 $X2=2.785
+ $Y2=0
r103 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=0.085
+ $X2=5.07 $Y2=0
r104 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.07 $Y=0.085
+ $X2=5.07 $Y2=0.38
r105 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r106 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.38
r107 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=0.085
+ $X2=2.785 $Y2=0
r108 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.785 $Y=0.085
+ $X2=2.785 $Y2=0.38
r109 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.945
+ $Y=0.235 $X2=5.08 $Y2=0.38
r110 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.38
r111 1 12 182 $w=1.7e-07 $l=6.28331e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.785 $Y2=0.38
.ends


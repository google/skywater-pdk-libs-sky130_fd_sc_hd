* File: sky130_fd_sc_hd__or4b_4.spice
* Created: Tue Sep  1 19:28:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or4b_4.pex.spice"
.subckt sky130_fd_sc_hd__or4b_4  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1017 N_A_109_93#_M1017_d N_D_N_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.10785 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_215_297#_M1003_d N_A_109_93#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1235 AS=0.16535 PD=1.03 PS=1.82 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_215_297#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=0 NRS=4.608 M=1 R=4.33333 SA=75000.7
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1006 N_A_215_297#_M1006_d N_B_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_215_297#_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.08775 PD=1.03 PS=0.92 NRD=17.532 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1004_d N_A_215_297#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.08775 PD=1.03 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_215_297#_M1008_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1008_d N_A_215_297#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_215_297#_M1011_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.08775 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_109_93#_M1010_d N_D_N_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_297_297# N_A_109_93#_M1002_g N_A_215_297#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.19 AS=0.26 PD=1.38 PS=2.52 NRD=26.5753 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.3 A=0.15 P=2.3 MULT=1
MM1014 A_403_297# N_C_M1014_g A_297_297# VPB PHIGHVT L=0.15 W=1 AD=0.135 AS=0.19
+ PD=1.27 PS=1.38 NRD=15.7403 NRS=26.5753 M=1 R=6.66667 SA=75000.7 SB=75002.8
+ A=0.15 P=2.3 MULT=1
MM1012 A_487_297# N_B_M1012_g A_403_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_487_297# VPB PHIGHVT L=0.15 W=1 AD=0.19
+ AS=0.135 PD=1.38 PS=1.27 NRD=9.8303 NRS=15.7403 M=1 R=6.66667 SA=75001.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1005_d N_A_215_297#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.19 AS=0.135 PD=1.38 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75002.1
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_215_297#_M1013_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1013_d N_A_215_297#_M1015_g N_X_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_A_215_297#_M1016_g N_X_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=8.7312 P=14.09
*
.include "sky130_fd_sc_hd__or4b_4.pxi.spice"
*
.ends
*
*

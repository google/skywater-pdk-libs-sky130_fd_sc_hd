* File: sky130_fd_sc_hd__o2bb2a_4.pex.spice
* Created: Tue Sep  1 19:23:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%B1 3 6 8 10 13 15 19 20 22 25 26 27
c80 26 0 1.22288e-19 $X=0.41 $Y=1.16
c81 19 0 1.20505e-19 $X=1.73 $Y=1.16
c82 8 0 1.14637e-19 $X=1.73 $Y=0.995
r83 25 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=1.325
r84 25 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=0.995
r85 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r86 22 34 8.29932 $w=4.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.33 $Y=1.19
+ $X2=0.33 $Y2=1.53
r87 22 26 0.732293 $w=4.88e-07 $l=3e-08 $layer=LI1_cond $X=0.33 $Y=1.19 $X2=0.33
+ $Y2=1.16
r88 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r89 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.73 $Y=1.445
+ $X2=1.73 $Y2=1.16
r90 16 34 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.575 $Y=1.53
+ $X2=0.33 $Y2=1.53
r91 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.53
+ $X2=1.73 $Y2=1.445
r92 15 16 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.565 $Y=1.53
+ $X2=0.575 $Y2=1.53
r93 11 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r94 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r95 8 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r96 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r97 6 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r98 3 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%B2 1 3 6 8 10 13 15 22
c48 6 0 1.22288e-19 $X=0.89 $Y=1.985
r49 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.31
+ $Y2=1.16
r50 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.89 $Y=1.16 $X2=1.1
+ $Y2=1.16
r51 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%A_415_21# 1 2 3 10 12 15 17 19 22 24 27 30
+ 32 34 35 36 37 41 42 48 49 52
c122 52 0 1.27834e-19 $X=4.56 $Y=1.96
c123 48 0 1.20878e-19 $X=4.14 $Y=0.73
c124 42 0 1.20678e-19 $X=3.72 $Y=1.875
c125 27 0 1.82667e-19 $X=2.78 $Y=1.16
c126 10 0 1.56657e-19 $X=2.15 $Y=0.995
r127 53 55 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r128 48 49 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0.775
+ $X2=3.975 $Y2=0.775
r129 42 45 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.875
+ $X2=3.72 $Y2=1.96
r130 38 42 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1.875
+ $X2=3.72 $Y2=1.875
r131 37 52 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=1.875
+ $X2=4.56 $Y2=1.875
r132 37 38 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=4.435 $Y=1.875
+ $X2=3.845 $Y2=1.875
r133 35 42 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.595 $Y=1.875
+ $X2=3.72 $Y2=1.875
r134 35 36 27.7273 $w=1.78e-07 $l=4.5e-07 $layer=LI1_cond $X=3.595 $Y=1.875
+ $X2=3.145 $Y2=1.875
r135 34 49 51.1414 $w=1.78e-07 $l=8.3e-07 $layer=LI1_cond $X=3.145 $Y=0.815
+ $X2=3.975 $Y2=0.815
r136 32 36 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.05 $Y=1.785
+ $X2=3.145 $Y2=1.875
r137 31 41 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=1.245
+ $X2=3.05 $Y2=1.16
r138 31 32 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=3.05 $Y=1.245
+ $X2=3.05 $Y2=1.785
r139 30 41 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=1.075
+ $X2=3.05 $Y2=1.16
r140 29 34 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.05 $Y=0.905
+ $X2=3.145 $Y2=0.815
r141 29 30 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.05 $Y=0.905
+ $X2=3.05 $Y2=1.075
r142 27 55 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.78 $Y=1.16
+ $X2=2.57 $Y2=1.16
r143 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.16 $X2=2.78 $Y2=1.16
r144 24 41 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.955 $Y=1.16
+ $X2=3.05 $Y2=1.16
r145 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.955 $Y=1.16
+ $X2=2.78 $Y2=1.16
r146 20 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r147 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r148 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r149 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r150 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r151 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r152 10 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r153 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
r154 3 52 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.96
r155 2 45 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=1.96
r156 1 48 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%A1_N 3 6 8 10 13 17 18 20 21 23 26 29
c90 29 0 5.08858e-19 $X=4.77 $Y=1.16
c91 18 0 1.20678e-19 $X=3.48 $Y=1.16
c92 17 0 1.82667e-19 $X=3.48 $Y=1.16
c93 13 0 1.48522e-19 $X=4.77 $Y=1.985
c94 8 0 2.18852e-19 $X=4.77 $Y=0.995
r95 23 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.16 $X2=4.77 $Y2=1.16
r96 22 23 9.12351 $w=3.58e-07 $l=2.85e-07 $layer=LI1_cond $X=4.785 $Y=1.445
+ $X2=4.785 $Y2=1.16
r97 20 22 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=4.605 $Y=1.53
+ $X2=4.785 $Y2=1.445
r98 20 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.605 $Y=1.53
+ $X2=3.645 $Y2=1.53
r99 18 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=3.48 $Y2=1.325
r100 18 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=3.48 $Y2=0.995
r101 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.48
+ $Y=1.16 $X2=3.48 $Y2=1.16
r102 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.48 $Y=1.445
+ $X2=3.645 $Y2=1.53
r103 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.48 $Y=1.445
+ $X2=3.48 $Y2=1.16
r104 11 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.16
r105 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.985
r106 8 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.16
r107 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r108 6 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.51 $Y=1.985
+ $X2=3.51 $Y2=1.325
r109 3 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.56
+ $X2=3.51 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%A2_N 1 3 6 8 10 13 15 21 22
c45 8 0 6.86556e-20 $X=4.35 $Y=0.995
r46 20 22 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.145 $Y=1.16
+ $X2=4.35 $Y2=1.16
r47 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=1.16 $X2=4.145 $Y2=1.16
r48 17 20 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.145 $Y2=1.16
r49 15 21 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=3.93 $Y=1.175
+ $X2=4.145 $Y2=1.175
r50 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.985
r52 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
r54 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=1.325
+ $X2=3.93 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.93 $Y=1.325 $X2=3.93
+ $Y2=1.985
r56 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995 $X2=3.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%A_193_297# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 38 41 44 49 52 58 62 63 69 70 78 86
c157 70 0 8.263e-20 $X=5.31 $Y=1.53
c158 69 0 1.48522e-19 $X=5.31 $Y=1.53
c159 63 0 1.20505e-19 $X=2.675 $Y=1.53
c160 58 0 8.53932e-20 $X=2.36 $Y=0.73
c161 44 0 1.74908e-19 $X=5.455 $Y=1.16
r162 84 86 2.27329 $w=4.83e-07 $l=9e-08 $layer=LI1_cond $X=2.34 $Y=1.87 $X2=2.34
+ $Y2=1.96
r163 75 76 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=6.03 $Y2=1.16
r164 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.31 $Y=1.53
+ $X2=5.31 $Y2=1.53
r165 66 84 8.58799 $w=4.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.34 $Y=1.53
+ $X2=2.34 $Y2=1.87
r166 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.53
+ $X2=2.53 $Y2=1.53
r167 63 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.53
+ $X2=2.53 $Y2=1.53
r168 62 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.165 $Y=1.53
+ $X2=5.31 $Y2=1.53
r169 62 63 3.08168 $w=1.4e-07 $l=2.49e-06 $layer=MET1_cond $X=5.165 $Y=1.53
+ $X2=2.675 $Y2=1.53
r170 61 70 11.3257 $w=2.88e-07 $l=2.85e-07 $layer=LI1_cond $X=5.31 $Y=1.245
+ $X2=5.31 $Y2=1.53
r171 58 60 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.73
+ $X2=2.36 $Y2=0.815
r172 52 55 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.1 $Y=1.87 $X2=1.1
+ $Y2=1.96
r173 50 78 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=6.21 $Y=1.16
+ $X2=6.45 $Y2=1.16
r174 50 76 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.21 $Y=1.16
+ $X2=6.03 $Y2=1.16
r175 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.21
+ $Y=1.16 $X2=6.21 $Y2=1.16
r176 47 75 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.53 $Y=1.16 $X2=5.61
+ $Y2=1.16
r177 47 72 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.53 $Y=1.16
+ $X2=5.19 $Y2=1.16
r178 46 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.53 $Y=1.16
+ $X2=6.21 $Y2=1.16
r179 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.16 $X2=5.53 $Y2=1.16
r180 44 61 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=5.455 $Y=1.16
+ $X2=5.31 $Y2=1.245
r181 44 46 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.455 $Y=1.16
+ $X2=5.53 $Y2=1.16
r182 41 66 14.3211 $w=4.83e-07 $l=4.64892e-07 $layer=LI1_cond $X=2.32 $Y=1.075
+ $X2=2.34 $Y2=1.53
r183 41 60 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.32 $Y=1.075
+ $X2=2.32 $Y2=0.815
r184 39 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=1.87
+ $X2=1.1 $Y2=1.87
r185 38 84 6.94006 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.065 $Y=1.87
+ $X2=2.34 $Y2=1.87
r186 38 39 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.065 $Y=1.87
+ $X2=1.225 $Y2=1.87
r187 34 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r188 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r189 31 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r190 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r191 27 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r192 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.985
r193 24 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r194 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=0.56
r195 20 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.16
r196 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.985
r197 17 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.16
r198 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r199 13 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.16
r200 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.985
r201 10 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.16
r202 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r203 3 86 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.96
r204 3 66 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.62
r205 2 55 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r206 1 58 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 38 42 46
+ 49 50 52 53 54 55 56 76 83 84 92 95 97 100
c120 36 0 1.23485e-19 $X=4.98 $Y=1.96
r121 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r122 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r123 94 95 9.89763 $w=6.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.3 $Y=2.47
+ $X2=3.425 $Y2=2.47
r124 90 94 5.53409 $w=6.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.99 $Y=2.47
+ $X2=3.3 $Y2=2.47
r125 90 92 12.9325 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=2.47
+ $X2=2.695 $Y2=2.47
r126 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r127 84 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r128 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r129 81 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=2.72
+ $X2=6.66 $Y2=2.72
r130 81 83 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.785 $Y=2.72
+ $X2=7.13 $Y2=2.72
r131 80 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r132 80 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r133 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r134 77 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=5.82 $Y2=2.72
r135 77 79 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=6.21 $Y2=2.72
r136 76 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.66 $Y2=2.72
r137 76 79 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.21 $Y2=2.72
r138 75 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r139 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r140 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r141 72 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r142 71 95 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=3.425 $Y2=2.72
r143 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r144 68 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r145 67 92 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.695 $Y2=2.72
r146 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r147 64 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r148 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r149 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r150 60 63 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r151 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r152 58 87 3.63617 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r153 58 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 56 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r155 56 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r156 54 74 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=4.83 $Y2=2.72
r157 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=4.98 $Y2=2.72
r158 52 71 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.91 $Y2=2.72
r159 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.14 $Y2=2.72
r160 51 74 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.265 $Y=2.72
+ $X2=4.83 $Y2=2.72
r161 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.265 $Y=2.72
+ $X2=4.14 $Y2=2.72
r162 49 63 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.61 $Y2=2.72
r163 49 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.94 $Y2=2.72
r164 48 67 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.53 $Y2=2.72
r165 48 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=1.94 $Y2=2.72
r166 44 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=2.72
r167 44 46 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=1.99
r168 40 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.72
r169 40 42 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.33
r170 39 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=4.98 $Y2=2.72
r171 38 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.82 $Y2=2.72
r172 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.105 $Y2=2.72
r173 34 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r174 34 36 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=1.96
r175 30 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.72
r176 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.3
r177 26 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r178 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.3
r179 22 87 3.25784 $w=2.05e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.172 $Y2=2.72
r180 22 24 36.5188 $w=2.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=1.96
r181 7 46 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=1.99
r182 6 42 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2.33
r183 5 36 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=1.96
r184 4 32 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2.3
r185 3 94 300 $w=1.7e-07 $l=1.09455e-06 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=3.3 $Y2=2.3
r186 2 28 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.3
r187 1 24 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%A_109_297# 1 2 9 11 12 14
r18 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.52 $Y=2.3 $X2=1.52
+ $Y2=2.38
r19 11 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.395 $Y=2.38
+ $X2=1.52 $Y2=2.38
r20 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.395 $Y=2.38
+ $X2=0.805 $Y2=2.38
r21 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.68 $Y=2.295
+ $X2=0.805 $Y2=2.38
r22 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=2.295
+ $X2=0.68 $Y2=1.96
r23 2 14 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.3
r24 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35 37
+ 38
c74 24 0 9.79736e-20 $X=5.565 $Y=0.815
r75 41 47 1.28267 $w=3.05e-07 $l=2.4e-07 $layer=LI1_cond $X=6.757 $Y=1.415
+ $X2=6.757 $Y2=1.655
r76 38 47 2.44731 $w=3.34e-07 $l=6.7e-08 $layer=LI1_cond $X=6.69 $Y=1.655
+ $X2=6.757 $Y2=1.655
r77 38 44 16.4371 $w=3.34e-07 $l=4.5e-07 $layer=LI1_cond $X=6.69 $Y=1.655
+ $X2=6.24 $Y2=1.655
r78 37 41 8.50163 $w=3.03e-07 $l=2.25e-07 $layer=LI1_cond $X=6.757 $Y=1.19
+ $X2=6.757 $Y2=1.415
r79 36 37 10.7687 $w=3.03e-07 $l=2.85e-07 $layer=LI1_cond $X=6.757 $Y=0.905
+ $X2=6.757 $Y2=1.19
r80 34 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=0.815
+ $X2=6.24 $Y2=0.815
r81 33 36 7.42255 $w=1.8e-07 $l=1.91792e-07 $layer=LI1_cond $X=6.605 $Y=0.815
+ $X2=6.757 $Y2=0.905
r82 33 34 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=6.605 $Y=0.815
+ $X2=6.405 $Y2=0.815
r83 29 44 2.43566 $w=2.5e-07 $l=3e-07 $layer=LI1_cond $X=6.24 $Y=1.955 $X2=6.24
+ $Y2=1.655
r84 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.24 $Y=1.955
+ $X2=6.24 $Y2=1.96
r85 25 35 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.24 $Y=0.725 $X2=6.24
+ $Y2=0.815
r86 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.24 $Y=0.725
+ $X2=6.24 $Y2=0.39
r87 23 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=6.24 $Y2=0.815
r88 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=5.565 $Y2=0.815
r89 21 44 7.50035 $w=3.34e-07 $l=2.7037e-07 $layer=LI1_cond $X=6.115 $Y=1.87
+ $X2=6.24 $Y2=1.655
r90 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.115 $Y=1.87
+ $X2=5.525 $Y2=1.87
r91 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.4 $Y=1.955
+ $X2=5.525 $Y2=1.87
r92 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.4 $Y=1.955 $X2=5.4
+ $Y2=1.96
r93 13 24 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.4 $Y=0.725
+ $X2=5.565 $Y2=0.815
r94 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.4 $Y=0.725 $X2=5.4
+ $Y2=0.39
r95 4 44 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.62
r96 4 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.96
r97 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.96
r98 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.39
r99 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%A_27_47# 1 2 3 4 15 17 18 21 23 25 28 31 33
c64 33 0 2.9244e-20 $X=1.1 $Y=0.815
c65 23 0 1.56657e-19 $X=1.775 $Y=0.82
r66 29 35 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=0.365
+ $X2=1.9 $Y2=0.365
r67 29 31 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.365
+ $X2=2.78 $Y2=0.365
r68 26 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.9 $Y=0.735 $X2=1.9
+ $Y2=0.73
r69 25 35 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.9 $Y=0.475 $X2=1.9
+ $Y2=0.365
r70 25 28 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.9 $Y=0.475
+ $X2=1.9 $Y2=0.73
r71 24 33 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.265 $Y=0.82
+ $X2=1.1 $Y2=0.815
r72 23 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.775 $Y=0.82
+ $X2=1.9 $Y2=0.735
r73 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=0.82
+ $X2=1.265 $Y2=0.82
r74 19 33 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.1 $Y=0.725 $X2=1.1
+ $Y2=0.815
r75 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=0.725 $X2=1.1
+ $Y2=0.39
r76 17 33 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.815
+ $X2=1.1 $Y2=0.815
r77 17 18 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.815
+ $X2=0.425 $Y2=0.815
r78 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.425 $Y2=0.815
r79 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.26 $Y2=0.39
r80 4 31 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.39
r81 3 35 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.39
r82 3 28 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.73
r83 2 21 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r84 1 15 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%VGND 1 2 3 4 5 6 21 25 29 33 35 39 43 46 47
+ 49 50 52 53 54 55 57 58 59 85 86 89
r118 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r119 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r120 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r121 83 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r122 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r123 80 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0 $X2=5.82
+ $Y2=0
r124 80 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.21 $Y2=0
r125 79 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r126 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r127 76 79 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.83 $Y2=0
r128 75 78 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=4.83
+ $Y2=0
r129 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r130 73 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r131 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r132 70 73 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.99 $Y2=0
r133 69 72 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r134 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r135 67 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r136 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r137 59 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r138 59 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r139 57 82 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.21 $Y2=0
r140 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0 $X2=6.66
+ $Y2=0
r141 56 85 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=7.13 $Y2=0
r142 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0 $X2=6.66
+ $Y2=0
r143 54 78 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.83
+ $Y2=0
r144 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.98
+ $Y2=0
r145 52 72 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=0
+ $X2=2.99 $Y2=0
r146 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.3
+ $Y2=0
r147 51 75 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.45
+ $Y2=0
r148 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.3
+ $Y2=0
r149 49 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0
+ $X2=1.15 $Y2=0
r150 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.52
+ $Y2=0
r151 48 69 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.61
+ $Y2=0
r152 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.52
+ $Y2=0
r153 46 62 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r154 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r155 45 66 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=1.15 $Y2=0
r156 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r157 41 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0
r158 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0.39
r159 37 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r160 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.39
r161 36 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r162 35 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.82
+ $Y2=0
r163 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.065 $Y2=0
r164 31 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r165 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.39
r166 27 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.085 $X2=3.3
+ $Y2=0
r167 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0.39
r168 23 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r169 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.39
r170 19 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r171 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.39
r172 6 43 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.39
r173 5 39 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.39
r174 4 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.39
r175 3 29 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.3 $Y2=0.39
r176 2 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r177 1 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2A_4%A_717_47# 1 2 7 11 13
c23 13 0 6.86556e-20 $X=4.56 $Y=0.73
r24 11 16 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=0.475 $X2=4.6
+ $Y2=0.39
r25 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.6 $Y=0.475
+ $X2=4.6 $Y2=0.73
r26 7 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.475 $Y=0.39 $X2=4.6
+ $Y2=0.39
r27 7 9 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.475 $Y=0.39
+ $X2=3.72 $Y2=0.39
r28 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.39
r29 2 13 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.73
r30 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.39
.ends


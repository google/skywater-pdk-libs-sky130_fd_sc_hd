* File: sky130_fd_sc_hd__or4_2.spice.SKY130_FD_SC_HD__OR4_2.pxi
* Created: Thu Aug 27 14:44:07 2020
* 
x_PM_SKY130_FD_SC_HD__OR4_2%D N_D_M1005_g N_D_M1009_g D D N_D_c_66_n
+ PM_SKY130_FD_SC_HD__OR4_2%D
x_PM_SKY130_FD_SC_HD__OR4_2%C N_C_M1011_g N_C_M1000_g C C N_C_c_94_n
+ PM_SKY130_FD_SC_HD__OR4_2%C
x_PM_SKY130_FD_SC_HD__OR4_2%B N_B_M1002_g N_B_M1004_g N_B_c_131_n N_B_c_132_n B
+ B B N_B_c_134_n N_B_c_135_n PM_SKY130_FD_SC_HD__OR4_2%B
x_PM_SKY130_FD_SC_HD__OR4_2%A N_A_M1003_g N_A_M1008_g A N_A_c_170_n N_A_c_171_n
+ PM_SKY130_FD_SC_HD__OR4_2%A
x_PM_SKY130_FD_SC_HD__OR4_2%A_27_297# N_A_27_297#_M1005_d N_A_27_297#_M1004_d
+ N_A_27_297#_M1009_s N_A_27_297#_c_211_n N_A_27_297#_M1006_g
+ N_A_27_297#_M1001_g N_A_27_297#_c_212_n N_A_27_297#_M1007_g
+ N_A_27_297#_M1010_g N_A_27_297#_c_222_n N_A_27_297#_c_305_p
+ N_A_27_297#_c_213_n N_A_27_297#_c_214_n N_A_27_297#_c_316_p
+ N_A_27_297#_c_215_n N_A_27_297#_c_250_n N_A_27_297#_c_223_n
+ N_A_27_297#_c_224_n N_A_27_297#_c_216_n N_A_27_297#_c_225_n
+ N_A_27_297#_c_217_n N_A_27_297#_c_218_n N_A_27_297#_c_219_n
+ PM_SKY130_FD_SC_HD__OR4_2%A_27_297#
x_PM_SKY130_FD_SC_HD__OR4_2%VPWR N_VPWR_M1008_d N_VPWR_M1010_s N_VPWR_c_334_n
+ N_VPWR_c_335_n N_VPWR_c_336_n VPWR N_VPWR_c_337_n N_VPWR_c_338_n
+ N_VPWR_c_339_n N_VPWR_c_333_n PM_SKY130_FD_SC_HD__OR4_2%VPWR
x_PM_SKY130_FD_SC_HD__OR4_2%X N_X_M1006_d N_X_M1001_d N_X_c_368_n N_X_c_370_n
+ N_X_c_366_n X PM_SKY130_FD_SC_HD__OR4_2%X
x_PM_SKY130_FD_SC_HD__OR4_2%VGND N_VGND_M1005_s N_VGND_M1011_d N_VGND_M1003_d
+ N_VGND_M1007_s N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n
+ N_VGND_c_395_n N_VGND_c_396_n VGND N_VGND_c_397_n N_VGND_c_398_n
+ N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n
+ PM_SKY130_FD_SC_HD__OR4_2%VGND
cc_1 VNB N_D_M1005_g 0.0343362f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB D 0.0237123f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_D_c_66_n 0.0355361f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_C_M1011_g 0.0257827f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_5 VNB C 0.00562839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_C_c_94_n 0.0180743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_M1002_g 0.0181193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B_c_131_n 0.013575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_c_132_n 0.0128829f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_10 VNB N_A_M1003_g 0.0266374f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_11 VNB N_A_c_170_n 0.0206834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_c_171_n 0.00322228f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_13 VNB N_A_27_297#_c_211_n 0.0164401f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_14 VNB N_A_27_297#_c_212_n 0.0187042f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_15 VNB N_A_27_297#_c_213_n 0.00394971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_297#_c_214_n 0.00296979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_215_n 0.00105916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_216_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_217_n 0.00185649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_297#_c_218_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_297#_c_219_n 0.0462852f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_333_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_366_n 7.68963e-19 $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_24 VNB N_VGND_c_391_n 0.0104794f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_25 VNB N_VGND_c_392_n 0.0170104f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_26 VNB N_VGND_c_393_n 8.05577e-19 $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=0.85
cc_27 VNB N_VGND_c_394_n 5.60747e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_395_n 0.0118506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_396_n 0.0118658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_397_n 0.014035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_398_n 0.0115649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_399_n 0.0171221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_400_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_401_n 0.0052385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_402_n 0.188966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_D_M1009_g 0.0267282f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_37 VPB D 0.00363927f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_38 VPB N_D_c_66_n 0.0095147f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_39 VPB N_C_M1000_g 0.01663f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_40 VPB C 0.0018547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_C_c_94_n 0.00440081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B_M1002_g 0.0243581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B_c_134_n 0.0369905f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_44 VPB N_B_c_135_n 0.0473847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_M1008_g 0.021674f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_46 VPB N_A_c_170_n 0.00401117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_c_171_n 0.00159111f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_48 VPB N_A_27_297#_M1001_g 0.0209283f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_A_27_297#_M1010_g 0.0245282f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.16
cc_50 VPB N_A_27_297#_c_222_n 0.00536076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_297#_c_223_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_297#_c_224_n 0.0211961f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_297#_c_225_n 0.00201186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_297#_c_219_n 0.00736414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_334_n 0.0121128f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_56 VPB N_VPWR_c_335_n 0.0118214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_336_n 0.00792914f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_58 VPB N_VPWR_c_337_n 0.0489433f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=0.85
cc_59 VPB N_VPWR_c_338_n 0.018077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_339_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_333_n 0.0629537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_X_c_366_n 0.00111849f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_63 N_D_M1005_g N_C_M1011_g 0.0171645f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_64 D N_C_M1011_g 8.90377e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_65 N_D_M1009_g N_C_M1000_g 0.0254979f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_66 D C 0.0279811f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_67 N_D_c_66_n C 0.00905747f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_68 D N_C_c_94_n 2.65642e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_69 N_D_c_66_n N_C_c_94_n 0.0207331f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_70 N_D_M1009_g N_B_c_135_n 0.00441071f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_71 N_D_M1009_g N_A_27_297#_c_222_n 0.0112539f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_72 D N_A_27_297#_c_222_n 9.67991e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_73 N_D_M1005_g N_A_27_297#_c_214_n 0.00368534f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_74 D N_A_27_297#_c_214_n 0.00556624f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_75 N_D_M1009_g N_A_27_297#_c_224_n 0.0068783f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_76 D N_A_27_297#_c_224_n 0.0247997f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_77 N_D_c_66_n N_A_27_297#_c_224_n 0.00190153f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_78 N_D_M1005_g N_VGND_c_392_n 0.0102216f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_79 D N_VGND_c_392_n 0.0264529f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_80 N_D_c_66_n N_VGND_c_392_n 0.00113138f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_81 N_D_M1005_g N_VGND_c_393_n 5.21337e-19 $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_82 N_D_M1005_g N_VGND_c_397_n 0.00430458f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_83 N_D_M1005_g N_VGND_c_402_n 0.00749122f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_84 D N_VGND_c_402_n 0.00188851f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_85 C N_B_M1002_g 0.0186858f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_86 N_C_c_94_n N_B_M1002_g 0.041154f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_87 N_C_M1011_g N_B_c_131_n 0.0136904f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_88 N_C_M1011_g N_B_c_132_n 0.041154f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_89 N_C_M1000_g N_B_c_135_n 0.00439246f $X=0.95 $Y=1.695 $X2=0 $Y2=0
cc_90 C N_A_M1008_g 8.9759e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_91 C N_A_c_170_n 2.87148e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_92 C N_A_c_171_n 0.0281805f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_93 N_C_M1000_g N_A_27_297#_c_222_n 0.00925462f $X=0.95 $Y=1.695 $X2=0 $Y2=0
cc_94 C N_A_27_297#_c_222_n 0.0421076f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_95 N_C_c_94_n N_A_27_297#_c_222_n 3.74254e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_96 N_C_M1011_g N_A_27_297#_c_213_n 0.0110261f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_97 C N_A_27_297#_c_213_n 0.0414766f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_98 N_C_c_94_n N_A_27_297#_c_213_n 0.00179145f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_99 C N_A_27_297#_c_214_n 0.0152593f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_100 N_C_c_94_n N_A_27_297#_c_214_n 9.23324e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_101 N_C_M1000_g N_A_27_297#_c_224_n 9.69353e-19 $X=0.95 $Y=1.695 $X2=0 $Y2=0
cc_102 C N_A_27_297#_c_224_n 0.00868841f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_103 C N_A_27_297#_c_225_n 0.00860775f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_104 C A_109_297# 0.00398871f $X=1.07 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_105 C A_205_297# 0.00106447f $X=1.07 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_106 N_C_M1011_g N_VGND_c_392_n 5.50776e-19 $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_107 N_C_M1011_g N_VGND_c_393_n 0.00712013f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_108 N_C_M1011_g N_VGND_c_397_n 0.00322006f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_109 N_C_M1011_g N_VGND_c_402_n 0.00401385f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_110 N_B_M1002_g N_A_M1003_g 0.0033853f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_111 N_B_c_131_n N_A_M1003_g 0.0187947f $X=1.34 $Y=0.76 $X2=0 $Y2=0
cc_112 N_B_M1002_g N_A_M1008_g 0.0231912f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_113 N_B_c_135_n N_A_M1008_g 9.99953e-19 $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_114 N_B_M1002_g N_A_c_170_n 0.0150712f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_115 N_B_M1002_g N_A_c_171_n 0.00214352f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_116 N_B_M1002_g N_A_27_297#_c_222_n 0.0112861f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_117 N_B_c_134_n N_A_27_297#_c_222_n 0.00103679f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_118 N_B_c_135_n N_A_27_297#_c_222_n 0.0815054f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_119 N_B_c_131_n N_A_27_297#_c_213_n 0.00683722f $X=1.34 $Y=0.76 $X2=0 $Y2=0
cc_120 N_B_c_132_n N_A_27_297#_c_213_n 0.00984378f $X=1.34 $Y=0.91 $X2=0 $Y2=0
cc_121 N_B_c_135_n N_A_27_297#_c_250_n 0.0017825f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_122 N_B_c_135_n N_A_27_297#_c_224_n 0.026488f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_123 N_B_M1002_g N_A_27_297#_c_225_n 0.00491229f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_124 N_B_c_135_n N_A_27_297#_c_225_n 0.0138062f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_125 N_B_M1002_g N_VPWR_c_334_n 0.00249809f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_126 N_B_c_134_n N_VPWR_c_334_n 7.14013e-19 $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_127 N_B_c_135_n N_VPWR_c_334_n 0.0251801f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_128 N_B_c_134_n N_VPWR_c_337_n 0.00736312f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_129 N_B_c_135_n N_VPWR_c_337_n 0.0835718f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_130 N_B_c_134_n N_VPWR_c_333_n 0.0106165f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_131 N_B_c_135_n N_VPWR_c_333_n 0.0605377f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_132 N_B_c_131_n N_VGND_c_393_n 0.00673662f $X=1.34 $Y=0.76 $X2=0 $Y2=0
cc_133 N_B_c_132_n N_VGND_c_393_n 2.19529e-19 $X=1.34 $Y=0.91 $X2=0 $Y2=0
cc_134 N_B_c_131_n N_VGND_c_394_n 5.25642e-19 $X=1.34 $Y=0.76 $X2=0 $Y2=0
cc_135 N_B_c_131_n N_VGND_c_398_n 0.00322006f $X=1.34 $Y=0.76 $X2=0 $Y2=0
cc_136 N_B_c_131_n N_VGND_c_402_n 0.00390029f $X=1.34 $Y=0.76 $X2=0 $Y2=0
cc_137 N_A_M1003_g N_A_27_297#_c_211_n 0.0172443f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_138 N_A_M1008_g N_A_27_297#_M1001_g 0.0190165f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_139 N_A_c_171_n N_A_27_297#_c_222_n 7.66792e-19 $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_c_171_n N_A_27_297#_c_213_n 3.58777e-19 $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_M1003_g N_A_27_297#_c_215_n 0.0116543f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_142 N_A_c_170_n N_A_27_297#_c_215_n 0.00220162f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_c_171_n N_A_27_297#_c_215_n 0.0166868f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_M1008_g N_A_27_297#_c_250_n 0.013079f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_145 N_A_c_171_n N_A_27_297#_c_250_n 0.0131508f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_M1008_g N_A_27_297#_c_223_n 0.0034529f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_147 N_A_c_170_n N_A_27_297#_c_216_n 5.77159e-19 $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_c_171_n N_A_27_297#_c_216_n 0.0146254f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_M1008_g N_A_27_297#_c_225_n 0.00166288f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_150 N_A_c_170_n N_A_27_297#_c_225_n 8.39213e-19 $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_c_171_n N_A_27_297#_c_225_n 0.0130897f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_c_170_n N_A_27_297#_c_217_n 0.00186332f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_c_171_n N_A_27_297#_c_217_n 0.0261029f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_M1003_g N_A_27_297#_c_218_n 0.0034529f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_155 N_A_c_170_n N_A_27_297#_c_219_n 0.0203649f $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_171_n N_A_27_297#_c_219_n 3.5395e-19 $X=1.775 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_M1008_g N_VPWR_c_334_n 0.00298728f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_158 N_A_M1008_g N_VPWR_c_337_n 0.00264561f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_159 N_A_M1008_g N_VPWR_c_333_n 0.00333991f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_160 N_A_M1003_g N_VGND_c_393_n 5.2354e-19 $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_161 N_A_M1003_g N_VGND_c_394_n 0.00709299f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_162 N_A_M1003_g N_VGND_c_398_n 0.00322006f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_163 N_A_M1003_g N_VGND_c_402_n 0.00390029f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_164 N_A_27_297#_c_222_n A_109_297# 0.00243923f $X=1.51 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_165 N_A_27_297#_c_222_n A_205_297# 0.00102299f $X=1.51 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_27_297#_c_222_n A_277_297# 0.00246778f $X=1.51 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_27_297#_c_225_n A_277_297# 0.00526734f $X=1.595 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_27_297#_c_250_n N_VPWR_M1008_d 0.00526233f $X=2.065 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_27_297#_M1001_g N_VPWR_c_334_n 0.00348231f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_27_297#_c_250_n N_VPWR_c_334_n 0.0190361f $X=2.065 $Y=1.58 $X2=0
+ $Y2=0
cc_171 N_A_27_297#_c_225_n N_VPWR_c_334_n 0.0030545f $X=1.595 $Y=1.58 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_c_219_n N_VPWR_c_334_n 2.11345e-19 $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_27_297#_M1010_g N_VPWR_c_336_n 0.00639159f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_27_297#_M1001_g N_VPWR_c_338_n 0.00585385f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_27_297#_M1010_g N_VPWR_c_338_n 0.00503406f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_M1001_g N_VPWR_c_333_n 0.0118387f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_M1010_g N_VPWR_c_333_n 0.00967739f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_c_212_n N_X_c_368_n 0.00536146f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_27_297#_c_219_n N_X_c_368_n 0.00259703f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_27_297#_M1010_g N_X_c_370_n 0.00294462f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_27_297#_c_219_n N_X_c_370_n 0.00288868f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_211_n N_X_c_366_n 0.00151661f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_27_297#_M1001_g N_X_c_366_n 0.00115345f $X=2.28 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_27_297#_c_212_n N_X_c_366_n 0.00462154f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_27_297#_M1010_g N_X_c_366_n 0.00707148f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_27_297#_c_215_n N_X_c_366_n 0.00352178f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A_27_297#_c_223_n N_X_c_366_n 0.00841218f $X=2.15 $Y=1.495 $X2=0 $Y2=0
cc_188 N_A_27_297#_c_217_n N_X_c_366_n 0.0232251f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_27_297#_c_218_n N_X_c_366_n 0.00836616f $X=2.202 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_27_297#_c_219_n N_X_c_366_n 0.0229104f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_27_297#_M1010_g X 0.0119134f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_27_297#_c_213_n N_VGND_M1011_d 0.00160115f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_27_297#_c_215_n N_VGND_M1003_d 0.00482895f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_218_n N_VGND_M1003_d 6.98847e-19 $X=2.202 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_27_297#_c_305_p N_VGND_c_392_n 0.0182596f $X=0.71 $Y=0.47 $X2=0 $Y2=0
cc_196 N_A_27_297#_c_305_p N_VGND_c_393_n 0.0117247f $X=0.71 $Y=0.47 $X2=0 $Y2=0
cc_197 N_A_27_297#_c_213_n N_VGND_c_393_n 0.0160613f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_c_211_n N_VGND_c_394_n 0.0079064f $X=2.28 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_c_212_n N_VGND_c_394_n 9.49203e-19 $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_27_297#_c_215_n N_VGND_c_394_n 0.020701f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_27_297#_c_219_n N_VGND_c_394_n 2.33671e-19 $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_27_297#_c_212_n N_VGND_c_396_n 0.00815799f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_c_305_p N_VGND_c_397_n 0.00876148f $X=0.71 $Y=0.47 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_c_213_n N_VGND_c_397_n 0.00276686f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_205 N_A_27_297#_c_213_n N_VGND_c_398_n 0.00232396f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_27_297#_c_316_p N_VGND_c_398_n 0.00846569f $X=1.58 $Y=0.47 $X2=0
+ $Y2=0
cc_207 N_A_27_297#_c_215_n N_VGND_c_398_n 0.00232396f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A_27_297#_c_211_n N_VGND_c_399_n 0.00524631f $X=2.28 $Y=0.995 $X2=0
+ $Y2=0
cc_209 N_A_27_297#_c_212_n N_VGND_c_399_n 0.00513402f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_27_297#_c_215_n N_VGND_c_399_n 3.34073e-19 $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_211 N_A_27_297#_c_211_n N_VGND_c_402_n 0.00851181f $X=2.28 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_27_297#_c_212_n N_VGND_c_402_n 0.00968535f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_27_297#_c_305_p N_VGND_c_402_n 0.00625722f $X=0.71 $Y=0.47 $X2=0
+ $Y2=0
cc_214 N_A_27_297#_c_213_n N_VGND_c_402_n 0.0105423f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_27_297#_c_316_p N_VGND_c_402_n 0.00625722f $X=1.58 $Y=0.47 $X2=0
+ $Y2=0
cc_216 N_A_27_297#_c_215_n N_VGND_c_402_n 0.00637905f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_333_n N_X_M1001_d 0.00393857f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_336_n N_X_c_366_n 0.0733959f $X=2.935 $Y=1.66 $X2=0 $Y2=0
cc_219 N_VPWR_c_338_n X 0.0168871f $X=2.85 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_c_333_n X 0.0102668f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_c_336_n N_VGND_c_396_n 0.0079302f $X=2.935 $Y=1.66 $X2=0 $Y2=0
cc_222 N_X_c_368_n N_VGND_c_396_n 0.0250997f $X=2.595 $Y=0.587 $X2=0 $Y2=0
cc_223 N_X_c_366_n N_VGND_c_396_n 0.0169659f $X=2.542 $Y=1.495 $X2=0 $Y2=0
cc_224 N_X_c_368_n N_VGND_c_399_n 0.00796253f $X=2.595 $Y=0.587 $X2=0 $Y2=0
cc_225 N_X_M1006_d N_VGND_c_402_n 0.00409985f $X=2.355 $Y=0.235 $X2=0 $Y2=0
cc_226 N_X_c_368_n N_VGND_c_402_n 0.00913686f $X=2.595 $Y=0.587 $X2=0 $Y2=0

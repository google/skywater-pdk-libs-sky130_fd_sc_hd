* File: sky130_fd_sc_hd__a211oi_4.pex.spice
* Created: Thu Aug 27 13:59:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A211OI_4%A2 3 7 11 15 19 23 25 27 30 32 36 37 39 51
+ 54 59 62
c123 37 0 1.77722e-19 $X=3.41 $Y=1.16
c124 30 0 1.03215e-19 $X=3.41 $Y=1.985
c125 19 0 1.41833e-19 $X=1.31 $Y=0.56
r126 54 59 1.31771 $w=5.88e-07 $l=6.5e-08 $layer=LI1_cond $X=1.09 $Y=1.33
+ $X2=1.155 $Y2=1.33
r127 50 62 9.68168 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=1.33
+ $X2=1.385 $Y2=1.33
r128 49 51 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.22 $Y=1.16 $X2=1.31
+ $Y2=1.16
r129 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.16 $X2=1.22 $Y2=1.16
r130 47 49 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.22 $Y2=1.16
r131 45 47 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=0.88 $Y=1.16 $X2=0.89
+ $Y2=1.16
r132 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.88
+ $Y=1.16 $X2=0.88 $Y2=1.16
r133 42 45 91.0912 $w=2.7e-07 $l=4.1e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.88 $Y2=1.16
r134 39 50 1.11499 $w=5.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.165 $Y=1.33
+ $X2=1.22 $Y2=1.33
r135 39 59 0.202725 $w=5.88e-07 $l=1e-08 $layer=LI1_cond $X=1.165 $Y=1.33
+ $X2=1.155 $Y2=1.33
r136 39 54 0.202725 $w=5.88e-07 $l=1e-08 $layer=LI1_cond $X=1.08 $Y=1.33
+ $X2=1.09 $Y2=1.33
r137 39 46 4.0545 $w=5.88e-07 $l=2e-07 $layer=LI1_cond $X=1.08 $Y=1.33 $X2=0.88
+ $Y2=1.33
r138 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.16 $X2=3.41 $Y2=1.16
r139 34 36 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.41 $Y=1.445
+ $X2=3.41 $Y2=1.16
r140 32 34 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.245 $Y=1.535
+ $X2=3.41 $Y2=1.445
r141 32 62 114.606 $w=1.78e-07 $l=1.86e-06 $layer=LI1_cond $X=3.245 $Y=1.535
+ $X2=1.385 $Y2=1.535
r142 28 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r143 28 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r144 25 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r145 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r146 21 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r147 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r148 17 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r149 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r150 13 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r151 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r152 9 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.16
r153 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r154 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r155 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.985
r156 1 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r157 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%A1 3 7 11 15 19 23 27 31 35 41 46 47
r73 45 47 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=2.84 $Y=1.16
+ $X2=2.99 $Y2=1.16
r74 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.84
+ $Y=1.16 $X2=2.84 $Y2=1.16
r75 43 45 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.84 $Y2=1.16
r76 42 43 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16 $X2=2.57
+ $Y2=1.16
r77 40 42 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=2.15 $Y2=1.16
r78 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.82
+ $Y=1.16 $X2=1.82 $Y2=1.16
r79 37 40 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.73 $Y=1.16 $X2=1.82
+ $Y2=1.16
r80 35 46 36.7341 $w=2.38e-07 $l=7.65e-07 $layer=LI1_cond $X=2.075 $Y=1.155
+ $X2=2.84 $Y2=1.155
r81 35 41 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=2.075 $Y=1.155
+ $X2=1.82 $Y2=1.155
r82 29 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r83 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r84 25 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r85 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r86 21 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r87 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r88 17 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r89 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r90 13 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r91 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r92 9 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r93 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r94 5 37 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r95 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295 $X2=1.73
+ $Y2=1.985
r96 1 37 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r97 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%B1 1 3 6 10 12 14 17 19 21 24 27 31 38 39
+ 41 42 44 45 47 57 60 69
c140 69 0 1.88781e-19 $X=4.46 $Y=1.325
c141 42 0 1.03215e-19 $X=4.06 $Y=1.53
c142 41 0 1.74717e-19 $X=6.53 $Y=1.53
c143 39 0 3.99932e-19 $X=6.85 $Y=1.16
c144 17 0 1.85098e-19 $X=4.67 $Y=1.985
r145 56 57 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=1.16
+ $X2=4.745 $Y2=1.16
r146 53 69 8.55056 $w=5.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.25 $Y=1.325
+ $X2=4.46 $Y2=1.325
r147 53 65 6.90838 $w=5.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.25 $Y=1.325
+ $X2=3.915 $Y2=1.325
r148 52 54 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=4.25 $Y=1.16
+ $X2=4.315 $Y2=1.16
r149 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.25
+ $Y=1.16 $X2=4.25 $Y2=1.16
r150 49 52 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.83 $Y=1.16
+ $X2=4.25 $Y2=1.16
r151 47 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.915 $Y=1.53
+ $X2=3.915 $Y2=1.53
r152 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.675 $Y=1.53
+ $X2=6.675 $Y2=1.53
r153 42 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.53
+ $X2=3.915 $Y2=1.53
r154 41 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.53 $Y=1.53
+ $X2=6.675 $Y2=1.53
r155 41 42 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=6.53 $Y=1.53
+ $X2=4.06 $Y2=1.53
r156 39 61 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.852 $Y=1.16
+ $X2=6.852 $Y2=1.325
r157 39 60 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.852 $Y=1.16
+ $X2=6.852 $Y2=0.995
r158 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.16 $X2=6.85 $Y2=1.16
r159 35 45 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.675 $Y=1.325
+ $X2=6.675 $Y2=1.53
r160 34 38 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=6.675 $Y=1.16
+ $X2=6.85 $Y2=1.16
r161 34 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=1.16
+ $X2=6.675 $Y2=1.325
r162 32 56 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=4.59 $Y=1.16 $X2=4.67
+ $Y2=1.16
r163 32 54 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=4.59 $Y=1.16
+ $X2=4.315 $Y2=1.16
r164 31 69 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=4.59 $Y=1.155
+ $X2=4.46 $Y2=1.155
r165 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.59
+ $Y=1.16 $X2=4.59 $Y2=1.16
r166 27 61 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.89 $Y=1.985
+ $X2=6.89 $Y2=1.325
r167 24 60 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.86 $Y=0.56
+ $X2=6.86 $Y2=0.995
r168 19 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=0.995
+ $X2=4.745 $Y2=1.16
r169 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.745 $Y=0.995
+ $X2=4.745 $Y2=0.56
r170 15 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=1.325
+ $X2=4.67 $Y2=1.16
r171 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.67 $Y=1.325
+ $X2=4.67 $Y2=1.985
r172 12 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=0.995
+ $X2=4.315 $Y2=1.16
r173 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.315 $Y=0.995
+ $X2=4.315 $Y2=0.56
r174 8 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=1.325
+ $X2=4.25 $Y2=1.16
r175 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.25 $Y=1.325
+ $X2=4.25 $Y2=1.985
r176 4 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.325
+ $X2=3.83 $Y2=1.16
r177 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.83 $Y=1.325
+ $X2=3.83 $Y2=1.985
r178 1 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=1.16
r179 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%C1 3 5 7 10 12 14 17 19 21 22 24 27 31 33
+ 35 48
c89 48 0 1.88781e-19 $X=6.43 $Y=1.16
c90 33 0 2.33752e-19 $X=6.185 $Y=1.16
r91 45 46 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.98 $Y=1.16 $X2=6.01
+ $Y2=1.16
r92 44 45 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=5.59 $Y=1.16
+ $X2=5.98 $Y2=1.16
r93 43 44 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=5.55 $Y=1.16 $X2=5.59
+ $Y2=1.16
r94 42 43 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=5.17 $Y=1.16
+ $X2=5.55 $Y2=1.16
r95 40 42 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=5.165 $Y=1.16
+ $X2=5.17 $Y2=1.16
r96 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.165
+ $Y=1.16 $X2=5.165 $Y2=1.16
r97 37 40 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=5.12 $Y=1.16
+ $X2=5.165 $Y2=1.16
r98 35 41 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=5.295 $Y=1.155
+ $X2=5.165 $Y2=1.155
r99 34 48 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=6.185 $Y=1.16
+ $X2=6.43 $Y2=1.16
r100 34 46 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.185 $Y=1.16
+ $X2=6.01 $Y2=1.16
r101 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.185
+ $Y=1.16 $X2=6.185 $Y2=1.16
r102 31 35 40.0954 $w=2.38e-07 $l=8.35e-07 $layer=LI1_cond $X=6.13 $Y=1.155
+ $X2=5.295 $Y2=1.155
r103 31 33 3.26808 $w=2.4e-07 $l=1.1e-07 $layer=LI1_cond $X=6.13 $Y=1.155
+ $X2=6.24 $Y2=1.155
r104 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.16
r105 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.325
+ $X2=6.43 $Y2=1.985
r106 22 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=1.16
r107 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=0.56
r108 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.01 $Y=0.995
+ $X2=6.01 $Y2=1.16
r109 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.01 $Y=0.995
+ $X2=6.01 $Y2=0.56
r110 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.98 $Y=1.325
+ $X2=5.98 $Y2=1.16
r111 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.98 $Y=1.325
+ $X2=5.98 $Y2=1.985
r112 12 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.59 $Y=0.995
+ $X2=5.59 $Y2=1.16
r113 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.59 $Y=0.995
+ $X2=5.59 $Y2=0.56
r114 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.55 $Y=1.325
+ $X2=5.55 $Y2=1.16
r115 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.55 $Y=1.325
+ $X2=5.55 $Y2=1.985
r116 5 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=1.16
r117 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=0.56
r118 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.12 $Y=1.325
+ $X2=5.12 $Y2=1.16
r119 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.12 $Y=1.325
+ $X2=5.12 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%noxref_7 1 2 3 4 5 6 7 22 24 26 30 32 36 38
+ 42 44 46 47 52 57 59 61
c94 46 0 2.91989e-20 $X=3.62 $Y=2.105
c95 44 0 1.48523e-19 $X=3.535 $Y=1.95
c96 7 0 1.30877e-19 $X=6.965 $Y=1.485
r97 50 52 139.429 $w=2.08e-07 $l=2.64e-06 $layer=LI1_cond $X=4.46 $Y=2.36
+ $X2=7.1 $Y2=2.36
r98 48 65 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=2.36
+ $X2=3.62 $Y2=2.36
r99 48 50 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=3.705 $Y=2.36
+ $X2=4.46 $Y2=2.36
r100 47 65 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.62 $Y=2.255
+ $X2=3.62 $Y2=2.36
r101 46 63 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.62 $Y=2.105
+ $X2=3.62 $Y2=1.95
r102 46 47 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.62 $Y=2.105
+ $X2=3.62 $Y2=2.255
r103 45 61 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.95
+ $X2=2.78 $Y2=1.95
r104 44 63 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=1.95
+ $X2=3.62 $Y2=1.95
r105 44 45 24.9076 $w=3.08e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=1.95
+ $X2=2.865 $Y2=1.95
r106 40 61 3.57226 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.78 $Y=2.105
+ $X2=2.78 $Y2=1.95
r107 40 42 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.78 $Y=2.105
+ $X2=2.78 $Y2=2.3
r108 39 59 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.95
+ $X2=1.94 $Y2=1.95
r109 38 61 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=1.95
+ $X2=2.78 $Y2=1.95
r110 38 39 24.9076 $w=3.08e-07 $l=6.7e-07 $layer=LI1_cond $X=2.695 $Y=1.95
+ $X2=2.025 $Y2=1.95
r111 34 59 3.57226 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.94 $Y=2.105
+ $X2=1.94 $Y2=1.95
r112 34 36 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.94 $Y=2.105
+ $X2=1.94 $Y2=2.3
r113 33 57 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.95 $X2=1.1
+ $Y2=1.95
r114 32 59 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=1.95
+ $X2=1.94 $Y2=1.95
r115 32 33 24.9076 $w=3.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=1.95
+ $X2=1.185 $Y2=1.95
r116 28 57 3.44808 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.1 $Y=2.105
+ $X2=1.1 $Y2=1.95
r117 28 30 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.1 $Y=2.105
+ $X2=1.1 $Y2=2.3
r118 27 55 3.17836 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=0.345 $Y=1.94
+ $X2=0.22 $Y2=1.94
r119 26 57 3.14896 $w=3e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.015 $Y=1.94
+ $X2=1.1 $Y2=1.95
r120 26 27 26.6254 $w=2.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=1.94
+ $X2=0.345 $Y2=1.94
r121 22 55 3.6869 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=0.22 $Y=2.085
+ $X2=0.22 $Y2=1.94
r122 22 24 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=0.22 $Y=2.085
+ $X2=0.22 $Y2=2.3
r123 7 52 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=2.34
r124 6 50 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=2.36
r125 5 65 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2.3
r126 5 63 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.96
r127 4 61 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.96
r128 4 42 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2.3
r129 3 59 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r130 3 36 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.3
r131 2 57 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r132 2 30 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.3
r133 1 55 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r134 1 24 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 59 60 63
c112 59 0 9.10281e-20 $X=7.13 $Y=2.72
r113 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 59 60 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r115 57 60 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=7.13 $Y2=2.72
r116 56 59 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=7.13 $Y2=2.72
r117 56 57 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r118 54 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r120 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r121 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r122 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r123 48 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r125 45 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r126 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r128 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r129 38 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r131 36 53 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=2.99 $Y2=2.72
r132 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=3.2 $Y2=2.72
r133 35 56 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=2.72
+ $X2=3.45 $Y2=2.72
r134 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=2.72
+ $X2=3.2 $Y2=2.72
r135 33 50 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.36 $Y2=2.72
r137 32 53 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.99 $Y2=2.72
r138 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.36 $Y2=2.72
r139 30 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.52 $Y2=2.72
r141 29 50 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.72
+ $X2=1.52 $Y2=2.72
r143 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635 $X2=3.2
+ $Y2=2.72
r144 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2.36
r145 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r146 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.36
r147 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r148 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.36
r149 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r150 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r151 4 27 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.36
r152 3 23 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.36
r153 2 19 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.36
r154 1 15 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%noxref_9 1 2 7 13 15
r45 15 17 15.0229 $w=2.78e-07 $l=3.65e-07 $layer=LI1_cond $X=4.77 $Y=1.57
+ $X2=4.77 $Y2=1.935
r46 11 15 1.39851 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=4.91 $Y=1.57 $X2=4.77
+ $Y2=1.57
r47 11 13 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=4.91 $Y=1.57
+ $X2=5.765 $Y2=1.57
r48 7 17 0.291325 $w=3e-07 $l=1.4e-07 $layer=LI1_cond $X=4.63 $Y=1.935 $X2=4.77
+ $Y2=1.935
r49 7 9 22.6647 $w=2.98e-07 $l=5.9e-07 $layer=LI1_cond $X=4.63 $Y=1.935 $X2=4.04
+ $Y2=1.935
r50 2 13 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=5.625
+ $Y=1.485 $X2=5.765 $Y2=1.61
r51 1 9 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%Y 1 2 3 4 5 6 7 8 25 31 35 37 41 43 45 53
+ 55 57 63 65 67 69 70 71 72 73 76
c142 76 0 9.10281e-20 $X=7.102 $Y=1.865
c143 72 0 1.30877e-19 $X=7.102 $Y=1.495
c144 70 0 1.74717e-19 $X=6.355 $Y=0.74
c145 57 0 1.06175e-19 $X=7.105 $Y=0.72
c146 45 0 3.51279e-19 $X=6.93 $Y=1.975
c147 25 0 1.41833e-19 $X=3.235 $Y=0.77
r148 73 76 2.83177 $w=3.45e-07 $l=1.1e-07 $layer=LI1_cond $X=7.102 $Y=1.975
+ $X2=7.102 $Y2=1.865
r149 73 76 1.33617 $w=3.43e-07 $l=4e-08 $layer=LI1_cond $X=7.102 $Y=1.825
+ $X2=7.102 $Y2=1.865
r150 71 73 5.27785 $w=3.43e-07 $l=1.58e-07 $layer=LI1_cond $X=7.102 $Y=1.667
+ $X2=7.102 $Y2=1.825
r151 71 72 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=7.102 $Y=1.667
+ $X2=7.102 $Y2=1.495
r152 61 72 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.19 $Y=0.825
+ $X2=7.19 $Y2=1.495
r153 60 70 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=6.65 $Y=0.72
+ $X2=6.355 $Y2=0.72
r154 57 61 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.105 $Y=0.72
+ $X2=7.19 $Y2=0.825
r155 57 60 24.0303 $w=2.08e-07 $l=4.55e-07 $layer=LI1_cond $X=7.105 $Y=0.72
+ $X2=6.65 $Y2=0.72
r156 56 69 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=0.74
+ $X2=5.8 $Y2=0.74
r157 55 70 6.09095 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.23 $Y=0.74
+ $X2=6.355 $Y2=0.74
r158 55 56 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=6.23 $Y=0.74
+ $X2=5.885 $Y2=0.74
r159 51 69 2.68609 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.8 $Y=0.615
+ $X2=5.8 $Y2=0.74
r160 51 53 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.8 $Y=0.615
+ $X2=5.8 $Y2=0.42
r161 47 50 46.0977 $w=2.18e-07 $l=8.8e-07 $layer=LI1_cond $X=5.335 $Y=1.975
+ $X2=6.215 $Y2=1.975
r162 45 73 4.42786 $w=2.2e-07 $l=1.72e-07 $layer=LI1_cond $X=6.93 $Y=1.975
+ $X2=7.102 $Y2=1.975
r163 45 50 37.4544 $w=2.18e-07 $l=7.15e-07 $layer=LI1_cond $X=6.93 $Y=1.975
+ $X2=6.215 $Y2=1.975
r164 44 67 3.77418 $w=2.45e-07 $l=8.74643e-08 $layer=LI1_cond $X=5.045 $Y=0.745
+ $X2=4.96 $Y2=0.74
r165 43 69 3.77418 $w=2.45e-07 $l=8.74643e-08 $layer=LI1_cond $X=5.715 $Y=0.745
+ $X2=5.8 $Y2=0.74
r166 43 44 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=5.715 $Y=0.745
+ $X2=5.045 $Y2=0.745
r167 39 67 2.68609 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.96 $Y=0.615
+ $X2=4.96 $Y2=0.74
r168 39 41 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.96 $Y=0.615
+ $X2=4.96 $Y2=0.42
r169 38 65 7.22005 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=4.195 $Y=0.74
+ $X2=4.035 $Y2=0.74
r170 37 67 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=0.74
+ $X2=4.96 $Y2=0.74
r171 37 38 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.875 $Y=0.74
+ $X2=4.195 $Y2=0.74
r172 33 65 0.120199 $w=3.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.035 $Y=0.615
+ $X2=4.035 $Y2=0.74
r173 33 35 7.0227 $w=3.18e-07 $l=1.95e-07 $layer=LI1_cond $X=4.035 $Y=0.615
+ $X2=4.035 $Y2=0.42
r174 31 65 7.22005 $w=2.1e-07 $l=1.78885e-07 $layer=LI1_cond $X=3.875 $Y=0.78
+ $X2=4.035 $Y2=0.74
r175 31 63 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.875 $Y=0.78
+ $X2=3.33 $Y2=0.78
r176 27 30 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=1.94 $Y=0.77
+ $X2=2.78 $Y2=0.77
r177 25 63 5.69365 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=3.235 $Y=0.77
+ $X2=3.33 $Y2=0.77
r178 25 30 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=3.235 $Y=0.77
+ $X2=2.78 $Y2=0.77
r179 8 50 600 $w=1.7e-07 $l=5.69408e-07 $layer=licon1_PDIFF $count=1 $X=6.055
+ $Y=1.485 $X2=6.215 $Y2=1.98
r180 7 47 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=5.195
+ $Y=1.485 $X2=5.335 $Y2=1.98
r181 6 60 182 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.65 $Y2=0.74
r182 5 69 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=5.665
+ $Y=0.235 $X2=5.8 $Y2=0.76
r183 5 53 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.665
+ $Y=0.235 $X2=5.8 $Y2=0.42
r184 4 67 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.235 $X2=4.96 $Y2=0.76
r185 4 41 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.235 $X2=4.96 $Y2=0.42
r186 3 65 182 $w=1.7e-07 $l=5.97495e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.06 $Y2=0.76
r187 3 35 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.06 $Y2=0.42
r188 2 30 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.76
r189 1 27 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%VGND 1 2 3 4 5 6 7 22 24 28 32 34 38 40 44
+ 48 50 52 54 55 56 58 67 72 81 84 87 90 94
c126 50 0 1.06175e-19 $X=7.092 $Y=0.085
r127 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r128 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r129 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r130 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r131 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r132 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r133 76 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r134 76 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r135 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r136 73 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=0 $X2=6.22
+ $Y2=0
r137 73 75 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.385 $Y=0
+ $X2=6.67 $Y2=0
r138 72 93 5.03279 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=7.137 $Y2=0
r139 72 75 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.67
+ $Y2=0
r140 71 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r141 71 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r142 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r143 68 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.545 $Y=0 $X2=5.38
+ $Y2=0
r144 68 70 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.545 $Y=0
+ $X2=5.75 $Y2=0
r145 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.055 $Y=0 $X2=6.22
+ $Y2=0
r146 67 70 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.055 $Y=0
+ $X2=5.75 $Y2=0
r147 66 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r148 66 82 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=1.15
+ $Y2=0
r149 65 66 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r150 63 81 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.067 $Y2=0
r151 63 65 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=3.45 $Y2=0
r152 62 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r153 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r154 59 78 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r155 59 61 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r156 58 81 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.067
+ $Y2=0
r157 58 61 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.69
+ $Y2=0
r158 56 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r159 56 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r160 54 65 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.45
+ $Y2=0
r161 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.62
+ $Y2=0
r162 50 93 2.94713 $w=3.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=7.092 $Y=0.085
+ $X2=7.137 $Y2=0
r163 50 52 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=7.092 $Y=0.085
+ $X2=7.092 $Y2=0.36
r164 46 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=0.085
+ $X2=6.22 $Y2=0
r165 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.22 $Y=0.085
+ $X2=6.22 $Y2=0.36
r166 42 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.38 $Y=0.085
+ $X2=5.38 $Y2=0
r167 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.38 $Y=0.085
+ $X2=5.38 $Y2=0.36
r168 41 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.695 $Y=0 $X2=4.53
+ $Y2=0
r169 40 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.38
+ $Y2=0
r170 40 41 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.215 $Y=0
+ $X2=4.695 $Y2=0
r171 36 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.085
+ $X2=4.53 $Y2=0
r172 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.53 $Y=0.085
+ $X2=4.53 $Y2=0.36
r173 35 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.62
+ $Y2=0
r174 34 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=0 $X2=4.53
+ $Y2=0
r175 34 35 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.365 $Y=0
+ $X2=3.705 $Y2=0
r176 30 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0
r177 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0.36
r178 26 81 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.067 $Y=0.085
+ $X2=1.067 $Y2=0
r179 26 28 13.486 $w=2.33e-07 $l=2.75e-07 $layer=LI1_cond $X=1.067 $Y=0.085
+ $X2=1.067 $Y2=0.36
r180 22 78 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.197 $Y2=0
r181 22 24 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.38
r182 7 52 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.935
+ $Y=0.235 $X2=7.08 $Y2=0.36
r183 6 48 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.235 $X2=6.22 $Y2=0.36
r184 5 44 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.38 $Y2=0.36
r185 4 38 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.235 $X2=4.53 $Y2=0.36
r186 3 32 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.36
r187 2 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.36
r188 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_4%A_109_47# 1 2 3 4 13 15 16 21 24
r39 24 26 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=0.67 $Y=0.7 $X2=0.67
+ $Y2=0.78
r40 19 21 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.38 $X2=3.2
+ $Y2=0.38
r41 17 29 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.605 $Y=0.38
+ $X2=1.48 $Y2=0.38
r42 17 19 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=1.605 $Y=0.38
+ $X2=2.36 $Y2=0.38
r43 15 29 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.48 $Y=0.505
+ $X2=1.48 $Y2=0.38
r44 15 16 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=1.48 $Y=0.505
+ $X2=1.48 $Y2=0.695
r45 14 26 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.775 $Y=0.78
+ $X2=0.67 $Y2=0.78
r46 13 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.355 $Y=0.78
+ $X2=1.48 $Y2=0.695
r47 13 14 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.355 $Y=0.78
+ $X2=0.775 $Y2=0.78
r48 4 21 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.36
r49 3 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.36
r50 2 29 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.36
r51 1 24 182 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.7
.ends


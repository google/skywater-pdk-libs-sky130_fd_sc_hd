# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.075000 4.975000 1.320000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 1.800000 1.275000 ;
    END
  END SLEEP
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.385000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 2.295000 0.905000 2.625000 1.445000 ;
        RECT 2.295000 1.445000 3.305000 1.745000 ;
        RECT 2.295000 1.745000 2.465000 2.125000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.135000 1.745000 3.305000 2.125000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.905000 ;
      RECT 0.085000  1.455000 2.125000 1.665000 ;
      RECT 0.085000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.465000 ;
      RECT 1.375000  1.835000 1.625000 2.635000 ;
      RECT 1.795000  1.665000 2.125000 2.295000 ;
      RECT 1.795000  2.295000 3.855000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.635000  1.935000 2.965000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 2.795000  1.075000 4.275000 1.275000 ;
      RECT 3.475000  1.575000 3.855000 2.295000 ;
      RECT 3.555000  0.085000 3.845000 0.905000 ;
      RECT 4.025000  0.255000 4.355000 0.815000 ;
      RECT 4.025000  0.815000 4.275000 1.075000 ;
      RECT 4.025000  1.275000 4.275000 1.575000 ;
      RECT 4.025000  1.575000 4.355000 2.465000 ;
      RECT 4.525000  0.085000 4.815000 0.905000 ;
      RECT 4.525000  1.495000 4.930000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_4
END LIBRARY

* File: sky130_fd_sc_hd__nand3b_4.pex.spice
* Created: Thu Aug 27 14:29:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND3B_4%A_N 3 7 9 12
c28 12 0 1.22725e-19 $X=0.595 $Y=1.16
r29 12 15 43.5052 $w=3.65e-07 $l=1.45e-07 $layer=POLY_cond $X=0.577 $Y=1.16
+ $X2=0.577 $Y2=1.305
r30 12 14 43.5052 $w=3.65e-07 $l=1.45e-07 $layer=POLY_cond $X=0.577 $Y=1.16
+ $X2=0.577 $Y2=1.015
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r32 9 13 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.595 $Y2=1.175
r33 7 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.305
r34 3 14 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 47 51 54 60 63 64 68 76
c113 60 0 1.47016e-19 $X=2.46 $Y=1.16
c114 33 0 1.99733e-19 $X=2.67 $Y=0.56
c115 9 0 1.22725e-19 $X=1.41 $Y=0.56
r116 73 74 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.83 $Y=1.16
+ $X2=2.25 $Y2=1.16
r117 68 71 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.41 $Y2=1.16
r118 67 68 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.335 $Y2=1.16
r119 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r120 61 76 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.46 $Y=1.16
+ $X2=2.67 $Y2=1.16
r121 61 74 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.46 $Y=1.16
+ $X2=2.25 $Y2=1.16
r122 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r123 58 73 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.62 $Y=1.16
+ $X2=1.83 $Y2=1.16
r124 58 71 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.62 $Y=1.16
+ $X2=1.41 $Y2=1.16
r125 57 60 46.5818 $w=1.98e-07 $l=8.4e-07 $layer=LI1_cond $X=1.62 $Y=1.175
+ $X2=2.46 $Y2=1.175
r126 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.16 $X2=1.62 $Y2=1.16
r127 55 66 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=1.285 $Y=1.175
+ $X2=1.145 $Y2=1.175
r128 55 57 18.5773 $w=1.98e-07 $l=3.35e-07 $layer=LI1_cond $X=1.285 $Y=1.175
+ $X2=1.62 $Y2=1.175
r129 54 66 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=1.145 $Y=1.075
+ $X2=1.145 $Y2=1.175
r130 53 54 6.99698 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.145 $Y=0.905
+ $X2=1.145 $Y2=1.075
r131 52 63 2.45687 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=0.425 $Y=0.81
+ $X2=0.255 $Y2=0.81
r132 51 53 7.1467 $w=1.9e-07 $l=1.81384e-07 $layer=LI1_cond $X=1.005 $Y=0.81
+ $X2=1.145 $Y2=0.905
r133 51 52 33.8565 $w=1.88e-07 $l=5.8e-07 $layer=LI1_cond $X=1.005 $Y=0.81
+ $X2=0.425 $Y2=0.81
r134 47 49 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=2.34
r135 45 64 8.46734 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=1.615
+ $X2=0.255 $Y2=1.445
r136 45 47 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.255 $Y=1.615
+ $X2=0.255 $Y2=1.66
r137 43 63 3.98378 $w=2.57e-07 $l=1.30038e-07 $layer=LI1_cond $X=0.172 $Y=0.905
+ $X2=0.255 $Y2=0.81
r138 43 64 34.2234 $w=1.73e-07 $l=5.4e-07 $layer=LI1_cond $X=0.172 $Y=0.905
+ $X2=0.172 $Y2=1.445
r139 39 63 3.98378 $w=2.57e-07 $l=9.5e-08 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.81
r140 39 41 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.38
r141 35 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.16
r142 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.985
r143 31 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=1.16
r144 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=0.56
r145 27 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.16
r146 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.985
r147 23 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=1.16
r148 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=0.56
r149 19 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.16
r150 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.985
r151 15 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=1.16
r152 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=0.56
r153 11 71 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.16
r154 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.985
r155 7 71 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.16
r156 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r157 2 49 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r158 2 47 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r159 1 41 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%B 3 7 11 15 19 23 27 31 33 34 35 46
c78 46 0 1.47016e-19 $X=4.35 $Y=1.16
r79 44 46 52.2108 $w=2.7e-07 $l=2.35e-07 $layer=POLY_cond $X=4.115 $Y=1.16
+ $X2=4.35 $Y2=1.16
r80 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.115
+ $Y=1.16 $X2=4.115 $Y2=1.16
r81 42 44 41.1021 $w=2.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.115 $Y2=1.16
r82 41 42 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.51 $Y=1.16 $X2=3.93
+ $Y2=1.16
r83 39 41 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.09 $Y=1.16 $X2=3.51
+ $Y2=1.16
r84 35 45 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.115 $Y2=1.175
r85 34 45 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=4.115 $Y2=1.175
r86 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.935 $Y2=1.175
r87 29 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.16
r88 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.985
r89 25 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=1.16
r90 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
r91 21 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.16
r92 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.985
r93 17 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=1.16
r94 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=0.56
r95 13 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.16
r96 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.985
r97 9 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=1.16
r98 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=0.56
r99 5 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.16
r100 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.985
r101 1 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=1.16
r102 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%C 3 7 11 15 19 23 27 31 33 34 35 36 41 52
r83 50 52 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=6.335 $Y=1.16
+ $X2=6.55 $Y2=1.16
r84 48 50 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=6.13 $Y=1.16
+ $X2=6.335 $Y2=1.16
r85 47 48 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.71 $Y=1.16 $X2=6.13
+ $Y2=1.16
r86 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.29 $Y=1.16 $X2=5.71
+ $Y2=1.16
r87 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.05
+ $Y=1.16 $X2=5.05 $Y2=1.16
r88 41 46 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.215 $Y=1.16
+ $X2=5.29 $Y2=1.16
r89 41 43 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.215 $Y=1.16
+ $X2=5.05 $Y2=1.16
r90 36 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.335
+ $Y=1.16 $X2=6.335 $Y2=1.16
r91 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=5.795 $Y=1.175
+ $X2=6.255 $Y2=1.175
r92 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=5.335 $Y=1.175
+ $X2=5.795 $Y2=1.175
r93 34 44 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=5.335 $Y=1.175
+ $X2=5.05 $Y2=1.175
r94 33 44 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=4.875 $Y=1.175
+ $X2=5.05 $Y2=1.175
r95 29 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.16
r96 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.985
r97 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.55 $Y=1.025
+ $X2=6.55 $Y2=1.16
r98 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.55 $Y=1.025
+ $X2=6.55 $Y2=0.56
r99 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.13 $Y=1.295
+ $X2=6.13 $Y2=1.16
r100 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.13 $Y=1.295
+ $X2=6.13 $Y2=1.985
r101 17 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.13 $Y=1.025
+ $X2=6.13 $Y2=1.16
r102 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.13 $Y=1.025
+ $X2=6.13 $Y2=0.56
r103 13 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.71 $Y=1.295
+ $X2=5.71 $Y2=1.16
r104 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.71 $Y=1.295
+ $X2=5.71 $Y2=1.985
r105 9 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.71 $Y=1.025
+ $X2=5.71 $Y2=1.16
r106 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.71 $Y=1.025
+ $X2=5.71 $Y2=0.56
r107 5 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.29 $Y=1.295
+ $X2=5.29 $Y2=1.16
r108 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.29 $Y=1.295
+ $X2=5.29 $Y2=1.985
r109 1 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.29 $Y=1.025
+ $X2=5.29 $Y2=1.16
r110 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.29 $Y=1.025
+ $X2=5.29 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%VPWR 1 2 3 4 5 6 7 8 9 30 38 42 46 50 55 59
+ 64 65 67 68 70 71 73 74 76 77 78 80 95 107 108 111 114
r107 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r108 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r109 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r110 105 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r111 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r112 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r113 102 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.83 $Y2=2.72
r114 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 99 114 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=5.165 $Y=2.72
+ $X2=4.82 $Y2=2.72
r116 99 101 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.165 $Y=2.72
+ $X2=5.75 $Y2=2.72
r117 98 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r118 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r119 95 114 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.475 $Y=2.72
+ $X2=4.82 $Y2=2.72
r120 95 97 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=2.72
+ $X2=4.37 $Y2=2.72
r121 94 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r122 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r123 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r124 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r125 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r126 88 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r128 85 111 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=0.94 $Y2=2.72
r129 85 87 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.61 $Y2=2.72
r130 80 111 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.94 $Y2=2.72
r131 80 82 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r132 78 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r133 78 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r134 76 104 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.67 $Y2=2.72
r135 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=2.72
+ $X2=6.84 $Y2=2.72
r136 75 107 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=7.13 $Y2=2.72
r137 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=2.72
+ $X2=6.84 $Y2=2.72
r138 73 101 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=2.72
+ $X2=5.75 $Y2=2.72
r139 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=2.72
+ $X2=5.92 $Y2=2.72
r140 72 104 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.005 $Y=2.72
+ $X2=6.67 $Y2=2.72
r141 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.72
+ $X2=5.92 $Y2=2.72
r142 70 93 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.45 $Y2=2.72
r143 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=2.72
+ $X2=3.72 $Y2=2.72
r144 69 97 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=4.37 $Y2=2.72
r145 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.72 $Y2=2.72
r146 67 90 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r147 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.88 $Y2=2.72
r148 66 93 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=3.45 $Y2=2.72
r149 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=2.88 $Y2=2.72
r150 64 87 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r151 64 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.04 $Y2=2.72
r152 63 90 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.53 $Y2=2.72
r153 63 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.04 $Y2=2.72
r154 59 62 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.84 $Y=1.66
+ $X2=6.84 $Y2=2.34
r155 57 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.72
r156 57 62 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.34
r157 53 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.635
+ $X2=5.92 $Y2=2.72
r158 53 55 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.92 $Y=2.635
+ $X2=5.92 $Y2=2
r159 48 114 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.82 $Y=2.635
+ $X2=4.82 $Y2=2.72
r160 48 50 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=4.82 $Y=2.635
+ $X2=4.82 $Y2=2
r161 44 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2.72
r162 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.72 $Y=2.635
+ $X2=3.72 $Y2=2
r163 40 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=2.635
+ $X2=2.88 $Y2=2.72
r164 40 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.88 $Y=2.635
+ $X2=2.88 $Y2=2.34
r165 36 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r166 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2
r167 30 34 11.7874 $w=6.88e-07 $l=6.8e-07 $layer=LI1_cond $X=0.94 $Y=1.66
+ $X2=0.94 $Y2=2.34
r168 28 111 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=2.635
+ $X2=0.94 $Y2=2.72
r169 28 34 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.94 $Y=2.635
+ $X2=0.94 $Y2=2.34
r170 9 62 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.485 $X2=6.84 $Y2=2.34
r171 9 59 400 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.485 $X2=6.84 $Y2=1.66
r172 8 55 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.785
+ $Y=1.485 $X2=5.92 $Y2=2
r173 7 50 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=4.955
+ $Y=1.485 $X2=5.08 $Y2=2
r174 6 50 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2
r175 5 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2
r176 4 42 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2.34
r177 3 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2
r178 2 34 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.34
r179 2 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.66
r180 1 34 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r181 1 30 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%Y 1 2 3 4 5 6 7 8 25 31 33 39 45 47 51 53
+ 57 59 61 63 68 70 73 74 86 88 91 98
c134 61 0 1.62628e-19 $X=6.34 $Y=1.665
r135 97 98 8.09507 $w=5.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=1.725
+ $X2=3.465 $Y2=1.725
r136 90 92 10.4016 $w=5.58e-07 $l=4.87e-07 $layer=LI1_cond $X=2.46 $Y=1.725
+ $X2=2.947 $Y2=1.725
r137 90 91 8.09507 $w=5.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=1.725
+ $X2=2.295 $Y2=1.725
r138 81 88 1.39805 $w=3.03e-07 $l=3.7e-08 $layer=LI1_cond $X=2.947 $Y=1.227
+ $X2=2.947 $Y2=1.19
r139 74 97 6.08718 $w=5.58e-07 $l=2.85e-07 $layer=LI1_cond $X=3.015 $Y=1.725
+ $X2=3.3 $Y2=1.725
r140 74 92 1.45238 $w=5.58e-07 $l=6.8e-08 $layer=LI1_cond $X=3.015 $Y=1.725
+ $X2=2.947 $Y2=1.725
r141 74 92 4.30533 $w=3.05e-07 $l=2.8e-07 $layer=LI1_cond $X=2.947 $Y=1.445
+ $X2=2.947 $Y2=1.725
r142 73 88 0.90684 $w=3.03e-07 $l=2.4e-08 $layer=LI1_cond $X=2.947 $Y=1.166
+ $X2=2.947 $Y2=1.19
r143 73 86 5.67849 $w=3.03e-07 $l=9.1e-08 $layer=LI1_cond $X=2.947 $Y=1.166
+ $X2=2.947 $Y2=1.075
r144 73 74 6.41267 $w=4.73e-07 $l=1.94e-07 $layer=LI1_cond $X=2.947 $Y=1.251
+ $X2=2.947 $Y2=1.445
r145 73 81 0.90684 $w=3.03e-07 $l=2.4e-08 $layer=LI1_cond $X=2.947 $Y=1.251
+ $X2=2.947 $Y2=1.227
r146 61 72 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.34 $Y=1.665
+ $X2=6.34 $Y2=1.555
r147 61 63 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.34 $Y=1.665
+ $X2=6.34 $Y2=2.34
r148 60 70 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=1.555
+ $X2=5.5 $Y2=1.555
r149 59 72 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=1.555
+ $X2=6.34 $Y2=1.555
r150 59 60 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=6.175 $Y=1.555
+ $X2=5.665 $Y2=1.555
r151 55 70 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=5.5 $Y=1.665
+ $X2=5.5 $Y2=1.555
r152 55 57 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.5 $Y=1.665
+ $X2=5.5 $Y2=2.34
r153 54 68 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=1.555
+ $X2=4.14 $Y2=1.555
r154 53 70 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=1.555
+ $X2=5.5 $Y2=1.555
r155 53 54 53.9553 $w=2.18e-07 $l=1.03e-06 $layer=LI1_cond $X=5.335 $Y=1.555
+ $X2=4.305 $Y2=1.555
r156 49 68 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.14 $Y=1.665
+ $X2=4.14 $Y2=1.555
r157 49 51 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.14 $Y=1.665
+ $X2=4.14 $Y2=2.34
r158 47 68 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=1.555
+ $X2=4.14 $Y2=1.555
r159 47 98 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=3.975 $Y=1.555
+ $X2=3.465 $Y2=1.555
r160 43 97 3.83127 $w=3.3e-07 $l=2.8e-07 $layer=LI1_cond $X=3.3 $Y=2.005 $X2=3.3
+ $Y2=1.725
r161 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.3 $Y=2.005
+ $X2=3.3 $Y2=2.34
r162 41 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.88 $Y=0.905
+ $X2=2.88 $Y2=1.075
r163 37 90 3.83127 $w=3.3e-07 $l=2.8e-07 $layer=LI1_cond $X=2.46 $Y=2.005
+ $X2=2.46 $Y2=1.725
r164 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.46 $Y=2.005
+ $X2=2.46 $Y2=2.34
r165 36 66 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=1.555
+ $X2=1.62 $Y2=1.555
r166 36 91 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=1.785 $Y=1.555
+ $X2=2.295 $Y2=1.555
r167 31 66 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.555
r168 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=2.34
r169 27 30 35.8538 $w=2.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.62 $Y=0.77
+ $X2=2.46 $Y2=0.77
r170 25 41 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.795 $Y=0.77
+ $X2=2.88 $Y2=0.905
r171 25 30 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.795 $Y=0.77
+ $X2=2.46 $Y2=0.77
r172 8 72 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=1.66
r173 8 63 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=2.34
r174 7 70 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.5 $Y2=1.66
r175 7 57 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.5 $Y2=2.34
r176 6 68 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=1.66
r177 6 51 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2.34
r178 5 97 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=1.66
r179 5 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=2.34
r180 4 90 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.66
r181 4 39 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.34
r182 3 66 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=1.66
r183 3 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=2.34
r184 2 30 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.72
r185 1 27 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 59 60 63
r86 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r87 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r88 57 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r89 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r90 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r91 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r92 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r93 50 51 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r94 48 51 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r95 48 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r96 47 50 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r97 47 48 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r98 45 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.72
+ $Y2=0
r99 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r100 40 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.72
+ $Y2=0
r101 40 42 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r102 38 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r103 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r104 36 56 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.67
+ $Y2=0
r105 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.84
+ $Y2=0
r106 35 59 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.13 $Y2=0
r107 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=6.84
+ $Y2=0
r108 33 53 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.75
+ $Y2=0
r109 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.92
+ $Y2=0
r110 32 56 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.005 $Y=0 $X2=6.67
+ $Y2=0
r111 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0 $X2=5.92
+ $Y2=0
r112 30 50 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0 $X2=4.83
+ $Y2=0
r113 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.915 $Y=0 $X2=5.04
+ $Y2=0
r114 29 53 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.75 $Y2=0
r115 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5.04
+ $Y2=0
r116 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0
r117 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0.38
r118 21 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r119 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.38
r120 17 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0
r121 17 19 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0.38
r122 13 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r123 13 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.38
r124 4 27 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=6.625
+ $Y=0.235 $X2=6.84 $Y2=0.38
r125 3 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.235 $X2=5.92 $Y2=0.38
r126 2 19 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.08 $Y2=0.38
r127 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%A_215_47# 1 2 3 4 5 26
r34 24 26 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=3.72 $Y=0.36
+ $X2=4.56 $Y2=0.36
r35 22 24 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=2.88 $Y=0.36
+ $X2=3.72 $Y2=0.36
r36 20 22 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=2.04 $Y=0.36
+ $X2=2.88 $Y2=0.36
r37 17 20 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=1.2 $Y=0.36 $X2=2.04
+ $Y2=0.36
r38 5 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.38
r39 4 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.38
r40 3 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.38
r41 2 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.38
r42 1 17 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_4%A_633_47# 1 2 3 4 13 19 23 25 29 31 32
c58 25 0 1.62628e-19 $X=6.175 $Y=0.81
c59 13 0 1.99733e-19 $X=4.59 $Y=0.77
r60 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.34 $Y=0.715
+ $X2=6.34 $Y2=0.38
r61 26 32 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0.81
+ $X2=5.5 $Y2=0.81
r62 25 27 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=6.175 $Y=0.81
+ $X2=6.34 $Y2=0.715
r63 25 26 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=6.175 $Y=0.81
+ $X2=5.665 $Y2=0.81
r64 21 32 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=5.5 $Y=0.715 $X2=5.5
+ $Y2=0.81
r65 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.5 $Y=0.715 $X2=5.5
+ $Y2=0.38
r66 19 32 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0.81
+ $X2=5.5 $Y2=0.81
r67 19 31 35.6077 $w=1.88e-07 $l=6.1e-07 $layer=LI1_cond $X=5.335 $Y=0.81
+ $X2=4.725 $Y2=0.81
r68 15 18 35.8538 $w=2.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.3 $Y=0.77 $X2=4.14
+ $Y2=0.77
r69 13 31 6.78806 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.59 $Y=0.77
+ $X2=4.725 $Y2=0.77
r70 13 18 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.59 $Y=0.77
+ $X2=4.14 $Y2=0.77
r71 4 29 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.205
+ $Y=0.235 $X2=6.34 $Y2=0.38
r72 3 23 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.365
+ $Y=0.235 $X2=5.5 $Y2=0.38
r73 2 18 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.72
r74 1 15 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.72
.ends


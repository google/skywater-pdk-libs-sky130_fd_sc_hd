* File: sky130_fd_sc_hd__bufinv_16.spice
* Created: Tue Sep  1 18:59:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__bufinv_16.pex.spice"
.subckt sky130_fd_sc_hd__bufinv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1023 N_A_27_47#_M1023_d N_A_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75010.3 A=0.0975 P=1.6 MULT=1
MM1030 N_A_27_47#_M1030_d N_A_M1030_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75009.8 A=0.0975 P=1.6 MULT=1
MM1045 N_A_27_47#_M1030_d N_A_M1045_g N_VGND_M1045_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75009.4 A=0.0975 P=1.6 MULT=1
MM1027 N_A_361_47#_M1027_d N_A_27_47#_M1027_g N_VGND_M1045_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75009 A=0.0975 P=1.6 MULT=1
MM1028 N_A_361_47#_M1027_d N_A_27_47#_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75008.6 A=0.0975 P=1.6 MULT=1
MM1033 N_A_361_47#_M1033_d N_A_27_47#_M1033_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75008.2 A=0.0975 P=1.6 MULT=1
MM1036 N_A_361_47#_M1033_d N_A_27_47#_M1036_g N_VGND_M1036_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75007.7 A=0.0975 P=1.6 MULT=1
MM1040 N_A_361_47#_M1040_d N_A_27_47#_M1040_g N_VGND_M1036_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1041 N_A_361_47#_M1040_d N_A_27_47#_M1041_g N_VGND_M1041_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A_361_47#_M1000_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75006.5 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1000_d N_A_361_47#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75006.1 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_A_361_47#_M1006_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.8
+ SB=75005.6 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1006_d N_A_361_47#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.2
+ SB=75005.2 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1009_d N_A_361_47#_M1009_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.6
+ SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1009_d N_A_361_47#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.1
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1014_d N_A_361_47#_M1014_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.5
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1014_d N_A_361_47#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.9
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1018_d N_A_361_47#_M1018_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.3
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1018_d N_A_361_47#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.7
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1021 N_Y_M1021_d N_A_361_47#_M1021_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1034 N_Y_M1021_d N_A_361_47#_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.6
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1037 N_Y_M1037_d N_A_361_47#_M1037_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1046 N_Y_M1037_d N_A_361_47#_M1046_g N_VGND_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1047 N_Y_M1047_d N_A_361_47#_M1047_g N_VGND_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1049 N_Y_M1047_d N_A_361_47#_M1049_g N_VGND_M1049_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75010.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_27_47#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75010.3 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1007_d N_A_M1012_g N_A_27_47#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75009.8 A=0.15 P=2.3 MULT=1
MM1031 N_VPWR_M1031_d N_A_M1031_g N_A_27_47#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75009.4 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1031_d N_A_27_47#_M1001_g N_A_361_47#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75009 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_27_47#_M1013_g N_A_361_47#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75008.6 A=0.15 P=2.3 MULT=1
MM1029 N_VPWR_M1013_d N_A_27_47#_M1029_g N_A_361_47#_M1029_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75008.2 A=0.15 P=2.3 MULT=1
MM1035 N_VPWR_M1035_d N_A_27_47#_M1035_g N_A_361_47#_M1029_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75007.7 A=0.15 P=2.3 MULT=1
MM1043 N_VPWR_M1035_d N_A_27_47#_M1043_g N_A_361_47#_M1043_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75007.3 A=0.15 P=2.3 MULT=1
MM1044 N_VPWR_M1044_d N_A_27_47#_M1044_g N_A_361_47#_M1043_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75006.9 A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1002_d N_A_361_47#_M1002_g N_VPWR_M1044_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75006.5 A=0.15 P=2.3 MULT=1
MM1003 N_Y_M1002_d N_A_361_47#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4
+ SB=75006.1 A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1004_d N_A_361_47#_M1004_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.8
+ SB=75005.6 A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1004_d N_A_361_47#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.2
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1016 N_Y_M1016_d N_A_361_47#_M1016_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.6
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1017 N_Y_M1016_d N_A_361_47#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.1
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1020 N_Y_M1020_d N_A_361_47#_M1020_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.5
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1022 N_Y_M1020_d N_A_361_47#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.9
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1024 N_Y_M1024_d N_A_361_47#_M1024_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.3
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1025 N_Y_M1024_d N_A_361_47#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.7
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1026 N_Y_M1026_d N_A_361_47#_M1026_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1032 N_Y_M1026_d N_A_361_47#_M1032_g N_VPWR_M1032_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1038 N_Y_M1038_d N_A_361_47#_M1038_g N_VPWR_M1032_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1039 N_Y_M1038_d N_A_361_47#_M1039_g N_VPWR_M1039_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1042 N_Y_M1042_d N_A_361_47#_M1042_g N_VPWR_M1039_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1048 N_Y_M1042_d N_A_361_47#_M1048_g N_VPWR_M1048_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75010.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX50_noxref VNB VPB NWDIODE A=18.3291 P=26.05
*
.include "sky130_fd_sc_hd__bufinv_16.pxi.spice"
*
.ends
*
*

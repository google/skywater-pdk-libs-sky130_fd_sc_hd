* NGSPICE file created from sky130_fd_sc_hd__nand3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=8.1e+11p pd=7.62e+06u as=1.36e+12p ps=1.272e+07u
M1001 VPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR C Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_47# A Y VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u
M1004 VGND C a_277_47# VNB nshort w=650000u l=150000u
+  ad=3.705e+11p pd=3.74e+06u as=3.51e+11p ps=3.68e+06u
M1005 a_277_47# C VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_47# B a_277_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_277_47# B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* NGSPICE file created from sky130_fd_sc_hd__o41a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_103_21# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.2e+11p pd=3.04e+06u as=5.5e+11p ps=5.1e+06u
M1001 a_511_297# A3 a_393_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.9e+11p pd=2.78e+06u as=4.4e+11p ps=2.88e+06u
M1002 VPWR a_103_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=4.25e+11p ps=2.85e+06u
M1003 a_321_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=6.24e+11p pd=5.82e+06u as=6.695e+11p ps=5.96e+06u
M1004 a_321_47# B1 a_103_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1005 a_321_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_619_297# A2 a_511_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.9e+11p pd=2.78e+06u as=0p ps=0u
M1007 VGND A4 a_321_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_393_297# A4 a_103_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_619_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_321_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_103_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.47e+11p ps=2.06e+06u
.ends


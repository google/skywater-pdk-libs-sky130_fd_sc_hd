* File: sky130_fd_sc_hd__fahcin_1.pxi.spice
* Created: Thu Aug 27 14:21:31 2020
* 
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_67_199# N_A_67_199#_M1018_d N_A_67_199#_M1028_s
+ N_A_67_199#_M1010_d N_A_67_199#_M1003_d N_A_67_199#_M1011_d
+ N_A_67_199#_M1007_g N_A_67_199#_M1013_g N_A_67_199#_c_210_n
+ N_A_67_199#_c_217_n N_A_67_199#_c_211_n N_A_67_199#_c_230_p
+ N_A_67_199#_c_326_p N_A_67_199#_c_225_p N_A_67_199#_c_226_p
+ N_A_67_199#_c_235_p N_A_67_199#_c_212_n N_A_67_199#_c_213_n
+ N_A_67_199#_c_219_n N_A_67_199#_c_243_p N_A_67_199#_c_245_p
+ N_A_67_199#_c_246_p N_A_67_199#_c_220_n N_A_67_199#_c_271_p
+ N_A_67_199#_c_221_n N_A_67_199#_c_222_n N_A_67_199#_c_250_p
+ N_A_67_199#_c_251_p N_A_67_199#_c_214_n PM_SKY130_FD_SC_HD__FAHCIN_1%A_67_199#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A N_A_c_398_n N_A_M1018_g N_A_M1010_g A
+ N_A_c_400_n PM_SKY130_FD_SC_HD__FAHCIN_1%A
x_PM_SKY130_FD_SC_HD__FAHCIN_1%B N_B_c_440_n N_B_M1005_g N_B_M1027_g N_B_M1011_g
+ N_B_M1012_g N_B_c_441_n N_B_M1015_g N_B_M1004_g N_B_c_442_n N_B_c_443_n
+ N_B_c_444_n N_B_c_445_n N_B_c_446_n N_B_c_447_n B N_B_c_449_n N_B_c_450_n B
+ N_B_c_451_n N_B_c_452_n PM_SKY130_FD_SC_HD__FAHCIN_1%B
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_489_21# N_A_489_21#_M1015_s N_A_489_21#_M1004_s
+ N_A_489_21#_c_598_n N_A_489_21#_M1026_g N_A_489_21#_M1003_g
+ N_A_489_21#_c_599_n N_A_489_21#_M1028_g N_A_489_21#_M1020_g
+ N_A_489_21#_M1024_g N_A_489_21#_M1006_g N_A_489_21#_c_600_n
+ N_A_489_21#_c_601_n N_A_489_21#_c_602_n N_A_489_21#_c_603_n
+ N_A_489_21#_c_604_n N_A_489_21#_c_605_n N_A_489_21#_c_628_n
+ N_A_489_21#_c_615_n N_A_489_21#_c_616_n N_A_489_21#_c_617_n
+ N_A_489_21#_c_675_p N_A_489_21#_c_618_n N_A_489_21#_c_606_n
+ PM_SKY130_FD_SC_HD__FAHCIN_1%A_489_21#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_434_49# N_A_434_49#_M1005_d N_A_434_49#_M1027_d
+ N_A_434_49#_M1030_g N_A_434_49#_c_756_n N_A_434_49#_M1031_g
+ N_A_434_49#_c_757_n N_A_434_49#_M1019_g N_A_434_49#_M1023_g
+ N_A_434_49#_c_779_n N_A_434_49#_c_758_n N_A_434_49#_c_770_n
+ N_A_434_49#_c_759_n N_A_434_49#_c_788_n N_A_434_49#_c_760_n
+ N_A_434_49#_c_761_n N_A_434_49#_c_762_n N_A_434_49#_c_763_n
+ N_A_434_49#_c_764_n N_A_434_49#_c_765_n N_A_434_49#_c_766_n
+ N_A_434_49#_c_767_n PM_SKY130_FD_SC_HD__FAHCIN_1%A_434_49#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_721_47# N_A_721_47#_M1028_d N_A_721_47#_M1020_d
+ N_A_721_47#_M1009_g N_A_721_47#_c_948_n N_A_721_47#_M1014_g
+ N_A_721_47#_M1029_g N_A_721_47#_c_956_n N_A_721_47#_c_957_n
+ N_A_721_47#_M1000_g N_A_721_47#_c_949_n N_A_721_47#_c_950_n
+ N_A_721_47#_c_951_n N_A_721_47#_c_960_n N_A_721_47#_c_961_n
+ N_A_721_47#_c_962_n N_A_721_47#_c_952_n N_A_721_47#_c_976_n
+ N_A_721_47#_c_991_n N_A_721_47#_c_977_n N_A_721_47#_c_1014_n
+ N_A_721_47#_c_963_n N_A_721_47#_c_1015_n N_A_721_47#_c_964_n
+ N_A_721_47#_c_953_n N_A_721_47#_c_954_n N_A_721_47#_c_967_n
+ PM_SKY130_FD_SC_HD__FAHCIN_1%A_721_47#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_1636_315# N_A_1636_315#_M1019_d
+ N_A_1636_315#_M1022_d N_A_1636_315#_M1000_s N_A_1636_315#_M1016_d
+ N_A_1636_315#_M1001_g N_A_1636_315#_M1002_g N_A_1636_315#_c_1161_n
+ N_A_1636_315#_c_1145_n N_A_1636_315#_c_1146_n N_A_1636_315#_c_1152_n
+ N_A_1636_315#_c_1138_n N_A_1636_315#_c_1159_n N_A_1636_315#_c_1184_p
+ N_A_1636_315#_c_1139_n N_A_1636_315#_c_1140_n N_A_1636_315#_c_1141_n
+ N_A_1636_315#_c_1149_n N_A_1636_315#_c_1160_n N_A_1636_315#_c_1142_n
+ N_A_1636_315#_c_1143_n PM_SKY130_FD_SC_HD__FAHCIN_1%A_1636_315#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%CIN N_CIN_M1016_g N_CIN_c_1262_n N_CIN_M1022_g
+ N_CIN_c_1263_n N_CIN_M1008_g N_CIN_M1021_g N_CIN_c_1264_n N_CIN_c_1265_n
+ N_CIN_c_1266_n CIN PM_SKY130_FD_SC_HD__FAHCIN_1%CIN
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_1647_49# N_A_1647_49#_M1029_d
+ N_A_1647_49#_M1000_d N_A_1647_49#_M1017_g N_A_1647_49#_M1025_g
+ N_A_1647_49#_c_1328_n N_A_1647_49#_c_1329_n N_A_1647_49#_c_1335_n
+ N_A_1647_49#_c_1336_n N_A_1647_49#_c_1337_n N_A_1647_49#_c_1330_n
+ N_A_1647_49#_c_1331_n N_A_1647_49#_c_1332_n N_A_1647_49#_c_1340_n
+ PM_SKY130_FD_SC_HD__FAHCIN_1%A_1647_49#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1026_d
+ N_A_27_47#_M1012_d N_A_27_47#_M1013_s N_A_27_47#_M1027_s N_A_27_47#_M1020_s
+ N_A_27_47#_c_1441_n N_A_27_47#_c_1434_n N_A_27_47#_c_1456_n
+ N_A_27_47#_c_1463_n N_A_27_47#_c_1503_n N_A_27_47#_c_1442_n
+ N_A_27_47#_c_1435_n N_A_27_47#_c_1436_n N_A_27_47#_c_1477_n
+ N_A_27_47#_c_1478_n N_A_27_47#_c_1437_n N_A_27_47#_c_1444_n
+ N_A_27_47#_c_1438_n N_A_27_47#_c_1446_n N_A_27_47#_c_1447_n
+ N_A_27_47#_c_1439_n N_A_27_47#_c_1448_n N_A_27_47#_c_1440_n
+ N_A_27_47#_c_1519_n PM_SKY130_FD_SC_HD__FAHCIN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%VPWR N_VPWR_M1013_d N_VPWR_M1004_d N_VPWR_M1002_d
+ N_VPWR_M1021_d N_VPWR_c_1602_n N_VPWR_c_1603_n N_VPWR_c_1604_n N_VPWR_c_1605_n
+ N_VPWR_c_1606_n VPWR N_VPWR_c_1607_n N_VPWR_c_1608_n N_VPWR_c_1609_n
+ N_VPWR_c_1610_n N_VPWR_c_1601_n N_VPWR_c_1612_n N_VPWR_c_1613_n
+ N_VPWR_c_1614_n N_VPWR_c_1615_n PM_SKY130_FD_SC_HD__FAHCIN_1%VPWR
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_1142_49# N_A_1142_49#_M1024_d
+ N_A_1142_49#_M1014_d N_A_1142_49#_M1006_d N_A_1142_49#_c_1729_n
+ N_A_1142_49#_c_1745_n N_A_1142_49#_c_1738_n N_A_1142_49#_c_1751_n
+ N_A_1142_49#_c_1730_n N_A_1142_49#_c_1732_n N_A_1142_49#_c_1739_n
+ N_A_1142_49#_c_1740_n PM_SKY130_FD_SC_HD__FAHCIN_1%A_1142_49#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%COUT N_COUT_M1031_d N_COUT_M1030_d COUT COUT
+ N_COUT_c_1802_n COUT PM_SKY130_FD_SC_HD__FAHCIN_1%COUT
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_1251_49# N_A_1251_49#_M1031_s
+ N_A_1251_49#_M1008_s N_A_1251_49#_M1009_d N_A_1251_49#_M1021_s
+ N_A_1251_49#_c_1829_n N_A_1251_49#_c_1861_n N_A_1251_49#_c_1834_n
+ N_A_1251_49#_c_1835_n N_A_1251_49#_c_1880_n N_A_1251_49#_c_1838_n
+ N_A_1251_49#_c_1836_n N_A_1251_49#_c_1881_n N_A_1251_49#_c_1830_n
+ N_A_1251_49#_c_1831_n N_A_1251_49#_c_1832_n N_A_1251_49#_c_1889_n
+ N_A_1251_49#_c_1833_n PM_SKY130_FD_SC_HD__FAHCIN_1%A_1251_49#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%A_1565_49# N_A_1565_49#_M1029_s
+ N_A_1565_49#_M1001_s N_A_1565_49#_M1023_d N_A_1565_49#_c_1971_n
+ N_A_1565_49#_c_1963_n N_A_1565_49#_c_2009_n N_A_1565_49#_c_1964_n
+ N_A_1565_49#_c_1965_n N_A_1565_49#_c_1966_n N_A_1565_49#_c_1967_n
+ N_A_1565_49#_c_1993_n PM_SKY130_FD_SC_HD__FAHCIN_1%A_1565_49#
x_PM_SKY130_FD_SC_HD__FAHCIN_1%SUM N_SUM_M1025_d N_SUM_M1017_d SUM SUM SUM SUM
+ SUM SUM N_SUM_c_2022_n PM_SKY130_FD_SC_HD__FAHCIN_1%SUM
x_PM_SKY130_FD_SC_HD__FAHCIN_1%VGND N_VGND_M1007_d N_VGND_M1015_d N_VGND_M1001_d
+ N_VGND_M1008_d N_VGND_c_2040_n N_VGND_c_2041_n N_VGND_c_2042_n N_VGND_c_2043_n
+ N_VGND_c_2044_n N_VGND_c_2045_n VGND N_VGND_c_2046_n N_VGND_c_2047_n
+ N_VGND_c_2048_n N_VGND_c_2049_n N_VGND_c_2050_n N_VGND_c_2051_n
+ N_VGND_c_2052_n PM_SKY130_FD_SC_HD__FAHCIN_1%VGND
cc_1 VNB N_A_67_199#_c_210_n 0.00625651f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.325
cc_2 VNB N_A_67_199#_c_211_n 0.00332932f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.82
cc_3 VNB N_A_67_199#_c_212_n 0.00601615f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.34
cc_4 VNB N_A_67_199#_c_213_n 0.026083f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_5 VNB N_A_67_199#_c_214_n 0.0205236f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_6 VNB N_A_c_398_n 0.020424f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.235
cc_7 VNB A 0.00181874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_c_400_n 0.0300339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_c_440_n 0.0202962f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.235
cc_10 VNB N_B_c_441_n 0.0201069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_c_442_n 0.0344872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_443_n 0.00898261f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.325
cc_13 VNB N_B_c_444_n 0.0181948f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.82
cc_14 VNB N_B_c_445_n 0.021911f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_15 VNB N_B_c_446_n 0.0487553f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.585
cc_16 VNB N_B_c_447_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.465
cc_17 VNB B 0.00417432f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.735
cc_18 VNB N_B_c_449_n 0.00613646f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_19 VNB N_B_c_450_n 0.0034327f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=0.36
cc_20 VNB N_B_c_451_n 8.74233e-19 $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_21 VNB N_B_c_452_n 7.72065e-19 $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_22 VNB N_A_489_21#_c_598_n 0.021145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_489_21#_c_599_n 0.0225157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_489_21#_c_600_n 0.0101537f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.465
cc_25 VNB N_A_489_21#_c_601_n 0.0443961f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.735
cc_26 VNB N_A_489_21#_c_602_n 0.0139301f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_27 VNB N_A_489_21#_c_603_n 0.00188997f $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=0.36
cc_28 VNB N_A_489_21#_c_604_n 0.0020237f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=0.34
cc_29 VNB N_A_489_21#_c_605_n 0.0253462f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_30 VNB N_A_489_21#_c_606_n 0.0203142f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.87
cc_31 VNB N_A_434_49#_c_756_n 0.0189404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_434_49#_c_757_n 0.0188417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_434_49#_c_758_n 0.00346469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_434_49#_c_759_n 0.00950118f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.465
cc_35 VNB N_A_434_49#_c_760_n 0.0076264f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_36 VNB N_A_434_49#_c_761_n 0.00285941f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_37 VNB N_A_434_49#_c_762_n 0.00119646f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.36
cc_38 VNB N_A_434_49#_c_763_n 0.00580264f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_39 VNB N_A_434_49#_c_764_n 0.00190842f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_40 VNB N_A_434_49#_c_765_n 0.0360602f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.87
cc_41 VNB N_A_434_49#_c_766_n 0.047595f $X=-0.19 $Y=-0.24 $X2=3.305 $Y2=0.42
cc_42 VNB N_A_434_49#_c_767_n 0.00151079f $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=1.87
cc_43 VNB N_A_721_47#_c_948_n 0.020289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_721_47#_c_949_n 0.0133977f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.325
cc_45 VNB N_A_721_47#_c_950_n 0.0667997f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.82
cc_46 VNB N_A_721_47#_c_951_n 0.020274f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.82
cc_47 VNB N_A_721_47#_c_952_n 0.00259038f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.34
cc_48 VNB N_A_721_47#_c_953_n 0.00107146f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=0.36
cc_49 VNB N_A_721_47#_c_954_n 0.00363645f $X=-0.19 $Y=-0.24 $X2=4.08 $Y2=1.87
cc_50 VNB N_A_1636_315#_c_1138_n 0.00860754f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_51 VNB N_A_1636_315#_c_1139_n 0.00310926f $X=-0.19 $Y=-0.24 $X2=1.885
+ $Y2=0.38
cc_52 VNB N_A_1636_315#_c_1140_n 0.00517348f $X=-0.19 $Y=-0.24 $X2=0.602
+ $Y2=1.16
cc_53 VNB N_A_1636_315#_c_1141_n 0.00423574f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_54 VNB N_A_1636_315#_c_1142_n 0.0224625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1636_315#_c_1143_n 0.0202796f $X=-0.19 $Y=-0.24 $X2=2.11 $Y2=1.87
cc_56 VNB N_CIN_c_1262_n 0.0207742f $X=-0.19 $Y=-0.24 $X2=4.145 $Y2=1.61
cc_57 VNB N_CIN_c_1263_n 0.0204768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_CIN_c_1264_n 0.0116244f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_59 VNB N_CIN_c_1265_n 0.0437832f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.555
cc_60 VNB N_CIN_c_1266_n 0.0101793f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.555
cc_61 VNB N_A_1647_49#_c_1328_n 0.00385467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1647_49#_c_1329_n 7.04441e-19 $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=1.325
cc_63 VNB N_A_1647_49#_c_1330_n 0.0226007f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=0.36
cc_64 VNB N_A_1647_49#_c_1331_n 0.00571475f $X=-0.19 $Y=-0.24 $X2=1.325 $Y2=0.36
cc_65 VNB N_A_1647_49#_c_1332_n 0.0201404f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.36
cc_66 VNB N_A_27_47#_c_1434_n 0.0187016f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.585
cc_67 VNB N_A_27_47#_c_1435_n 0.0013204f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.34
cc_68 VNB N_A_27_47#_c_1436_n 0.00104233f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.38
cc_69 VNB N_A_27_47#_c_1437_n 0.00295877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_27_47#_c_1438_n 0.0227289f $X=-0.19 $Y=-0.24 $X2=3.305 $Y2=0.42
cc_71 VNB N_A_27_47#_c_1439_n 0.00824219f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.87
cc_72 VNB N_A_27_47#_c_1440_n 0.00372324f $X=-0.19 $Y=-0.24 $X2=4.225 $Y2=1.87
cc_73 VNB N_VPWR_c_1601_n 0.516438f $X=-0.19 $Y=-0.24 $X2=2.51 $Y2=1.87
cc_74 VNB N_A_1142_49#_c_1729_n 0.00685453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1142_49#_c_1730_n 0.00120965f $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=0.555
cc_76 VNB COUT 0.00193947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_COUT_c_1802_n 8.43544e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1251_49#_c_1829_n 0.00597029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1251_49#_c_1830_n 0.0200172f $X=-0.19 $Y=-0.24 $X2=0.602 $Y2=1.16
cc_80 VNB N_A_1251_49#_c_1831_n 0.00443263f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_81 VNB N_A_1251_49#_c_1832_n 0.0110757f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.38
cc_82 VNB N_A_1251_49#_c_1833_n 0.00135949f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.87
cc_83 VNB N_A_1565_49#_c_1963_n 0.00587953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1565_49#_c_1964_n 6.78455e-19 $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=0.995
cc_85 VNB N_A_1565_49#_c_1965_n 0.00734551f $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=0.555
cc_86 VNB N_A_1565_49#_c_1966_n 0.00862893f $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=1.325
cc_87 VNB N_A_1565_49#_c_1967_n 0.00180358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB SUM 0.0297243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_SUM_c_2022_n 0.0160045f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.5
cc_90 VNB N_VGND_c_2040_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.555
cc_91 VNB N_VGND_c_2041_n 0.00294634f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_92 VNB N_VGND_c_2042_n 0.00485258f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.82
cc_93 VNB N_VGND_c_2043_n 0.00288927f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.465
cc_94 VNB N_VGND_c_2044_n 0.111916f $X=-0.19 $Y=-0.24 $X2=1.16 $Y2=0.72
cc_95 VNB N_VGND_c_2045_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=0.36
cc_96 VNB N_VGND_c_2046_n 0.103307f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=0.38
cc_97 VNB N_VGND_c_2047_n 0.0295045f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=0.36
cc_98 VNB N_VGND_c_2048_n 0.0177665f $X=-0.19 $Y=-0.24 $X2=1.965 $Y2=1.87
cc_99 VNB N_VGND_c_2049_n 0.621019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_2050_n 0.0220858f $X=-0.19 $Y=-0.24 $X2=2.655 $Y2=1.87
cc_101 VNB N_VGND_c_2051_n 0.0051639f $X=-0.19 $Y=-0.24 $X2=4.225 $Y2=1.87
cc_102 VNB N_VGND_c_2052_n 0.00514867f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.995
cc_103 VPB N_A_67_199#_M1013_g 0.023979f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_104 VPB N_A_67_199#_c_210_n 0.00109618f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_105 VPB N_A_67_199#_c_217_n 0.00272323f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.5
cc_106 VPB N_A_67_199#_c_213_n 0.00620175f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_107 VPB N_A_67_199#_c_219_n 0.00386384f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.665
cc_108 VPB N_A_67_199#_c_220_n 0.00351091f $X=-0.19 $Y=1.305 $X2=4.08 $Y2=1.87
cc_109 VPB N_A_67_199#_c_221_n 0.00890077f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.87
cc_110 VPB N_A_67_199#_c_222_n 0.00332655f $X=-0.19 $Y=1.305 $X2=2.655 $Y2=1.87
cc_111 VPB N_A_M1010_g 0.0270986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_c_400_n 0.00852415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_B_M1027_g 0.0241329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_B_M1011_g 0.0348198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_B_M1004_g 0.0242935f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_116 VPB N_B_c_442_n 0.0158127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_B_c_443_n 5.80369e-19 $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_118 VPB N_B_c_444_n 0.00229037f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.82
cc_119 VPB N_B_c_446_n 0.0220588f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.585
cc_120 VPB N_B_c_447_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.465
cc_121 VPB B 0.0034641f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.735
cc_122 VPB N_B_c_452_n 0.00255216f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_123 VPB N_A_489_21#_M1003_g 0.0212549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_489_21#_M1020_g 0.0218106f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_125 VPB N_A_489_21#_M1006_g 0.0229057f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_126 VPB N_A_489_21#_c_600_n 7.08375e-19 $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.465
cc_127 VPB N_A_489_21#_c_601_n 0.0246268f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.735
cc_128 VPB N_A_489_21#_c_602_n 8.40309e-19 $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_129 VPB N_A_489_21#_c_604_n 0.00329861f $X=-0.19 $Y=1.305 $X2=2.1 $Y2=0.34
cc_130 VPB N_A_489_21#_c_605_n 0.00613509f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_131 VPB N_A_489_21#_c_615_n 0.0160478f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_489_21#_c_616_n 0.00558812f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.665
cc_133 VPB N_A_489_21#_c_617_n 0.00676255f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_489_21#_c_618_n 0.00842032f $X=-0.19 $Y=1.305 $X2=2.51 $Y2=1.87
cc_135 VPB N_A_434_49#_M1030_g 0.0208531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_434_49#_M1023_g 0.0284423f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_137 VPB N_A_434_49#_c_770_n 0.00251074f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.82
cc_138 VPB N_A_434_49#_c_761_n 4.7406e-19 $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_139 VPB N_A_434_49#_c_762_n 0.00272473f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=0.36
cc_140 VPB N_A_434_49#_c_763_n 8.12858e-19 $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.82
cc_141 VPB N_A_434_49#_c_764_n 4.66358e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_142 VPB N_A_434_49#_c_765_n 0.0115302f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.87
cc_143 VPB N_A_434_49#_c_766_n 0.00534447f $X=-0.19 $Y=1.305 $X2=3.305 $Y2=0.42
cc_144 VPB N_A_721_47#_M1009_g 0.0216864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_721_47#_c_956_n 0.0230178f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_146 VPB N_A_721_47#_c_957_n 0.017473f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_147 VPB N_A_721_47#_c_949_n 0.00248297f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_148 VPB N_A_721_47#_c_950_n 0.0566748f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.82
cc_149 VPB N_A_721_47#_c_960_n 0.00358583f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.72
cc_150 VPB N_A_721_47#_c_961_n 0.0161847f $X=-0.19 $Y=1.305 $X2=1.995 $Y2=0.36
cc_151 VPB N_A_721_47#_c_962_n 0.00224654f $X=-0.19 $Y=1.305 $X2=1.325 $Y2=0.36
cc_152 VPB N_A_721_47#_c_963_n 0.0165276f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.585
cc_153 VPB N_A_721_47#_c_964_n 0.00625617f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.87
cc_154 VPB N_A_721_47#_c_953_n 0.00206858f $X=-0.19 $Y=1.305 $X2=2.1 $Y2=0.36
cc_155 VPB N_A_721_47#_c_954_n 0.00167678f $X=-0.19 $Y=1.305 $X2=4.08 $Y2=1.87
cc_156 VPB N_A_721_47#_c_967_n 0.00498551f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.87
cc_157 VPB N_A_1636_315#_M1002_g 0.0225f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_158 VPB N_A_1636_315#_c_1145_n 0.00634436f $X=-0.19 $Y=1.305 $X2=0.695
+ $Y2=1.5
cc_159 VPB N_A_1636_315#_c_1146_n 0.00184985f $X=-0.19 $Y=1.305 $X2=0.995
+ $Y2=0.82
cc_160 VPB N_A_1636_315#_c_1138_n 0.00555891f $X=-0.19 $Y=1.305 $X2=1.16
+ $Y2=0.72
cc_161 VPB N_A_1636_315#_c_1141_n 0.0105395f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_162 VPB N_A_1636_315#_c_1149_n 0.00466989f $X=-0.19 $Y=1.305 $X2=1.16
+ $Y2=0.38
cc_163 VPB N_A_1636_315#_c_1142_n 0.00451844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_CIN_M1016_g 0.0232402f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.485
cc_165 VPB N_CIN_M1021_g 0.023149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_CIN_c_1264_n 7.09285e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_167 VPB N_CIN_c_1265_n 0.019685f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_168 VPB N_CIN_c_1266_n 6.56727e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_169 VPB N_A_1647_49#_M1017_g 0.0220957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1647_49#_c_1328_n 7.47965e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_1647_49#_c_1335_n 0.0199045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1647_49#_c_1336_n 0.00101562f $X=-0.19 $Y=1.305 $X2=0.695
+ $Y2=1.325
cc_173 VPB N_A_1647_49#_c_1337_n 0.00131607f $X=-0.19 $Y=1.305 $X2=1.16
+ $Y2=0.465
cc_174 VPB N_A_1647_49#_c_1330_n 0.00600825f $X=-0.19 $Y=1.305 $X2=1.995
+ $Y2=0.36
cc_175 VPB N_A_1647_49#_c_1331_n 0.00253093f $X=-0.19 $Y=1.305 $X2=1.325
+ $Y2=0.36
cc_176 VPB N_A_1647_49#_c_1340_n 0.00490459f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_177 VPB N_A_27_47#_c_1441_n 0.0181919f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.325
cc_178 VPB N_A_27_47#_c_1442_n 0.0148626f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=0.36
cc_179 VPB N_A_27_47#_c_1436_n 0.00206094f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.38
cc_180 VPB N_A_27_47#_c_1444_n 0.020102f $X=-0.19 $Y=1.305 $X2=3.305 $Y2=0.42
cc_181 VPB N_A_27_47#_c_1438_n 0.00898713f $X=-0.19 $Y=1.305 $X2=3.305 $Y2=0.42
cc_182 VPB N_A_27_47#_c_1446_n 0.00880588f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.87
cc_183 VPB N_A_27_47#_c_1447_n 0.00224823f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.87
cc_184 VPB N_A_27_47#_c_1448_n 7.93366e-19 $X=-0.19 $Y=1.305 $X2=2.655 $Y2=1.87
cc_185 VPB N_VPWR_c_1602_n 0.00465796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1603_n 0.105493f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.555
cc_187 VPB N_VPWR_c_1604_n 0.00281836f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_188 VPB N_VPWR_c_1605_n 0.00469901f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.82
cc_189 VPB N_VPWR_c_1606_n 0.00231609f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=0.465
cc_190 VPB N_VPWR_c_1607_n 0.0172154f $X=-0.19 $Y=1.305 $X2=1.995 $Y2=0.36
cc_191 VPB N_VPWR_c_1608_n 0.109665f $X=-0.19 $Y=1.305 $X2=2.1 $Y2=0.34
cc_192 VPB N_VPWR_c_1609_n 0.0312887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1610_n 0.0167387f $X=-0.19 $Y=1.305 $X2=3.305 $Y2=0.42
cc_194 VPB N_VPWR_c_1601_n 0.110293f $X=-0.19 $Y=1.305 $X2=2.51 $Y2=1.87
cc_195 VPB N_VPWR_c_1612_n 0.00323923f $X=-0.19 $Y=1.305 $X2=2.8 $Y2=1.87
cc_196 VPB N_VPWR_c_1613_n 0.00507288f $X=-0.19 $Y=1.305 $X2=1.965 $Y2=1.87
cc_197 VPB N_VPWR_c_1614_n 0.00324066f $X=-0.19 $Y=1.305 $X2=2.655 $Y2=1.87
cc_198 VPB N_VPWR_c_1615_n 0.0036033f $X=-0.19 $Y=1.305 $X2=4.225 $Y2=1.87
cc_199 VPB N_A_1142_49#_c_1729_n 0.00438008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1142_49#_c_1732_n 0.00150393f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.325
cc_201 VPB COUT 0.00104353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_1251_49#_c_1834_n 0.00129808f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.325
cc_203 VPB N_A_1251_49#_c_1835_n 0.00787825f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.985
cc_204 VPB N_A_1251_49#_c_1836_n 0.00249994f $X=-0.19 $Y=1.305 $X2=1.325
+ $Y2=0.36
cc_205 VPB N_A_1251_49#_c_1833_n 0.00183316f $X=-0.19 $Y=1.305 $X2=1.365
+ $Y2=1.87
cc_206 VPB N_A_1565_49#_c_1966_n 0.00380247f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.325
cc_207 VPB SUM 0.0206533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB SUM 0.0287211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 N_A_67_199#_c_210_n N_A_c_398_n 0.0068634f $X=0.695 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_210 N_A_67_199#_c_211_n N_A_c_398_n 0.0105647f $X=0.995 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_67_199#_c_225_p N_A_c_398_n 0.00258977f $X=1.16 $Y=0.465 $X2=-0.19
+ $Y2=-0.24
cc_212 N_A_67_199#_c_226_p N_A_c_398_n 0.00439001f $X=1.16 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_213 N_A_67_199#_c_214_n N_A_c_398_n 0.0190131f $X=0.5 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_67_199#_M1013_g N_A_M1010_g 0.0350328f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_67_199#_c_217_n N_A_M1010_g 0.00394699f $X=0.695 $Y=1.5 $X2=0 $Y2=0
cc_216 N_A_67_199#_c_230_p N_A_M1010_g 0.0125067f $X=1.28 $Y=1.585 $X2=0 $Y2=0
cc_217 N_A_67_199#_c_219_n N_A_M1010_g 0.00744116f $X=1.365 $Y=1.665 $X2=0 $Y2=0
cc_218 N_A_67_199#_c_210_n A 0.0161919f $X=0.695 $Y=1.325 $X2=0 $Y2=0
cc_219 N_A_67_199#_c_211_n A 0.0298669f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_220 N_A_67_199#_c_230_p A 0.0169989f $X=1.28 $Y=1.585 $X2=0 $Y2=0
cc_221 N_A_67_199#_c_235_p A 4.10315e-19 $X=1.995 $Y=0.36 $X2=0 $Y2=0
cc_222 N_A_67_199#_c_219_n A 0.00379181f $X=1.365 $Y=1.665 $X2=0 $Y2=0
cc_223 N_A_67_199#_c_211_n N_A_c_400_n 0.00739621f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_224 N_A_67_199#_c_230_p N_A_c_400_n 0.00511078f $X=1.28 $Y=1.585 $X2=0 $Y2=0
cc_225 N_A_67_199#_c_213_n N_A_c_400_n 0.0208492f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_67_199#_c_219_n N_A_c_400_n 6.89875e-19 $X=1.365 $Y=1.665 $X2=0 $Y2=0
cc_227 N_A_67_199#_c_226_p N_B_c_440_n 0.00324097f $X=1.16 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_228 N_A_67_199#_c_212_n N_B_c_440_n 0.00487626f $X=2.515 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_229 N_A_67_199#_c_243_p N_B_c_440_n 0.00387065f $X=2.1 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_230 N_A_67_199#_c_219_n N_B_M1027_g 0.00857993f $X=1.365 $Y=1.665 $X2=0 $Y2=0
cc_231 N_A_67_199#_c_245_p N_B_M1027_g 0.00207742f $X=2.51 $Y=1.87 $X2=0 $Y2=0
cc_232 N_A_67_199#_c_246_p N_B_M1027_g 0.00279765f $X=2.11 $Y=1.87 $X2=0 $Y2=0
cc_233 N_A_67_199#_c_221_n N_B_M1027_g 0.00700985f $X=1.965 $Y=1.87 $X2=0 $Y2=0
cc_234 N_A_67_199#_c_222_n N_B_M1027_g 0.00108364f $X=2.655 $Y=1.87 $X2=0 $Y2=0
cc_235 N_A_67_199#_c_220_n N_B_M1011_g 0.00258135f $X=4.08 $Y=1.87 $X2=0 $Y2=0
cc_236 N_A_67_199#_c_250_p N_B_M1011_g 7.63489e-19 $X=4.225 $Y=1.87 $X2=0 $Y2=0
cc_237 N_A_67_199#_c_251_p N_B_M1011_g 0.00865293f $X=4.225 $Y=1.87 $X2=0 $Y2=0
cc_238 N_A_67_199#_c_251_p N_B_M1004_g 0.00387974f $X=4.225 $Y=1.87 $X2=0 $Y2=0
cc_239 N_A_67_199#_c_235_p N_B_c_442_n 0.00700393f $X=1.995 $Y=0.36 $X2=0 $Y2=0
cc_240 N_A_67_199#_c_246_p N_B_c_442_n 0.0032044f $X=2.11 $Y=1.87 $X2=0 $Y2=0
cc_241 N_A_67_199#_c_221_n N_B_c_442_n 0.00731952f $X=1.965 $Y=1.87 $X2=0 $Y2=0
cc_242 N_A_67_199#_c_251_p N_B_c_444_n 0.00156571f $X=4.225 $Y=1.87 $X2=0 $Y2=0
cc_243 N_A_67_199#_M1018_d B 0.0077132f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_244 N_A_67_199#_c_211_n B 0.0110561f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_245 N_A_67_199#_c_226_p B 0.00509683f $X=1.16 $Y=0.72 $X2=0 $Y2=0
cc_246 N_A_67_199#_c_235_p B 0.0139594f $X=1.995 $Y=0.36 $X2=0 $Y2=0
cc_247 N_A_67_199#_c_221_n B 0.00861067f $X=1.965 $Y=1.87 $X2=0 $Y2=0
cc_248 N_A_67_199#_M1018_d N_B_c_449_n 0.00199924f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_249 N_A_67_199#_c_235_p N_B_c_449_n 0.00656416f $X=1.995 $Y=0.36 $X2=0 $Y2=0
cc_250 N_A_67_199#_c_212_n N_B_c_449_n 0.00926564f $X=2.515 $Y=0.34 $X2=0 $Y2=0
cc_251 N_A_67_199#_M1018_d N_B_c_450_n 0.00215729f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_252 N_A_67_199#_c_211_n N_B_c_450_n 0.00585767f $X=0.995 $Y=0.82 $X2=0 $Y2=0
cc_253 N_A_67_199#_c_235_p N_B_c_450_n 0.00266787f $X=1.995 $Y=0.36 $X2=0 $Y2=0
cc_254 N_A_67_199#_c_251_p N_B_c_452_n 0.00484475f $X=4.225 $Y=1.87 $X2=0 $Y2=0
cc_255 N_A_67_199#_c_212_n N_A_489_21#_c_598_n 0.0163725f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_256 N_A_67_199#_c_245_p N_A_489_21#_M1003_g 0.00252506f $X=2.51 $Y=1.87 $X2=0
+ $Y2=0
cc_257 N_A_67_199#_c_271_p N_A_489_21#_M1003_g 0.00243281f $X=2.8 $Y=1.87 $X2=0
+ $Y2=0
cc_258 N_A_67_199#_c_221_n N_A_489_21#_M1003_g 5.35429e-19 $X=1.965 $Y=1.87
+ $X2=0 $Y2=0
cc_259 N_A_67_199#_c_222_n N_A_489_21#_M1003_g 0.0051368f $X=2.655 $Y=1.87 $X2=0
+ $Y2=0
cc_260 N_A_67_199#_c_220_n N_A_489_21#_M1020_g 0.0058639f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_261 N_A_67_199#_c_212_n N_A_489_21#_c_601_n 4.57112e-19 $X=2.515 $Y=0.34
+ $X2=0 $Y2=0
cc_262 N_A_67_199#_c_271_p N_A_489_21#_c_601_n 0.00167015f $X=2.8 $Y=1.87 $X2=0
+ $Y2=0
cc_263 N_A_67_199#_c_222_n N_A_489_21#_c_601_n 0.00376167f $X=2.655 $Y=1.87
+ $X2=0 $Y2=0
cc_264 N_A_67_199#_c_220_n N_A_489_21#_c_628_n 3.63034e-19 $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_265 N_A_67_199#_c_271_p N_A_489_21#_c_628_n 0.00105951f $X=2.8 $Y=1.87 $X2=0
+ $Y2=0
cc_266 N_A_67_199#_c_222_n N_A_489_21#_c_628_n 0.00419843f $X=2.655 $Y=1.87
+ $X2=0 $Y2=0
cc_267 N_A_67_199#_c_220_n N_A_489_21#_c_615_n 0.0705151f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_268 N_A_67_199#_c_250_p N_A_489_21#_c_615_n 0.0261743f $X=4.225 $Y=1.87 $X2=0
+ $Y2=0
cc_269 N_A_67_199#_c_251_p N_A_489_21#_c_615_n 0.00878124f $X=4.225 $Y=1.87
+ $X2=0 $Y2=0
cc_270 N_A_67_199#_c_220_n N_A_489_21#_c_616_n 0.0279447f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_271 N_A_67_199#_c_220_n N_A_489_21#_c_617_n 0.00113365f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_272 N_A_67_199#_c_251_p N_A_489_21#_c_618_n 0.00196374f $X=4.225 $Y=1.87
+ $X2=0 $Y2=0
cc_273 N_A_67_199#_c_212_n N_A_434_49#_M1005_d 0.00314538f $X=2.515 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_274 N_A_67_199#_c_245_p N_A_434_49#_M1027_d 0.00460449f $X=2.51 $Y=1.87 $X2=0
+ $Y2=0
cc_275 N_A_67_199#_c_212_n N_A_434_49#_c_779_n 0.0146467f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_276 N_A_67_199#_c_243_p N_A_434_49#_c_779_n 0.00433984f $X=2.1 $Y=0.36 $X2=0
+ $Y2=0
cc_277 N_A_67_199#_c_245_p N_A_434_49#_c_770_n 0.00398041f $X=2.51 $Y=1.87 $X2=0
+ $Y2=0
cc_278 N_A_67_199#_c_246_p N_A_434_49#_c_770_n 9.36352e-19 $X=2.11 $Y=1.87 $X2=0
+ $Y2=0
cc_279 N_A_67_199#_c_271_p N_A_434_49#_c_770_n 9.24792e-19 $X=2.8 $Y=1.87 $X2=0
+ $Y2=0
cc_280 N_A_67_199#_c_245_p N_A_434_49#_c_759_n 0.0129408f $X=2.51 $Y=1.87 $X2=0
+ $Y2=0
cc_281 N_A_67_199#_c_220_n N_A_434_49#_c_759_n 0.00340191f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_282 N_A_67_199#_c_271_p N_A_434_49#_c_759_n 0.0147845f $X=2.8 $Y=1.87 $X2=0
+ $Y2=0
cc_283 N_A_67_199#_c_222_n N_A_434_49#_c_759_n 0.00164718f $X=2.655 $Y=1.87
+ $X2=0 $Y2=0
cc_284 N_A_67_199#_c_245_p N_A_434_49#_c_788_n 0.00481091f $X=2.51 $Y=1.87 $X2=0
+ $Y2=0
cc_285 N_A_67_199#_c_246_p N_A_434_49#_c_788_n 0.00980484f $X=2.11 $Y=1.87 $X2=0
+ $Y2=0
cc_286 N_A_67_199#_c_221_n N_A_434_49#_c_788_n 4.62044e-19 $X=1.965 $Y=1.87
+ $X2=0 $Y2=0
cc_287 N_A_67_199#_c_245_p N_A_434_49#_c_762_n 0.00273443f $X=2.51 $Y=1.87 $X2=0
+ $Y2=0
cc_288 N_A_67_199#_c_246_p N_A_434_49#_c_762_n 0.00207713f $X=2.11 $Y=1.87 $X2=0
+ $Y2=0
cc_289 N_A_67_199#_c_221_n N_A_434_49#_c_762_n 0.00137144f $X=1.965 $Y=1.87
+ $X2=0 $Y2=0
cc_290 N_A_67_199#_c_220_n N_A_721_47#_M1020_d 0.00281165f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_291 N_A_67_199#_c_220_n N_A_721_47#_c_960_n 0.0133801f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_292 N_A_67_199#_c_250_p N_A_721_47#_c_960_n 0.00218435f $X=4.225 $Y=1.87
+ $X2=0 $Y2=0
cc_293 N_A_67_199#_c_251_p N_A_721_47#_c_960_n 0.0253803f $X=4.225 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_67_199#_M1011_d N_A_721_47#_c_961_n 0.00520868f $X=4.145 $Y=1.61
+ $X2=0 $Y2=0
cc_295 N_A_67_199#_c_220_n N_A_721_47#_c_961_n 0.00458634f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_67_199#_c_250_p N_A_721_47#_c_961_n 8.96902e-19 $X=4.225 $Y=1.87
+ $X2=0 $Y2=0
cc_297 N_A_67_199#_c_251_p N_A_721_47#_c_961_n 0.0210702f $X=4.225 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_67_199#_c_251_p N_A_721_47#_c_976_n 0.00243682f $X=4.225 $Y=1.87
+ $X2=0 $Y2=0
cc_299 N_A_67_199#_c_250_p N_A_721_47#_c_977_n 6.37902e-19 $X=4.225 $Y=1.87
+ $X2=0 $Y2=0
cc_300 N_A_67_199#_c_251_p N_A_721_47#_c_977_n 0.00748065f $X=4.225 $Y=1.87
+ $X2=0 $Y2=0
cc_301 N_A_67_199#_c_212_n N_A_27_47#_M1026_d 0.00632791f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_302 N_A_67_199#_c_246_p N_A_27_47#_M1027_s 0.00495068f $X=2.11 $Y=1.87 $X2=0
+ $Y2=0
cc_303 N_A_67_199#_c_221_n N_A_27_47#_M1027_s 0.00546515f $X=1.965 $Y=1.87 $X2=0
+ $Y2=0
cc_304 N_A_67_199#_c_220_n N_A_27_47#_M1020_s 0.00292858f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_305 N_A_67_199#_M1013_g N_A_27_47#_c_1441_n 0.00625347f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_306 N_A_67_199#_c_226_p N_A_27_47#_c_1434_n 0.00527756f $X=1.16 $Y=0.72 $X2=0
+ $Y2=0
cc_307 N_A_67_199#_c_214_n N_A_27_47#_c_1434_n 0.00700681f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_67_199#_M1010_d N_A_27_47#_c_1456_n 0.00186286f $X=1.05 $Y=1.485
+ $X2=0 $Y2=0
cc_309 N_A_67_199#_M1013_g N_A_27_47#_c_1456_n 0.0101197f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_310 N_A_67_199#_c_210_n N_A_27_47#_c_1456_n 0.00414367f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_311 N_A_67_199#_c_230_p N_A_27_47#_c_1456_n 0.0156825f $X=1.28 $Y=1.585 $X2=0
+ $Y2=0
cc_312 N_A_67_199#_c_326_p N_A_27_47#_c_1456_n 0.0137412f $X=0.78 $Y=1.585 $X2=0
+ $Y2=0
cc_313 N_A_67_199#_c_213_n N_A_27_47#_c_1456_n 3.28412e-19 $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_314 N_A_67_199#_c_219_n N_A_27_47#_c_1456_n 0.0138143f $X=1.365 $Y=1.665
+ $X2=0 $Y2=0
cc_315 N_A_67_199#_M1010_d N_A_27_47#_c_1463_n 0.0068106f $X=1.05 $Y=1.485 $X2=0
+ $Y2=0
cc_316 N_A_67_199#_M1013_g N_A_27_47#_c_1463_n 5.25648e-19 $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_317 N_A_67_199#_c_219_n N_A_27_47#_c_1463_n 0.00250582f $X=1.365 $Y=1.665
+ $X2=0 $Y2=0
cc_318 N_A_67_199#_M1003_d N_A_27_47#_c_1442_n 0.00253023f $X=2.595 $Y=1.485
+ $X2=0 $Y2=0
cc_319 N_A_67_199#_c_245_p N_A_27_47#_c_1442_n 0.00706323f $X=2.51 $Y=1.87 $X2=0
+ $Y2=0
cc_320 N_A_67_199#_c_246_p N_A_27_47#_c_1442_n 0.00207268f $X=2.11 $Y=1.87 $X2=0
+ $Y2=0
cc_321 N_A_67_199#_c_220_n N_A_27_47#_c_1442_n 0.00908299f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_322 N_A_67_199#_c_271_p N_A_27_47#_c_1442_n 0.00215819f $X=2.8 $Y=1.87 $X2=0
+ $Y2=0
cc_323 N_A_67_199#_c_221_n N_A_27_47#_c_1442_n 0.00124299f $X=1.965 $Y=1.87
+ $X2=0 $Y2=0
cc_324 N_A_67_199#_c_222_n N_A_27_47#_c_1442_n 0.0119898f $X=2.655 $Y=1.87 $X2=0
+ $Y2=0
cc_325 N_A_67_199#_c_212_n N_A_27_47#_c_1435_n 0.0149451f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_326 N_A_67_199#_c_220_n N_A_27_47#_c_1436_n 0.0145428f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_327 N_A_67_199#_c_271_p N_A_27_47#_c_1436_n 0.00142508f $X=2.8 $Y=1.87 $X2=0
+ $Y2=0
cc_328 N_A_67_199#_c_222_n N_A_27_47#_c_1436_n 0.00881385f $X=2.655 $Y=1.87
+ $X2=0 $Y2=0
cc_329 N_A_67_199#_c_212_n N_A_27_47#_c_1477_n 0.0116127f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_330 N_A_67_199#_c_212_n N_A_27_47#_c_1478_n 0.0148585f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_331 N_A_67_199#_c_210_n N_A_27_47#_c_1437_n 0.00556977f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_332 N_A_67_199#_c_213_n N_A_27_47#_c_1437_n 0.00146618f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_A_67_199#_c_214_n N_A_27_47#_c_1437_n 0.00216178f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_67_199#_M1013_g N_A_27_47#_c_1444_n 0.00819617f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_335 N_A_67_199#_c_210_n N_A_27_47#_c_1444_n 0.0010813f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_336 N_A_67_199#_c_326_p N_A_27_47#_c_1444_n 0.0140939f $X=0.78 $Y=1.585 $X2=0
+ $Y2=0
cc_337 N_A_67_199#_c_213_n N_A_27_47#_c_1444_n 0.00150157f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_A_67_199#_M1013_g N_A_27_47#_c_1438_n 0.00270966f $X=0.475 $Y=1.985
+ $X2=0 $Y2=0
cc_339 N_A_67_199#_c_210_n N_A_27_47#_c_1438_n 0.0315979f $X=0.695 $Y=1.325
+ $X2=0 $Y2=0
cc_340 N_A_67_199#_c_217_n N_A_27_47#_c_1438_n 0.00561378f $X=0.695 $Y=1.5 $X2=0
+ $Y2=0
cc_341 N_A_67_199#_c_213_n N_A_27_47#_c_1438_n 0.00822704f $X=0.51 $Y=1.16 $X2=0
+ $Y2=0
cc_342 N_A_67_199#_c_214_n N_A_27_47#_c_1438_n 0.00268818f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A_67_199#_M1010_d N_A_27_47#_c_1446_n 0.00614173f $X=1.05 $Y=1.485
+ $X2=0 $Y2=0
cc_344 N_A_67_199#_c_230_p N_A_27_47#_c_1446_n 0.00517777f $X=1.28 $Y=1.585
+ $X2=0 $Y2=0
cc_345 N_A_67_199#_c_219_n N_A_27_47#_c_1446_n 0.0132101f $X=1.365 $Y=1.665
+ $X2=0 $Y2=0
cc_346 N_A_67_199#_c_221_n N_A_27_47#_c_1446_n 0.0249023f $X=1.965 $Y=1.87 $X2=0
+ $Y2=0
cc_347 N_A_67_199#_c_246_p N_A_27_47#_c_1447_n 0.00169077f $X=2.11 $Y=1.87 $X2=0
+ $Y2=0
cc_348 N_A_67_199#_M1028_s N_A_27_47#_c_1439_n 0.00239272f $X=3.18 $Y=0.235
+ $X2=0 $Y2=0
cc_349 N_A_67_199#_c_212_n N_A_27_47#_c_1439_n 0.0283951f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_350 N_A_67_199#_c_220_n N_A_27_47#_c_1448_n 0.00289643f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_351 N_A_67_199#_c_217_n N_VPWR_M1013_d 3.11669e-19 $X=0.695 $Y=1.5 $X2=-0.19
+ $Y2=-0.24
cc_352 N_A_67_199#_c_230_p N_VPWR_M1013_d 0.0018145f $X=1.28 $Y=1.585 $X2=-0.19
+ $Y2=-0.24
cc_353 N_A_67_199#_c_326_p N_VPWR_M1013_d 0.00415932f $X=0.78 $Y=1.585 $X2=-0.19
+ $Y2=-0.24
cc_354 N_A_67_199#_M1013_g N_VPWR_c_1602_n 0.00280412f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A_67_199#_M1013_g N_VPWR_c_1607_n 0.0042268f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A_67_199#_M1010_d N_VPWR_c_1601_n 0.00208741f $X=1.05 $Y=1.485 $X2=0
+ $Y2=0
cc_357 N_A_67_199#_M1013_g N_VPWR_c_1601_n 0.00684251f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_358 N_A_67_199#_c_245_p N_VPWR_c_1601_n 0.020224f $X=2.51 $Y=1.87 $X2=0 $Y2=0
cc_359 N_A_67_199#_c_246_p N_VPWR_c_1601_n 0.0160351f $X=2.11 $Y=1.87 $X2=0
+ $Y2=0
cc_360 N_A_67_199#_c_220_n N_VPWR_c_1601_n 0.0630331f $X=4.08 $Y=1.87 $X2=0
+ $Y2=0
cc_361 N_A_67_199#_c_271_p N_VPWR_c_1601_n 0.0149228f $X=2.8 $Y=1.87 $X2=0 $Y2=0
cc_362 N_A_67_199#_c_250_p N_VPWR_c_1601_n 0.0145846f $X=4.225 $Y=1.87 $X2=0
+ $Y2=0
cc_363 N_A_67_199#_c_210_n N_VGND_M1007_d 0.00396202f $X=0.695 $Y=1.325
+ $X2=-0.19 $Y2=-0.24
cc_364 N_A_67_199#_c_211_n N_VGND_M1007_d 5.44633e-19 $X=0.995 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_365 N_A_67_199#_c_210_n N_VGND_c_2040_n 0.0117147f $X=0.695 $Y=1.325 $X2=0
+ $Y2=0
cc_366 N_A_67_199#_c_211_n N_VGND_c_2040_n 0.00132365f $X=0.995 $Y=0.82 $X2=0
+ $Y2=0
cc_367 N_A_67_199#_c_225_p N_VGND_c_2040_n 0.0148348f $X=1.16 $Y=0.465 $X2=0
+ $Y2=0
cc_368 N_A_67_199#_c_226_p N_VGND_c_2040_n 0.00527979f $X=1.16 $Y=0.72 $X2=0
+ $Y2=0
cc_369 N_A_67_199#_c_214_n N_VGND_c_2040_n 0.00383303f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_67_199#_c_211_n N_VGND_c_2046_n 0.00224601f $X=0.995 $Y=0.82 $X2=0
+ $Y2=0
cc_371 N_A_67_199#_c_225_p N_VGND_c_2046_n 0.0210601f $X=1.16 $Y=0.465 $X2=0
+ $Y2=0
cc_372 N_A_67_199#_c_235_p N_VGND_c_2046_n 0.0707535f $X=1.995 $Y=0.36 $X2=0
+ $Y2=0
cc_373 N_A_67_199#_c_212_n N_VGND_c_2046_n 0.0554858f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_374 N_A_67_199#_M1018_d N_VGND_c_2049_n 0.00438671f $X=1.025 $Y=0.235 $X2=0
+ $Y2=0
cc_375 N_A_67_199#_M1028_s N_VGND_c_2049_n 0.00202171f $X=3.18 $Y=0.235 $X2=0
+ $Y2=0
cc_376 N_A_67_199#_c_210_n N_VGND_c_2049_n 0.00127085f $X=0.695 $Y=1.325 $X2=0
+ $Y2=0
cc_377 N_A_67_199#_c_211_n N_VGND_c_2049_n 0.00458421f $X=0.995 $Y=0.82 $X2=0
+ $Y2=0
cc_378 N_A_67_199#_c_225_p N_VGND_c_2049_n 0.0124843f $X=1.16 $Y=0.465 $X2=0
+ $Y2=0
cc_379 N_A_67_199#_c_235_p N_VGND_c_2049_n 0.022547f $X=1.995 $Y=0.36 $X2=0
+ $Y2=0
cc_380 N_A_67_199#_c_212_n N_VGND_c_2049_n 0.0150136f $X=2.515 $Y=0.34 $X2=0
+ $Y2=0
cc_381 N_A_67_199#_c_214_n N_VGND_c_2049_n 0.0106925f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_382 N_A_67_199#_c_210_n N_VGND_c_2050_n 3.07438e-19 $X=0.695 $Y=1.325 $X2=0
+ $Y2=0
cc_383 N_A_67_199#_c_214_n N_VGND_c_2050_n 0.00541359f $X=0.5 $Y=0.995 $X2=0
+ $Y2=0
cc_384 A N_B_c_442_n 6.60282e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_385 N_A_c_400_n N_B_c_442_n 0.0214042f $X=1.175 $Y=1.16 $X2=0 $Y2=0
cc_386 N_A_c_398_n B 0.00226237f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_387 A B 0.0159767f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_388 N_A_c_400_n B 0.00331525f $X=1.175 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_c_398_n N_B_c_450_n 0.00127453f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_390 N_A_M1010_g N_A_27_47#_c_1441_n 5.78297e-19 $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_391 N_A_c_398_n N_A_27_47#_c_1434_n 5.98586e-19 $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_392 N_A_M1010_g N_A_27_47#_c_1456_n 0.0104009f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A_M1010_g N_A_27_47#_c_1463_n 0.0075453f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A_M1010_g N_A_27_47#_c_1503_n 0.00814033f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_395 N_A_M1010_g N_A_27_47#_c_1444_n 0.00103455f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_396 N_A_M1010_g N_A_27_47#_c_1447_n 0.00194926f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A_M1010_g N_VPWR_c_1602_n 0.0059862f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_398 N_A_M1010_g N_VPWR_c_1603_n 0.00390371f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_399 N_A_M1010_g N_VPWR_c_1601_n 0.00710619f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A_c_398_n N_VGND_c_2040_n 0.00384648f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_c_398_n N_VGND_c_2046_n 0.00422898f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_402 N_A_c_398_n N_VGND_c_2049_n 0.0072906f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_403 N_B_c_440_n N_A_489_21#_c_598_n 0.0265904f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_404 N_B_c_449_n N_A_489_21#_c_598_n 0.00401801f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_405 N_B_M1027_g N_A_489_21#_M1003_g 0.0265904f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_406 N_B_c_445_n N_A_489_21#_c_599_n 0.0137472f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_407 N_B_M1011_g N_A_489_21#_M1020_g 0.0289737f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_408 N_B_M1004_g N_A_489_21#_M1006_g 0.0356525f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_409 N_B_c_443_n N_A_489_21#_c_600_n 0.0265904f $X=2.095 $Y=1.16 $X2=0 $Y2=0
cc_410 N_B_c_449_n N_A_489_21#_c_601_n 0.00601333f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_411 N_B_c_444_n N_A_489_21#_c_602_n 0.0129182f $X=4.27 $Y=1.16 $X2=0 $Y2=0
cc_412 N_B_c_441_n N_A_489_21#_c_603_n 0.00490819f $X=5.125 $Y=0.995 $X2=0 $Y2=0
cc_413 N_B_c_445_n N_A_489_21#_c_603_n 0.00367982f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_414 N_B_c_451_n N_A_489_21#_c_603_n 0.00665271f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_415 N_B_c_452_n N_A_489_21#_c_603_n 0.0126697f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_416 N_B_c_447_n N_A_489_21#_c_604_n 0.00546111f $X=5.125 $Y=1.16 $X2=0 $Y2=0
cc_417 N_B_c_447_n N_A_489_21#_c_605_n 0.021509f $X=5.125 $Y=1.16 $X2=0 $Y2=0
cc_418 N_B_c_443_n N_A_489_21#_c_628_n 2.01375e-19 $X=2.095 $Y=1.16 $X2=0 $Y2=0
cc_419 N_B_c_449_n N_A_489_21#_c_628_n 0.00277067f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_420 N_B_M1011_g N_A_489_21#_c_615_n 0.0065988f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_421 N_B_c_444_n N_A_489_21#_c_615_n 0.00339751f $X=4.27 $Y=1.16 $X2=0 $Y2=0
cc_422 N_B_c_452_n N_A_489_21#_c_615_n 0.0035358f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_423 N_B_M1011_g N_A_489_21#_c_618_n 0.00800906f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_424 N_B_M1004_g N_A_489_21#_c_618_n 0.0147854f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_425 N_B_c_446_n N_A_489_21#_c_618_n 0.0274104f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_426 N_B_c_447_n N_A_489_21#_c_618_n 0.00995875f $X=5.125 $Y=1.16 $X2=0 $Y2=0
cc_427 N_B_c_452_n N_A_489_21#_c_618_n 0.0125603f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_428 N_B_c_441_n N_A_489_21#_c_606_n 0.0157995f $X=5.125 $Y=0.995 $X2=0 $Y2=0
cc_429 N_B_c_449_n N_A_434_49#_M1005_d 4.43088e-19 $X=4.225 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_430 N_B_c_440_n N_A_434_49#_c_779_n 0.00828913f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_431 B N_A_434_49#_c_779_n 0.0063676f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_432 N_B_c_449_n N_A_434_49#_c_779_n 0.0140059f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_433 N_B_c_450_n N_A_434_49#_c_779_n 0.00128472f $X=1.755 $Y=0.85 $X2=0 $Y2=0
cc_434 N_B_c_440_n N_A_434_49#_c_758_n 0.00428791f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_435 N_B_c_442_n N_A_434_49#_c_758_n 0.0032583f $X=2.02 $Y=1.16 $X2=0 $Y2=0
cc_436 N_B_c_443_n N_A_434_49#_c_758_n 0.00349007f $X=2.095 $Y=1.16 $X2=0 $Y2=0
cc_437 B N_A_434_49#_c_758_n 0.0208669f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_438 N_B_c_449_n N_A_434_49#_c_758_n 0.00906427f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_439 N_B_c_450_n N_A_434_49#_c_758_n 0.00128381f $X=1.755 $Y=0.85 $X2=0 $Y2=0
cc_440 N_B_M1027_g N_A_434_49#_c_770_n 0.00319381f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_441 N_B_c_444_n N_A_434_49#_c_759_n 0.00274495f $X=4.27 $Y=1.16 $X2=0 $Y2=0
cc_442 N_B_c_446_n N_A_434_49#_c_759_n 0.0136654f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_443 N_B_c_449_n N_A_434_49#_c_759_n 0.156786f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_444 N_B_c_451_n N_A_434_49#_c_759_n 0.0253176f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_445 N_B_c_452_n N_A_434_49#_c_759_n 0.0128416f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_446 N_B_c_442_n N_A_434_49#_c_788_n 0.00265654f $X=2.02 $Y=1.16 $X2=0 $Y2=0
cc_447 B N_A_434_49#_c_788_n 0.00635599f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_448 N_B_c_449_n N_A_434_49#_c_788_n 0.0255037f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_449 N_B_M1027_g N_A_434_49#_c_762_n 0.00450435f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_450 N_B_c_442_n N_A_434_49#_c_762_n 0.00304094f $X=2.02 $Y=1.16 $X2=0 $Y2=0
cc_451 N_B_c_443_n N_A_434_49#_c_762_n 0.00406409f $X=2.095 $Y=1.16 $X2=0 $Y2=0
cc_452 N_B_c_449_n N_A_721_47#_M1028_d 0.00183087f $X=4.225 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_453 N_B_M1011_g N_A_721_47#_c_960_n 0.0145753f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_454 N_B_c_452_n N_A_721_47#_c_960_n 2.10079e-19 $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_455 N_B_M1011_g N_A_721_47#_c_961_n 0.0118658f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_456 N_B_M1004_g N_A_721_47#_c_961_n 0.00597424f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_457 N_B_c_444_n N_A_721_47#_c_952_n 0.00599801f $X=4.27 $Y=1.16 $X2=0 $Y2=0
cc_458 N_B_c_445_n N_A_721_47#_c_952_n 0.00115759f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_459 N_B_c_449_n N_A_721_47#_c_952_n 0.010847f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_460 N_B_c_451_n N_A_721_47#_c_952_n 0.00226876f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_461 N_B_c_452_n N_A_721_47#_c_952_n 0.0280077f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_462 N_B_M1011_g N_A_721_47#_c_976_n 0.00307394f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_463 N_B_M1004_g N_A_721_47#_c_976_n 0.00787832f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_464 N_B_M1004_g N_A_721_47#_c_991_n 0.00986772f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_465 N_B_M1004_g N_A_721_47#_c_977_n 0.00369168f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_466 N_B_c_446_n N_A_721_47#_c_977_n 4.43504e-19 $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_467 N_B_c_444_n N_A_721_47#_c_954_n 0.00609207f $X=4.27 $Y=1.16 $X2=0 $Y2=0
cc_468 N_B_c_449_n N_A_721_47#_c_954_n 0.00129243f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_469 N_B_c_452_n N_A_721_47#_c_954_n 0.0115417f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_470 N_B_c_451_n N_A_27_47#_M1012_d 0.00177119f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_471 N_B_c_452_n N_A_27_47#_M1012_d 0.00459504f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_472 N_B_M1027_g N_A_27_47#_c_1442_n 0.0125333f $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_473 N_B_c_449_n N_A_27_47#_c_1435_n 0.0109361f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_474 N_B_c_444_n N_A_27_47#_c_1436_n 3.10296e-19 $X=4.27 $Y=1.16 $X2=0 $Y2=0
cc_475 N_B_c_445_n N_A_27_47#_c_1477_n 0.00260871f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_476 N_B_c_449_n N_A_27_47#_c_1439_n 0.0356614f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_477 N_B_M1011_g N_A_27_47#_c_1448_n 2.74497e-19 $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_478 N_B_c_441_n N_A_27_47#_c_1440_n 0.0037945f $X=5.125 $Y=0.995 $X2=0 $Y2=0
cc_479 N_B_c_445_n N_A_27_47#_c_1440_n 0.00198465f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_480 N_B_c_446_n N_A_27_47#_c_1440_n 0.0026102f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_481 N_B_c_451_n N_A_27_47#_c_1440_n 0.00164354f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_482 N_B_c_452_n N_A_27_47#_c_1440_n 0.0137147f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_483 N_B_c_444_n N_A_27_47#_c_1519_n 2.49317e-19 $X=4.27 $Y=1.16 $X2=0 $Y2=0
cc_484 N_B_c_445_n N_A_27_47#_c_1519_n 0.00813469f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_485 N_B_c_449_n N_A_27_47#_c_1519_n 0.008106f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_486 N_B_c_451_n N_A_27_47#_c_1519_n 3.07703e-19 $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_487 N_B_M1027_g N_VPWR_c_1603_n 9.44495e-19 $X=2.095 $Y=1.905 $X2=0 $Y2=0
cc_488 N_B_M1011_g N_VPWR_c_1603_n 0.00336115f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_489 N_B_M1004_g N_VPWR_c_1603_n 0.00421091f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_490 N_B_M1004_g N_VPWR_c_1604_n 0.00556491f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_491 N_B_M1011_g N_VPWR_c_1601_n 0.00685129f $X=4.07 $Y=2.03 $X2=0 $Y2=0
cc_492 N_B_M1004_g N_VPWR_c_1601_n 0.00738011f $X=5.125 $Y=1.985 $X2=0 $Y2=0
cc_493 N_B_M1004_g N_A_1142_49#_c_1729_n 5.46172e-19 $X=5.125 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_B_c_441_n N_VGND_c_2041_n 0.0150187f $X=5.125 $Y=0.995 $X2=0 $Y2=0
cc_495 N_B_c_440_n N_VGND_c_2046_n 0.00357877f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_496 N_B_c_441_n N_VGND_c_2046_n 0.00505556f $X=5.125 $Y=0.995 $X2=0 $Y2=0
cc_497 N_B_c_445_n N_VGND_c_2046_n 0.00351226f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_498 N_B_c_440_n N_VGND_c_2049_n 0.00662925f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_499 N_B_c_441_n N_VGND_c_2049_n 0.00995901f $X=5.125 $Y=0.995 $X2=0 $Y2=0
cc_500 N_B_c_445_n N_VGND_c_2049_n 0.00686244f $X=4.127 $Y=0.995 $X2=0 $Y2=0
cc_501 N_B_c_449_n N_VGND_c_2049_n 0.116256f $X=4.225 $Y=0.85 $X2=0 $Y2=0
cc_502 N_B_c_450_n N_VGND_c_2049_n 0.0149427f $X=1.755 $Y=0.85 $X2=0 $Y2=0
cc_503 N_B_c_451_n N_VGND_c_2049_n 0.0148223f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_504 N_A_489_21#_c_598_n N_A_434_49#_c_758_n 0.00310513f $X=2.52 $Y=0.995
+ $X2=0 $Y2=0
cc_505 N_A_489_21#_c_628_n N_A_434_49#_c_758_n 0.00827314f $X=2.805 $Y=1.16
+ $X2=0 $Y2=0
cc_506 N_A_489_21#_M1003_g N_A_434_49#_c_770_n 0.00310513f $X=2.52 $Y=1.905
+ $X2=0 $Y2=0
cc_507 N_A_489_21#_c_616_n N_A_434_49#_c_770_n 0.00624624f $X=3.18 $Y=1.53 $X2=0
+ $Y2=0
cc_508 N_A_489_21#_c_600_n N_A_434_49#_c_759_n 0.00500331f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_509 N_A_489_21#_c_601_n N_A_434_49#_c_759_n 0.00361395f $X=3.455 $Y=1.16
+ $X2=0 $Y2=0
cc_510 N_A_489_21#_c_602_n N_A_434_49#_c_759_n 0.00442392f $X=3.557 $Y=1.16
+ $X2=0 $Y2=0
cc_511 N_A_489_21#_c_604_n N_A_434_49#_c_759_n 0.0383848f $X=5.545 $Y=1.16 $X2=0
+ $Y2=0
cc_512 N_A_489_21#_c_605_n N_A_434_49#_c_759_n 0.004742f $X=5.545 $Y=1.16 $X2=0
+ $Y2=0
cc_513 N_A_489_21#_c_628_n N_A_434_49#_c_759_n 0.0190202f $X=2.805 $Y=1.16 $X2=0
+ $Y2=0
cc_514 N_A_489_21#_c_615_n N_A_434_49#_c_759_n 0.120229f $X=4.7 $Y=1.53 $X2=0
+ $Y2=0
cc_515 N_A_489_21#_c_616_n N_A_434_49#_c_759_n 0.0258328f $X=3.18 $Y=1.53 $X2=0
+ $Y2=0
cc_516 N_A_489_21#_c_675_p N_A_434_49#_c_759_n 0.025437f $X=4.845 $Y=1.53 $X2=0
+ $Y2=0
cc_517 N_A_489_21#_c_618_n N_A_434_49#_c_759_n 0.0394641f $X=4.845 $Y=1.53 $X2=0
+ $Y2=0
cc_518 N_A_489_21#_c_628_n N_A_434_49#_c_788_n 2.50543e-19 $X=2.805 $Y=1.16
+ $X2=0 $Y2=0
cc_519 N_A_489_21#_c_600_n N_A_434_49#_c_762_n 0.00310513f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_520 N_A_489_21#_c_628_n N_A_434_49#_c_762_n 5.67894e-19 $X=2.805 $Y=1.16
+ $X2=0 $Y2=0
cc_521 N_A_489_21#_c_617_n N_A_434_49#_c_762_n 0.00736909f $X=3.035 $Y=1.53
+ $X2=0 $Y2=0
cc_522 N_A_489_21#_c_606_n N_A_434_49#_c_763_n 0.00149902f $X=5.56 $Y=0.995
+ $X2=0 $Y2=0
cc_523 N_A_489_21#_c_605_n N_A_434_49#_c_765_n 0.00665199f $X=5.545 $Y=1.16
+ $X2=0 $Y2=0
cc_524 N_A_489_21#_c_615_n N_A_721_47#_M1020_d 8.14763e-19 $X=4.7 $Y=1.53 $X2=0
+ $Y2=0
cc_525 N_A_489_21#_c_602_n N_A_721_47#_c_960_n 0.00386403f $X=3.557 $Y=1.16
+ $X2=0 $Y2=0
cc_526 N_A_489_21#_c_615_n N_A_721_47#_c_960_n 0.0131883f $X=4.7 $Y=1.53 $X2=0
+ $Y2=0
cc_527 N_A_489_21#_M1004_s N_A_721_47#_c_961_n 0.00318137f $X=4.79 $Y=1.485
+ $X2=0 $Y2=0
cc_528 N_A_489_21#_c_618_n N_A_721_47#_c_961_n 0.00422939f $X=4.845 $Y=1.53
+ $X2=0 $Y2=0
cc_529 N_A_489_21#_M1020_g N_A_721_47#_c_962_n 0.0013897f $X=3.585 $Y=1.905
+ $X2=0 $Y2=0
cc_530 N_A_489_21#_c_599_n N_A_721_47#_c_952_n 0.00144563f $X=3.53 $Y=0.995
+ $X2=0 $Y2=0
cc_531 N_A_489_21#_c_602_n N_A_721_47#_c_952_n 0.00134715f $X=3.557 $Y=1.16
+ $X2=0 $Y2=0
cc_532 N_A_489_21#_M1004_s N_A_721_47#_c_976_n 0.0045681f $X=4.79 $Y=1.485 $X2=0
+ $Y2=0
cc_533 N_A_489_21#_M1006_g N_A_721_47#_c_976_n 5.30718e-19 $X=5.635 $Y=1.985
+ $X2=0 $Y2=0
cc_534 N_A_489_21#_M1006_g N_A_721_47#_c_991_n 0.0144138f $X=5.635 $Y=1.985
+ $X2=0 $Y2=0
cc_535 N_A_489_21#_c_604_n N_A_721_47#_c_991_n 0.0121036f $X=5.545 $Y=1.16 $X2=0
+ $Y2=0
cc_536 N_A_489_21#_c_605_n N_A_721_47#_c_991_n 0.00229431f $X=5.545 $Y=1.16
+ $X2=0 $Y2=0
cc_537 N_A_489_21#_c_618_n N_A_721_47#_c_991_n 0.00796435f $X=4.845 $Y=1.53
+ $X2=0 $Y2=0
cc_538 N_A_489_21#_M1004_s N_A_721_47#_c_977_n 0.00458918f $X=4.79 $Y=1.485
+ $X2=0 $Y2=0
cc_539 N_A_489_21#_c_675_p N_A_721_47#_c_977_n 0.00119591f $X=4.845 $Y=1.53
+ $X2=0 $Y2=0
cc_540 N_A_489_21#_c_618_n N_A_721_47#_c_977_n 0.0157891f $X=4.845 $Y=1.53 $X2=0
+ $Y2=0
cc_541 N_A_489_21#_M1006_g N_A_721_47#_c_1014_n 0.00743023f $X=5.635 $Y=1.985
+ $X2=0 $Y2=0
cc_542 N_A_489_21#_M1006_g N_A_721_47#_c_1015_n 0.00383087f $X=5.635 $Y=1.985
+ $X2=0 $Y2=0
cc_543 N_A_489_21#_c_602_n N_A_721_47#_c_954_n 0.0016475f $X=3.557 $Y=1.16 $X2=0
+ $Y2=0
cc_544 N_A_489_21#_c_615_n N_A_721_47#_c_954_n 0.00496925f $X=4.7 $Y=1.53 $X2=0
+ $Y2=0
cc_545 N_A_489_21#_c_615_n N_A_27_47#_M1020_s 0.00130271f $X=4.7 $Y=1.53 $X2=0
+ $Y2=0
cc_546 N_A_489_21#_c_616_n N_A_27_47#_M1020_s 4.85103e-19 $X=3.18 $Y=1.53 $X2=0
+ $Y2=0
cc_547 N_A_489_21#_M1003_g N_A_27_47#_c_1442_n 0.0127243f $X=2.52 $Y=1.905 $X2=0
+ $Y2=0
cc_548 N_A_489_21#_c_598_n N_A_27_47#_c_1435_n 6.16041e-19 $X=2.52 $Y=0.995
+ $X2=0 $Y2=0
cc_549 N_A_489_21#_c_601_n N_A_27_47#_c_1435_n 0.00522283f $X=3.455 $Y=1.16
+ $X2=0 $Y2=0
cc_550 N_A_489_21#_c_628_n N_A_27_47#_c_1435_n 0.0165044f $X=2.805 $Y=1.16 $X2=0
+ $Y2=0
cc_551 N_A_489_21#_c_598_n N_A_27_47#_c_1436_n 0.00137727f $X=2.52 $Y=0.995
+ $X2=0 $Y2=0
cc_552 N_A_489_21#_M1003_g N_A_27_47#_c_1436_n 0.00334557f $X=2.52 $Y=1.905
+ $X2=0 $Y2=0
cc_553 N_A_489_21#_c_599_n N_A_27_47#_c_1436_n 0.00224671f $X=3.53 $Y=0.995
+ $X2=0 $Y2=0
cc_554 N_A_489_21#_M1020_g N_A_27_47#_c_1436_n 0.00940077f $X=3.585 $Y=1.905
+ $X2=0 $Y2=0
cc_555 N_A_489_21#_c_601_n N_A_27_47#_c_1436_n 0.0158901f $X=3.455 $Y=1.16 $X2=0
+ $Y2=0
cc_556 N_A_489_21#_c_602_n N_A_27_47#_c_1436_n 0.00407852f $X=3.557 $Y=1.16
+ $X2=0 $Y2=0
cc_557 N_A_489_21#_c_628_n N_A_27_47#_c_1436_n 0.0122547f $X=2.805 $Y=1.16 $X2=0
+ $Y2=0
cc_558 N_A_489_21#_c_615_n N_A_27_47#_c_1436_n 0.0111716f $X=4.7 $Y=1.53 $X2=0
+ $Y2=0
cc_559 N_A_489_21#_c_616_n N_A_27_47#_c_1436_n 0.00339232f $X=3.18 $Y=1.53 $X2=0
+ $Y2=0
cc_560 N_A_489_21#_c_617_n N_A_27_47#_c_1436_n 0.024478f $X=3.035 $Y=1.53 $X2=0
+ $Y2=0
cc_561 N_A_489_21#_c_599_n N_A_27_47#_c_1477_n 0.0105455f $X=3.53 $Y=0.995 $X2=0
+ $Y2=0
cc_562 N_A_489_21#_c_599_n N_A_27_47#_c_1478_n 0.00548278f $X=3.53 $Y=0.995
+ $X2=0 $Y2=0
cc_563 N_A_489_21#_c_598_n N_A_27_47#_c_1439_n 2.62007e-19 $X=2.52 $Y=0.995
+ $X2=0 $Y2=0
cc_564 N_A_489_21#_c_599_n N_A_27_47#_c_1439_n 0.0153035f $X=3.53 $Y=0.995 $X2=0
+ $Y2=0
cc_565 N_A_489_21#_c_601_n N_A_27_47#_c_1439_n 0.0125787f $X=3.455 $Y=1.16 $X2=0
+ $Y2=0
cc_566 N_A_489_21#_c_602_n N_A_27_47#_c_1439_n 0.00294337f $X=3.557 $Y=1.16
+ $X2=0 $Y2=0
cc_567 N_A_489_21#_c_628_n N_A_27_47#_c_1439_n 0.0140232f $X=2.805 $Y=1.16 $X2=0
+ $Y2=0
cc_568 N_A_489_21#_M1003_g N_A_27_47#_c_1448_n 0.00351169f $X=2.52 $Y=1.905
+ $X2=0 $Y2=0
cc_569 N_A_489_21#_M1020_g N_A_27_47#_c_1448_n 0.00554289f $X=3.585 $Y=1.905
+ $X2=0 $Y2=0
cc_570 N_A_489_21#_M1003_g N_VPWR_c_1603_n 9.44495e-19 $X=2.52 $Y=1.905 $X2=0
+ $Y2=0
cc_571 N_A_489_21#_M1020_g N_VPWR_c_1603_n 0.00544188f $X=3.585 $Y=1.905 $X2=0
+ $Y2=0
cc_572 N_A_489_21#_M1006_g N_VPWR_c_1604_n 0.00902456f $X=5.635 $Y=1.985 $X2=0
+ $Y2=0
cc_573 N_A_489_21#_M1006_g N_VPWR_c_1608_n 0.00341689f $X=5.635 $Y=1.985 $X2=0
+ $Y2=0
cc_574 N_A_489_21#_M1004_s N_VPWR_c_1601_n 0.00210267f $X=4.79 $Y=1.485 $X2=0
+ $Y2=0
cc_575 N_A_489_21#_M1020_g N_VPWR_c_1601_n 0.00369216f $X=3.585 $Y=1.905 $X2=0
+ $Y2=0
cc_576 N_A_489_21#_M1006_g N_VPWR_c_1601_n 0.00540327f $X=5.635 $Y=1.985 $X2=0
+ $Y2=0
cc_577 N_A_489_21#_M1006_g N_A_1142_49#_c_1729_n 0.00573282f $X=5.635 $Y=1.985
+ $X2=0 $Y2=0
cc_578 N_A_489_21#_c_604_n N_A_1142_49#_c_1729_n 0.0242985f $X=5.545 $Y=1.16
+ $X2=0 $Y2=0
cc_579 N_A_489_21#_c_618_n N_A_1142_49#_c_1729_n 0.0111642f $X=4.845 $Y=1.53
+ $X2=0 $Y2=0
cc_580 N_A_489_21#_c_606_n N_A_1142_49#_c_1729_n 0.0122311f $X=5.56 $Y=0.995
+ $X2=0 $Y2=0
cc_581 N_A_489_21#_M1006_g N_A_1142_49#_c_1738_n 0.00281901f $X=5.635 $Y=1.985
+ $X2=0 $Y2=0
cc_582 N_A_489_21#_c_606_n N_A_1142_49#_c_1739_n 0.00655158f $X=5.56 $Y=0.995
+ $X2=0 $Y2=0
cc_583 N_A_489_21#_M1006_g N_A_1142_49#_c_1740_n 8.4745e-19 $X=5.635 $Y=1.985
+ $X2=0 $Y2=0
cc_584 N_A_489_21#_c_606_n N_A_1251_49#_c_1838_n 0.00354077f $X=5.56 $Y=0.995
+ $X2=0 $Y2=0
cc_585 N_A_489_21#_c_604_n N_VGND_c_2041_n 0.0212879f $X=5.545 $Y=1.16 $X2=0
+ $Y2=0
cc_586 N_A_489_21#_c_605_n N_VGND_c_2041_n 0.00226374f $X=5.545 $Y=1.16 $X2=0
+ $Y2=0
cc_587 N_A_489_21#_c_606_n N_VGND_c_2041_n 0.00593607f $X=5.56 $Y=0.995 $X2=0
+ $Y2=0
cc_588 N_A_489_21#_c_606_n N_VGND_c_2044_n 0.00536492f $X=5.56 $Y=0.995 $X2=0
+ $Y2=0
cc_589 N_A_489_21#_c_598_n N_VGND_c_2046_n 0.00357766f $X=2.52 $Y=0.995 $X2=0
+ $Y2=0
cc_590 N_A_489_21#_c_599_n N_VGND_c_2046_n 0.0041652f $X=3.53 $Y=0.995 $X2=0
+ $Y2=0
cc_591 N_A_489_21#_c_603_n N_VGND_c_2046_n 0.00429232f $X=4.915 $Y=0.74 $X2=0
+ $Y2=0
cc_592 N_A_489_21#_M1015_s N_VGND_c_2049_n 0.0051911f $X=4.79 $Y=0.605 $X2=0
+ $Y2=0
cc_593 N_A_489_21#_c_598_n N_VGND_c_2049_n 0.00662918f $X=2.52 $Y=0.995 $X2=0
+ $Y2=0
cc_594 N_A_489_21#_c_599_n N_VGND_c_2049_n 0.00747617f $X=3.53 $Y=0.995 $X2=0
+ $Y2=0
cc_595 N_A_489_21#_c_603_n N_VGND_c_2049_n 0.00553188f $X=4.915 $Y=0.74 $X2=0
+ $Y2=0
cc_596 N_A_489_21#_c_606_n N_VGND_c_2049_n 0.0110279f $X=5.56 $Y=0.995 $X2=0
+ $Y2=0
cc_597 N_A_434_49#_M1030_g N_A_721_47#_M1009_g 0.0371801f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_598 N_A_434_49#_c_756_n N_A_721_47#_c_948_n 0.0260017f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_599 N_A_434_49#_M1023_g N_A_721_47#_c_956_n 0.0257608f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_600 N_A_434_49#_c_760_n N_A_721_47#_c_956_n 0.00329127f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_601 N_A_434_49#_c_766_n N_A_721_47#_c_956_n 0.00395049f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_602 N_A_434_49#_c_760_n N_A_721_47#_c_949_n 0.0101614f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_603 N_A_434_49#_c_765_n N_A_721_47#_c_949_n 0.0214585f $X=6.63 $Y=1.16 $X2=0
+ $Y2=0
cc_604 N_A_434_49#_M1023_g N_A_721_47#_c_950_n 2.73351e-19 $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_605 N_A_434_49#_c_760_n N_A_721_47#_c_950_n 0.0265382f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_606 N_A_434_49#_c_766_n N_A_721_47#_c_950_n 0.0190701f $X=8.935 $Y=1.16 $X2=0
+ $Y2=0
cc_607 N_A_434_49#_c_757_n N_A_721_47#_c_951_n 0.0149133f $X=8.6 $Y=0.96 $X2=0
+ $Y2=0
cc_608 N_A_434_49#_c_759_n N_A_721_47#_c_960_n 2.63373e-19 $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_609 N_A_434_49#_c_759_n N_A_721_47#_c_952_n 0.00409089f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_610 N_A_434_49#_M1030_g N_A_721_47#_c_1014_n 0.00350227f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_611 N_A_434_49#_M1030_g N_A_721_47#_c_963_n 0.0119433f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_612 N_A_434_49#_c_760_n N_A_721_47#_c_953_n 0.0164128f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_613 N_A_434_49#_c_759_n N_A_721_47#_c_954_n 0.0130466f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_614 N_A_434_49#_c_760_n N_A_721_47#_c_967_n 0.00362829f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_615 N_A_434_49#_M1023_g N_A_1636_315#_c_1145_n 0.0146628f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_616 N_A_434_49#_c_766_n N_A_1636_315#_c_1152_n 0.00954492f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_617 N_A_434_49#_c_767_n N_A_1636_315#_c_1152_n 0.00925003f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_618 N_A_434_49#_c_757_n N_A_1636_315#_c_1138_n 0.00311679f $X=8.6 $Y=0.96
+ $X2=0 $Y2=0
cc_619 N_A_434_49#_M1023_g N_A_1636_315#_c_1138_n 0.0117267f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_620 N_A_434_49#_c_764_n N_A_1636_315#_c_1138_n 0.00772348f $X=8.985 $Y=1.19
+ $X2=0 $Y2=0
cc_621 N_A_434_49#_c_766_n N_A_1636_315#_c_1138_n 0.00368376f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_622 N_A_434_49#_c_767_n N_A_1636_315#_c_1138_n 0.0216383f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_623 N_A_434_49#_M1023_g N_A_1636_315#_c_1159_n 0.00700327f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_624 N_A_434_49#_M1023_g N_A_1636_315#_c_1160_n 0.00358172f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_625 N_A_434_49#_c_757_n N_A_1647_49#_c_1328_n 0.00160562f $X=8.6 $Y=0.96
+ $X2=0 $Y2=0
cc_626 N_A_434_49#_M1023_g N_A_1647_49#_c_1328_n 0.00116952f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_627 N_A_434_49#_c_760_n N_A_1647_49#_c_1328_n 0.0124451f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_628 N_A_434_49#_c_764_n N_A_1647_49#_c_1328_n 6.1128e-19 $X=8.985 $Y=1.19
+ $X2=0 $Y2=0
cc_629 N_A_434_49#_c_766_n N_A_1647_49#_c_1328_n 0.00695756f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_630 N_A_434_49#_c_767_n N_A_1647_49#_c_1328_n 0.0140666f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_631 N_A_434_49#_c_757_n N_A_1647_49#_c_1329_n 0.00655441f $X=8.6 $Y=0.96
+ $X2=0 $Y2=0
cc_632 N_A_434_49#_c_760_n N_A_1647_49#_c_1329_n 0.001989f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_633 N_A_434_49#_M1023_g N_A_1647_49#_c_1335_n 0.0085344f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_634 N_A_434_49#_c_760_n N_A_1647_49#_c_1335_n 0.0140421f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_635 N_A_434_49#_c_764_n N_A_1647_49#_c_1335_n 0.0265246f $X=8.985 $Y=1.19
+ $X2=0 $Y2=0
cc_636 N_A_434_49#_c_766_n N_A_1647_49#_c_1335_n 0.00188533f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_637 N_A_434_49#_c_767_n N_A_1647_49#_c_1335_n 0.00498177f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_638 N_A_434_49#_M1023_g N_A_1647_49#_c_1336_n 4.4878e-19 $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_639 N_A_434_49#_c_760_n N_A_1647_49#_c_1336_n 0.026091f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_640 N_A_434_49#_M1023_g N_A_1647_49#_c_1340_n 0.0107283f $X=8.935 $Y=1.995
+ $X2=0 $Y2=0
cc_641 N_A_434_49#_c_760_n N_A_1647_49#_c_1340_n 0.0021315f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_642 N_A_434_49#_c_766_n N_A_1647_49#_c_1340_n 0.00780225f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_643 N_A_434_49#_c_767_n N_A_1647_49#_c_1340_n 0.00288506f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_644 N_A_434_49#_M1027_d N_A_27_47#_c_1442_n 0.00267395f $X=2.17 $Y=1.485
+ $X2=0 $Y2=0
cc_645 N_A_434_49#_c_770_n N_A_27_47#_c_1442_n 0.002595f $X=2.305 $Y=1.62 $X2=0
+ $Y2=0
cc_646 N_A_434_49#_c_779_n N_A_27_47#_c_1435_n 0.00265835f $X=2.187 $Y=0.877
+ $X2=0 $Y2=0
cc_647 N_A_434_49#_c_758_n N_A_27_47#_c_1435_n 0.0012144f $X=2.187 $Y=1.148
+ $X2=0 $Y2=0
cc_648 N_A_434_49#_c_759_n N_A_27_47#_c_1435_n 4.0994e-19 $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_649 N_A_434_49#_c_759_n N_A_27_47#_c_1436_n 0.0111296f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_650 N_A_434_49#_c_758_n N_A_27_47#_c_1439_n 3.9727e-19 $X=2.187 $Y=1.148
+ $X2=0 $Y2=0
cc_651 N_A_434_49#_c_759_n N_A_27_47#_c_1439_n 0.0116483f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_652 N_A_434_49#_M1030_g N_VPWR_c_1608_n 9.44495e-19 $X=6.575 $Y=1.905 $X2=0
+ $Y2=0
cc_653 N_A_434_49#_M1023_g N_VPWR_c_1608_n 0.00313972f $X=8.935 $Y=1.995 $X2=0
+ $Y2=0
cc_654 N_A_434_49#_M1023_g N_VPWR_c_1601_n 0.00519382f $X=8.935 $Y=1.995 $X2=0
+ $Y2=0
cc_655 N_A_434_49#_M1030_g N_A_1142_49#_c_1729_n 0.00356489f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_656 N_A_434_49#_c_759_n N_A_1142_49#_c_1729_n 0.0286752f $X=6.08 $Y=1.19
+ $X2=0 $Y2=0
cc_657 N_A_434_49#_c_761_n N_A_1142_49#_c_1729_n 0.00275249f $X=6.37 $Y=1.19
+ $X2=0 $Y2=0
cc_658 N_A_434_49#_c_765_n N_A_1142_49#_c_1729_n 9.64063e-19 $X=6.63 $Y=1.16
+ $X2=0 $Y2=0
cc_659 N_A_434_49#_M1030_g N_A_1142_49#_c_1745_n 0.00382305f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_660 N_A_434_49#_c_759_n N_A_1142_49#_c_1745_n 0.00437461f $X=6.08 $Y=1.19
+ $X2=0 $Y2=0
cc_661 N_A_434_49#_c_761_n N_A_1142_49#_c_1745_n 0.00433012f $X=6.37 $Y=1.19
+ $X2=0 $Y2=0
cc_662 N_A_434_49#_c_763_n N_A_1142_49#_c_1745_n 0.013108f $X=6.225 $Y=1.19
+ $X2=0 $Y2=0
cc_663 N_A_434_49#_c_765_n N_A_1142_49#_c_1745_n 0.00363059f $X=6.63 $Y=1.16
+ $X2=0 $Y2=0
cc_664 N_A_434_49#_M1030_g N_A_1142_49#_c_1738_n 0.00215498f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_665 N_A_434_49#_M1030_g N_A_1142_49#_c_1751_n 0.00931505f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_666 N_A_434_49#_c_760_n N_A_1142_49#_c_1730_n 0.0201739f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_667 N_A_434_49#_M1030_g N_A_1142_49#_c_1732_n 6.70022e-19 $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_668 N_A_434_49#_c_760_n N_A_1142_49#_c_1732_n 0.0101391f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_669 N_A_434_49#_c_756_n N_A_1142_49#_c_1739_n 0.00313733f $X=6.63 $Y=0.995
+ $X2=0 $Y2=0
cc_670 N_A_434_49#_c_759_n N_A_1142_49#_c_1739_n 0.00500613f $X=6.08 $Y=1.19
+ $X2=0 $Y2=0
cc_671 N_A_434_49#_c_763_n N_A_1142_49#_c_1739_n 0.0441632f $X=6.225 $Y=1.19
+ $X2=0 $Y2=0
cc_672 N_A_434_49#_M1030_g N_A_1142_49#_c_1740_n 0.00321587f $X=6.575 $Y=1.905
+ $X2=0 $Y2=0
cc_673 N_A_434_49#_c_763_n N_A_1142_49#_c_1740_n 0.00169815f $X=6.225 $Y=1.19
+ $X2=0 $Y2=0
cc_674 N_A_434_49#_c_765_n N_A_1142_49#_c_1740_n 0.00214523f $X=6.63 $Y=1.16
+ $X2=0 $Y2=0
cc_675 N_A_434_49#_M1030_g COUT 0.00635668f $X=6.575 $Y=1.905 $X2=0 $Y2=0
cc_676 N_A_434_49#_c_756_n COUT 0.00161643f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_677 N_A_434_49#_c_760_n COUT 0.0330527f $X=8.84 $Y=1.19 $X2=0 $Y2=0
cc_678 N_A_434_49#_c_761_n COUT 5.6439e-19 $X=6.37 $Y=1.19 $X2=0 $Y2=0
cc_679 N_A_434_49#_c_763_n COUT 0.0271315f $X=6.225 $Y=1.19 $X2=0 $Y2=0
cc_680 N_A_434_49#_c_765_n COUT 0.0101219f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_681 N_A_434_49#_M1030_g COUT 0.00293392f $X=6.575 $Y=1.905 $X2=0 $Y2=0
cc_682 N_A_434_49#_c_756_n N_COUT_c_1802_n 0.00522673f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_683 N_A_434_49#_c_760_n N_COUT_c_1802_n 0.002594f $X=8.84 $Y=1.19 $X2=0 $Y2=0
cc_684 N_A_434_49#_c_763_n N_COUT_c_1802_n 0.0129305f $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_685 N_A_434_49#_c_763_n N_A_1251_49#_M1031_s 0.00373082f $X=6.225 $Y=1.19
+ $X2=-0.19 $Y2=-0.24
cc_686 N_A_434_49#_c_756_n N_A_1251_49#_c_1829_n 0.00808644f $X=6.63 $Y=0.995
+ $X2=0 $Y2=0
cc_687 N_A_434_49#_c_756_n N_A_1251_49#_c_1838_n 0.00530807f $X=6.63 $Y=0.995
+ $X2=0 $Y2=0
cc_688 N_A_434_49#_c_760_n N_A_1251_49#_c_1838_n 0.00490782f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_689 N_A_434_49#_c_761_n N_A_1251_49#_c_1838_n 4.57094e-19 $X=6.37 $Y=1.19
+ $X2=0 $Y2=0
cc_690 N_A_434_49#_c_763_n N_A_1251_49#_c_1838_n 0.0132225f $X=6.225 $Y=1.19
+ $X2=0 $Y2=0
cc_691 N_A_434_49#_c_765_n N_A_1251_49#_c_1838_n 0.00400012f $X=6.63 $Y=1.16
+ $X2=0 $Y2=0
cc_692 N_A_434_49#_c_760_n N_A_1251_49#_c_1836_n 0.025635f $X=8.84 $Y=1.19 $X2=0
+ $Y2=0
cc_693 N_A_434_49#_c_757_n N_A_1251_49#_c_1830_n 0.00426885f $X=8.6 $Y=0.96
+ $X2=0 $Y2=0
cc_694 N_A_434_49#_c_760_n N_A_1251_49#_c_1830_n 0.0872966f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_695 N_A_434_49#_c_764_n N_A_1251_49#_c_1830_n 0.0266205f $X=8.985 $Y=1.19
+ $X2=0 $Y2=0
cc_696 N_A_434_49#_c_766_n N_A_1251_49#_c_1830_n 0.00672159f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_697 N_A_434_49#_c_767_n N_A_1251_49#_c_1830_n 0.00180356f $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_698 N_A_434_49#_c_760_n N_A_1251_49#_c_1831_n 0.0257857f $X=8.84 $Y=1.19
+ $X2=0 $Y2=0
cc_699 N_A_434_49#_c_757_n N_A_1565_49#_c_1963_n 0.0124254f $X=8.6 $Y=0.96 $X2=0
+ $Y2=0
cc_700 N_A_434_49#_c_766_n N_A_1565_49#_c_1963_n 9.39927e-19 $X=8.935 $Y=1.16
+ $X2=0 $Y2=0
cc_701 N_A_434_49#_c_759_n N_VGND_c_2041_n 0.00211029f $X=6.08 $Y=1.19 $X2=0
+ $Y2=0
cc_702 N_A_434_49#_c_756_n N_VGND_c_2044_n 0.00352679f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_703 N_A_434_49#_c_757_n N_VGND_c_2044_n 0.00357877f $X=8.6 $Y=0.96 $X2=0
+ $Y2=0
cc_704 N_A_434_49#_c_763_n N_VGND_c_2044_n 0.00189245f $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_705 N_A_434_49#_c_756_n N_VGND_c_2049_n 0.00646238f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_706 N_A_434_49#_c_757_n N_VGND_c_2049_n 0.00676309f $X=8.6 $Y=0.96 $X2=0
+ $Y2=0
cc_707 N_A_434_49#_c_763_n N_VGND_c_2049_n 0.00355378f $X=6.225 $Y=1.19 $X2=0
+ $Y2=0
cc_708 N_A_721_47#_c_950_n N_A_1636_315#_c_1161_n 0.00454307f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_709 N_A_721_47#_c_964_n N_A_1636_315#_c_1161_n 0.0180111f $X=7.865 $Y=2.295
+ $X2=0 $Y2=0
cc_710 N_A_721_47#_c_957_n N_A_1636_315#_c_1145_n 0.01147f $X=8.515 $Y=1.5 $X2=0
+ $Y2=0
cc_711 N_A_721_47#_c_963_n N_A_1636_315#_c_1146_n 0.0112831f $X=7.78 $Y=2.38
+ $X2=0 $Y2=0
cc_712 N_A_721_47#_c_956_n N_A_1647_49#_c_1328_n 0.0087759f $X=8.44 $Y=1.425
+ $X2=0 $Y2=0
cc_713 N_A_721_47#_c_951_n N_A_1647_49#_c_1328_n 0.00530648f $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_714 N_A_721_47#_c_953_n N_A_1647_49#_c_1328_n 0.0171951f $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_715 N_A_721_47#_c_956_n N_A_1647_49#_c_1329_n 0.00195876f $X=8.44 $Y=1.425
+ $X2=0 $Y2=0
cc_716 N_A_721_47#_c_951_n N_A_1647_49#_c_1329_n 0.00217451f $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_717 N_A_721_47#_c_953_n N_A_1647_49#_c_1336_n 0.00151468f $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_718 N_A_721_47#_c_956_n N_A_1647_49#_c_1340_n 0.00443311f $X=8.44 $Y=1.425
+ $X2=0 $Y2=0
cc_719 N_A_721_47#_c_957_n N_A_1647_49#_c_1340_n 0.0181141f $X=8.515 $Y=1.5
+ $X2=0 $Y2=0
cc_720 N_A_721_47#_c_964_n N_A_1647_49#_c_1340_n 0.00752892f $X=7.865 $Y=2.295
+ $X2=0 $Y2=0
cc_721 N_A_721_47#_c_953_n N_A_1647_49#_c_1340_n 0.011786f $X=7.95 $Y=1.16 $X2=0
+ $Y2=0
cc_722 N_A_721_47#_c_960_n N_A_27_47#_c_1436_n 0.0151785f $X=3.795 $Y=1.99 $X2=0
+ $Y2=0
cc_723 N_A_721_47#_c_952_n N_A_27_47#_c_1436_n 0.00750846f $X=3.985 $Y=0.76
+ $X2=0 $Y2=0
cc_724 N_A_721_47#_c_954_n N_A_27_47#_c_1436_n 0.00839475f $X=3.985 $Y=1.235
+ $X2=0 $Y2=0
cc_725 N_A_721_47#_M1028_d N_A_27_47#_c_1477_n 0.00378275f $X=3.605 $Y=0.235
+ $X2=0 $Y2=0
cc_726 N_A_721_47#_c_952_n N_A_27_47#_c_1477_n 0.0115352f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_727 N_A_721_47#_M1028_d N_A_27_47#_c_1478_n 6.64705e-19 $X=3.605 $Y=0.235
+ $X2=0 $Y2=0
cc_728 N_A_721_47#_M1028_d N_A_27_47#_c_1439_n 6.80925e-19 $X=3.605 $Y=0.235
+ $X2=0 $Y2=0
cc_729 N_A_721_47#_c_952_n N_A_27_47#_c_1439_n 0.0122849f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_730 N_A_721_47#_c_954_n N_A_27_47#_c_1439_n 0.00109524f $X=3.985 $Y=1.235
+ $X2=0 $Y2=0
cc_731 N_A_721_47#_c_962_n N_A_27_47#_c_1448_n 0.0119613f $X=3.88 $Y=2.375 $X2=0
+ $Y2=0
cc_732 N_A_721_47#_M1028_d N_A_27_47#_c_1519_n 0.00882466f $X=3.605 $Y=0.235
+ $X2=0 $Y2=0
cc_733 N_A_721_47#_c_952_n N_A_27_47#_c_1519_n 0.0114751f $X=3.985 $Y=0.76 $X2=0
+ $Y2=0
cc_734 N_A_721_47#_c_991_n N_VPWR_M1004_d 0.00699141f $X=5.825 $Y=1.98 $X2=0
+ $Y2=0
cc_735 N_A_721_47#_c_961_n N_VPWR_c_1603_n 0.0728111f $X=4.815 $Y=2.375 $X2=0
+ $Y2=0
cc_736 N_A_721_47#_c_962_n N_VPWR_c_1603_n 0.0118156f $X=3.88 $Y=2.375 $X2=0
+ $Y2=0
cc_737 N_A_721_47#_c_991_n N_VPWR_c_1603_n 0.00267364f $X=5.825 $Y=1.98 $X2=0
+ $Y2=0
cc_738 N_A_721_47#_c_961_n N_VPWR_c_1604_n 0.012593f $X=4.815 $Y=2.375 $X2=0
+ $Y2=0
cc_739 N_A_721_47#_c_976_n N_VPWR_c_1604_n 0.00373191f $X=4.94 $Y=2.29 $X2=0
+ $Y2=0
cc_740 N_A_721_47#_c_991_n N_VPWR_c_1604_n 0.0206205f $X=5.825 $Y=1.98 $X2=0
+ $Y2=0
cc_741 N_A_721_47#_c_1014_n N_VPWR_c_1604_n 0.003425f $X=5.91 $Y=2.295 $X2=0
+ $Y2=0
cc_742 N_A_721_47#_c_1015_n N_VPWR_c_1604_n 0.0109407f $X=5.995 $Y=2.38 $X2=0
+ $Y2=0
cc_743 N_A_721_47#_M1009_g N_VPWR_c_1608_n 9.44495e-19 $X=6.995 $Y=1.905 $X2=0
+ $Y2=0
cc_744 N_A_721_47#_c_957_n N_VPWR_c_1608_n 0.00313972f $X=8.515 $Y=1.5 $X2=0
+ $Y2=0
cc_745 N_A_721_47#_c_991_n N_VPWR_c_1608_n 0.00335963f $X=5.825 $Y=1.98 $X2=0
+ $Y2=0
cc_746 N_A_721_47#_c_963_n N_VPWR_c_1608_n 0.126769f $X=7.78 $Y=2.38 $X2=0 $Y2=0
cc_747 N_A_721_47#_c_1015_n N_VPWR_c_1608_n 0.0118015f $X=5.995 $Y=2.38 $X2=0
+ $Y2=0
cc_748 N_A_721_47#_c_957_n N_VPWR_c_1601_n 0.00519382f $X=8.515 $Y=1.5 $X2=0
+ $Y2=0
cc_749 N_A_721_47#_c_961_n N_VPWR_c_1601_n 0.0337884f $X=4.815 $Y=2.375 $X2=0
+ $Y2=0
cc_750 N_A_721_47#_c_962_n N_VPWR_c_1601_n 0.00311148f $X=3.88 $Y=2.375 $X2=0
+ $Y2=0
cc_751 N_A_721_47#_c_991_n N_VPWR_c_1601_n 0.0121802f $X=5.825 $Y=1.98 $X2=0
+ $Y2=0
cc_752 N_A_721_47#_c_963_n N_VPWR_c_1601_n 0.0730221f $X=7.78 $Y=2.38 $X2=0
+ $Y2=0
cc_753 N_A_721_47#_c_1015_n N_VPWR_c_1601_n 0.00651702f $X=5.995 $Y=2.38 $X2=0
+ $Y2=0
cc_754 N_A_721_47#_c_991_n N_A_1142_49#_M1006_d 0.00626813f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_755 N_A_721_47#_c_1014_n N_A_1142_49#_M1006_d 0.00716186f $X=5.91 $Y=2.295
+ $X2=0 $Y2=0
cc_756 N_A_721_47#_c_963_n N_A_1142_49#_M1006_d 0.0128212f $X=7.78 $Y=2.38 $X2=0
+ $Y2=0
cc_757 N_A_721_47#_c_1015_n N_A_1142_49#_M1006_d 0.00490995f $X=5.995 $Y=2.38
+ $X2=0 $Y2=0
cc_758 N_A_721_47#_c_991_n N_A_1142_49#_c_1729_n 0.0223447f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_759 N_A_721_47#_c_991_n N_A_1142_49#_c_1745_n 0.0019685f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_760 N_A_721_47#_c_963_n N_A_1142_49#_c_1745_n 0.00601442f $X=7.78 $Y=2.38
+ $X2=0 $Y2=0
cc_761 N_A_721_47#_M1009_g N_A_1142_49#_c_1751_n 0.01446f $X=6.995 $Y=1.905
+ $X2=0 $Y2=0
cc_762 N_A_721_47#_c_963_n N_A_1142_49#_c_1751_n 0.0083871f $X=7.78 $Y=2.38
+ $X2=0 $Y2=0
cc_763 N_A_721_47#_c_948_n N_A_1142_49#_c_1730_n 0.00664727f $X=7.055 $Y=0.995
+ $X2=0 $Y2=0
cc_764 N_A_721_47#_c_949_n N_A_1142_49#_c_1730_n 0.00505614f $X=7.025 $Y=1.16
+ $X2=0 $Y2=0
cc_765 N_A_721_47#_c_950_n N_A_1142_49#_c_1730_n 0.0117706f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_766 N_A_721_47#_M1009_g N_A_1142_49#_c_1732_n 0.0187858f $X=6.995 $Y=1.905
+ $X2=0 $Y2=0
cc_767 N_A_721_47#_c_949_n N_A_1142_49#_c_1732_n 0.00292034f $X=7.025 $Y=1.16
+ $X2=0 $Y2=0
cc_768 N_A_721_47#_c_950_n N_A_1142_49#_c_1732_n 0.00398638f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_769 N_A_721_47#_c_991_n N_A_1142_49#_c_1740_n 0.0130086f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_770 N_A_721_47#_c_1014_n N_A_1142_49#_c_1740_n 0.00414373f $X=5.91 $Y=2.295
+ $X2=0 $Y2=0
cc_771 N_A_721_47#_c_963_n N_A_1142_49#_c_1740_n 0.0448489f $X=7.78 $Y=2.38
+ $X2=0 $Y2=0
cc_772 N_A_721_47#_c_963_n N_COUT_M1030_d 0.00166235f $X=7.78 $Y=2.38 $X2=0
+ $Y2=0
cc_773 N_A_721_47#_c_948_n COUT 5.04756e-19 $X=7.055 $Y=0.995 $X2=0 $Y2=0
cc_774 N_A_721_47#_c_949_n COUT 0.00356487f $X=7.025 $Y=1.16 $X2=0 $Y2=0
cc_775 N_A_721_47#_c_948_n N_COUT_c_1802_n 2.94306e-19 $X=7.055 $Y=0.995 $X2=0
+ $Y2=0
cc_776 N_A_721_47#_c_949_n N_COUT_c_1802_n 2.47785e-19 $X=7.025 $Y=1.16 $X2=0
+ $Y2=0
cc_777 N_A_721_47#_c_963_n N_A_1251_49#_M1009_d 0.0189848f $X=7.78 $Y=2.38 $X2=0
+ $Y2=0
cc_778 N_A_721_47#_c_964_n N_A_1251_49#_M1009_d 0.0154561f $X=7.865 $Y=2.295
+ $X2=0 $Y2=0
cc_779 N_A_721_47#_c_953_n N_A_1251_49#_M1009_d 8.43292e-19 $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_780 N_A_721_47#_c_967_n N_A_1251_49#_M1009_d 0.00306849f $X=7.907 $Y=1.72
+ $X2=0 $Y2=0
cc_781 N_A_721_47#_c_948_n N_A_1251_49#_c_1829_n 0.0141786f $X=7.055 $Y=0.995
+ $X2=0 $Y2=0
cc_782 N_A_721_47#_c_949_n N_A_1251_49#_c_1829_n 8.79554e-19 $X=7.025 $Y=1.16
+ $X2=0 $Y2=0
cc_783 N_A_721_47#_c_950_n N_A_1251_49#_c_1829_n 0.00443758f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_784 N_A_721_47#_c_951_n N_A_1251_49#_c_1829_n 5.47211e-19 $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_785 N_A_721_47#_M1009_g N_A_1251_49#_c_1861_n 0.00301685f $X=6.995 $Y=1.905
+ $X2=0 $Y2=0
cc_786 N_A_721_47#_c_963_n N_A_1251_49#_c_1861_n 0.0128008f $X=7.78 $Y=2.38
+ $X2=0 $Y2=0
cc_787 N_A_721_47#_c_953_n N_A_1251_49#_c_1861_n 8.7702e-19 $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_788 N_A_721_47#_c_967_n N_A_1251_49#_c_1861_n 0.0336903f $X=7.907 $Y=1.72
+ $X2=0 $Y2=0
cc_789 N_A_721_47#_c_948_n N_A_1251_49#_c_1838_n 7.8676e-19 $X=7.055 $Y=0.995
+ $X2=0 $Y2=0
cc_790 N_A_721_47#_M1009_g N_A_1251_49#_c_1836_n 0.00105176f $X=6.995 $Y=1.905
+ $X2=0 $Y2=0
cc_791 N_A_721_47#_c_950_n N_A_1251_49#_c_1836_n 0.0229067f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_792 N_A_721_47#_c_953_n N_A_1251_49#_c_1836_n 0.0258205f $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_793 N_A_721_47#_c_950_n N_A_1251_49#_c_1830_n 0.00187896f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_794 N_A_721_47#_c_951_n N_A_1251_49#_c_1830_n 0.00611779f $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_795 N_A_721_47#_c_953_n N_A_1251_49#_c_1830_n 0.00163363f $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_796 N_A_721_47#_c_950_n N_A_1251_49#_c_1831_n 0.00194076f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_797 N_A_721_47#_c_951_n N_A_1251_49#_c_1831_n 0.00183791f $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_798 N_A_721_47#_c_948_n N_A_1251_49#_c_1832_n 0.00502701f $X=7.055 $Y=0.995
+ $X2=0 $Y2=0
cc_799 N_A_721_47#_c_950_n N_A_1251_49#_c_1832_n 0.00935867f $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_800 N_A_721_47#_c_951_n N_A_1251_49#_c_1832_n 0.00460812f $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_801 N_A_721_47#_c_953_n N_A_1251_49#_c_1832_n 0.00743847f $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_802 N_A_721_47#_c_950_n N_A_1565_49#_c_1971_n 9.26558e-19 $X=7.995 $Y=1.16
+ $X2=0 $Y2=0
cc_803 N_A_721_47#_c_953_n N_A_1565_49#_c_1971_n 0.00653698f $X=7.95 $Y=1.16
+ $X2=0 $Y2=0
cc_804 N_A_721_47#_c_951_n N_A_1565_49#_c_1963_n 0.00986682f $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_805 N_A_721_47#_c_948_n N_VGND_c_2044_n 0.00351226f $X=7.055 $Y=0.995 $X2=0
+ $Y2=0
cc_806 N_A_721_47#_c_951_n N_VGND_c_2044_n 0.00351226f $X=8.115 $Y=0.995 $X2=0
+ $Y2=0
cc_807 N_A_721_47#_M1028_d N_VGND_c_2049_n 0.00240414f $X=3.605 $Y=0.235 $X2=0
+ $Y2=0
cc_808 N_A_721_47#_c_948_n N_VGND_c_2049_n 0.00647149f $X=7.055 $Y=0.995 $X2=0
+ $Y2=0
cc_809 N_A_721_47#_c_951_n N_VGND_c_2049_n 0.00645346f $X=8.115 $Y=0.995 $X2=0
+ $Y2=0
cc_810 N_A_1636_315#_M1002_g N_CIN_M1016_g 0.0442256f $X=10.065 $Y=1.985 $X2=0
+ $Y2=0
cc_811 N_A_1636_315#_c_1141_n N_CIN_M1016_g 0.0208549f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_812 N_A_1636_315#_c_1149_n N_CIN_M1016_g 0.00592601f $X=10.7 $Y=2.31 $X2=0
+ $Y2=0
cc_813 N_A_1636_315#_c_1139_n N_CIN_c_1262_n 0.0089675f $X=10.53 $Y=0.82 $X2=0
+ $Y2=0
cc_814 N_A_1636_315#_c_1140_n N_CIN_c_1262_n 0.00739176f $X=10.72 $Y=0.4 $X2=0
+ $Y2=0
cc_815 N_A_1636_315#_c_1141_n N_CIN_c_1262_n 9.635e-19 $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_816 N_A_1636_315#_c_1143_n N_CIN_c_1262_n 0.0193376f $X=10.065 $Y=0.995 $X2=0
+ $Y2=0
cc_817 N_A_1636_315#_c_1139_n N_CIN_c_1263_n 6.87385e-19 $X=10.53 $Y=0.82 $X2=0
+ $Y2=0
cc_818 N_A_1636_315#_c_1141_n N_CIN_M1021_g 0.00107298f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_819 N_A_1636_315#_c_1139_n N_CIN_c_1264_n 8.04291e-19 $X=10.53 $Y=0.82 $X2=0
+ $Y2=0
cc_820 N_A_1636_315#_c_1141_n N_CIN_c_1264_n 0.0069139f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_821 N_A_1636_315#_c_1142_n N_CIN_c_1264_n 0.0215662f $X=10.065 $Y=1.16 $X2=0
+ $Y2=0
cc_822 N_A_1636_315#_c_1139_n N_CIN_c_1265_n 0.00578114f $X=10.53 $Y=0.82 $X2=0
+ $Y2=0
cc_823 N_A_1636_315#_c_1141_n N_CIN_c_1265_n 0.00592002f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_824 N_A_1636_315#_c_1139_n CIN 0.0250787f $X=10.53 $Y=0.82 $X2=0 $Y2=0
cc_825 N_A_1636_315#_c_1141_n CIN 0.0424662f $X=10.71 $Y=2.025 $X2=0 $Y2=0
cc_826 N_A_1636_315#_c_1145_n N_A_1647_49#_M1000_d 0.00165831f $X=9.24 $Y=2.38
+ $X2=0 $Y2=0
cc_827 N_A_1636_315#_M1002_g N_A_1647_49#_c_1335_n 0.00385016f $X=10.065
+ $Y=1.985 $X2=0 $Y2=0
cc_828 N_A_1636_315#_c_1138_n N_A_1647_49#_c_1335_n 0.0210222f $X=9.325 $Y=1.875
+ $X2=0 $Y2=0
cc_829 N_A_1636_315#_c_1184_p N_A_1647_49#_c_1335_n 0.0125749f $X=10.055 $Y=1.96
+ $X2=0 $Y2=0
cc_830 N_A_1636_315#_c_1139_n N_A_1647_49#_c_1335_n 3.12387e-19 $X=10.53 $Y=0.82
+ $X2=0 $Y2=0
cc_831 N_A_1636_315#_c_1141_n N_A_1647_49#_c_1335_n 0.0640764f $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_832 N_A_1636_315#_c_1142_n N_A_1647_49#_c_1335_n 9.6356e-19 $X=10.065 $Y=1.16
+ $X2=0 $Y2=0
cc_833 N_A_1636_315#_c_1138_n N_A_1647_49#_c_1336_n 0.00131308f $X=9.325
+ $Y=1.875 $X2=0 $Y2=0
cc_834 N_A_1636_315#_M1000_s N_A_1647_49#_c_1340_n 0.00341774f $X=8.18 $Y=1.575
+ $X2=0 $Y2=0
cc_835 N_A_1636_315#_c_1161_n N_A_1647_49#_c_1340_n 6.89312e-19 $X=8.305 $Y=2.12
+ $X2=0 $Y2=0
cc_836 N_A_1636_315#_c_1145_n N_A_1647_49#_c_1340_n 0.0195185f $X=9.24 $Y=2.38
+ $X2=0 $Y2=0
cc_837 N_A_1636_315#_c_1138_n N_A_1647_49#_c_1340_n 0.0154191f $X=9.325 $Y=1.875
+ $X2=0 $Y2=0
cc_838 N_A_1636_315#_c_1159_n N_A_1647_49#_c_1340_n 0.00336848f $X=9.325
+ $Y=2.295 $X2=0 $Y2=0
cc_839 N_A_1636_315#_c_1160_n N_A_1647_49#_c_1340_n 0.00805744f $X=9.325 $Y=1.96
+ $X2=0 $Y2=0
cc_840 N_A_1636_315#_c_1141_n N_VPWR_M1002_d 0.00195566f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_841 N_A_1636_315#_M1002_g N_VPWR_c_1605_n 0.00268723f $X=10.065 $Y=1.985
+ $X2=0 $Y2=0
cc_842 N_A_1636_315#_c_1141_n N_VPWR_c_1605_n 0.0130469f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_843 N_A_1636_315#_M1002_g N_VPWR_c_1608_n 0.00431122f $X=10.065 $Y=1.985
+ $X2=0 $Y2=0
cc_844 N_A_1636_315#_c_1145_n N_VPWR_c_1608_n 0.0659458f $X=9.24 $Y=2.38 $X2=0
+ $Y2=0
cc_845 N_A_1636_315#_c_1146_n N_VPWR_c_1608_n 0.0119306f $X=8.39 $Y=2.38 $X2=0
+ $Y2=0
cc_846 N_A_1636_315#_c_1184_p N_VPWR_c_1608_n 0.00985633f $X=10.055 $Y=1.96
+ $X2=0 $Y2=0
cc_847 N_A_1636_315#_c_1141_n N_VPWR_c_1608_n 0.00131017f $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_848 N_A_1636_315#_c_1141_n N_VPWR_c_1609_n 0.00235518f $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_849 N_A_1636_315#_c_1149_n N_VPWR_c_1609_n 0.0224828f $X=10.7 $Y=2.31 $X2=0
+ $Y2=0
cc_850 N_A_1636_315#_M1016_d N_VPWR_c_1601_n 0.00213418f $X=10.56 $Y=1.485 $X2=0
+ $Y2=0
cc_851 N_A_1636_315#_M1002_g N_VPWR_c_1601_n 0.00721611f $X=10.065 $Y=1.985
+ $X2=0 $Y2=0
cc_852 N_A_1636_315#_c_1145_n N_VPWR_c_1601_n 0.036823f $X=9.24 $Y=2.38 $X2=0
+ $Y2=0
cc_853 N_A_1636_315#_c_1146_n N_VPWR_c_1601_n 0.00649922f $X=8.39 $Y=2.38 $X2=0
+ $Y2=0
cc_854 N_A_1636_315#_c_1184_p N_VPWR_c_1601_n 0.0173811f $X=10.055 $Y=1.96 $X2=0
+ $Y2=0
cc_855 N_A_1636_315#_c_1141_n N_VPWR_c_1601_n 0.00832204f $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_856 N_A_1636_315#_c_1149_n N_VPWR_c_1601_n 0.0132199f $X=10.7 $Y=2.31 $X2=0
+ $Y2=0
cc_857 N_A_1636_315#_c_1141_n N_A_1251_49#_c_1834_n 0.0443688f $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_858 N_A_1636_315#_c_1149_n N_A_1251_49#_c_1835_n 0.0339937f $X=10.7 $Y=2.31
+ $X2=0 $Y2=0
cc_859 N_A_1636_315#_c_1140_n N_A_1251_49#_c_1880_n 0.0273464f $X=10.72 $Y=0.4
+ $X2=0 $Y2=0
cc_860 N_A_1636_315#_c_1139_n N_A_1251_49#_c_1881_n 0.00872264f $X=10.53 $Y=0.82
+ $X2=0 $Y2=0
cc_861 N_A_1636_315#_M1019_d N_A_1251_49#_c_1830_n 0.0048766f $X=8.675 $Y=0.245
+ $X2=0 $Y2=0
cc_862 N_A_1636_315#_c_1152_n N_A_1251_49#_c_1830_n 0.0141024f $X=9.24 $Y=0.68
+ $X2=0 $Y2=0
cc_863 N_A_1636_315#_c_1138_n N_A_1251_49#_c_1830_n 0.0166729f $X=9.325 $Y=1.875
+ $X2=0 $Y2=0
cc_864 N_A_1636_315#_c_1139_n N_A_1251_49#_c_1830_n 0.0253325f $X=10.53 $Y=0.82
+ $X2=0 $Y2=0
cc_865 N_A_1636_315#_c_1141_n N_A_1251_49#_c_1830_n 0.0210222f $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_866 N_A_1636_315#_c_1142_n N_A_1251_49#_c_1830_n 5.57837e-19 $X=10.065
+ $Y=1.16 $X2=0 $Y2=0
cc_867 N_A_1636_315#_c_1143_n N_A_1251_49#_c_1830_n 0.00503235f $X=10.065
+ $Y=0.995 $X2=0 $Y2=0
cc_868 N_A_1636_315#_c_1139_n N_A_1251_49#_c_1889_n 3.70194e-19 $X=10.53 $Y=0.82
+ $X2=0 $Y2=0
cc_869 N_A_1636_315#_c_1141_n N_A_1251_49#_c_1833_n 6.0064e-19 $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_870 N_A_1636_315#_c_1145_n N_A_1565_49#_M1023_d 0.0103526f $X=9.24 $Y=2.38
+ $X2=0 $Y2=0
cc_871 N_A_1636_315#_c_1138_n N_A_1565_49#_M1023_d 0.0101884f $X=9.325 $Y=1.875
+ $X2=0 $Y2=0
cc_872 N_A_1636_315#_c_1159_n N_A_1565_49#_M1023_d 0.00935662f $X=9.325 $Y=2.295
+ $X2=0 $Y2=0
cc_873 N_A_1636_315#_c_1184_p N_A_1565_49#_M1023_d 0.0194298f $X=10.055 $Y=1.96
+ $X2=0 $Y2=0
cc_874 N_A_1636_315#_c_1160_n N_A_1565_49#_M1023_d 0.00364924f $X=9.325 $Y=1.96
+ $X2=0 $Y2=0
cc_875 N_A_1636_315#_M1019_d N_A_1565_49#_c_1963_n 0.0183955f $X=8.675 $Y=0.245
+ $X2=0 $Y2=0
cc_876 N_A_1636_315#_c_1152_n N_A_1565_49#_c_1963_n 0.0448229f $X=9.24 $Y=0.68
+ $X2=0 $Y2=0
cc_877 N_A_1636_315#_c_1143_n N_A_1565_49#_c_1964_n 0.00194921f $X=10.065
+ $Y=0.995 $X2=0 $Y2=0
cc_878 N_A_1636_315#_c_1152_n N_A_1565_49#_c_1965_n 0.011843f $X=9.24 $Y=0.68
+ $X2=0 $Y2=0
cc_879 N_A_1636_315#_c_1140_n N_A_1565_49#_c_1965_n 0.00489878f $X=10.72 $Y=0.4
+ $X2=0 $Y2=0
cc_880 N_A_1636_315#_c_1143_n N_A_1565_49#_c_1965_n 0.00303692f $X=10.065
+ $Y=0.995 $X2=0 $Y2=0
cc_881 N_A_1636_315#_M1002_g N_A_1565_49#_c_1966_n 0.00340389f $X=10.065
+ $Y=1.985 $X2=0 $Y2=0
cc_882 N_A_1636_315#_c_1141_n N_A_1565_49#_c_1966_n 0.039819f $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_883 N_A_1636_315#_c_1142_n N_A_1565_49#_c_1966_n 0.00752814f $X=10.065
+ $Y=1.16 $X2=0 $Y2=0
cc_884 N_A_1636_315#_c_1143_n N_A_1565_49#_c_1966_n 0.00244964f $X=10.065
+ $Y=0.995 $X2=0 $Y2=0
cc_885 N_A_1636_315#_c_1138_n N_A_1565_49#_c_1967_n 0.043999f $X=9.325 $Y=1.875
+ $X2=0 $Y2=0
cc_886 N_A_1636_315#_c_1141_n N_A_1565_49#_c_1967_n 0.00586752f $X=10.71
+ $Y=2.025 $X2=0 $Y2=0
cc_887 N_A_1636_315#_c_1142_n N_A_1565_49#_c_1967_n 8.53648e-19 $X=10.065
+ $Y=1.16 $X2=0 $Y2=0
cc_888 N_A_1636_315#_c_1143_n N_A_1565_49#_c_1967_n 0.00260688f $X=10.065
+ $Y=0.995 $X2=0 $Y2=0
cc_889 N_A_1636_315#_M1002_g N_A_1565_49#_c_1993_n 0.00187515f $X=10.065
+ $Y=1.985 $X2=0 $Y2=0
cc_890 N_A_1636_315#_c_1138_n N_A_1565_49#_c_1993_n 0.00974348f $X=9.325
+ $Y=1.875 $X2=0 $Y2=0
cc_891 N_A_1636_315#_c_1184_p N_A_1565_49#_c_1993_n 0.0208998f $X=10.055 $Y=1.96
+ $X2=0 $Y2=0
cc_892 N_A_1636_315#_c_1141_n N_A_1565_49#_c_1993_n 0.00869812f $X=10.71
+ $Y=2.025 $X2=0 $Y2=0
cc_893 N_A_1636_315#_c_1142_n N_A_1565_49#_c_1993_n 0.00143352f $X=10.065
+ $Y=1.16 $X2=0 $Y2=0
cc_894 N_A_1636_315#_c_1139_n N_VGND_M1001_d 5.2343e-19 $X=10.53 $Y=0.82 $X2=0
+ $Y2=0
cc_895 N_A_1636_315#_c_1141_n N_VGND_M1001_d 0.0033195f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_896 N_A_1636_315#_c_1140_n N_VGND_c_2042_n 0.0199993f $X=10.72 $Y=0.4 $X2=0
+ $Y2=0
cc_897 N_A_1636_315#_c_1141_n N_VGND_c_2042_n 0.013297f $X=10.71 $Y=2.025 $X2=0
+ $Y2=0
cc_898 N_A_1636_315#_c_1143_n N_VGND_c_2042_n 0.00380764f $X=10.065 $Y=0.995
+ $X2=0 $Y2=0
cc_899 N_A_1636_315#_c_1143_n N_VGND_c_2044_n 0.00545275f $X=10.065 $Y=0.995
+ $X2=0 $Y2=0
cc_900 N_A_1636_315#_c_1139_n N_VGND_c_2047_n 0.00205365f $X=10.53 $Y=0.82 $X2=0
+ $Y2=0
cc_901 N_A_1636_315#_c_1140_n N_VGND_c_2047_n 0.0204614f $X=10.72 $Y=0.4 $X2=0
+ $Y2=0
cc_902 N_A_1636_315#_M1022_d N_VGND_c_2049_n 0.0017338f $X=10.585 $Y=0.235 $X2=0
+ $Y2=0
cc_903 N_A_1636_315#_c_1139_n N_VGND_c_2049_n 0.00178463f $X=10.53 $Y=0.82 $X2=0
+ $Y2=0
cc_904 N_A_1636_315#_c_1140_n N_VGND_c_2049_n 0.00664209f $X=10.72 $Y=0.4 $X2=0
+ $Y2=0
cc_905 N_A_1636_315#_c_1141_n N_VGND_c_2049_n 4.58187e-19 $X=10.71 $Y=2.025
+ $X2=0 $Y2=0
cc_906 N_A_1636_315#_c_1143_n N_VGND_c_2049_n 0.00752144f $X=10.065 $Y=0.995
+ $X2=0 $Y2=0
cc_907 N_CIN_M1021_g N_A_1647_49#_M1017_g 0.0261027f $X=11.45 $Y=1.985 $X2=0
+ $Y2=0
cc_908 N_CIN_M1021_g N_A_1647_49#_c_1335_n 0.00976642f $X=11.45 $Y=1.985 $X2=0
+ $Y2=0
cc_909 N_CIN_c_1265_n N_A_1647_49#_c_1335_n 0.00340455f $X=11.375 $Y=1.16 $X2=0
+ $Y2=0
cc_910 CIN N_A_1647_49#_c_1335_n 0.00365164f $X=10.74 $Y=1.105 $X2=0 $Y2=0
cc_911 N_CIN_M1021_g N_A_1647_49#_c_1337_n 0.00144107f $X=11.45 $Y=1.985 $X2=0
+ $Y2=0
cc_912 N_CIN_c_1266_n N_A_1647_49#_c_1330_n 0.0216941f $X=11.45 $Y=1.16 $X2=0
+ $Y2=0
cc_913 N_CIN_c_1266_n N_A_1647_49#_c_1331_n 0.00446904f $X=11.45 $Y=1.16 $X2=0
+ $Y2=0
cc_914 N_CIN_c_1263_n N_A_1647_49#_c_1332_n 0.0193354f $X=11.45 $Y=0.995 $X2=0
+ $Y2=0
cc_915 N_CIN_M1016_g N_VPWR_c_1605_n 0.00268723f $X=10.485 $Y=1.985 $X2=0 $Y2=0
cc_916 N_CIN_M1021_g N_VPWR_c_1606_n 0.00280208f $X=11.45 $Y=1.985 $X2=0 $Y2=0
cc_917 N_CIN_M1016_g N_VPWR_c_1609_n 0.00422443f $X=10.485 $Y=1.985 $X2=0 $Y2=0
cc_918 N_CIN_M1021_g N_VPWR_c_1609_n 0.00541359f $X=11.45 $Y=1.985 $X2=0 $Y2=0
cc_919 N_CIN_M1016_g N_VPWR_c_1601_n 0.00703375f $X=10.485 $Y=1.985 $X2=0 $Y2=0
cc_920 N_CIN_M1021_g N_VPWR_c_1601_n 0.0108548f $X=11.45 $Y=1.985 $X2=0 $Y2=0
cc_921 N_CIN_M1016_g N_A_1251_49#_c_1834_n 0.0014909f $X=10.485 $Y=1.985 $X2=0
+ $Y2=0
cc_922 N_CIN_M1021_g N_A_1251_49#_c_1834_n 0.00203012f $X=11.45 $Y=1.985 $X2=0
+ $Y2=0
cc_923 N_CIN_c_1265_n N_A_1251_49#_c_1834_n 0.00366648f $X=11.375 $Y=1.16 $X2=0
+ $Y2=0
cc_924 N_CIN_M1021_g N_A_1251_49#_c_1835_n 0.0101256f $X=11.45 $Y=1.985 $X2=0
+ $Y2=0
cc_925 N_CIN_c_1262_n N_A_1251_49#_c_1880_n 9.04978e-19 $X=10.51 $Y=0.995 $X2=0
+ $Y2=0
cc_926 N_CIN_c_1263_n N_A_1251_49#_c_1881_n 0.00384601f $X=11.45 $Y=0.995 $X2=0
+ $Y2=0
cc_927 N_CIN_c_1262_n N_A_1251_49#_c_1830_n 0.00197973f $X=10.51 $Y=0.995 $X2=0
+ $Y2=0
cc_928 N_CIN_c_1264_n N_A_1251_49#_c_1830_n 5.63257e-19 $X=10.497 $Y=1.16 $X2=0
+ $Y2=0
cc_929 N_CIN_c_1265_n N_A_1251_49#_c_1830_n 0.00894399f $X=11.375 $Y=1.16 $X2=0
+ $Y2=0
cc_930 CIN N_A_1251_49#_c_1830_n 0.00558207f $X=10.74 $Y=1.105 $X2=0 $Y2=0
cc_931 N_CIN_c_1263_n N_A_1251_49#_c_1889_n 0.00516076f $X=11.45 $Y=0.995 $X2=0
+ $Y2=0
cc_932 N_CIN_M1016_g N_A_1251_49#_c_1833_n 0.00279091f $X=10.485 $Y=1.985 $X2=0
+ $Y2=0
cc_933 N_CIN_c_1262_n N_A_1251_49#_c_1833_n 0.00196745f $X=10.51 $Y=0.995 $X2=0
+ $Y2=0
cc_934 N_CIN_c_1263_n N_A_1251_49#_c_1833_n 0.00741274f $X=11.45 $Y=0.995 $X2=0
+ $Y2=0
cc_935 N_CIN_M1021_g N_A_1251_49#_c_1833_n 0.00393605f $X=11.45 $Y=1.985 $X2=0
+ $Y2=0
cc_936 N_CIN_c_1265_n N_A_1251_49#_c_1833_n 0.0220421f $X=11.375 $Y=1.16 $X2=0
+ $Y2=0
cc_937 N_CIN_c_1266_n N_A_1251_49#_c_1833_n 0.00395206f $X=11.45 $Y=1.16 $X2=0
+ $Y2=0
cc_938 CIN N_A_1251_49#_c_1833_n 0.0136896f $X=10.74 $Y=1.105 $X2=0 $Y2=0
cc_939 N_CIN_c_1262_n N_A_1565_49#_c_1965_n 4.80288e-19 $X=10.51 $Y=0.995 $X2=0
+ $Y2=0
cc_940 N_CIN_c_1263_n N_SUM_c_2022_n 7.72042e-19 $X=11.45 $Y=0.995 $X2=0 $Y2=0
cc_941 N_CIN_c_1262_n N_VGND_c_2042_n 0.00437781f $X=10.51 $Y=0.995 $X2=0 $Y2=0
cc_942 N_CIN_c_1263_n N_VGND_c_2043_n 0.0101282f $X=11.45 $Y=0.995 $X2=0 $Y2=0
cc_943 N_CIN_c_1262_n N_VGND_c_2047_n 0.00413062f $X=10.51 $Y=0.995 $X2=0 $Y2=0
cc_944 N_CIN_c_1263_n N_VGND_c_2047_n 0.00428962f $X=11.45 $Y=0.995 $X2=0 $Y2=0
cc_945 N_CIN_c_1262_n N_VGND_c_2049_n 0.00699361f $X=10.51 $Y=0.995 $X2=0 $Y2=0
cc_946 N_CIN_c_1263_n N_VGND_c_2049_n 0.00680675f $X=11.45 $Y=0.995 $X2=0 $Y2=0
cc_947 N_A_1647_49#_c_1335_n N_VPWR_M1002_d 3.3943e-19 $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_948 N_A_1647_49#_c_1335_n N_VPWR_M1021_d 0.00228444f $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_949 N_A_1647_49#_c_1337_n N_VPWR_M1021_d 0.00180492f $X=11.765 $Y=1.53 $X2=0
+ $Y2=0
cc_950 N_A_1647_49#_c_1331_n N_VPWR_M1021_d 0.00128737f $X=11.87 $Y=1.16 $X2=0
+ $Y2=0
cc_951 N_A_1647_49#_c_1335_n N_VPWR_c_1605_n 6.3305e-19 $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_952 N_A_1647_49#_M1017_g N_VPWR_c_1606_n 0.0135622f $X=11.87 $Y=1.985 $X2=0
+ $Y2=0
cc_953 N_A_1647_49#_c_1335_n N_VPWR_c_1606_n 0.00226154f $X=11.62 $Y=1.53 $X2=0
+ $Y2=0
cc_954 N_A_1647_49#_c_1337_n N_VPWR_c_1606_n 0.00669312f $X=11.765 $Y=1.53 $X2=0
+ $Y2=0
cc_955 N_A_1647_49#_c_1331_n N_VPWR_c_1606_n 0.00992907f $X=11.87 $Y=1.16 $X2=0
+ $Y2=0
cc_956 N_A_1647_49#_M1017_g N_VPWR_c_1610_n 0.00447018f $X=11.87 $Y=1.985 $X2=0
+ $Y2=0
cc_957 N_A_1647_49#_M1017_g N_VPWR_c_1601_n 0.00860724f $X=11.87 $Y=1.985 $X2=0
+ $Y2=0
cc_958 N_A_1647_49#_M1017_g N_A_1251_49#_c_1834_n 7.52739e-19 $X=11.87 $Y=1.985
+ $X2=0 $Y2=0
cc_959 N_A_1647_49#_c_1335_n N_A_1251_49#_c_1834_n 0.0339216f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_960 N_A_1647_49#_c_1337_n N_A_1251_49#_c_1834_n 0.00177524f $X=11.765 $Y=1.53
+ $X2=0 $Y2=0
cc_961 N_A_1647_49#_c_1332_n N_A_1251_49#_c_1881_n 0.00179054f $X=11.87 $Y=0.995
+ $X2=0 $Y2=0
cc_962 N_A_1647_49#_M1029_d N_A_1251_49#_c_1830_n 5.85211e-19 $X=8.235 $Y=0.245
+ $X2=0 $Y2=0
cc_963 N_A_1647_49#_c_1329_n N_A_1251_49#_c_1830_n 0.0188099f $X=8.39 $Y=0.76
+ $X2=0 $Y2=0
cc_964 N_A_1647_49#_c_1335_n N_A_1251_49#_c_1830_n 0.0893135f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_965 N_A_1647_49#_c_1329_n N_A_1251_49#_c_1831_n 0.001045f $X=8.39 $Y=0.76
+ $X2=0 $Y2=0
cc_966 N_A_1647_49#_c_1329_n N_A_1251_49#_c_1832_n 0.00295833f $X=8.39 $Y=0.76
+ $X2=0 $Y2=0
cc_967 N_A_1647_49#_c_1335_n N_A_1251_49#_c_1889_n 0.0126255f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_968 N_A_1647_49#_c_1332_n N_A_1251_49#_c_1889_n 0.00112497f $X=11.87 $Y=0.995
+ $X2=0 $Y2=0
cc_969 N_A_1647_49#_M1017_g N_A_1251_49#_c_1833_n 3.23024e-19 $X=11.87 $Y=1.985
+ $X2=0 $Y2=0
cc_970 N_A_1647_49#_c_1337_n N_A_1251_49#_c_1833_n 0.00125324f $X=11.765 $Y=1.53
+ $X2=0 $Y2=0
cc_971 N_A_1647_49#_c_1330_n N_A_1251_49#_c_1833_n 2.99878e-19 $X=11.87 $Y=1.16
+ $X2=0 $Y2=0
cc_972 N_A_1647_49#_c_1331_n N_A_1251_49#_c_1833_n 0.0342796f $X=11.87 $Y=1.16
+ $X2=0 $Y2=0
cc_973 N_A_1647_49#_c_1335_n N_A_1565_49#_M1023_d 0.0109275f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_974 N_A_1647_49#_M1029_d N_A_1565_49#_c_1963_n 0.00351836f $X=8.235 $Y=0.245
+ $X2=0 $Y2=0
cc_975 N_A_1647_49#_c_1329_n N_A_1565_49#_c_1963_n 0.0133054f $X=8.39 $Y=0.76
+ $X2=0 $Y2=0
cc_976 N_A_1647_49#_c_1335_n N_A_1565_49#_c_1966_n 0.00845622f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_977 N_A_1647_49#_c_1335_n N_A_1565_49#_c_1993_n 0.0123644f $X=11.62 $Y=1.53
+ $X2=0 $Y2=0
cc_978 N_A_1647_49#_M1017_g SUM 0.00620927f $X=11.87 $Y=1.985 $X2=0 $Y2=0
cc_979 N_A_1647_49#_c_1337_n SUM 0.00263862f $X=11.765 $Y=1.53 $X2=0 $Y2=0
cc_980 N_A_1647_49#_c_1330_n SUM 0.00757246f $X=11.87 $Y=1.16 $X2=0 $Y2=0
cc_981 N_A_1647_49#_c_1331_n SUM 0.0414319f $X=11.87 $Y=1.16 $X2=0 $Y2=0
cc_982 N_A_1647_49#_c_1332_n SUM 0.00715959f $X=11.87 $Y=0.995 $X2=0 $Y2=0
cc_983 N_A_1647_49#_c_1332_n N_SUM_c_2022_n 0.00490295f $X=11.87 $Y=0.995 $X2=0
+ $Y2=0
cc_984 N_A_1647_49#_c_1330_n N_VGND_c_2043_n 4.51599e-19 $X=11.87 $Y=1.16 $X2=0
+ $Y2=0
cc_985 N_A_1647_49#_c_1331_n N_VGND_c_2043_n 0.0065286f $X=11.87 $Y=1.16 $X2=0
+ $Y2=0
cc_986 N_A_1647_49#_c_1332_n N_VGND_c_2043_n 0.00323533f $X=11.87 $Y=0.995 $X2=0
+ $Y2=0
cc_987 N_A_1647_49#_c_1332_n N_VGND_c_2048_n 0.00579312f $X=11.87 $Y=0.995 $X2=0
+ $Y2=0
cc_988 N_A_1647_49#_c_1332_n N_VGND_c_2049_n 0.0115602f $X=11.87 $Y=0.995 $X2=0
+ $Y2=0
cc_989 N_A_27_47#_c_1456_n N_VPWR_M1013_d 0.00541207f $X=0.94 $Y=1.925 $X2=-0.19
+ $Y2=-0.24
cc_990 N_A_27_47#_c_1456_n N_VPWR_c_1602_n 0.0126308f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_991 N_A_27_47#_c_1463_n N_VPWR_c_1602_n 0.00242328f $X=1.025 $Y=2.215 $X2=0
+ $Y2=0
cc_992 N_A_27_47#_c_1503_n N_VPWR_c_1602_n 0.0133618f $X=1.11 $Y=2.3 $X2=0 $Y2=0
cc_993 N_A_27_47#_c_1456_n N_VPWR_c_1603_n 0.00208831f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_994 N_A_27_47#_c_1503_n N_VPWR_c_1603_n 0.00633644f $X=1.11 $Y=2.3 $X2=0
+ $Y2=0
cc_995 N_A_27_47#_c_1446_n N_VPWR_c_1603_n 0.025708f $X=1.715 $Y=2.34 $X2=0
+ $Y2=0
cc_996 N_A_27_47#_c_1447_n N_VPWR_c_1603_n 0.0988797f $X=1.97 $Y=2.34 $X2=0
+ $Y2=0
cc_997 N_A_27_47#_c_1448_n N_VPWR_c_1603_n 0.0186052f $X=3.29 $Y=2.38 $X2=0
+ $Y2=0
cc_998 N_A_27_47#_c_1441_n N_VPWR_c_1607_n 0.0221067f $X=0.265 $Y=2.31 $X2=0
+ $Y2=0
cc_999 N_A_27_47#_c_1456_n N_VPWR_c_1607_n 0.00191602f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_1000 N_A_27_47#_M1013_s N_VPWR_c_1601_n 0.00213418f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_1001 N_A_27_47#_M1020_s N_VPWR_c_1601_n 0.00202962f $X=3.165 $Y=1.485 $X2=0
+ $Y2=0
cc_1002 N_A_27_47#_c_1441_n N_VPWR_c_1601_n 0.0130045f $X=0.265 $Y=2.31 $X2=0
+ $Y2=0
cc_1003 N_A_27_47#_c_1456_n N_VPWR_c_1601_n 0.00872069f $X=0.94 $Y=1.925 $X2=0
+ $Y2=0
cc_1004 N_A_27_47#_c_1503_n N_VPWR_c_1601_n 0.00570549f $X=1.11 $Y=2.3 $X2=0
+ $Y2=0
cc_1005 N_A_27_47#_c_1444_n N_VPWR_c_1601_n 2.06696e-19 $X=0.265 $Y=1.63 $X2=0
+ $Y2=0
cc_1006 N_A_27_47#_c_1446_n N_VPWR_c_1601_n 0.0214051f $X=1.715 $Y=2.34 $X2=0
+ $Y2=0
cc_1007 N_A_27_47#_c_1447_n N_VPWR_c_1601_n 0.0278358f $X=1.97 $Y=2.34 $X2=0
+ $Y2=0
cc_1008 N_A_27_47#_c_1448_n N_VPWR_c_1601_n 0.0048573f $X=3.29 $Y=2.38 $X2=0
+ $Y2=0
cc_1009 N_A_27_47#_c_1434_n N_VGND_c_2040_n 0.0188898f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_1010 N_A_27_47#_c_1440_n N_VGND_c_2041_n 0.00690613f $X=4.405 $Y=0.39 $X2=0
+ $Y2=0
cc_1011 N_A_27_47#_c_1478_n N_VGND_c_2046_n 0.00986382f $X=3.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1012 N_A_27_47#_c_1439_n N_VGND_c_2046_n 0.00186133f $X=3.375 $Y=0.79 $X2=0
+ $Y2=0
cc_1013 N_A_27_47#_c_1519_n N_VGND_c_2046_n 0.0500253f $X=4.24 $Y=0.365 $X2=0
+ $Y2=0
cc_1014 N_A_27_47#_M1007_s N_VGND_c_2049_n 0.00213418f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_1015 N_A_27_47#_c_1434_n N_VGND_c_2049_n 0.0123905f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_1016 N_A_27_47#_c_1478_n N_VGND_c_2049_n 0.00301895f $X=3.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1017 N_A_27_47#_c_1437_n N_VGND_c_2049_n 3.91258e-19 $X=0.257 $Y=0.805 $X2=0
+ $Y2=0
cc_1018 N_A_27_47#_c_1439_n N_VGND_c_2049_n 0.00228493f $X=3.375 $Y=0.79 $X2=0
+ $Y2=0
cc_1019 N_A_27_47#_c_1519_n N_VGND_c_2049_n 0.0149518f $X=4.24 $Y=0.365 $X2=0
+ $Y2=0
cc_1020 N_A_27_47#_c_1434_n N_VGND_c_2050_n 0.0209072f $X=0.265 $Y=0.38 $X2=0
+ $Y2=0
cc_1021 N_A_27_47#_c_1437_n N_VGND_c_2050_n 2.33971e-19 $X=0.257 $Y=0.805 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1601_n N_A_1142_49#_M1006_d 0.00562065f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1601_n N_A_1251_49#_M1021_s 0.00209319f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1024 N_VPWR_c_1609_n N_A_1251_49#_c_1835_n 0.0210382f $X=11.575 $Y=2.72 $X2=0
+ $Y2=0
cc_1025 N_VPWR_c_1601_n N_A_1251_49#_c_1835_n 0.0124268f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1026 N_VPWR_c_1601_n N_A_1565_49#_M1023_d 0.00581128f $X=12.19 $Y=2.72 $X2=0
+ $Y2=0
cc_1027 N_VPWR_c_1601_n N_SUM_M1017_d 0.0042075f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1028 N_VPWR_c_1610_n SUM 0.0235249f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1029 N_VPWR_c_1601_n SUM 0.0128192f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_1030 N_A_1142_49#_c_1751_n N_COUT_M1030_d 0.00324451f $X=7.04 $Y=2.04 $X2=0
+ $Y2=0
cc_1031 N_A_1142_49#_c_1729_n COUT 0.00590902f $X=5.885 $Y=1.555 $X2=0 $Y2=0
cc_1032 N_A_1142_49#_c_1730_n COUT 0.0199735f $X=7.125 $Y=1.23 $X2=0 $Y2=0
cc_1033 N_A_1142_49#_c_1732_n COUT 0.0205108f $X=7.125 $Y=1.955 $X2=0 $Y2=0
cc_1034 N_A_1142_49#_c_1729_n COUT 4.18687e-19 $X=5.885 $Y=1.555 $X2=0 $Y2=0
cc_1035 N_A_1142_49#_c_1745_n COUT 0.00777354f $X=6.2 $Y=1.64 $X2=0 $Y2=0
cc_1036 N_A_1142_49#_c_1751_n COUT 0.015187f $X=7.04 $Y=2.04 $X2=0 $Y2=0
cc_1037 N_A_1142_49#_c_1730_n N_COUT_c_1802_n 0.013211f $X=7.125 $Y=1.23 $X2=0
+ $Y2=0
cc_1038 N_A_1142_49#_c_1751_n N_A_1251_49#_M1009_d 0.0027538f $X=7.04 $Y=2.04
+ $X2=0 $Y2=0
cc_1039 N_A_1142_49#_c_1732_n N_A_1251_49#_M1009_d 0.00499655f $X=7.125 $Y=1.955
+ $X2=0 $Y2=0
cc_1040 N_A_1142_49#_M1014_d N_A_1251_49#_c_1829_n 0.00561037f $X=7.13 $Y=0.245
+ $X2=0 $Y2=0
cc_1041 N_A_1142_49#_c_1730_n N_A_1251_49#_c_1829_n 0.0156983f $X=7.125 $Y=1.23
+ $X2=0 $Y2=0
cc_1042 N_A_1142_49#_c_1751_n N_A_1251_49#_c_1861_n 0.0138309f $X=7.04 $Y=2.04
+ $X2=0 $Y2=0
cc_1043 N_A_1142_49#_c_1732_n N_A_1251_49#_c_1861_n 0.0307964f $X=7.125 $Y=1.955
+ $X2=0 $Y2=0
cc_1044 N_A_1142_49#_c_1739_n N_A_1251_49#_c_1838_n 0.0103218f $X=5.845 $Y=0.58
+ $X2=0 $Y2=0
cc_1045 N_A_1142_49#_c_1730_n N_A_1251_49#_c_1836_n 0.00834029f $X=7.125 $Y=1.23
+ $X2=0 $Y2=0
cc_1046 N_A_1142_49#_c_1732_n N_A_1251_49#_c_1836_n 0.0200856f $X=7.125 $Y=1.955
+ $X2=0 $Y2=0
cc_1047 N_A_1142_49#_c_1730_n N_A_1251_49#_c_1831_n 0.00772608f $X=7.125 $Y=1.23
+ $X2=0 $Y2=0
cc_1048 N_A_1142_49#_c_1730_n N_A_1251_49#_c_1832_n 0.0323983f $X=7.125 $Y=1.23
+ $X2=0 $Y2=0
cc_1049 N_A_1142_49#_c_1739_n N_VGND_c_2044_n 0.00999822f $X=5.845 $Y=0.58 $X2=0
+ $Y2=0
cc_1050 N_A_1142_49#_c_1739_n N_VGND_c_2049_n 0.0101398f $X=5.845 $Y=0.58 $X2=0
+ $Y2=0
cc_1051 N_COUT_M1031_d N_A_1251_49#_c_1829_n 0.0031917f $X=6.705 $Y=0.245 $X2=0
+ $Y2=0
cc_1052 N_COUT_c_1802_n N_A_1251_49#_c_1829_n 0.0160879f $X=6.735 $Y=0.925 $X2=0
+ $Y2=0
cc_1053 N_A_1251_49#_c_1830_n N_A_1565_49#_M1029_s 0.00238205f $X=11.16 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1054 N_A_1251_49#_c_1830_n N_A_1565_49#_c_1971_n 0.00277415f $X=11.16 $Y=0.85
+ $X2=0 $Y2=0
cc_1055 N_A_1251_49#_c_1832_n N_A_1565_49#_c_1971_n 0.0232269f $X=7.605 $Y=0.85
+ $X2=0 $Y2=0
cc_1056 N_A_1251_49#_c_1830_n N_A_1565_49#_c_1963_n 0.0176987f $X=11.16 $Y=0.85
+ $X2=0 $Y2=0
cc_1057 N_A_1251_49#_c_1829_n N_A_1565_49#_c_2009_n 0.0156276f $X=7.52 $Y=0.34
+ $X2=0 $Y2=0
cc_1058 N_A_1251_49#_c_1830_n N_A_1565_49#_c_1966_n 0.00917535f $X=11.16 $Y=0.85
+ $X2=0 $Y2=0
cc_1059 N_A_1251_49#_c_1830_n N_A_1565_49#_c_1967_n 0.0160105f $X=11.16 $Y=0.85
+ $X2=0 $Y2=0
cc_1060 N_A_1251_49#_c_1830_n N_A_1565_49#_c_1993_n 0.00104887f $X=11.16 $Y=0.85
+ $X2=0 $Y2=0
cc_1061 N_A_1251_49#_c_1881_n SUM 0.00262228f $X=11.28 $Y=0.805 $X2=0 $Y2=0
cc_1062 N_A_1251_49#_c_1889_n SUM 0.00181067f $X=11.305 $Y=0.85 $X2=0 $Y2=0
cc_1063 N_A_1251_49#_c_1830_n N_VGND_M1001_d 9.93578e-19 $X=11.16 $Y=0.85 $X2=0
+ $Y2=0
cc_1064 N_A_1251_49#_c_1830_n N_VGND_c_2042_n 8.18814e-19 $X=11.16 $Y=0.85 $X2=0
+ $Y2=0
cc_1065 N_A_1251_49#_c_1829_n N_VGND_c_2044_n 0.0665874f $X=7.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1066 N_A_1251_49#_c_1838_n N_VGND_c_2044_n 0.0200031f $X=6.42 $Y=0.34 $X2=0
+ $Y2=0
cc_1067 N_A_1251_49#_c_1880_n N_VGND_c_2047_n 0.0105862f $X=11.24 $Y=0.55 $X2=0
+ $Y2=0
cc_1068 N_A_1251_49#_c_1881_n N_VGND_c_2047_n 8.99889e-19 $X=11.28 $Y=0.805
+ $X2=0 $Y2=0
cc_1069 N_A_1251_49#_c_1829_n N_VGND_c_2049_n 0.0353917f $X=7.52 $Y=0.34 $X2=0
+ $Y2=0
cc_1070 N_A_1251_49#_c_1880_n N_VGND_c_2049_n 0.00292257f $X=11.24 $Y=0.55 $X2=0
+ $Y2=0
cc_1071 N_A_1251_49#_c_1838_n N_VGND_c_2049_n 0.0122613f $X=6.42 $Y=0.34 $X2=0
+ $Y2=0
cc_1072 N_A_1251_49#_c_1881_n N_VGND_c_2049_n 9.51601e-19 $X=11.28 $Y=0.805
+ $X2=0 $Y2=0
cc_1073 N_A_1251_49#_c_1830_n N_VGND_c_2049_n 0.165116f $X=11.16 $Y=0.85 $X2=0
+ $Y2=0
cc_1074 N_A_1251_49#_c_1831_n N_VGND_c_2049_n 0.0154677f $X=7.75 $Y=0.85 $X2=0
+ $Y2=0
cc_1075 N_A_1251_49#_c_1889_n N_VGND_c_2049_n 0.0149084f $X=11.305 $Y=0.85 $X2=0
+ $Y2=0
cc_1076 N_A_1565_49#_c_1964_n N_VGND_c_2042_n 0.0117758f $X=9.81 $Y=0.425 $X2=0
+ $Y2=0
cc_1077 N_A_1565_49#_c_1965_n N_VGND_c_2042_n 0.0091072f $X=9.81 $Y=0.655 $X2=0
+ $Y2=0
cc_1078 N_A_1565_49#_c_1963_n N_VGND_c_2044_n 0.0951651f $X=9.64 $Y=0.34 $X2=0
+ $Y2=0
cc_1079 N_A_1565_49#_c_2009_n N_VGND_c_2044_n 0.0114347f $X=8.035 $Y=0.34 $X2=0
+ $Y2=0
cc_1080 N_A_1565_49#_c_1964_n N_VGND_c_2044_n 0.0218171f $X=9.81 $Y=0.425 $X2=0
+ $Y2=0
cc_1081 N_A_1565_49#_c_1963_n N_VGND_c_2049_n 0.0267792f $X=9.64 $Y=0.34 $X2=0
+ $Y2=0
cc_1082 N_A_1565_49#_c_2009_n N_VGND_c_2049_n 0.0030628f $X=8.035 $Y=0.34 $X2=0
+ $Y2=0
cc_1083 N_A_1565_49#_c_1964_n N_VGND_c_2049_n 0.00615485f $X=9.81 $Y=0.425 $X2=0
+ $Y2=0
cc_1084 N_SUM_c_2022_n N_VGND_c_2048_n 0.0217448f $X=12.16 $Y=0.39 $X2=0 $Y2=0
cc_1085 N_SUM_M1025_d N_VGND_c_2049_n 0.00229814f $X=12 $Y=0.235 $X2=0 $Y2=0
cc_1086 N_SUM_c_2022_n N_VGND_c_2049_n 0.0129038f $X=12.16 $Y=0.39 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nand4bb_2.spice.pex
* Created: Thu Aug 27 14:30:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%B_N 4 5 7 10 14 18 20 21 25 27
c40 20 0 1.9583e-19 $X=0.235 $Y=1.19
c41 18 0 2.62595e-20 $X=0.47 $Y=1.86
c42 10 0 6.73268e-20 $X=0.47 $Y=2.275
r43 25 28 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r44 25 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r45 20 21 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r46 20 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r47 16 18 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.86
+ $X2=0.47 $Y2=1.86
r48 12 14 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r49 8 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.935
+ $X2=0.47 $Y2=1.86
r50 8 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.47 $Y=1.935 $X2=0.47
+ $Y2=2.275
r51 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r52 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r53 4 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.785
+ $X2=0.305 $Y2=1.86
r54 4 28 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.305 $Y=1.785
+ $X2=0.305 $Y2=1.4
r55 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r56 1 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%A_N 3 7 9 10 14
c38 7 0 1.7806e-19 $X=0.89 $Y=2.275
c39 3 0 1.60458e-19 $X=0.89 $Y=0.445
r40 14 17 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.777 $Y=1.255
+ $X2=0.777 $Y2=1.42
r41 14 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.777 $Y=1.255
+ $X2=0.777 $Y2=1.09
r42 9 10 14.061 $w=2.95e-07 $l=3.4e-07 $layer=LI1_cond $X=0.725 $Y=1.19
+ $X2=0.725 $Y2=1.53
r43 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.255 $X2=0.725 $Y2=1.255
r44 7 17 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.89 $Y=2.275
+ $X2=0.89 $Y2=1.42
r45 3 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%A_193_47# 1 2 7 9 12 14 16 20 22 25 29 35
+ 38 41 42 43
c79 38 0 1.42688e-19 $X=1.495 $Y=1.16
c80 29 0 6.73268e-20 $X=1.4 $Y=2.307
r81 41 43 46.8987 $w=1.73e-07 $l=7.4e-07 $layer=LI1_cond $X=1.487 $Y=2.15
+ $X2=1.487 $Y2=1.41
r82 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r83 36 43 5.54545 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=1.49 $Y=1.32 $X2=1.49
+ $Y2=1.41
r84 36 38 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=1.49 $Y=1.32
+ $X2=1.49 $Y2=1.16
r85 35 42 5.54545 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=1.49 $Y=0.805 $X2=1.49
+ $Y2=0.715
r86 35 38 21.8737 $w=1.78e-07 $l=3.55e-07 $layer=LI1_cond $X=1.49 $Y=0.805
+ $X2=1.49 $Y2=1.16
r87 33 42 9.82338 $w=1.73e-07 $l=1.55e-07 $layer=LI1_cond $X=1.487 $Y=0.56
+ $X2=1.487 $Y2=0.715
r88 29 41 7.5664 $w=3.15e-07 $l=1.95724e-07 $layer=LI1_cond $X=1.4 $Y=2.307
+ $X2=1.487 $Y2=2.15
r89 29 31 10.9756 $w=3.13e-07 $l=3e-07 $layer=LI1_cond $X=1.4 $Y=2.307 $X2=1.1
+ $Y2=2.307
r90 25 33 7.48781 $w=3.05e-07 $l=1.91625e-07 $layer=LI1_cond $X=1.4 $Y=0.407
+ $X2=1.487 $Y2=0.56
r91 25 27 11.3355 $w=3.03e-07 $l=3e-07 $layer=LI1_cond $X=1.4 $Y=0.407 $X2=1.1
+ $Y2=0.407
r92 22 39 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=1.965 $Y=1.16
+ $X2=1.495 $Y2=1.16
r93 22 23 11.9831 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.965 $Y=1.16
+ $X2=2.04 $Y2=1.16
r94 14 23 71.0316 $w=2.85e-07 $l=4.2e-07 $layer=POLY_cond $X=2.46 $Y=1.16
+ $X2=2.04 $Y2=1.16
r95 14 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.46 $Y=1.295
+ $X2=2.46 $Y2=1.985
r96 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.46 $Y=1.025
+ $X2=2.46 $Y2=0.56
r97 10 23 17.7656 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.325
+ $X2=2.04 $Y2=1.16
r98 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.04 $Y=1.325
+ $X2=2.04 $Y2=1.985
r99 7 23 17.7656 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=0.995
+ $X2=2.04 $Y2=1.16
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.04 $Y=0.995
+ $X2=2.04 $Y2=0.56
r101 2 31 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=2.065 $X2=1.1 $Y2=2.33
r102 1 27 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%A_27_47# 1 2 9 13 17 21 25 29 31 32 33 34
+ 39 42 49 50
r113 48 50 86.6477 $w=2.7e-07 $l=3.9e-07 $layer=POLY_cond $X=2.91 $Y=1.16
+ $X2=3.3 $Y2=1.16
r114 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.16 $X2=2.91 $Y2=1.16
r115 45 48 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.88 $Y=1.16 $X2=2.91
+ $Y2=1.16
r116 42 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.19
+ $X2=2.99 $Y2=1.19
r117 38 42 1.18376 $w=2.3e-07 $l=1.845e-06 $layer=MET1_cond $X=1.145 $Y=1.19
+ $X2=2.99 $Y2=1.19
r118 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.145 $Y=1.19
+ $X2=1.145 $Y2=1.19
r119 36 39 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.145 $Y=1.785
+ $X2=1.145 $Y2=1.19
r120 35 39 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.145 $Y=0.9
+ $X2=1.145 $Y2=1.19
r121 33 36 6.85817 $w=1.95e-07 $l=1.32868e-07 $layer=LI1_cond $X=1.06 $Y=1.882
+ $X2=1.145 $Y2=1.785
r122 33 34 39.2448 $w=1.93e-07 $l=6.9e-07 $layer=LI1_cond $X=1.06 $Y=1.882
+ $X2=0.37 $Y2=1.882
r123 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=0.815
+ $X2=1.145 $Y2=0.9
r124 31 32 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.06 $Y=0.815
+ $X2=0.345 $Y2=0.815
r125 27 34 7.13288 $w=1.95e-07 $l=1.85642e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.37 $Y2=1.882
r126 27 29 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.227 $Y2=2.275
r127 23 32 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.73
+ $X2=0.345 $Y2=0.815
r128 23 25 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=0.215 $Y=0.73
+ $X2=0.215 $Y2=0.46
r129 19 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.3 $Y=1.295
+ $X2=3.3 $Y2=1.16
r130 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.3 $Y=1.295
+ $X2=3.3 $Y2=1.985
r131 15 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.3 $Y=1.025
+ $X2=3.3 $Y2=1.16
r132 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.3 $Y=1.025
+ $X2=3.3 $Y2=0.56
r133 11 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.88 $Y=1.295
+ $X2=2.88 $Y2=1.16
r134 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.88 $Y=1.295
+ $X2=2.88 $Y2=1.985
r135 7 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.88 $Y=1.025
+ $X2=2.88 $Y2=1.16
r136 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.88 $Y=1.025
+ $X2=2.88 $Y2=0.56
r137 2 29 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.275
r138 1 25 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%C 5 9 13 17 19 20 23 27
c48 13 0 1.79953e-19 $X=4.66 $Y=0.56
r49 25 27 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.45 $Y=1.16
+ $X2=4.66 $Y2=1.16
r50 23 25 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.24 $Y=1.16
+ $X2=4.45 $Y2=1.16
r51 20 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.45
+ $Y=1.16 $X2=4.45 $Y2=1.16
r52 19 20 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.93 $Y=1.175
+ $X2=4.39 $Y2=1.175
r53 15 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.66 $Y=1.295
+ $X2=4.66 $Y2=1.16
r54 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.66 $Y=1.295
+ $X2=4.66 $Y2=1.985
r55 11 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.66 $Y=1.025
+ $X2=4.66 $Y2=1.16
r56 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.66 $Y=1.025
+ $X2=4.66 $Y2=0.56
r57 7 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.24 $Y=1.295
+ $X2=4.24 $Y2=1.16
r58 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.24 $Y=1.295 $X2=4.24
+ $Y2=1.985
r59 3 23 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.24 $Y=1.025
+ $X2=4.24 $Y2=1.16
r60 3 5 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.24 $Y=1.025
+ $X2=4.24 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%D 3 7 11 15 17 20 21 25
c51 3 0 7.99167e-20 $X=5.08 $Y=0.56
r52 21 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.71
+ $Y=1.16 $X2=5.71 $Y2=1.16
r53 20 21 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=5.31 $Y=1.175 $X2=5.71
+ $Y2=1.175
r54 17 25 27.9249 $w=2.9e-07 $l=1.35e-07 $layer=POLY_cond $X=5.575 $Y=1.16
+ $X2=5.71 $Y2=1.16
r55 17 19 12.6663 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=5.575 $Y=1.16
+ $X2=5.5 $Y2=1.16
r56 13 19 16.847 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.5 $Y=1.305 $X2=5.5
+ $Y2=1.16
r57 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.5 $Y=1.305 $X2=5.5
+ $Y2=1.985
r58 9 19 16.847 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.5 $Y=1.015 $X2=5.5
+ $Y2=1.16
r59 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.5 $Y=1.015 $X2=5.5
+ $Y2=0.56
r60 1 19 73.8832 $w=2.74e-07 $l=4.2e-07 $layer=POLY_cond $X=5.08 $Y=1.16 $X2=5.5
+ $Y2=1.16
r61 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.08 $Y=1.295 $X2=5.08
+ $Y2=1.985
r62 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.08 $Y=1.025
+ $X2=5.08 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%VPWR 1 2 3 4 5 6 21 25 29 33 35 39 41 45
+ 47 49 53 54 55 57 66 72 75 78 83 87
c88 87 0 2.62595e-20 $X=5.75 $Y=2.72
r89 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r90 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r91 79 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r92 79 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r93 78 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r94 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r95 76 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r96 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r97 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r98 70 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r99 70 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r100 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r101 67 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=4.87 $Y2=2.72
r102 67 69 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=5.29 $Y2=2.72
r103 66 86 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=5.625 $Y=2.72
+ $X2=5.802 $Y2=2.72
r104 66 69 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.625 $Y=2.72
+ $X2=5.29 $Y2=2.72
r105 65 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r106 65 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r107 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r108 62 72 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.652 $Y2=2.72
r109 62 64 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=1.61 $Y2=2.72
r110 57 72 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.652 $Y2=2.72
r111 57 59 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r112 55 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 55 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r114 53 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=2.72
+ $X2=1.61 $Y2=2.72
r115 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=2.72
+ $X2=1.83 $Y2=2.72
r116 49 52 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.76 $Y=1.66
+ $X2=5.76 $Y2=2.34
r117 47 86 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.76 $Y=2.635
+ $X2=5.802 $Y2=2.72
r118 47 52 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.76 $Y=2.635
+ $X2=5.76 $Y2=2.34
r119 43 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=2.635
+ $X2=4.87 $Y2=2.72
r120 43 45 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.87 $Y=2.635
+ $X2=4.87 $Y2=2
r121 42 78 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.115 $Y=2.72
+ $X2=3.77 $Y2=2.72
r122 41 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.72
+ $X2=4.87 $Y2=2.72
r123 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.785 $Y=2.72
+ $X2=4.115 $Y2=2.72
r124 37 78 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=2.635
+ $X2=3.77 $Y2=2.72
r125 37 39 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=3.77 $Y=2.635
+ $X2=3.77 $Y2=2
r126 36 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.63 $Y2=2.72
r127 35 78 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=3.77 $Y2=2.72
r128 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=2.755 $Y2=2.72
r129 31 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=2.72
r130 31 33 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=2
r131 30 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.83 $Y2=2.72
r132 29 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.63 $Y2=2.72
r133 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=1.915 $Y2=2.72
r134 25 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.83 $Y=1.66
+ $X2=1.83 $Y2=2.34
r135 23 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.72
r136 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.34
r137 19 72 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.652 $Y=2.635
+ $X2=0.652 $Y2=2.72
r138 19 21 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=0.652 $Y=2.635
+ $X2=0.652 $Y2=2.36
r139 6 52 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.575
+ $Y=1.485 $X2=5.71 $Y2=2.34
r140 6 49 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.575
+ $Y=1.485 $X2=5.71 $Y2=1.66
r141 5 45 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.735
+ $Y=1.485 $X2=4.87 $Y2=2
r142 4 39 150 $w=1.7e-07 $l=7.91675e-07 $layer=licon1_PDIFF $count=4 $X=3.375
+ $Y=1.485 $X2=3.95 $Y2=2
r143 3 33 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.485 $X2=2.67 $Y2=2
r144 2 28 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=1.485 $X2=1.83 $Y2=2.34
r145 2 25 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=1.485 $X2=1.83 $Y2=1.66
r146 1 21 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%Y 1 2 3 4 5 18 22 24 28 30 31 34 36 38 40
+ 42 44 47 48
r92 48 58 16.0818 $w=2.18e-07 $l=3.07e-07 $layer=LI1_cond $X=3.397 $Y=1.555
+ $X2=3.09 $Y2=1.555
r93 47 48 7.94868 $w=4.73e-07 $l=2.55e-07 $layer=LI1_cond $X=3.397 $Y=1.19
+ $X2=3.397 $Y2=1.445
r94 38 46 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=5.29 $Y=1.665
+ $X2=5.29 $Y2=1.555
r95 38 40 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.29 $Y=1.665
+ $X2=5.29 $Y2=2.34
r96 37 44 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=1.555
+ $X2=4.45 $Y2=1.555
r97 36 46 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=1.555
+ $X2=5.29 $Y2=1.555
r98 36 37 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=5.125 $Y=1.555
+ $X2=4.615 $Y2=1.555
r99 32 44 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.45 $Y=1.665
+ $X2=4.45 $Y2=1.555
r100 32 34 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.45 $Y=1.665
+ $X2=4.45 $Y2=2.34
r101 31 48 5.23838 $w=2.18e-07 $l=1e-07 $layer=LI1_cond $X=3.55 $Y=1.555
+ $X2=3.45 $Y2=1.555
r102 30 44 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=1.555
+ $X2=4.45 $Y2=1.555
r103 30 31 38.5021 $w=2.18e-07 $l=7.35e-07 $layer=LI1_cond $X=4.285 $Y=1.555
+ $X2=3.55 $Y2=1.555
r104 28 58 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.09 $Y=2.34
+ $X2=3.09 $Y2=1.665
r105 25 42 2.35378 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=1.555
+ $X2=2.25 $Y2=1.555
r106 24 58 8.64332 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=1.555
+ $X2=3.09 $Y2=1.555
r107 24 25 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=2.925 $Y=1.555
+ $X2=2.415 $Y2=1.555
r108 20 42 4.08154 $w=2.9e-07 $l=1.28452e-07 $layer=LI1_cond $X=2.21 $Y=1.665
+ $X2=2.25 $Y2=1.555
r109 20 22 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=2.21 $Y=1.665
+ $X2=2.21 $Y2=1.785
r110 16 42 4.08154 $w=2.9e-07 $l=1.1e-07 $layer=LI1_cond $X=2.25 $Y=1.445
+ $X2=2.25 $Y2=1.555
r111 16 18 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=2.25 $Y=1.445
+ $X2=2.25 $Y2=0.74
r112 5 46 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.155
+ $Y=1.485 $X2=5.29 $Y2=1.66
r113 5 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.155
+ $Y=1.485 $X2=5.29 $Y2=2.34
r114 4 44 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.485 $X2=4.45 $Y2=1.66
r115 4 34 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.485 $X2=4.45 $Y2=2.34
r116 3 58 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.09 $Y2=1.66
r117 3 28 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.485 $X2=3.09 $Y2=2.34
r118 2 22 300 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_PDIFF $count=2 $X=2.115
+ $Y=1.485 $X2=2.25 $Y2=1.785
r119 1 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.25 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%VGND 1 2 9 13 15 17 22 29 30 33 36
r68 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r69 33 34 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r70 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r71 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r72 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0 $X2=5.29
+ $Y2=0
r73 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.375 $Y=0 $X2=5.75
+ $Y2=0
r74 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r75 26 34 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.83 $Y=0 $X2=0.69
+ $Y2=0
r76 25 26 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r77 23 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.64
+ $Y2=0
r78 23 25 265.203 $w=1.68e-07 $l=4.065e-06 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=4.83 $Y2=0
r79 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=0 $X2=5.29
+ $Y2=0
r80 22 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.205 $Y=0 $X2=4.83
+ $Y2=0
r81 17 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.64
+ $Y2=0
r82 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r83 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r84 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r85 11 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0
r86 11 13 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0.4
r87 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=0.085
+ $X2=0.64 $Y2=0
r88 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.64 $Y=0.085
+ $X2=0.64 $Y2=0.38
r89 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.155
+ $Y=0.235 $X2=5.29 $Y2=0.4
r90 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%A_341_47# 1 2 3 14 19
r24 17 19 4.03881 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=0.42
+ $X2=1.915 $Y2=0.42
r25 12 14 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.67 $Y=0.37
+ $X2=3.51 $Y2=0.37
r26 12 19 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=2.67 $Y=0.37
+ $X2=1.915 $Y2=0.37
r27 3 14 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.235 $X2=3.51 $Y2=0.4
r28 2 12 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.235 $X2=2.67 $Y2=0.4
r29 1 17 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.235 $X2=1.83 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%A_591_47# 1 2 11
c26 11 0 7.99167e-20 $X=4.45 $Y=0.74
r27 8 11 62.6929 $w=2.48e-07 $l=1.36e-06 $layer=LI1_cond $X=3.09 $Y=0.78
+ $X2=4.45 $Y2=0.78
r28 2 11 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.315
+ $Y=0.235 $X2=4.45 $Y2=0.74
r29 1 8 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.09 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_2%A_781_47# 1 2 3 10 14 15 16 20
c39 15 0 1.79953e-19 $X=4.91 $Y=0.735
r40 18 20 11.0305 $w=3.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.72 $Y=0.735
+ $X2=5.72 $Y2=0.4
r41 17 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.035 $Y=0.82
+ $X2=4.91 $Y2=0.82
r42 16 18 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.545 $Y=0.82
+ $X2=5.72 $Y2=0.735
r43 16 17 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.545 $Y=0.82
+ $X2=5.035 $Y2=0.82
r44 15 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=0.735
+ $X2=4.91 $Y2=0.82
r45 14 23 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=4.91 $Y=0.485
+ $X2=4.91 $Y2=0.37
r46 14 15 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=4.91 $Y=0.485
+ $X2=4.91 $Y2=0.735
r47 10 23 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=4.785 $Y=0.37
+ $X2=4.91 $Y2=0.37
r48 10 12 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=4.785 $Y=0.37
+ $X2=4.03 $Y2=0.37
r49 3 20 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.4
r50 2 25 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.735
+ $Y=0.235 $X2=4.87 $Y2=0.74
r51 2 23 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.735
+ $Y=0.235 $X2=4.87 $Y2=0.4
r52 1 12 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.03 $Y2=0.4
.ends


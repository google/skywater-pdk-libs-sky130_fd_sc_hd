* NGSPICE file created from sky130_fd_sc_hd__fa_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_1014_47# B VGND VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=1.482e+12p ps=1.557e+07u
M1001 VGND CIN a_1014_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR a_1271_47# SUM VPB phighvt w=1e+06u l=150000u
+  ad=2.2815e+12p pd=2.109e+07u as=5.4e+11p ps=5.08e+06u
M1003 VGND A a_1451_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1004 a_1014_369# A VPWR VPB phighvt w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=0p ps=0u
M1005 COUT a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1006 a_79_21# B a_456_371# VPB phighvt w=630000u l=150000u
+  ad=2.644e+11p pd=2.11e+06u as=1.8585e+11p ps=1.85e+06u
M1007 a_1451_371# B a_1356_369# VPB phighvt w=630000u l=150000u
+  ad=2.457e+11p pd=2.04e+06u as=2.0725e+11p ps=1.93e+06u
M1008 SUM a_1271_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1356_369# CIN a_1271_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1010 a_79_21# B a_461_47# VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=1.365e+11p ps=1.49e+06u
M1011 VPWR a_79_21# COUT VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 SUM a_1271_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR CIN a_1014_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_658_47# B VGND VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=0p ps=0u
M1015 VGND a_1271_47# SUM VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.03e+11p ps=3.84e+06u
M1016 a_1271_47# a_79_21# a_1014_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1271_47# a_79_21# a_1014_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1018 VGND A a_658_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_658_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.392e+11p ps=3.62e+06u
M1020 VGND a_79_21# COUT VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.51e+11p ps=3.68e+06u
M1021 a_658_47# CIN a_79_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1271_47# SUM VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1014_369# B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_461_47# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1271_47# SUM VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A a_1451_371# VPB phighvt w=630000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 SUM a_1271_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_79_21# COUT VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 COUT a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1451_47# B a_1379_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1031 COUT a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_658_369# CIN a_79_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 SUM a_1271_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_456_371# A VPWR VPB phighvt w=630000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_79_21# COUT VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 COUT a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1379_47# CIN a_1271_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_658_369# B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1014_47# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__a2111o_4.pex.spice
* Created: Tue Sep  1 18:50:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2111O_4%D1 3 5 7 10 12 14 15 16 24
c39 24 0 1.34048e-19 $X=0.92 $Y=1.16
c40 5 0 1.31746e-20 $X=0.56 $Y=0.995
r41 24 25 10.6772 $w=3.16e-07 $l=7e-08 $layer=POLY_cond $X=0.92 $Y=1.16 $X2=0.99
+ $Y2=1.16
r42 23 24 54.9114 $w=3.16e-07 $l=3.6e-07 $layer=POLY_cond $X=0.56 $Y=1.16
+ $X2=0.92 $Y2=1.16
r43 22 23 10.6772 $w=3.16e-07 $l=7e-08 $layer=POLY_cond $X=0.49 $Y=1.16 $X2=0.56
+ $Y2=1.16
r44 20 22 33.557 $w=3.16e-07 $l=2.2e-07 $layer=POLY_cond $X=0.27 $Y=1.16
+ $X2=0.49 $Y2=1.16
r45 15 16 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.227 $Y=1.16
+ $X2=0.227 $Y2=1.53
r46 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r47 12 25 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.16
r48 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r49 8 24 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=1.16
r50 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=1.985
r51 5 23 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=0.995
+ $X2=0.56 $Y2=1.16
r52 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.56 $Y=0.995 $X2=0.56
+ $Y2=0.56
r53 1 22 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r54 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%C1 3 5 7 10 12 14 15 16 17
c49 17 0 1.31746e-20 $X=2.07 $Y=1.19
c50 12 0 1.90293e-19 $X=1.885 $Y=0.995
r51 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.85
+ $Y=1.16 $X2=1.85 $Y2=1.16
r52 24 26 12.4286 $w=3.25e-07 $l=7e-08 $layer=POLY_cond $X=1.78 $Y=1.157
+ $X2=1.85 $Y2=1.157
r53 17 27 8.17863 $w=3.08e-07 $l=2.2e-07 $layer=LI1_cond $X=2.07 $Y=1.13
+ $X2=1.85 $Y2=1.13
r54 16 27 8.92214 $w=3.08e-07 $l=2.4e-07 $layer=LI1_cond $X=1.61 $Y=1.13
+ $X2=1.85 $Y2=1.13
r55 15 16 17.1008 $w=3.08e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=1.13
+ $X2=1.61 $Y2=1.13
r56 12 26 6.2143 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=1.885 $Y=1.157
+ $X2=1.85 $Y2=1.157
r57 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.885 $Y=0.995
+ $X2=1.885 $Y2=0.56
r58 8 24 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=1.78 $Y=1.32 $X2=1.78
+ $Y2=1.157
r59 8 10 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.78 $Y=1.32
+ $X2=1.78 $Y2=1.985
r60 5 24 63.9185 $w=3.25e-07 $l=3.6e-07 $layer=POLY_cond $X=1.42 $Y=1.157
+ $X2=1.78 $Y2=1.157
r61 5 21 12.4286 $w=3.25e-07 $l=7e-08 $layer=POLY_cond $X=1.42 $Y=1.157 $X2=1.35
+ $Y2=1.157
r62 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.42 $Y=0.995 $X2=1.42
+ $Y2=0.56
r63 1 21 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=1.35 $Y=1.32 $X2=1.35
+ $Y2=1.157
r64 1 3 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.35 $Y=1.32 $X2=1.35
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%B1 1 3 6 10 12 14 15 16 24
c48 24 0 1.90293e-19 $X=3.09 $Y=1.16
r49 23 25 10.6531 $w=3.25e-07 $l=6e-08 $layer=POLY_cond $X=3.09 $Y=1.157
+ $X2=3.15 $Y2=1.157
r50 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.16 $X2=3.09 $Y2=1.16
r51 21 23 65.694 $w=3.25e-07 $l=3.7e-07 $layer=POLY_cond $X=2.72 $Y=1.157
+ $X2=3.09 $Y2=1.157
r52 16 24 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=3 $Y=1.13 $X2=3.09
+ $Y2=1.13
r53 15 16 17.1008 $w=3.08e-07 $l=4.6e-07 $layer=LI1_cond $X=2.54 $Y=1.13 $X2=3
+ $Y2=1.13
r54 12 25 33.7348 $w=3.25e-07 $l=1.9e-07 $layer=POLY_cond $X=3.34 $Y=1.157
+ $X2=3.15 $Y2=1.157
r55 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.56
r56 8 25 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=3.15 $Y=1.32 $X2=3.15
+ $Y2=1.157
r57 8 10 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.15 $Y=1.32
+ $X2=3.15 $Y2=1.985
r58 4 21 20.86 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=2.72 $Y=1.32 $X2=2.72
+ $Y2=1.157
r59 4 6 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.72 $Y=1.32 $X2=2.72
+ $Y2=1.985
r60 1 21 62.143 $w=3.25e-07 $l=3.5e-07 $layer=POLY_cond $X=2.37 $Y=1.157
+ $X2=2.72 $Y2=1.157
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=0.995 $X2=2.37
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%A1 1 3 6 8 10 13 15 16 25
c45 16 0 1.66891e-19 $X=4.38 $Y=1.19
c46 6 0 1.29441e-19 $X=3.815 $Y=1.985
r47 23 25 14.4261 $w=3.4e-07 $l=8.5e-08 $layer=POLY_cond $X=4.245 $Y=1.165
+ $X2=4.33 $Y2=1.165
r48 22 23 6.78873 $w=3.4e-07 $l=4e-08 $layer=POLY_cond $X=4.205 $Y=1.165
+ $X2=4.245 $Y2=1.165
r49 21 22 66.1901 $w=3.4e-07 $l=3.9e-07 $layer=POLY_cond $X=3.815 $Y=1.165
+ $X2=4.205 $Y2=1.165
r50 19 21 6.78873 $w=3.4e-07 $l=4e-08 $layer=POLY_cond $X=3.775 $Y=1.165
+ $X2=3.815 $Y2=1.165
r51 16 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.33
+ $Y=1.16 $X2=4.33 $Y2=1.16
r52 15 16 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.92 $Y=1.175
+ $X2=4.33 $Y2=1.175
r53 11 23 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.245 $Y=1.335
+ $X2=4.245 $Y2=1.165
r54 11 13 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.245 $Y=1.335
+ $X2=4.245 $Y2=1.985
r55 8 22 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.205 $Y=0.995
+ $X2=4.205 $Y2=1.165
r56 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.205 $Y=0.995
+ $X2=4.205 $Y2=0.56
r57 4 21 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.815 $Y=1.335
+ $X2=3.815 $Y2=1.165
r58 4 6 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.815 $Y=1.335
+ $X2=3.815 $Y2=1.985
r59 1 19 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.775 $Y=0.995
+ $X2=3.775 $Y2=1.165
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.775 $Y=0.995
+ $X2=3.775 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%A2 1 3 6 8 10 13 15 16 22 23 25
c42 23 0 1.66891e-19 $X=5.615 $Y=1.16
c43 22 0 1.69924e-19 $X=5.46 $Y=1.16
r44 21 23 23.5678 $w=3.17e-07 $l=1.55e-07 $layer=POLY_cond $X=5.46 $Y=1.16
+ $X2=5.615 $Y2=1.16
r45 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.46
+ $Y=1.16 $X2=5.46 $Y2=1.16
r46 19 21 41.8139 $w=3.17e-07 $l=2.75e-07 $layer=POLY_cond $X=5.185 $Y=1.16
+ $X2=5.46 $Y2=1.16
r47 16 22 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=5.31 $Y=1.175
+ $X2=5.46 $Y2=1.175
r48 15 16 25.7864 $w=1.98e-07 $l=4.65e-07 $layer=LI1_cond $X=4.845 $Y=1.175
+ $X2=5.31 $Y2=1.175
r49 15 25 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=4.845 $Y=1.175
+ $X2=4.84 $Y2=1.175
r50 11 23 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.615 $Y=1.325
+ $X2=5.615 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.615 $Y=1.325
+ $X2=5.615 $Y2=1.985
r52 8 23 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.615 $Y=0.995
+ $X2=5.615 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.615 $Y=0.995
+ $X2=5.615 $Y2=0.56
r54 4 19 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.185 $Y=1.325
+ $X2=5.185 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.185 $Y=1.325
+ $X2=5.185 $Y2=1.985
r56 1 19 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.185 $Y=0.995
+ $X2=5.185 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.185 $Y=0.995
+ $X2=5.185 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%A_44_47# 1 2 3 4 5 6 19 21 24 26 28 31 33
+ 35 38 40 42 45 49 53 55 56 59 61 65 67 69 72 75 77 78 80 81 86 92 93 104
c183 104 0 1.69924e-19 $X=7.335 $Y=1.16
r184 101 102 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.475 $Y=1.16
+ $X2=6.905 $Y2=1.16
r185 87 104 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.155 $Y=1.16
+ $X2=7.335 $Y2=1.16
r186 87 102 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.155 $Y=1.16
+ $X2=6.905 $Y2=1.16
r187 86 87 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.155
+ $Y=1.16 $X2=7.155 $Y2=1.16
r188 84 101 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.135 $Y=1.16
+ $X2=6.475 $Y2=1.16
r189 84 98 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.135 $Y=1.16
+ $X2=6.045 $Y2=1.16
r190 83 86 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.135 $Y=1.16
+ $X2=7.155 $Y2=1.16
r191 83 84 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.135
+ $Y=1.16 $X2=6.135 $Y2=1.16
r192 81 83 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.975 $Y=1.16
+ $X2=6.135 $Y2=1.16
r193 79 81 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.885 $Y=1.245
+ $X2=5.975 $Y2=1.16
r194 79 80 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=5.885 $Y=1.245
+ $X2=5.885 $Y2=1.445
r195 77 80 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=5.795 $Y=1.535
+ $X2=5.885 $Y2=1.445
r196 77 78 131.859 $w=1.78e-07 $l=2.14e-06 $layer=LI1_cond $X=5.795 $Y=1.535
+ $X2=3.655 $Y2=1.535
r197 73 95 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.655 $Y=0.35
+ $X2=3.56 $Y2=0.35
r198 73 75 44.3636 $w=1.88e-07 $l=7.6e-07 $layer=LI1_cond $X=3.655 $Y=0.35
+ $X2=4.415 $Y2=0.35
r199 72 78 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.56 $Y=1.445
+ $X2=3.655 $Y2=1.535
r200 71 97 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.56 $Y=0.805
+ $X2=3.56 $Y2=0.71
r201 71 72 37.3589 $w=1.88e-07 $l=6.4e-07 $layer=LI1_cond $X=3.56 $Y=0.805
+ $X2=3.56 $Y2=1.445
r202 70 97 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.56 $Y=0.615
+ $X2=3.56 $Y2=0.71
r203 69 95 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.56 $Y=0.445
+ $X2=3.56 $Y2=0.35
r204 69 70 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.56 $Y=0.445
+ $X2=3.56 $Y2=0.615
r205 68 93 5.93234 $w=1.9e-07 $l=1.13e-07 $layer=LI1_cond $X=2.24 $Y=0.71
+ $X2=2.127 $Y2=0.71
r206 67 97 1.34256 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.465 $Y=0.71
+ $X2=3.56 $Y2=0.71
r207 67 68 71.5072 $w=1.88e-07 $l=1.225e-06 $layer=LI1_cond $X=3.465 $Y=0.71
+ $X2=2.24 $Y2=0.71
r208 63 93 0.741404 $w=2.25e-07 $l=9.5e-08 $layer=LI1_cond $X=2.127 $Y=0.615
+ $X2=2.127 $Y2=0.71
r209 63 65 9.98784 $w=2.23e-07 $l=1.95e-07 $layer=LI1_cond $X=2.127 $Y=0.615
+ $X2=2.127 $Y2=0.42
r210 62 92 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=1.34 $Y=0.71
+ $X2=1.225 $Y2=0.71
r211 61 93 5.93234 $w=1.9e-07 $l=1.12e-07 $layer=LI1_cond $X=2.015 $Y=0.71
+ $X2=2.127 $Y2=0.71
r212 61 62 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=2.015 $Y=0.71
+ $X2=1.34 $Y2=0.71
r213 57 92 0.47666 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=1.225 $Y=0.615
+ $X2=1.225 $Y2=0.71
r214 57 59 9.77071 $w=2.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.225 $Y=0.615
+ $X2=1.225 $Y2=0.42
r215 55 92 6.30264 $w=1.8e-07 $l=1.19896e-07 $layer=LI1_cond $X=1.11 $Y=0.72
+ $X2=1.225 $Y2=0.71
r216 55 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.11 $Y=0.72
+ $X2=0.87 $Y2=0.72
r217 51 56 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=0.72
+ $X2=0.87 $Y2=0.72
r218 51 53 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.705 $Y=0.805
+ $X2=0.705 $Y2=1.67
r219 47 51 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.31 $Y=0.72
+ $X2=0.705 $Y2=0.72
r220 47 49 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.31 $Y=0.635
+ $X2=0.31 $Y2=0.42
r221 43 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.335 $Y=1.325
+ $X2=7.335 $Y2=1.16
r222 43 45 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.335 $Y=1.325
+ $X2=7.335 $Y2=1.985
r223 40 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.335 $Y=0.995
+ $X2=7.335 $Y2=1.16
r224 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.335 $Y=0.995
+ $X2=7.335 $Y2=0.56
r225 36 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.325
+ $X2=6.905 $Y2=1.16
r226 36 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.905 $Y=1.325
+ $X2=6.905 $Y2=1.985
r227 33 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=0.995
+ $X2=6.905 $Y2=1.16
r228 33 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.905 $Y=0.995
+ $X2=6.905 $Y2=0.56
r229 29 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.475 $Y=1.325
+ $X2=6.475 $Y2=1.16
r230 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.475 $Y=1.325
+ $X2=6.475 $Y2=1.985
r231 26 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.475 $Y=0.995
+ $X2=6.475 $Y2=1.16
r232 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.475 $Y=0.995
+ $X2=6.475 $Y2=0.56
r233 22 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.325
+ $X2=6.045 $Y2=1.16
r234 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.045 $Y=1.325
+ $X2=6.045 $Y2=1.985
r235 19 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=0.995
+ $X2=6.045 $Y2=1.16
r236 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.045 $Y=0.995
+ $X2=6.045 $Y2=0.56
r237 6 53 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.705 $Y2=1.67
r238 5 75 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.28
+ $Y=0.235 $X2=4.415 $Y2=0.36
r239 4 97 182 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.56 $Y2=0.76
r240 4 95 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.56 $Y2=0.42
r241 3 65 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.235 $X2=2.1 $Y2=0.42
r242 2 59 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.205 $Y2=0.42
r243 1 49 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.22
+ $Y=0.235 $X2=0.345 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%A_30_297# 1 2 3 12 14 15 18 20 24 27
c38 18 0 1.34048e-19 $X=1.135 $Y=1.62
r39 22 24 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.03 $Y=2.295
+ $X2=2.03 $Y2=1.96
r40 21 27 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.23 $Y=2.38
+ $X2=1.135 $Y2=2.38
r41 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.9 $Y=2.38
+ $X2=2.03 $Y2=2.295
r42 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.9 $Y=2.38 $X2=1.23
+ $Y2=2.38
r43 16 27 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=2.295
+ $X2=1.135 $Y2=2.38
r44 16 18 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=1.135 $Y=2.295
+ $X2=1.135 $Y2=1.62
r45 14 27 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.04 $Y=2.38
+ $X2=1.135 $Y2=2.38
r46 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.04 $Y=2.38
+ $X2=0.37 $Y2=2.38
r47 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.24 $Y=2.295
+ $X2=0.37 $Y2=2.38
r48 10 12 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=2.295
+ $X2=0.24 $Y2=1.96
r49 3 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.855
+ $Y=1.485 $X2=1.99 $Y2=1.96
r50 2 27 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.135 $Y2=2.3
r51 2 18 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.485 $X2=1.135 $Y2=1.62
r52 1 12 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=1.485 $X2=0.275 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%A_285_297# 1 2 9 11 12 16
c36 16 0 1.29441e-19 $X=2.935 $Y=1.62
r37 11 16 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.845 $Y=1.54
+ $X2=2.972 $Y2=1.54
r38 11 12 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.845 $Y=1.54
+ $X2=1.73 $Y2=1.54
r39 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.625
+ $X2=1.73 $Y2=1.54
r40 7 9 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.565 $Y=1.625
+ $X2=1.565 $Y2=1.67
r41 2 16 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=2.795
+ $Y=1.485 $X2=2.935 $Y2=1.62
r42 1 9 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=1.425
+ $Y=1.485 $X2=1.565 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%A_477_297# 1 2 3 4 15 17 18 19 22 23 27 29
+ 36 38
r63 30 36 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.625 $Y=1.895 $X2=4.495
+ $Y2=1.895
r64 29 38 3.27269 $w=2e-07 $l=9.2e-08 $layer=LI1_cond $X=5.31 $Y=1.895 $X2=5.402
+ $Y2=1.895
r65 29 30 37.9864 $w=1.98e-07 $l=6.85e-07 $layer=LI1_cond $X=5.31 $Y=1.895
+ $X2=4.625 $Y2=1.895
r66 25 36 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=4.495 $Y=1.995
+ $X2=4.495 $Y2=1.895
r67 25 27 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=4.495 $Y=1.995
+ $X2=4.495 $Y2=2.25
r68 24 34 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.65 $Y=1.895
+ $X2=3.485 $Y2=1.895
r69 23 36 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.365 $Y=1.895 $X2=4.495
+ $Y2=1.895
r70 23 24 39.65 $w=1.98e-07 $l=7.15e-07 $layer=LI1_cond $X=4.365 $Y=1.895
+ $X2=3.65 $Y2=1.895
r71 20 22 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=3.485 $Y=2.295
+ $X2=3.485 $Y2=2.24
r72 19 34 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=3.485 $Y=1.995
+ $X2=3.485 $Y2=1.895
r73 19 22 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.485 $Y=1.995
+ $X2=3.485 $Y2=2.24
r74 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.32 $Y=2.38
+ $X2=3.485 $Y2=2.295
r75 17 18 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.32 $Y=2.38
+ $X2=2.675 $Y2=2.38
r76 13 18 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=2.507 $Y=2.295
+ $X2=2.675 $Y2=2.38
r77 13 15 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=2.507 $Y=2.295
+ $X2=2.507 $Y2=1.88
r78 4 38 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=5.26
+ $Y=1.485 $X2=5.4 $Y2=1.96
r79 3 36 600 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.485 $X2=4.455 $Y2=1.91
r80 3 27 600 $w=1.7e-07 $l=8.29759e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.485 $X2=4.455 $Y2=2.25
r81 2 34 600 $w=1.7e-07 $l=5.29268e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.485 $Y2=1.9
r82 2 22 600 $w=1.7e-07 $l=8.754e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.485 $Y2=2.24
r83 1 15 300 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=2 $X=2.385
+ $Y=1.485 $X2=2.51 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%VPWR 1 2 3 4 5 18 20 24 28 32 34 36 38 40
+ 45 50 55 61 64 67 70 74
r117 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r118 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r119 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r121 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r122 61 62 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r123 59 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r124 59 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r125 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r126 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.855 $Y=2.72
+ $X2=6.69 $Y2=2.72
r127 56 58 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.855 $Y=2.72
+ $X2=7.13 $Y2=2.72
r128 55 73 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=7.385 $Y=2.72
+ $X2=7.602 $Y2=2.72
r129 55 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.385 $Y=2.72
+ $X2=7.13 $Y2=2.72
r130 54 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r131 54 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r132 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r133 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.995 $Y=2.72
+ $X2=5.83 $Y2=2.72
r134 51 53 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.995 $Y=2.72
+ $X2=6.21 $Y2=2.72
r135 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.525 $Y=2.72
+ $X2=6.69 $Y2=2.72
r136 50 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.525 $Y=2.72
+ $X2=6.21 $Y2=2.72
r137 49 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r138 49 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r139 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r140 46 64 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=5.14 $Y=2.72
+ $X2=4.972 $Y2=2.72
r141 46 48 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.14 $Y=2.72
+ $X2=5.29 $Y2=2.72
r142 45 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=2.72
+ $X2=5.83 $Y2=2.72
r143 45 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.665 $Y=2.72
+ $X2=5.29 $Y2=2.72
r144 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=2.72
+ $X2=4.03 $Y2=2.72
r145 40 42 237.15 $w=1.68e-07 $l=3.635e-06 $layer=LI1_cond $X=3.865 $Y=2.72
+ $X2=0.23 $Y2=2.72
r146 38 62 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r147 38 42 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r148 34 73 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.55 $Y=2.635
+ $X2=7.602 $Y2=2.72
r149 34 36 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=7.55 $Y=2.635
+ $X2=7.55 $Y2=1.97
r150 30 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.69 $Y=2.635
+ $X2=6.69 $Y2=2.72
r151 30 32 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=6.69 $Y=2.635
+ $X2=6.69 $Y2=1.97
r152 26 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=2.635
+ $X2=5.83 $Y2=2.72
r153 26 28 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=5.83 $Y=2.635
+ $X2=5.83 $Y2=1.885
r154 22 64 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.972 $Y=2.635
+ $X2=4.972 $Y2=2.72
r155 22 24 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=4.972 $Y=2.635
+ $X2=4.972 $Y2=2.34
r156 21 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=2.72
+ $X2=4.03 $Y2=2.72
r157 20 64 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.805 $Y=2.72
+ $X2=4.972 $Y2=2.72
r158 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.805 $Y=2.72
+ $X2=4.195 $Y2=2.72
r159 16 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.635
+ $X2=4.03 $Y2=2.72
r160 16 18 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.03 $Y=2.635
+ $X2=4.03 $Y2=2.25
r161 5 36 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=7.41
+ $Y=1.485 $X2=7.55 $Y2=1.97
r162 4 32 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=6.55
+ $Y=1.485 $X2=6.69 $Y2=1.97
r163 3 28 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=5.69
+ $Y=1.485 $X2=5.83 $Y2=1.885
r164 2 24 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.485 $X2=4.975 $Y2=2.34
r165 1 18 600 $w=1.7e-07 $l=8.32061e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.485 $X2=4.03 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35 37
+ 38 39 40 41 47 48 50
r64 47 50 2.11673 $w=2.43e-07 $l=4.5e-08 $layer=LI1_cond $X=7.612 $Y=0.805
+ $X2=7.612 $Y2=0.85
r65 41 48 2.91961 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=7.612 $Y=1.55
+ $X2=7.612 $Y2=1.465
r66 41 48 0.470385 $w=2.43e-07 $l=1e-08 $layer=LI1_cond $X=7.612 $Y=1.455
+ $X2=7.612 $Y2=1.465
r67 40 41 12.4652 $w=2.43e-07 $l=2.65e-07 $layer=LI1_cond $X=7.612 $Y=1.19
+ $X2=7.612 $Y2=1.455
r68 39 47 2.91961 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=7.612 $Y=0.72
+ $X2=7.612 $Y2=0.805
r69 39 40 15.0523 $w=2.43e-07 $l=3.2e-07 $layer=LI1_cond $X=7.612 $Y=0.87
+ $X2=7.612 $Y2=1.19
r70 39 50 0.94077 $w=2.43e-07 $l=2e-08 $layer=LI1_cond $X=7.612 $Y=0.87
+ $X2=7.612 $Y2=0.85
r71 36 38 4.74942 $w=2.1e-07 $l=1.13248e-07 $layer=LI1_cond $X=7.215 $Y=1.55
+ $X2=7.12 $Y2=1.59
r72 35 41 4.1905 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=7.49 $Y=1.55
+ $X2=7.612 $Y2=1.55
r73 35 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.49 $Y=1.55
+ $X2=7.215 $Y2=1.55
r74 34 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.215 $Y=0.72
+ $X2=7.12 $Y2=0.72
r75 33 39 4.1905 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=7.49 $Y=0.72
+ $X2=7.612 $Y2=0.72
r76 33 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.49 $Y=0.72
+ $X2=7.215 $Y2=0.72
r77 29 38 1.70532 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=7.12 $Y=1.715
+ $X2=7.12 $Y2=1.59
r78 29 31 7.00478 $w=1.88e-07 $l=1.2e-07 $layer=LI1_cond $X=7.12 $Y=1.715
+ $X2=7.12 $Y2=1.835
r79 25 37 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.12 $Y=0.635
+ $X2=7.12 $Y2=0.72
r80 25 27 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=7.12 $Y=0.635
+ $X2=7.12 $Y2=0.42
r81 23 38 4.74942 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=7.025 $Y=1.59
+ $X2=7.12 $Y2=1.59
r82 23 24 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.025 $Y=1.59
+ $X2=6.355 $Y2=1.59
r83 21 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.025 $Y=0.72
+ $X2=7.12 $Y2=0.72
r84 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.025 $Y=0.72
+ $X2=6.355 $Y2=0.72
r85 17 24 6.98266 $w=2.5e-07 $l=1.65831e-07 $layer=LI1_cond $X=6.26 $Y=1.715
+ $X2=6.355 $Y2=1.59
r86 17 19 7.00478 $w=1.88e-07 $l=1.2e-07 $layer=LI1_cond $X=6.26 $Y=1.715
+ $X2=6.26 $Y2=1.835
r87 13 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.26 $Y=0.635
+ $X2=6.355 $Y2=0.72
r88 13 15 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=6.26 $Y=0.635
+ $X2=6.26 $Y2=0.42
r89 4 31 300 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=2 $X=6.98
+ $Y=1.485 $X2=7.12 $Y2=1.835
r90 3 19 300 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=2 $X=6.12
+ $Y=1.485 $X2=6.26 $Y2=1.835
r91 2 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.98
+ $Y=0.235 $X2=7.12 $Y2=0.42
r92 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.235 $X2=6.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%VGND 1 2 3 4 5 6 7 26 30 34 38 42 44 46 48
+ 50 60 65 70 75 81 84 89 95 97 100 103 107
r135 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r136 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r137 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r138 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r139 94 95 10.2686 $w=5.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.105 $Y=0.18
+ $X2=3.295 $Y2=0.18
r140 91 94 2.59526 $w=5.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.99 $Y=0.18
+ $X2=3.105 $Y2=0.18
r141 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r142 88 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r143 87 91 10.3811 $w=5.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=0.18
+ $X2=2.99 $Y2=0.18
r144 87 89 8.46316 $w=5.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.53 $Y=0.18
+ $X2=2.42 $Y2=0.18
r145 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r146 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r147 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r148 79 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r149 79 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.67 $Y2=0
r150 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r151 76 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.855 $Y=0
+ $X2=6.69 $Y2=0
r152 76 78 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.855 $Y=0
+ $X2=7.13 $Y2=0
r153 75 106 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=7.385 $Y=0
+ $X2=7.602 $Y2=0
r154 75 78 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.385 $Y=0
+ $X2=7.13 $Y2=0
r155 74 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r156 74 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r157 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r158 71 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.995 $Y=0
+ $X2=5.83 $Y2=0
r159 71 73 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.995 $Y=0
+ $X2=6.21 $Y2=0
r160 70 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.525 $Y=0
+ $X2=6.69 $Y2=0
r161 70 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.525 $Y=0
+ $X2=6.21 $Y2=0
r162 69 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r163 69 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r164 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r165 66 97 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=4.972
+ $Y2=0
r166 66 68 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.29
+ $Y2=0
r167 65 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0
+ $X2=5.83 $Y2=0
r168 65 68 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.665 $Y=0
+ $X2=5.29 $Y2=0
r169 64 98 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.83 $Y2=0
r170 64 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r171 63 95 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=3.295 $Y2=0
r172 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r173 60 97 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.805 $Y=0
+ $X2=4.972 $Y2=0
r174 60 63 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=4.805 $Y=0
+ $X2=3.45 $Y2=0
r175 59 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r176 59 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r177 58 89 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.42
+ $Y2=0
r178 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r179 56 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.675
+ $Y2=0
r180 56 58 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=2.07
+ $Y2=0
r181 54 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r182 54 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r183 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r184 51 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=0.775
+ $Y2=0
r185 51 53 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=1.15
+ $Y2=0
r186 50 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.675
+ $Y2=0
r187 50 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.15
+ $Y2=0
r188 48 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r189 44 106 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.55 $Y=0.085
+ $X2=7.602 $Y2=0
r190 44 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.55 $Y=0.085
+ $X2=7.55 $Y2=0.38
r191 40 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.69 $Y=0.085
+ $X2=6.69 $Y2=0
r192 40 42 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.69 $Y=0.085
+ $X2=6.69 $Y2=0.36
r193 36 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=0.085
+ $X2=5.83 $Y2=0
r194 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.83 $Y=0.085
+ $X2=5.83 $Y2=0.36
r195 32 97 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.972 $Y=0.085
+ $X2=4.972 $Y2=0
r196 32 34 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=4.972 $Y=0.085
+ $X2=4.972 $Y2=0.36
r197 28 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0
r198 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0.36
r199 24 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.085
+ $X2=0.775 $Y2=0
r200 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.775 $Y=0.085
+ $X2=0.775 $Y2=0.38
r201 7 46 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.235 $X2=7.55 $Y2=0.38
r202 6 42 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=6.55
+ $Y=0.235 $X2=6.69 $Y2=0.36
r203 5 38 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.69
+ $Y=0.235 $X2=5.83 $Y2=0.36
r204 4 34 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.83
+ $Y=0.235 $X2=4.975 $Y2=0.36
r205 3 94 91 $w=1.7e-07 $l=7.19792e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.235 $X2=3.105 $Y2=0.36
r206 2 30 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.675 $Y2=0.36
r207 1 26 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.235 $X2=0.775 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_4%A_770_47# 1 2 7 13
r21 11 13 11.6904 $w=1.83e-07 $l=1.95e-07 $layer=LI1_cond $X=5.402 $Y=0.615
+ $X2=5.402 $Y2=0.42
r22 7 11 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=5.31 $Y=0.7
+ $X2=5.402 $Y2=0.615
r23 7 9 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=5.31 $Y=0.7 $X2=3.99
+ $Y2=0.7
r24 2 13 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.26
+ $Y=0.235 $X2=5.4 $Y2=0.42
r25 1 9 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=3.85
+ $Y=0.235 $X2=3.99 $Y2=0.7
.ends


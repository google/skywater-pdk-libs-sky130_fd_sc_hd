* File: sky130_fd_sc_hd__or4b_2.spice
* Created: Tue Sep  1 19:28:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or4b_2.pex.spice"
.subckt sky130_fd_sc_hd__or4b_2  VNB VPB D_N A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_D_N_M1001_g N_A_27_53#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=8.568 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1001_d N_A_176_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_176_21#_M1004_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1006 N_A_176_21#_M1006_d N_A_M1006_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0787009 PD=0.75 PS=0.773271 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75001.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_A_176_21#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0693 PD=0.69 PS=0.75 NRD=0 NRS=15.708 M=1 R=2.8 SA=75002.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1000 N_A_176_21#_M1000_d N_C_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_27_53#_M1012_g N_A_176_21#_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_D_N_M1007_g N_A_27_53#_M1007_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.100149 AS=0.1092 PD=0.887324 PS=1.36 NRD=86.0299 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1007_d N_A_176_21#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.238451 AS=0.135 PD=2.11268 PS=1.27 NRD=12.7853 NRS=0 M=1 R=6.66667
+ SA=75000.4 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_176_21#_M1011_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.237113 AS=0.135 PD=2.10563 PS=1.27 NRD=12.7853 NRS=0 M=1 R=6.66667
+ SA=75000.8 SB=75001 A=0.15 P=2.3 MULT=1
MM1002 A_387_297# N_A_M1002_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0693
+ AS=0.0995873 PD=0.75 PS=0.884366 NRD=51.5943 NRS=85.4192 M=1 R=2.8 SA=75001.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1010 A_483_297# N_B_M1010_g A_387_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0693 PD=0.63 PS=0.75 NRD=23.443 NRS=51.5943 M=1 R=2.8 SA=75002.1 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1013 A_555_297# N_C_M1013_g A_483_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.0693
+ AS=0.0441 PD=0.75 PS=0.63 NRD=51.5943 NRS=23.443 M=1 R=2.8 SA=75002.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_176_21#_M1005_d N_A_27_53#_M1005_g A_555_297# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0693 PD=1.36 PS=0.75 NRD=0 NRS=51.5943 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
DX14_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__or4b_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nand2_4.pex.spice
* Created: Tue Sep  1 19:15:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND2_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 47
r90 45 47 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.73 $Y2=1.16
r91 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r92 43 45 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r93 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r94 41 42 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r95 38 41 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r96 32 46 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.2
+ $X2=1.52 $Y2=1.2
r97 31 46 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.2
+ $X2=1.52 $Y2=1.2
r98 30 31 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.2
+ $X2=1.155 $Y2=1.2
r99 29 30 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.2
+ $X2=0.695 $Y2=1.2
r100 29 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r101 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r102 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r103 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r104 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r105 18 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r106 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r107 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r108 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r109 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r110 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r111 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r112 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r113 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r114 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r115 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r116 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 42
c72 1 0 1.56657e-19 $X=2.15 $Y=0.995
r73 40 42 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.2 $Y=1.16 $X2=3.41
+ $Y2=1.16
r74 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.2 $Y=1.16
+ $X2=3.2 $Y2=1.16
r75 38 40 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.99 $Y=1.16 $X2=3.2
+ $Y2=1.16
r76 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r77 35 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r78 30 31 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=3.455 $Y=1.2
+ $X2=3.915 $Y2=1.2
r79 30 41 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.455 $Y=1.2
+ $X2=3.2 $Y2=1.2
r80 29 41 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=2.995 $Y=1.2
+ $X2=3.2 $Y2=1.2
r81 25 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r82 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r83 22 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r84 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r85 18 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r86 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r87 15 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r88 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r89 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r90 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r91 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r92 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r93 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r94 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
r95 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r96 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995 $X2=2.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_4%VPWR 1 2 3 4 5 16 18 24 28 32 36 39 40 42 43
+ 45 46 48 49 50 66 67
r65 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r66 64 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r69 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r74 52 70 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r75 52 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 50 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 50 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 48 63 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.45 $Y2=2.72
r79 48 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.66 $Y2=2.72
r80 47 66 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.91 $Y2=2.72
r81 47 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.66 $Y2=2.72
r82 45 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.53 $Y2=2.72
r83 45 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.78 $Y2=2.72
r84 44 63 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 44 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.78 $Y2=2.72
r86 42 57 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r87 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.94 $Y2=2.72
r88 41 60 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.94 $Y2=2.72
r90 39 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72 $X2=1.1
+ $Y2=2.72
r92 38 57 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72 $X2=1.1
+ $Y2=2.72
r94 34 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=2.635
+ $X2=3.66 $Y2=2.72
r95 34 36 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.66 $Y=2.635
+ $X2=3.66 $Y2=2
r96 30 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r97 30 32 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r98 26 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r99 26 28 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r100 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r101 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r102 18 21 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r103 16 70 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r104 16 21 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r105 5 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2
r106 4 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r107 3 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r108 2 24 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r109 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r110 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_4%Y 1 2 3 4 5 6 19 21 23 27 29 31 32 35 39 41
+ 42 43 45 50 55
r87 62 64 0.91215 $w=5.35e-07 $l=4e-08 $layer=LI1_cond $X=2.32 $Y=1.37 $X2=2.36
+ $Y2=1.37
r88 55 62 5.58692 $w=5.35e-07 $l=2.45e-07 $layer=LI1_cond $X=2.075 $Y=1.37
+ $X2=2.32 $Y2=1.37
r89 43 54 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=1.665 $X2=3.2
+ $Y2=1.58
r90 43 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.2 $Y=1.665
+ $X2=3.2 $Y2=2.34
r91 42 64 9.93083 $w=5.35e-07 $l=2.80624e-07 $layer=LI1_cond $X=2.525 $Y=1.58
+ $X2=2.36 $Y2=1.37
r92 41 54 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=1.58
+ $X2=3.2 $Y2=1.58
r93 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.035 $Y=1.58
+ $X2=2.525 $Y2=1.58
r94 37 52 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.445 $Y=0.72
+ $X2=2.32 $Y2=0.72
r95 37 39 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.445 $Y=0.72
+ $X2=3.2 $Y2=0.72
r96 33 64 3.564 $w=3.3e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=1.665 $X2=2.36
+ $Y2=1.37
r97 33 35 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=2.34
r98 32 62 5.20553 $w=2.5e-07 $l=2.95e-07 $layer=LI1_cond $X=2.32 $Y=1.075
+ $X2=2.32 $Y2=1.37
r99 31 52 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=0.805
+ $X2=2.32 $Y2=0.72
r100 31 32 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.32 $Y=0.805
+ $X2=2.32 $Y2=1.075
r101 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.58
+ $X2=1.52 $Y2=1.58
r102 29 55 9.93083 $w=5.35e-07 $l=2.80624e-07 $layer=LI1_cond $X=1.91 $Y=1.58
+ $X2=2.075 $Y2=1.37
r103 29 30 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.91 $Y=1.58
+ $X2=1.685 $Y2=1.58
r104 25 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.58
r105 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r106 24 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.58
+ $X2=0.68 $Y2=1.58
r107 23 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.58
+ $X2=1.52 $Y2=1.58
r108 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.58
+ $X2=0.845 $Y2=1.58
r109 19 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.58
r110 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r111 6 54 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.66
r112 6 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.34
r113 5 64 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.66
r114 5 35 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.34
r115 4 50 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r116 4 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r117 3 48 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r118 3 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r119 2 39 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.72
r120 1 52 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 28 29 30
+ 34 36 38
c75 29 0 1.56657e-19 $X=1.9 $Y=0.715
r76 34 44 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.66 $Y=0.465
+ $X2=3.66 $Y2=0.36
r77 34 36 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.66 $Y=0.465
+ $X2=3.66 $Y2=0.72
r78 31 40 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=0.36
+ $X2=1.9 $Y2=0.36
r79 31 33 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.36
+ $X2=2.78 $Y2=0.36
r80 30 44 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.535 $Y=0.36
+ $X2=3.66 $Y2=0.36
r81 30 33 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=3.535 $Y=0.36
+ $X2=2.78 $Y2=0.36
r82 29 42 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=1.9 $Y=0.715 $X2=1.9
+ $Y2=0.81
r83 28 40 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.9 $Y=0.465 $X2=1.9
+ $Y2=0.36
r84 28 29 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.9 $Y=0.465 $X2=1.9
+ $Y2=0.715
r85 27 38 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0.81
+ $X2=1.1 $Y2=0.81
r86 26 42 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=1.775 $Y=0.81
+ $X2=1.9 $Y2=0.81
r87 26 27 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=0.81
+ $X2=1.265 $Y2=0.81
r88 22 38 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=1.1 $Y=0.715 $X2=1.1
+ $Y2=0.81
r89 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=0.715 $X2=1.1
+ $Y2=0.38
r90 20 38 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.81
+ $X2=1.1 $Y2=0.81
r91 20 21 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.81
+ $X2=0.425 $Y2=0.81
r92 16 21 7.51555 $w=1.9e-07 $l=2.102e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.425 $Y2=0.81
r93 16 18 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.257 $Y2=0.38
r94 5 44 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.38
r95 5 36 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.72
r96 4 33 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.38
r97 3 42 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.72
r98 3 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r99 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r100 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_4%VGND 1 2 9 13 16 17 19 20 21 34 35
r55 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r56 32 35 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r57 31 34 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r58 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r59 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r60 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 21 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r62 21 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r63 19 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.15
+ $Y2=0
r64 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.52
+ $Y2=0
r65 18 31 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.61
+ $Y2=0
r66 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.52
+ $Y2=0
r67 16 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r68 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r69 15 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=1.15
+ $Y2=0
r70 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r71 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r72 11 13 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.38
r73 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r74 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0.38
r75 2 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r76 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


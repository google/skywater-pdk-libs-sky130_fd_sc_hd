# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlxbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.955000 1.785000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 0.415000 5.480000 0.745000 ;
        RECT 5.140000 1.670000 5.480000 2.465000 ;
        RECT 5.310000 0.745000 5.480000 1.670000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555000 0.255000 6.815000 0.825000 ;
        RECT 6.555000 1.505000 6.815000 2.465000 ;
        RECT 6.625000 0.825000 6.815000 1.505000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.900000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.875000  0.085000 2.230000 0.445000 ;
        RECT 3.765000  0.085000 4.095000 0.610000 ;
        RECT 4.640000  0.085000 4.970000 0.495000 ;
        RECT 6.090000  0.085000 6.385000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.900000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.980000 1.835000 2.295000 2.635000 ;
        RECT 3.780000 2.175000 3.950000 2.635000 ;
        RECT 4.720000 1.830000 4.970000 2.635000 ;
        RECT 6.090000 1.835000 6.385000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.780000 0.805000 ;
      RECT 0.175000 1.795000 0.780000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.610000 0.805000 0.780000 1.070000 ;
      RECT 0.610000 1.070000 0.840000 1.400000 ;
      RECT 0.610000 1.400000 0.780000 1.795000 ;
      RECT 1.015000 0.345000 1.185000 1.685000 ;
      RECT 1.015000 1.685000 1.240000 2.465000 ;
      RECT 1.480000 1.495000 2.165000 1.665000 ;
      RECT 1.480000 1.665000 1.810000 2.415000 ;
      RECT 1.535000 0.345000 1.705000 0.615000 ;
      RECT 1.535000 0.615000 2.165000 0.785000 ;
      RECT 1.995000 0.785000 2.165000 0.905000 ;
      RECT 1.995000 0.905000 2.365000 1.235000 ;
      RECT 1.995000 1.235000 2.165000 1.495000 ;
      RECT 2.495000 1.355000 2.780000 2.005000 ;
      RECT 2.565000 0.705000 3.120000 1.035000 ;
      RECT 2.790000 0.365000 3.525000 0.535000 ;
      RECT 2.920000 2.105000 3.620000 2.115000 ;
      RECT 2.920000 2.115000 3.615000 2.130000 ;
      RECT 2.920000 2.130000 3.610000 2.275000 ;
      RECT 2.950000 1.035000 3.120000 1.415000 ;
      RECT 2.950000 1.415000 3.290000 1.910000 ;
      RECT 3.355000 0.535000 3.525000 0.995000 ;
      RECT 3.355000 0.995000 4.225000 1.165000 ;
      RECT 3.360000 2.075000 3.630000 2.090000 ;
      RECT 3.360000 2.090000 3.625000 2.105000 ;
      RECT 3.375000 2.060000 3.630000 2.075000 ;
      RECT 3.420000 2.030000 3.630000 2.060000 ;
      RECT 3.430000 2.015000 3.630000 2.030000 ;
      RECT 3.460000 1.165000 4.225000 1.325000 ;
      RECT 3.460000 1.325000 3.630000 2.015000 ;
      RECT 3.800000 1.535000 4.580000 1.620000 ;
      RECT 3.800000 1.620000 4.550000 1.865000 ;
      RECT 4.300000 0.415000 4.470000 0.660000 ;
      RECT 4.300000 0.660000 4.580000 0.840000 ;
      RECT 4.300000 1.865000 4.550000 2.435000 ;
      RECT 4.395000 0.840000 4.580000 0.995000 ;
      RECT 4.395000 0.995000 5.140000 1.325000 ;
      RECT 4.395000 1.325000 4.580000 1.535000 ;
      RECT 5.660000 0.255000 5.910000 0.995000 ;
      RECT 5.660000 0.995000 6.455000 1.325000 ;
      RECT 5.660000 1.325000 5.910000 2.465000 ;
    LAYER mcon ;
      RECT 0.610000 1.445000 0.780000 1.615000 ;
      RECT 1.070000 1.785000 1.240000 1.955000 ;
      RECT 2.495000 1.785000 2.665000 1.955000 ;
      RECT 2.955000 1.445000 3.125000 1.615000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.185000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.725000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.435000 1.755000 2.725000 1.800000 ;
      RECT 2.435000 1.940000 2.725000 1.985000 ;
      RECT 2.895000 1.415000 3.185000 1.460000 ;
      RECT 2.895000 1.600000 3.185000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxbn_1

* File: sky130_fd_sc_hd__dlygate4sd2_1.pex.spice
* Created: Tue Sep  1 19:06:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A 3 7 9 10 15 17
c32 17 0 7.45863e-20 $X=0.58 $Y=1.16
r33 14 17 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=0.32 $Y=1.16
+ $X2=0.58 $Y2=1.16
r34 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.16 $X2=0.32 $Y2=1.16
r35 9 10 7.53086 $w=5.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.355 $Y=1.19
+ $X2=0.355 $Y2=1.53
r36 9 15 0.664488 $w=5.38e-07 $l=3e-08 $layer=LI1_cond $X=0.355 $Y=1.19
+ $X2=0.355 $Y2=1.16
r37 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.325
+ $X2=0.58 $Y2=1.16
r38 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.58 $Y=1.325 $X2=0.58
+ $Y2=2.275
r39 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.58 $Y2=1.16
r40 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.58 $Y=0.995 $X2=0.58
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_49_47# 1 2 9 13 17 21 23 24 25 26 27
+ 28 32
c66 32 0 1.52587e-19 $X=1 $Y=1.16
c67 27 0 1.19506e-19 $X=0.912 $Y=1.325
c68 25 0 7.45863e-20 $X=0.795 $Y=1.895
r69 32 35 43.3395 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.16 $X2=1
+ $Y2=1.325
r70 32 34 43.3395 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.16 $X2=1
+ $Y2=0.995
r71 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r72 29 31 16.6364 $w=2.64e-07 $l=3.6e-07 $layer=LI1_cond $X=0.94 $Y=0.8 $X2=0.94
+ $Y2=1.16
r73 27 31 7.80106 $w=2.64e-07 $l=1.78452e-07 $layer=LI1_cond $X=0.912 $Y=1.325
+ $X2=0.94 $Y2=1.16
r74 27 28 22.5585 $w=2.33e-07 $l=4.6e-07 $layer=LI1_cond $X=0.912 $Y=1.325
+ $X2=0.912 $Y2=1.785
r75 25 28 6.82613 $w=2.2e-07 $l=1.62969e-07 $layer=LI1_cond $X=0.795 $Y=1.895
+ $X2=0.912 $Y2=1.785
r76 25 26 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=0.795 $Y=1.895
+ $X2=0.485 $Y2=1.895
r77 23 29 3.3128 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.795 $Y=0.8 $X2=0.94
+ $Y2=0.8
r78 23 24 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.795 $Y=0.8
+ $X2=0.485 $Y2=0.8
r79 19 26 7.59172 $w=2.2e-07 $l=2.48998e-07 $layer=LI1_cond $X=0.285 $Y=2.005
+ $X2=0.485 $Y2=1.895
r80 19 21 5.90627 $w=3.98e-07 $l=2.05e-07 $layer=LI1_cond $X=0.285 $Y=2.005
+ $X2=0.285 $Y2=2.21
r81 15 24 8.37092 $w=1.7e-07 $l=2.38747e-07 $layer=LI1_cond $X=0.285 $Y=0.715
+ $X2=0.485 $Y2=0.8
r82 15 17 5.90627 $w=3.98e-07 $l=2.05e-07 $layer=LI1_cond $X=0.285 $Y=0.715
+ $X2=0.285 $Y2=0.51
r83 13 35 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=1.015 $Y=2.275
+ $X2=1.015 $Y2=1.325
r84 9 34 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=1.015 $Y=0.445
+ $X2=1.015 $Y2=0.995
r85 2 21 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=2.065 $X2=0.37 $Y2=2.21
r86 1 17 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_221_47# 1 2 9 13 16 18 21 27 32 34
+ 37
c61 37 0 7.47284e-20 $X=1.985 $Y=1.16
r62 30 32 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.24 $Y=2.3 $X2=1.34
+ $Y2=2.3
r63 25 27 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.24 $Y=0.42 $X2=1.34
+ $Y2=0.42
r64 22 37 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.76 $Y=1.16
+ $X2=1.985 $Y2=1.16
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.76
+ $Y=1.16 $X2=1.76 $Y2=1.16
r66 19 34 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.425 $Y=1.335
+ $X2=1.34 $Y2=1.335
r67 19 21 7.15511 $w=5.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.425 $Y=1.335
+ $X2=1.76 $Y2=1.335
r68 18 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=2.135
+ $X2=1.34 $Y2=2.3
r69 17 34 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=1.34 $Y=1.615
+ $X2=1.34 $Y2=1.335
r70 17 18 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.34 $Y=1.615
+ $X2=1.34 $Y2=2.135
r71 16 34 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=1.34 $Y=1.055
+ $X2=1.34 $Y2=1.335
r72 15 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=0.585
+ $X2=1.34 $Y2=0.42
r73 15 16 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.34 $Y=0.585
+ $X2=1.34 $Y2=1.055
r74 11 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.325
+ $X2=1.985 $Y2=1.16
r75 11 13 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=1.985 $Y=1.325
+ $X2=1.985 $Y2=2.275
r76 7 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.985 $Y2=1.16
r77 7 9 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.985 $Y2=0.445
r78 2 30 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=2.065 $X2=1.24 $Y2=2.3
r79 1 25 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.235 $X2=1.24 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_327_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c67 26 0 1.18733e-19 $X=2.3 $Y=1.325
c68 24 0 7.47284e-20 $X=2.2 $Y=1.895
r69 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.16
+ $X2=2.42 $Y2=1.325
r70 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.16
+ $X2=2.42 $Y2=0.995
r71 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.16 $X2=2.42 $Y2=1.16
r72 28 30 17.1562 $w=2.56e-07 $l=3.6e-07 $layer=LI1_cond $X=2.352 $Y=0.8
+ $X2=2.352 $Y2=1.16
r73 26 30 8.48013 $w=2.56e-07 $l=1.89222e-07 $layer=LI1_cond $X=2.3 $Y=1.325
+ $X2=2.352 $Y2=1.16
r74 26 27 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.3 $Y=1.325 $X2=2.3
+ $Y2=1.785
r75 24 27 6.83662 $w=2.2e-07 $l=1.51987e-07 $layer=LI1_cond $X=2.2 $Y=1.895
+ $X2=2.3 $Y2=1.785
r76 24 25 17.0247 $w=2.18e-07 $l=3.25e-07 $layer=LI1_cond $X=2.2 $Y=1.895
+ $X2=1.875 $Y2=1.895
r77 22 28 3.13337 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.2 $Y=0.8 $X2=2.352
+ $Y2=0.8
r78 22 23 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.2 $Y=0.8
+ $X2=1.875 $Y2=0.8
r79 18 25 6.87824 $w=2.2e-07 $l=1.76635e-07 $layer=LI1_cond $X=1.745 $Y=2.005
+ $X2=1.875 $Y2=1.895
r80 18 20 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=1.745 $Y=2.005
+ $X2=1.745 $Y2=2.21
r81 14 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.745 $Y=0.715
+ $X2=1.875 $Y2=0.8
r82 14 16 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=1.745 $Y=0.715
+ $X2=1.745 $Y2=0.51
r83 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.475 $Y=1.985
+ $X2=2.475 $Y2=1.325
r84 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.475 $Y=0.56
+ $X2=2.475 $Y2=0.995
r85 2 20 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.635
+ $Y=2.065 $X2=1.76 $Y2=2.21
r86 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.235 $X2=1.76 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%VPWR 1 2 11 15 18 19 20 30 31 34
r41 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 25 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 24 27 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r48 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 22 34 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.79 $Y2=2.72
r50 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 18 27 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 18 19 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=2.237 $Y2=2.72
r54 17 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.4 $Y=2.72 $X2=2.99
+ $Y2=2.72
r55 17 19 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=2.4 $Y=2.72 $X2=2.237
+ $Y2=2.72
r56 13 19 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.237 $Y=2.635
+ $X2=2.237 $Y2=2.72
r57 13 15 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=2.237 $Y=2.635
+ $X2=2.237 $Y2=2.34
r58 9 34 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=2.635
+ $X2=0.79 $Y2=2.72
r59 9 11 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.79 $Y=2.635
+ $X2=0.79 $Y2=2.34
r60 2 15 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.075
+ $Y=2.065 $X2=2.235 $Y2=2.34
r61 1 11 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=2.065 $X2=0.79 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%X 1 2 7 8 9 10 11 12 24 43
r16 43 44 1.18924 $w=5.63e-07 $l=3.5e-08 $layer=LI1_cond $X=2.852 $Y=1.53
+ $X2=2.852 $Y2=1.495
r17 24 41 0.650043 $w=4.58e-07 $l=2.5e-08 $layer=LI1_cond $X=2.905 $Y=0.85
+ $X2=2.905 $Y2=0.825
r18 11 12 7.19764 $w=5.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.852 $Y=1.87
+ $X2=2.852 $Y2=2.21
r19 11 29 1.96877 $w=5.63e-07 $l=9.3e-08 $layer=LI1_cond $X=2.852 $Y=1.87
+ $X2=2.852 $Y2=1.777
r20 10 29 4.69964 $w=5.63e-07 $l=2.22e-07 $layer=LI1_cond $X=2.852 $Y=1.555
+ $X2=2.852 $Y2=1.777
r21 10 43 0.529238 $w=5.63e-07 $l=2.5e-08 $layer=LI1_cond $X=2.852 $Y=1.555
+ $X2=2.852 $Y2=1.53
r22 10 44 0.650043 $w=4.58e-07 $l=2.5e-08 $layer=LI1_cond $X=2.905 $Y=1.47
+ $X2=2.905 $Y2=1.495
r23 9 10 7.28048 $w=4.58e-07 $l=2.8e-07 $layer=LI1_cond $X=2.905 $Y=1.19
+ $X2=2.905 $Y2=1.47
r24 8 41 1.0834 $w=5.63e-07 $l=3e-08 $layer=LI1_cond $X=2.852 $Y=0.795 $X2=2.852
+ $Y2=0.825
r25 8 9 8.06053 $w=4.58e-07 $l=3.1e-07 $layer=LI1_cond $X=2.905 $Y=0.88
+ $X2=2.905 $Y2=1.19
r26 8 24 0.780051 $w=4.58e-07 $l=3e-08 $layer=LI1_cond $X=2.905 $Y=0.88
+ $X2=2.905 $Y2=0.85
r27 7 8 6.03332 $w=5.63e-07 $l=2.85e-07 $layer=LI1_cond $X=2.852 $Y=0.51
+ $X2=2.852 $Y2=0.795
r28 2 11 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=1.485 $X2=2.685 $Y2=1.87
r29 1 7 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.235 $X2=2.685 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%VGND 1 2 11 15 18 19 20 30 31 34
c45 11 0 1.52587e-19 $X=0.79 $Y=0.38
r46 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r48 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r49 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r50 25 28 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r51 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r52 24 27 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r53 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 22 34 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.79
+ $Y2=0
r55 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.15
+ $Y2=0
r56 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r57 18 27 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r58 18 19 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.237
+ $Y2=0
r59 17 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.99
+ $Y2=0
r60 17 19 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.237
+ $Y2=0
r61 13 19 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.237 $Y=0.085
+ $X2=2.237 $Y2=0
r62 13 15 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=2.237 $Y=0.085
+ $X2=2.237 $Y2=0.38
r63 9 34 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r64 9 11 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.38
r65 2 15 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.235 $X2=2.235 $Y2=0.38
r66 1 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.655
+ $Y=0.235 $X2=0.79 $Y2=0.38
.ends


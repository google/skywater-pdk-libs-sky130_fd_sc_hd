* File: sky130_fd_sc_hd__o21a_4.pxi.spice
* Created: Tue Sep  1 19:21:18 2020
* 
x_PM_SKY130_FD_SC_HD__O21A_4%A_80_21# N_A_80_21#_M1012_d N_A_80_21#_M1008_s
+ N_A_80_21#_M1015_d N_A_80_21#_c_83_n N_A_80_21#_M1005_g N_A_80_21#_M1000_g
+ N_A_80_21#_c_84_n N_A_80_21#_M1007_g N_A_80_21#_M1002_g N_A_80_21#_c_85_n
+ N_A_80_21#_M1009_g N_A_80_21#_M1006_g N_A_80_21#_c_86_n N_A_80_21#_M1018_g
+ N_A_80_21#_M1013_g N_A_80_21#_c_94_n N_A_80_21#_c_95_n N_A_80_21#_c_87_n
+ N_A_80_21#_c_99_p N_A_80_21#_c_129_p N_A_80_21#_c_149_p N_A_80_21#_c_102_p
+ N_A_80_21#_c_88_n N_A_80_21#_c_109_p N_A_80_21#_c_117_p N_A_80_21#_c_89_n
+ PM_SKY130_FD_SC_HD__O21A_4%A_80_21#
x_PM_SKY130_FD_SC_HD__O21A_4%B1 N_B1_M1008_g N_B1_c_212_n N_B1_M1012_g
+ N_B1_M1014_g N_B1_c_213_n N_B1_M1019_g B1 N_B1_c_217_n N_B1_c_214_n
+ PM_SKY130_FD_SC_HD__O21A_4%B1
x_PM_SKY130_FD_SC_HD__O21A_4%A1 N_A1_M1003_g N_A1_M1001_g N_A1_M1017_g
+ N_A1_M1011_g N_A1_c_265_n N_A1_c_266_n N_A1_c_282_n N_A1_c_285_n A1
+ N_A1_c_267_n N_A1_c_268_n N_A1_c_269_n N_A1_c_270_n N_A1_c_277_n
+ PM_SKY130_FD_SC_HD__O21A_4%A1
x_PM_SKY130_FD_SC_HD__O21A_4%A2 N_A2_c_340_n N_A2_M1010_g N_A2_M1015_g
+ N_A2_c_341_n N_A2_M1016_g N_A2_M1004_g A2 N_A2_c_342_n N_A2_c_343_n
+ PM_SKY130_FD_SC_HD__O21A_4%A2
x_PM_SKY130_FD_SC_HD__O21A_4%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1013_d
+ N_VPWR_M1014_d N_VPWR_M1011_s N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_390_n
+ N_VPWR_c_391_n N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n
+ N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n VPWR N_VPWR_c_399_n
+ N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_387_n PM_SKY130_FD_SC_HD__O21A_4%VPWR
x_PM_SKY130_FD_SC_HD__O21A_4%X N_X_M1005_d N_X_M1009_d N_X_M1000_s N_X_M1006_s
+ N_X_c_479_n N_X_c_480_n N_X_c_485_n N_X_c_486_n N_X_c_506_n N_X_c_491_n
+ N_X_c_510_n N_X_c_495_n N_X_c_497_n X N_X_c_477_n X
+ PM_SKY130_FD_SC_HD__O21A_4%X
x_PM_SKY130_FD_SC_HD__O21A_4%VGND N_VGND_M1005_s N_VGND_M1007_s N_VGND_M1018_s
+ N_VGND_M1003_d N_VGND_M1016_s N_VGND_c_533_n N_VGND_c_534_n N_VGND_c_535_n
+ N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n VGND N_VGND_c_539_n
+ N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n
+ N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n
+ PM_SKY130_FD_SC_HD__O21A_4%VGND
x_PM_SKY130_FD_SC_HD__O21A_4%A_475_47# N_A_475_47#_M1012_s N_A_475_47#_M1019_s
+ N_A_475_47#_M1010_d N_A_475_47#_M1017_s N_A_475_47#_c_625_n
+ N_A_475_47#_c_626_n N_A_475_47#_c_639_n PM_SKY130_FD_SC_HD__O21A_4%A_475_47#
cc_1 VNB N_A_80_21#_c_83_n 0.0184169f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_84_n 0.0160024f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_A_80_21#_c_85_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.995
cc_4 VNB N_A_80_21#_c_86_n 0.0186877f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.995
cc_5 VNB N_A_80_21#_c_87_n 0.00362584f $X=-0.19 $Y=-0.24 $X2=2.93 $Y2=0.76
cc_6 VNB N_A_80_21#_c_88_n 0.0110211f $X=-0.19 $Y=-0.24 $X2=2.215 $Y2=0.762
cc_7 VNB N_A_80_21#_c_89_n 0.0882322f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=1.16
cc_8 VNB N_B1_c_212_n 0.0195826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_213_n 0.0170566f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_10 VNB N_B1_c_214_n 0.0438359f $X=-0.19 $Y=-0.24 $X2=1.655 $Y2=1.325
cc_11 VNB N_A1_c_265_n 0.00164747f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_12 VNB N_A1_c_266_n 0.0298551f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_13 VNB N_A1_c_267_n 0.0179078f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.56
cc_14 VNB N_A1_c_268_n 0.0300205f $X=-0.19 $Y=-0.24 $X2=1.655 $Y2=1.985
cc_15 VNB N_A1_c_269_n 0.0147456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_270_n 0.022077f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.995
cc_17 VNB N_A2_c_340_n 0.0168121f $X=-0.19 $Y=-0.24 $X2=2.79 $Y2=0.235
cc_18 VNB N_A2_c_341_n 0.016201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_342_n 0.0374603f $X=-0.19 $Y=-0.24 $X2=1.225 $Y2=1.985
cc_20 VNB N_A2_c_343_n 0.00118947f $X=-0.19 $Y=-0.24 $X2=1.225 $Y2=1.985
cc_21 VNB N_VPWR_c_387_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_22 VNB N_X_c_477_n 0.00760135f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.165
cc_23 VNB X 0.0238419f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_24 VNB N_VGND_c_533_n 0.0103103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_534_n 0.0119016f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_26 VNB N_VGND_c_535_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=1.225 $Y2=1.985
cc_27 VNB N_VGND_c_536_n 0.00526464f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.56
cc_28 VNB N_VGND_c_537_n 0.00275439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_538_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=1.325
cc_30 VNB N_VGND_c_539_n 0.0122979f $X=-0.19 $Y=-0.24 $X2=2.115 $Y2=1.165
cc_31 VNB N_VGND_c_540_n 0.0127251f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=1.165
cc_32 VNB N_VGND_c_541_n 0.0378687f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=0.762
cc_33 VNB N_VGND_c_542_n 0.0122674f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=1.957
cc_34 VNB N_VGND_c_543_n 0.0164562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_544_n 0.279007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_545_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=2.75 $Y2=1.96
cc_37 VNB N_VGND_c_546_n 0.00510127f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.16
cc_38 VNB N_VGND_c_547_n 0.00528879f $X=-0.19 $Y=-0.24 $X2=0.795 $Y2=1.16
cc_39 VNB N_VGND_c_548_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.16
cc_40 VNB N_A_475_47#_c_625_n 0.00286189f $X=-0.19 $Y=-0.24 $X2=0.795 $Y2=1.325
cc_41 VNB N_A_475_47#_c_626_n 0.00813518f $X=-0.19 $Y=-0.24 $X2=1.225 $Y2=1.985
cc_42 VPB N_A_80_21#_M1000_g 0.0219111f $X=-0.19 $Y=1.305 $X2=0.795 $Y2=1.985
cc_43 VPB N_A_80_21#_M1002_g 0.0184823f $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.985
cc_44 VPB N_A_80_21#_M1006_g 0.0184531f $X=-0.19 $Y=1.305 $X2=1.655 $Y2=1.985
cc_45 VPB N_A_80_21#_M1013_g 0.0180704f $X=-0.19 $Y=1.305 $X2=2.085 $Y2=1.985
cc_46 VPB N_A_80_21#_c_94_n 0.012031f $X=-0.19 $Y=1.305 $X2=2.115 $Y2=1.165
cc_47 VPB N_A_80_21#_c_95_n 8.87389e-19 $X=-0.19 $Y=1.305 $X2=2.22 $Y2=1.83
cc_48 VPB N_A_80_21#_c_89_n 0.0220601f $X=-0.19 $Y=1.305 $X2=2.085 $Y2=1.16
cc_49 VPB N_B1_M1008_g 0.0183085f $X=-0.19 $Y=1.305 $X2=4.24 $Y2=1.485
cc_50 VPB N_B1_M1014_g 0.0198754f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_51 VPB N_B1_c_217_n 0.00148153f $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.985
cc_52 VPB N_B1_c_214_n 0.0107386f $X=-0.19 $Y=1.305 $X2=1.655 $Y2=1.325
cc_53 VPB N_A1_M1001_g 0.0208794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A1_M1011_g 0.0225929f $X=-0.19 $Y=1.305 $X2=0.795 $Y2=1.325
cc_55 VPB N_A1_c_265_n 0.00140938f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.995
cc_56 VPB N_A1_c_266_n 0.00809547f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.56
cc_57 VPB N_A1_c_268_n 0.00675079f $X=-0.19 $Y=1.305 $X2=1.655 $Y2=1.985
cc_58 VPB N_A1_c_269_n 0.00714312f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A1_c_277_n 0.00881036f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=0.56
cc_60 VPB N_A2_M1015_g 0.0190486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A2_M1004_g 0.0190548f $X=-0.19 $Y=1.305 $X2=0.795 $Y2=1.325
cc_62 VPB N_A2_c_342_n 0.00675039f $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.985
cc_63 VPB N_A2_c_343_n 0.00110374f $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.985
cc_64 VPB N_VPWR_c_388_n 0.026733f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.56
cc_65 VPB N_VPWR_c_389_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=1.225 $Y2=1.985
cc_66 VPB N_VPWR_c_390_n 3.08929e-19 $X=-0.19 $Y=1.305 $X2=1.335 $Y2=0.56
cc_67 VPB N_VPWR_c_391_n 0.0105978f $X=-0.19 $Y=1.305 $X2=1.655 $Y2=1.985
cc_68 VPB N_VPWR_c_392_n 0.0261341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_393_n 0.0153494f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=0.56
cc_70 VPB N_VPWR_c_394_n 0.00510842f $X=-0.19 $Y=1.305 $X2=2.085 $Y2=1.325
cc_71 VPB N_VPWR_c_395_n 0.0129398f $X=-0.19 $Y=1.305 $X2=2.085 $Y2=1.985
cc_72 VPB N_VPWR_c_396_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_397_n 0.0129938f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.165
cc_74 VPB N_VPWR_c_398_n 0.00462744f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_75 VPB N_VPWR_c_399_n 0.0366436f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_400_n 0.0113761f $X=-0.19 $Y=1.305 $X2=4.38 $Y2=1.99
cc_77 VPB N_VPWR_c_401_n 0.0122827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_387_n 0.0562047f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_79 VPB N_X_c_479_n 0.00770909f $X=-0.19 $Y=1.305 $X2=0.795 $Y2=1.325
cc_80 VPB N_X_c_480_n 0.0176557f $X=-0.19 $Y=1.305 $X2=0.795 $Y2=1.985
cc_81 VPB X 0.0123549f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_82 N_A_80_21#_M1013_g N_B1_M1008_g 0.0252208f $X=2.085 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_95_n N_B1_M1008_g 0.00515707f $X=2.22 $Y=1.83 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_99_p N_B1_M1008_g 0.012959f $X=2.655 $Y=1.957 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_87_n N_B1_c_212_n 0.011662f $X=2.93 $Y=0.76 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_88_n N_B1_c_212_n 0.00441186f $X=2.215 $Y=0.762 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_102_p N_B1_M1014_g 0.0133664f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_87_n N_B1_c_213_n 0.00381045f $X=2.93 $Y=0.76 $X2=0 $Y2=0
cc_89 N_A_80_21#_M1008_s N_B1_c_217_n 0.00202214f $X=2.61 $Y=1.485 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_87_n N_B1_c_217_n 0.0352021f $X=2.93 $Y=0.76 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_99_p N_B1_c_217_n 0.00786612f $X=2.655 $Y=1.957 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_102_p N_B1_c_217_n 0.01151f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_88_n N_B1_c_217_n 0.0430685f $X=2.215 $Y=0.762 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_109_p N_B1_c_217_n 0.0122818f $X=2.75 $Y=1.96 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_89_n N_B1_c_217_n 5.10896e-19 $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_87_n N_B1_c_214_n 0.00819502f $X=2.93 $Y=0.76 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_102_p N_B1_c_214_n 0.00223133f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_88_n N_B1_c_214_n 0.00515707f $X=2.215 $Y=0.762 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_109_p N_B1_c_214_n 4.19987e-19 $X=2.75 $Y=1.96 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_89_n N_B1_c_214_n 0.0252208f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_102_p N_A1_M1001_g 0.0155419f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_117_p N_A1_M1001_g 0.00132842f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_117_p N_A1_M1011_g 0.0017887f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_102_p N_A1_c_266_n 0.00170362f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_105 N_A_80_21#_M1015_d N_A1_c_282_n 0.00332286f $X=4.24 $Y=1.485 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_102_p N_A1_c_282_n 0.0230368f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_117_p N_A1_c_282_n 0.0172374f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_102_p N_A1_c_285_n 0.0199333f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_102_p N_A2_M1015_g 0.00980579f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_117_p N_A2_M1015_g 0.00712025f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_117_p N_A2_M1004_g 0.0106248f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_95_n N_VPWR_M1013_d 0.00355959f $X=2.22 $Y=1.83 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_99_p N_VPWR_M1013_d 0.00438728f $X=2.655 $Y=1.957 $X2=0
+ $Y2=0
cc_114 N_A_80_21#_c_129_p N_VPWR_M1013_d 0.00103261f $X=2.315 $Y=1.957 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_c_102_p N_VPWR_M1014_d 0.0206981f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_116 N_A_80_21#_M1000_g N_VPWR_c_388_n 0.0114143f $X=0.795 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_80_21#_M1002_g N_VPWR_c_388_n 6.1315e-19 $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_80_21#_M1000_g N_VPWR_c_389_n 6.1315e-19 $X=0.795 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_80_21#_M1002_g N_VPWR_c_389_n 0.0103509f $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_80_21#_M1006_g N_VPWR_c_389_n 0.0103509f $X=1.655 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_80_21#_M1013_g N_VPWR_c_389_n 6.1315e-19 $X=2.085 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_80_21#_M1006_g N_VPWR_c_390_n 5.08691e-19 $X=1.655 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_80_21#_M1013_g N_VPWR_c_390_n 0.00655764f $X=2.085 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_80_21#_c_99_p N_VPWR_c_390_n 0.0085803f $X=2.655 $Y=1.957 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_129_p N_VPWR_c_390_n 0.0100754f $X=2.315 $Y=1.957 $X2=0
+ $Y2=0
cc_126 N_A_80_21#_c_117_p N_VPWR_c_392_n 0.0154707f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_127 N_A_80_21#_M1000_g N_VPWR_c_395_n 0.00486043f $X=0.795 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_M1002_g N_VPWR_c_395_n 0.00486043f $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_A_80_21#_M1006_g N_VPWR_c_397_n 0.00486043f $X=1.655 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_80_21#_M1013_g N_VPWR_c_397_n 0.00476417f $X=2.085 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_c_102_p N_VPWR_c_399_n 0.00862733f $X=4.215 $Y=1.99 $X2=0
+ $Y2=0
cc_132 N_A_80_21#_c_117_p N_VPWR_c_399_n 0.0166316f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_99_p N_VPWR_c_400_n 0.00252184f $X=2.655 $Y=1.957 $X2=0
+ $Y2=0
cc_134 N_A_80_21#_c_149_p N_VPWR_c_400_n 0.0123954f $X=2.75 $Y=2.3 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_102_p N_VPWR_c_400_n 0.00263122f $X=4.215 $Y=1.99 $X2=0
+ $Y2=0
cc_136 N_A_80_21#_c_102_p N_VPWR_c_401_n 0.0424296f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_117_p N_VPWR_c_401_n 0.00529302f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_138 N_A_80_21#_M1008_s N_VPWR_c_387_n 0.00252469f $X=2.61 $Y=1.485 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_M1015_d N_VPWR_c_387_n 0.00224096f $X=4.24 $Y=1.485 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_M1000_g N_VPWR_c_387_n 0.00822531f $X=0.795 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_80_21#_M1002_g N_VPWR_c_387_n 0.00822531f $X=1.225 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_80_21#_M1006_g N_VPWR_c_387_n 0.00822531f $X=1.655 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_M1013_g N_VPWR_c_387_n 0.00786326f $X=2.085 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_c_99_p N_VPWR_c_387_n 0.00500811f $X=2.655 $Y=1.957 $X2=0
+ $Y2=0
cc_145 N_A_80_21#_c_129_p N_VPWR_c_387_n 0.0011786f $X=2.315 $Y=1.957 $X2=0
+ $Y2=0
cc_146 N_A_80_21#_c_149_p N_VPWR_c_387_n 0.00722721f $X=2.75 $Y=2.3 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_102_p N_VPWR_c_387_n 0.0215892f $X=4.215 $Y=1.99 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_117_p N_VPWR_c_387_n 0.0120843f $X=4.38 $Y=2.02 $X2=0 $Y2=0
cc_149 N_A_80_21#_M1000_g N_X_c_479_n 0.0157301f $X=0.795 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_94_n N_X_c_479_n 0.0257396f $X=2.115 $Y=1.165 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_89_n N_X_c_479_n 0.00498754f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_80_21#_c_89_n N_X_c_485_n 0.0022939f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_84_n N_X_c_486_n 0.0101429f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_80_21#_c_85_n N_X_c_486_n 0.0101376f $X=1.335 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_80_21#_c_86_n N_X_c_486_n 0.005173f $X=1.765 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_80_21#_c_88_n N_X_c_486_n 0.00632392f $X=2.215 $Y=0.762 $X2=0 $Y2=0
cc_157 N_A_80_21#_c_89_n N_X_c_486_n 0.00520952f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_80_21#_M1002_g N_X_c_491_n 0.0137508f $X=1.225 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_80_21#_M1006_g N_X_c_491_n 0.0134702f $X=1.655 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_80_21#_c_94_n N_X_c_491_n 0.0523251f $X=2.115 $Y=1.165 $X2=0 $Y2=0
cc_161 N_A_80_21#_c_89_n N_X_c_491_n 0.00141679f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_80_21#_c_83_n N_X_c_495_n 0.0135536f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_80_21#_c_94_n N_X_c_495_n 0.0711211f $X=2.115 $Y=1.165 $X2=0 $Y2=0
cc_164 N_A_80_21#_c_94_n N_X_c_497_n 0.0139676f $X=2.115 $Y=1.165 $X2=0 $Y2=0
cc_165 N_A_80_21#_c_89_n N_X_c_497_n 7.50945e-19 $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_80_21#_c_83_n X 0.0171386f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_80_21#_M1000_g X 0.0054738f $X=0.795 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_80_21#_c_94_n X 0.0276497f $X=2.115 $Y=1.165 $X2=0 $Y2=0
cc_169 N_A_80_21#_c_102_p A_934_297# 0.00464299f $X=4.215 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_80_21#_c_83_n N_VGND_c_534_n 0.00907946f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_80_21#_c_84_n N_VGND_c_534_n 0.00114137f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_80_21#_c_83_n N_VGND_c_535_n 0.00104385f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A_80_21#_c_84_n N_VGND_c_535_n 0.00765006f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_174 N_A_80_21#_c_85_n N_VGND_c_535_n 0.00765006f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_A_80_21#_c_86_n N_VGND_c_535_n 0.00104385f $X=1.765 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_80_21#_c_85_n N_VGND_c_536_n 0.00114137f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_80_21#_c_86_n N_VGND_c_536_n 0.00936889f $X=1.765 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_80_21#_c_94_n N_VGND_c_536_n 0.00889986f $X=2.115 $Y=1.165 $X2=0
+ $Y2=0
cc_179 N_A_80_21#_c_88_n N_VGND_c_536_n 0.00224089f $X=2.215 $Y=0.762 $X2=0
+ $Y2=0
cc_180 N_A_80_21#_c_89_n N_VGND_c_536_n 0.0053922f $X=2.085 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_80_21#_c_83_n N_VGND_c_539_n 0.00353537f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_80_21#_c_84_n N_VGND_c_539_n 0.00351072f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_80_21#_c_85_n N_VGND_c_540_n 0.00351072f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_80_21#_c_86_n N_VGND_c_540_n 0.00458831f $X=1.765 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_80_21#_c_87_n N_VGND_c_541_n 3.56478e-19 $X=2.93 $Y=0.76 $X2=0 $Y2=0
cc_186 N_A_80_21#_c_88_n N_VGND_c_541_n 0.0032847f $X=2.215 $Y=0.762 $X2=0 $Y2=0
cc_187 N_A_80_21#_M1012_d N_VGND_c_544_n 0.00224864f $X=2.79 $Y=0.235 $X2=0
+ $Y2=0
cc_188 N_A_80_21#_c_83_n N_VGND_c_544_n 0.00415708f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_80_21#_c_84_n N_VGND_c_544_n 0.00411677f $X=0.905 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_80_21#_c_85_n N_VGND_c_544_n 0.00411677f $X=1.335 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_80_21#_c_86_n N_VGND_c_544_n 0.00747175f $X=1.765 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_80_21#_c_87_n N_VGND_c_544_n 0.00198975f $X=2.93 $Y=0.76 $X2=0 $Y2=0
cc_193 N_A_80_21#_c_88_n N_VGND_c_544_n 0.00520079f $X=2.215 $Y=0.762 $X2=0
+ $Y2=0
cc_194 N_A_80_21#_c_87_n N_A_475_47#_M1012_s 0.00766144f $X=2.93 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_195 N_A_80_21#_M1012_d N_A_475_47#_c_625_n 0.00324248f $X=2.79 $Y=0.235 $X2=0
+ $Y2=0
cc_196 N_A_80_21#_c_87_n N_A_475_47#_c_625_n 0.0416037f $X=2.93 $Y=0.76 $X2=0
+ $Y2=0
cc_197 N_B1_M1014_g N_A1_M1001_g 0.0150016f $X=2.965 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B1_c_217_n N_A1_M1001_g 0.00106089f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_M1014_g N_A1_c_265_n 6.04418e-19 $X=2.965 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B1_c_217_n N_A1_c_265_n 0.0211699f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B1_c_214_n N_A1_c_265_n 0.00153946f $X=3.145 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_c_217_n N_A1_c_266_n 8.36424e-19 $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B1_c_214_n N_A1_c_266_n 0.0218769f $X=3.145 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B1_M1014_g N_A1_c_285_n 0.00250544f $X=2.965 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B1_c_217_n N_A1_c_285_n 0.00666698f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B1_c_213_n N_A1_c_267_n 0.0189724f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B1_c_217_n N_VPWR_M1014_d 0.00246039f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B1_M1008_g N_VPWR_c_390_n 0.00650804f $X=2.535 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1014_g N_VPWR_c_390_n 5.05034e-19 $X=2.965 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_M1008_g N_VPWR_c_400_n 0.00353537f $X=2.535 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1014_g N_VPWR_c_400_n 0.00351072f $X=2.965 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1008_g N_VPWR_c_401_n 5.14256e-19 $X=2.535 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1014_g N_VPWR_c_401_n 0.00728383f $X=2.965 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1008_g N_VPWR_c_387_n 0.00411309f $X=2.535 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1014_g N_VPWR_c_387_n 0.0040578f $X=2.965 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B1_c_212_n N_VGND_c_536_n 0.00234448f $X=2.715 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_212_n N_VGND_c_541_n 0.00357877f $X=2.715 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_213_n N_VGND_c_541_n 0.00357877f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_212_n N_VGND_c_544_n 0.00657863f $X=2.715 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B1_c_213_n N_VGND_c_544_n 0.00553294f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B1_c_212_n N_A_475_47#_c_625_n 0.00920885f $X=2.715 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_B1_c_213_n N_A_475_47#_c_625_n 0.0136954f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B1_c_217_n N_A_475_47#_c_625_n 0.0016068f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A1_c_267_n N_A2_c_340_n 0.0253749f $X=3.622 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_225 N_A1_M1001_g N_A2_M1015_g 0.0371745f $X=3.735 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A1_c_282_n N_A2_M1015_g 0.0135953f $X=5.03 $Y=1.6 $X2=0 $Y2=0
cc_227 N_A1_c_270_n N_A2_c_341_n 0.0271828f $X=5.115 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A1_M1011_g N_A2_M1004_g 0.0574807f $X=5.025 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A1_c_282_n N_A2_M1004_g 0.015925f $X=5.03 $Y=1.6 $X2=0 $Y2=0
cc_230 N_A1_c_269_n N_A2_M1004_g 8.93695e-19 $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A1_c_265_n N_A2_c_342_n 0.00243785f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A1_c_266_n N_A2_c_342_n 0.0371745f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A1_c_282_n N_A2_c_342_n 0.00198407f $X=5.03 $Y=1.6 $X2=0 $Y2=0
cc_234 N_A1_c_268_n N_A2_c_342_n 0.0217057f $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A1_c_269_n N_A2_c_342_n 0.00118629f $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A1_c_265_n N_A2_c_343_n 0.0141901f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A1_c_266_n N_A2_c_343_n 0.00122759f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A1_c_282_n N_A2_c_343_n 0.0356877f $X=5.03 $Y=1.6 $X2=0 $Y2=0
cc_239 N_A1_c_268_n N_A2_c_343_n 0.00112056f $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A1_c_269_n N_A2_c_343_n 0.0149099f $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A1_c_285_n N_VPWR_M1014_d 0.00443886f $X=3.785 $Y=1.6 $X2=0 $Y2=0
cc_242 N_A1_c_277_n N_VPWR_M1011_s 0.00405261f $X=5.215 $Y=1.495 $X2=0 $Y2=0
cc_243 N_A1_M1011_g N_VPWR_c_392_n 0.0159381f $X=5.025 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A1_c_268_n N_VPWR_c_392_n 5.66234e-19 $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A1_c_277_n N_VPWR_c_392_n 0.0191225f $X=5.215 $Y=1.495 $X2=0 $Y2=0
cc_246 N_A1_M1001_g N_VPWR_c_399_n 0.00351072f $X=3.735 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A1_M1011_g N_VPWR_c_399_n 0.00486043f $X=5.025 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A1_M1001_g N_VPWR_c_401_n 0.0098987f $X=3.735 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A1_M1001_g N_VPWR_c_387_n 0.00412777f $X=3.735 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A1_M1011_g N_VPWR_c_387_n 0.0083285f $X=5.025 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A1_c_282_n A_934_297# 0.0082784f $X=5.03 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_252 N_A1_c_282_n A_762_297# 0.0126417f $X=5.03 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_253 N_A1_c_267_n N_VGND_c_537_n 0.004165f $X=3.622 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_270_n N_VGND_c_538_n 0.0140643f $X=5.115 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_267_n N_VGND_c_541_n 0.0041289f $X=3.622 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A1_c_270_n N_VGND_c_543_n 0.00351072f $X=5.115 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A1_c_267_n N_VGND_c_544_n 0.00602536f $X=3.622 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A1_c_270_n N_VGND_c_544_n 0.00510435f $X=5.115 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_c_265_n N_A_475_47#_c_626_n 0.0104494f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A1_c_266_n N_A_475_47#_c_626_n 9.83838e-19 $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A1_c_267_n N_A_475_47#_c_626_n 0.00953887f $X=3.622 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A1_c_268_n N_A_475_47#_c_626_n 0.00107332f $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A1_c_269_n N_A_475_47#_c_626_n 0.0232666f $X=5.115 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A1_c_270_n N_A_475_47#_c_626_n 0.012024f $X=5.115 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A1_c_265_n N_A_475_47#_c_639_n 0.00736299f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A1_c_266_n N_A_475_47#_c_639_n 0.00244243f $X=3.6 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A1_c_267_n N_A_475_47#_c_639_n 0.00670959f $X=3.622 $Y=0.995 $X2=0
+ $Y2=0
cc_268 N_A2_M1004_g N_VPWR_c_392_n 0.00271859f $X=4.595 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A2_M1015_g N_VPWR_c_399_n 0.00413555f $X=4.165 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A2_M1004_g N_VPWR_c_399_n 0.00549615f $X=4.595 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A2_M1015_g N_VPWR_c_401_n 0.00176586f $X=4.165 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A2_M1015_g N_VPWR_c_387_n 0.00576772f $X=4.165 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A2_M1004_g N_VPWR_c_387_n 0.00996598f $X=4.595 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A2_c_340_n N_VGND_c_537_n 0.00770381f $X=4.165 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_c_341_n N_VGND_c_537_n 0.00104439f $X=4.595 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A2_c_340_n N_VGND_c_538_n 0.00104385f $X=4.165 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A2_c_341_n N_VGND_c_538_n 0.0076143f $X=4.595 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A2_c_340_n N_VGND_c_542_n 0.00351072f $X=4.165 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A2_c_341_n N_VGND_c_542_n 0.00351072f $X=4.595 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A2_c_340_n N_VGND_c_544_n 0.00411677f $X=4.165 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A2_c_341_n N_VGND_c_544_n 0.00411677f $X=4.595 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A2_c_340_n N_A_475_47#_c_626_n 0.0115826f $X=4.165 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A2_c_341_n N_A_475_47#_c_626_n 0.00967692f $X=4.595 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A2_c_342_n N_A_475_47#_c_626_n 0.0018779f $X=4.605 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A2_c_343_n N_A_475_47#_c_626_n 0.0297167f $X=4.605 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A2_c_340_n N_A_475_47#_c_639_n 6.22612e-19 $X=4.165 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_387_n N_X_M1000_s 0.00535672f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_387_n N_X_M1006_s 0.00570388f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_M1000_d N_X_c_479_n 0.0049628f $X=0.455 $Y=1.485 $X2=0 $Y2=0
cc_290 N_VPWR_c_388_n N_X_c_479_n 0.0220026f $X=0.58 $Y=1.955 $X2=0 $Y2=0
cc_291 N_VPWR_c_395_n N_X_c_506_n 0.0124538f $X=1.275 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_387_n N_X_c_506_n 0.00724021f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_M1002_d N_X_c_491_n 0.00340337f $X=1.3 $Y=1.485 $X2=0 $Y2=0
cc_294 N_VPWR_c_389_n N_X_c_491_n 0.0170777f $X=1.44 $Y=1.955 $X2=0 $Y2=0
cc_295 N_VPWR_c_397_n N_X_c_510_n 0.012099f $X=2.135 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_c_387_n N_X_c_510_n 0.00684987f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_c_387_n A_934_297# 0.00318969f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_298 N_VPWR_c_387_n A_762_297# 0.0119688f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_299 N_X_c_495_n N_VGND_M1005_s 0.00106441f $X=0.595 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_300 N_X_c_477_n N_VGND_M1005_s 0.00276922f $X=0.205 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_301 X N_VGND_M1005_s 0.0012787f $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_302 N_X_c_486_n N_VGND_M1007_s 0.00331894f $X=1.55 $Y=0.71 $X2=0 $Y2=0
cc_303 N_X_c_495_n N_VGND_c_534_n 0.00339507f $X=0.595 $Y=0.71 $X2=0 $Y2=0
cc_304 N_X_c_477_n N_VGND_c_534_n 0.0190055f $X=0.205 $Y=0.805 $X2=0 $Y2=0
cc_305 N_X_c_486_n N_VGND_c_535_n 0.0160246f $X=1.55 $Y=0.71 $X2=0 $Y2=0
cc_306 N_X_c_485_n N_VGND_c_539_n 0.00590569f $X=0.69 $Y=0.72 $X2=0 $Y2=0
cc_307 N_X_c_495_n N_VGND_c_539_n 0.0024694f $X=0.595 $Y=0.71 $X2=0 $Y2=0
cc_308 N_X_c_486_n N_VGND_c_540_n 0.00680276f $X=1.55 $Y=0.71 $X2=0 $Y2=0
cc_309 N_X_M1005_d N_VGND_c_544_n 0.00320258f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_310 N_X_M1009_d N_VGND_c_544_n 0.00318969f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_311 N_X_c_485_n N_VGND_c_544_n 0.00979563f $X=0.69 $Y=0.72 $X2=0 $Y2=0
cc_312 N_X_c_486_n N_VGND_c_544_n 0.013196f $X=1.55 $Y=0.71 $X2=0 $Y2=0
cc_313 N_X_c_495_n N_VGND_c_544_n 0.00466137f $X=0.595 $Y=0.71 $X2=0 $Y2=0
cc_314 N_X_c_477_n N_VGND_c_544_n 0.00132683f $X=0.205 $Y=0.805 $X2=0 $Y2=0
cc_315 N_VGND_c_544_n N_A_475_47#_M1012_s 0.00213443f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_316 N_VGND_c_544_n N_A_475_47#_M1019_s 0.00287475f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_544_n N_A_475_47#_M1010_d 0.00318969f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_c_544_n N_A_475_47#_M1017_s 0.0030331f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_536_n N_A_475_47#_c_625_n 0.0170888f $X=1.98 $Y=0.38 $X2=0 $Y2=0
cc_320 N_VGND_c_541_n N_A_475_47#_c_625_n 0.0536006f $X=3.775 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_544_n N_A_475_47#_c_625_n 0.0338032f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_M1003_d N_A_475_47#_c_626_n 0.0112892f $X=3.73 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_VGND_M1016_s N_A_475_47#_c_626_n 0.00768399f $X=4.67 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_VGND_c_537_n N_A_475_47#_c_626_n 0.020311f $X=3.94 $Y=0.36 $X2=0 $Y2=0
cc_325 N_VGND_c_538_n N_A_475_47#_c_626_n 0.0159085f $X=4.81 $Y=0.36 $X2=0 $Y2=0
cc_326 N_VGND_c_541_n N_A_475_47#_c_626_n 0.00259773f $X=3.775 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_542_n N_A_475_47#_c_626_n 0.00846777f $X=4.645 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_543_n N_A_475_47#_c_626_n 0.00728503f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_544_n N_A_475_47#_c_626_n 0.0331269f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_330 N_VGND_c_541_n N_A_475_47#_c_639_n 0.0206214f $X=3.775 $Y=0 $X2=0 $Y2=0
cc_331 N_VGND_c_544_n N_A_475_47#_c_639_n 0.0123641f $X=5.29 $Y=0 $X2=0 $Y2=0

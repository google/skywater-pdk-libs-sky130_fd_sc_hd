* File: sky130_fd_sc_hd__a2111oi_1.pex.spice
* Created: Tue Sep  1 18:50:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2111OI_1%D1 3 6 8 9 10 11 17 18 19
r30 17 20 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.16
+ $X2=0.935 $Y2=1.325
r31 17 19 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.16
+ $X2=0.935 $Y2=0.995
r32 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.16 $X2=0.95 $Y2=1.16
r33 10 11 9.03704 $w=4.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.01 $Y=1.87
+ $X2=1.01 $Y2=2.21
r34 9 10 9.03704 $w=4.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.01 $Y=1.53 $X2=1.01
+ $Y2=1.87
r35 8 9 9.03704 $w=4.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.01 $Y=1.19 $X2=1.01
+ $Y2=1.53
r36 8 18 0.797386 $w=4.48e-07 $l=3e-08 $layer=LI1_cond $X=1.01 $Y=1.19 $X2=1.01
+ $Y2=1.16
r37 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.01 $Y=1.985
+ $X2=1.01 $Y2=1.325
r38 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.97 $Y=0.56 $X2=0.97
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%C1 3 6 7 8 9 10 16 18 19
r31 16 19 56.3675 $w=3.1e-07 $l=2.2e-07 $layer=POLY_cond $X=1.585 $Y=1.16
+ $X2=1.585 $Y2=1.38
r32 16 18 50.7832 $w=3.1e-07 $l=1.9e-07 $layer=POLY_cond $X=1.585 $Y=1.16
+ $X2=1.585 $Y2=0.97
r33 9 10 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.602 $Y=1.87
+ $X2=1.602 $Y2=2.21
r34 8 9 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.602 $Y=1.53
+ $X2=1.602 $Y2=1.87
r35 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.602 $Y=1.16
+ $X2=1.602 $Y2=1.53
r36 7 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.605
+ $Y=1.16 $X2=1.605 $Y2=1.16
r37 6 19 194.407 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=1.505 $Y=1.985
+ $X2=1.505 $Y2=1.38
r38 3 18 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.505 $Y=0.56
+ $X2=1.505 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%B1 3 6 8 9 10 11 17 19
c38 17 0 1.34745e-19 $X=2.105 $Y=1.16
c39 8 0 1.92208e-19 $X=2.07 $Y=1.19
c40 6 0 1.92762e-19 $X=2.025 $Y=1.985
r41 17 20 49.0286 $w=2.95e-07 $l=1.7e-07 $layer=POLY_cond $X=2.097 $Y=1.16
+ $X2=2.097 $Y2=1.33
r42 17 19 55.129 $w=2.95e-07 $l=2e-07 $layer=POLY_cond $X=2.097 $Y=1.16
+ $X2=2.097 $Y2=0.96
r43 10 11 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=2.077 $Y=1.87
+ $X2=2.077 $Y2=2.21
r44 9 10 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=2.077 $Y=1.53
+ $X2=2.077 $Y2=1.87
r45 9 32 5.44791 $w=2.73e-07 $l=1.3e-07 $layer=LI1_cond $X=2.077 $Y=1.53
+ $X2=2.077 $Y2=1.4
r46 8 32 8.7355 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.105 $Y=1.16
+ $X2=2.105 $Y2=1.4
r47 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.105
+ $Y=1.16 $X2=2.105 $Y2=1.16
r48 6 20 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.025 $Y=1.985
+ $X2=2.025 $Y2=1.33
r49 3 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.025 $Y=0.56 $X2=2.025
+ $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%A1 1 3 5 7 8 12
c34 12 0 1.92762e-19 $X=2.62 $Y=1.16
c35 5 0 1.34745e-19 $X=2.765 $Y=0.965
c36 3 0 1.92208e-19 $X=2.755 $Y=1.985
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.16 $X2=2.62 $Y2=1.16
r38 8 12 2.56098 $w=4.03e-07 $l=9e-08 $layer=LI1_cond $X=2.53 $Y=1.197 $X2=2.62
+ $Y2=1.197
r39 5 11 43.0453 $w=3.83e-07 $l=2.47053e-07 $layer=POLY_cond $X=2.765 $Y=0.965
+ $X2=2.647 $Y2=1.16
r40 5 7 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.765 $Y=0.965
+ $X2=2.765 $Y2=0.56
r41 1 11 38.6406 $w=3.83e-07 $l=2.07075e-07 $layer=POLY_cond $X=2.755 $Y=1.32
+ $X2=2.647 $Y2=1.16
r42 1 3 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.755 $Y=1.32
+ $X2=2.755 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%A2 3 6 8 10 11 12 17 19
r33 17 20 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.16
+ $X2=3.27 $Y2=1.325
r34 17 19 51.398 $w=3.4e-07 $l=1.95e-07 $layer=POLY_cond $X=3.27 $Y=1.16
+ $X2=3.27 $Y2=0.965
r35 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.16 $X2=3.26 $Y2=1.16
r36 12 18 8.10978 $w=2.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.45 $Y=1.155
+ $X2=3.26 $Y2=1.155
r37 10 11 20.3833 $w=1.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.997 $Y=0.51
+ $X2=2.997 $Y2=0.85
r38 9 11 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=2.997 $Y=1.02
+ $X2=2.997 $Y2=0.85
r39 8 18 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.09 $Y=1.155
+ $X2=3.26 $Y2=1.155
r40 8 9 7.13053 $w=2.7e-07 $l=1.75442e-07 $layer=LI1_cond $X=3.09 $Y=1.155
+ $X2=2.997 $Y2=1.02
r41 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.18 $Y=1.985
+ $X2=3.18 $Y2=1.325
r42 3 19 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.175 $Y=0.56
+ $X2=3.175 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%Y 1 2 3 10 14 16 20 22 23 24 25 26 27 34
c48 23 0 8.2804e-20 $X=0.23 $Y=0.85
r49 27 47 2.54435 $w=3.83e-07 $l=8.5e-08 $layer=LI1_cond $X=0.337 $Y=2.21
+ $X2=0.337 $Y2=2.295
r50 26 27 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.337 $Y=1.87
+ $X2=0.337 $Y2=2.21
r51 26 41 7.78273 $w=3.83e-07 $l=2.6e-07 $layer=LI1_cond $X=0.337 $Y=1.87
+ $X2=0.337 $Y2=1.61
r52 25 41 2.39469 $w=3.83e-07 $l=8e-08 $layer=LI1_cond $X=0.337 $Y=1.53
+ $X2=0.337 $Y2=1.61
r53 24 25 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.337 $Y=1.19
+ $X2=0.337 $Y2=1.53
r54 23 34 2.56146 $w=3.85e-07 $l=9e-08 $layer=LI1_cond $X=0.337 $Y=0.79
+ $X2=0.337 $Y2=0.88
r55 23 24 8.4712 $w=3.83e-07 $l=2.83e-07 $layer=LI1_cond $X=0.337 $Y=0.907
+ $X2=0.337 $Y2=1.19
r56 23 34 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=0.337 $Y=0.907
+ $X2=0.337 $Y2=0.88
r57 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.255 $Y=0.705
+ $X2=2.255 $Y2=0.39
r58 17 22 8.35232 $w=1.77e-07 $l=1.65997e-07 $layer=LI1_cond $X=1.375 $Y=0.792
+ $X2=1.21 $Y2=0.79
r59 16 18 16.7588 $w=1.15e-07 $l=2.03912e-07 $layer=LI1_cond $X=2.09 $Y=0.792
+ $X2=2.255 $Y2=0.705
r60 16 17 45.3143 $w=1.73e-07 $l=7.15e-07 $layer=LI1_cond $X=2.09 $Y=0.792
+ $X2=1.375 $Y2=0.792
r61 12 22 0.762005 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.21 $Y=0.7 $X2=1.21
+ $Y2=0.79
r62 12 14 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.21 $Y=0.7 $X2=1.21
+ $Y2=0.39
r63 11 23 5.4929 $w=1.8e-07 $l=1.93e-07 $layer=LI1_cond $X=0.53 $Y=0.79
+ $X2=0.337 $Y2=0.79
r64 10 22 8.35232 $w=1.77e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.79
+ $X2=1.21 $Y2=0.79
r65 10 11 31.7323 $w=1.78e-07 $l=5.15e-07 $layer=LI1_cond $X=1.045 $Y=0.79
+ $X2=0.53 $Y2=0.79
r66 3 47 400 $w=1.7e-07 $l=9.3314e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.485 $X2=0.445 $Y2=2.295
r67 3 41 400 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.485 $X2=0.445 $Y2=1.61
r68 2 20 91 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_NDIFF $count=2 $X=2.1
+ $Y=0.235 $X2=2.255 $Y2=0.39
r69 1 14 91 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.235 $X2=1.21 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%A_420_297# 1 2 9 11 12 15
r21 13 15 7.9627 $w=1.93e-07 $l=1.4e-07 $layer=LI1_cond $X=3.407 $Y=1.75
+ $X2=3.407 $Y2=1.89
r22 11 13 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=3.31 $Y=1.665
+ $X2=3.407 $Y2=1.75
r23 11 12 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.31 $Y=1.665
+ $X2=2.625 $Y2=1.665
r24 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.51 $Y=1.75
+ $X2=2.625 $Y2=1.665
r25 7 9 4.50956 $w=2.28e-07 $l=9e-08 $layer=LI1_cond $X=2.51 $Y=1.75 $X2=2.51
+ $Y2=1.84
r26 2 15 300 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=2 $X=3.255
+ $Y=1.485 $X2=3.395 $Y2=1.89
r27 1 9 300 $w=1.7e-07 $l=5.91439e-07 $layer=licon1_PDIFF $count=2 $X=2.1
+ $Y=1.485 $X2=2.54 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%VPWR 1 6 8 10 20 21 24
r37 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r38 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r39 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r40 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=2.72
+ $X2=2.965 $Y2=2.72
r41 18 20 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.13 $Y=2.72 $X2=3.45
+ $Y2=2.72
r42 17 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 16 17 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 12 16 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=2.72
+ $X2=2.965 $Y2=2.72
r46 10 16 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.8 $Y=2.72 $X2=2.53
+ $Y2=2.72
r47 8 17 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 8 12 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r49 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=2.635
+ $X2=2.965 $Y2=2.72
r50 4 6 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.965 $Y=2.635
+ $X2=2.965 $Y2=2.005
r51 1 6 300 $w=1.7e-07 $l=5.83609e-07 $layer=licon1_PDIFF $count=2 $X=2.83
+ $Y=1.485 $X2=2.965 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_HD__A2111OI_1%VGND 1 2 3 12 16 18 20 23 24 25 31 35 44
+ 48
c51 1 0 8.2804e-20 $X=0.155 $Y=0.235
r52 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r53 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r54 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r55 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r56 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r57 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r58 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r59 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r60 36 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.715
+ $Y2=0
r61 36 38 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.07
+ $Y2=0
r62 35 47 3.86939 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.475
+ $Y2=0
r63 35 41 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=2.99
+ $Y2=0
r64 34 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r65 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r66 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.715
+ $Y2=0
r67 31 33 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=0.69
+ $Y2=0
r68 25 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 25 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 23 28 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.315 $Y=0 $X2=0.23
+ $Y2=0
r71 23 24 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=0.315 $Y=0 $X2=0.472
+ $Y2=0
r72 22 33 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.69
+ $Y2=0
r73 22 24 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.472
+ $Y2=0
r74 18 47 3.20876 $w=2.4e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.475 $Y2=0
r75 18 20 18.7272 $w=2.38e-07 $l=3.9e-07 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0.475
r76 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=0.085
+ $X2=1.715 $Y2=0
r77 14 16 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.715 $Y=0.085
+ $X2=1.715 $Y2=0.37
r78 10 24 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.472 $Y=0.085
+ $X2=0.472 $Y2=0
r79 10 12 10.061 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=0.472 $Y=0.085
+ $X2=0.472 $Y2=0.36
r80 3 20 182 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.235 $X2=3.395 $Y2=0.475
r81 2 16 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.235 $X2=1.715 $Y2=0.37
r82 1 12 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.235 $X2=0.48 $Y2=0.36
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VGND D1 a_44_47# VNB nshort w=650000u l=150000u
+  ad=1.638e+12p pd=1.414e+07u as=9.3925e+11p ps=9.39e+06u
M1001 a_44_47# D1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR A1 a_477_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.365e+12p pd=1.273e+07u as=1.315e+12p ps=1.063e+07u
M1003 a_477_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_477_297# B1 a_285_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1005 a_44_47# D1 a_30_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.8e+11p pd=2.56e+06u as=8.05e+11p ps=7.61e+06u
M1006 a_285_297# C1 a_30_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_44_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1008 a_44_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_44_47# VGND VNB nshort w=650000u l=150000u
+  ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1010 a_770_47# A1 a_44_47# VNB nshort w=650000u l=150000u
+  ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1011 VGND A2 a_770_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_44_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_44_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_285_297# B1 a_477_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND C1 a_44_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_44_47# C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_477_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_30_297# D1 a_44_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND B1 a_44_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_44_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_44_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_770_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A2 a_477_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_30_297# C1 a_285_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_44_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_44_47# A1 a_770_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_44_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

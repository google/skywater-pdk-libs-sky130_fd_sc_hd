# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__clkdlybuf4s25_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.485000 1.320000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.702900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015000 0.255000 3.595000 0.640000 ;
        RECT 3.035000 1.565000 3.595000 2.465000 ;
        RECT 3.230000 0.640000 3.595000 1.565000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.580000  0.085000 0.910000 0.565000 ;
        RECT 2.240000  0.085000 2.845000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.600000 1.830000 0.925000 2.635000 ;
        RECT 2.235000 1.835000 2.845000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.410000 0.735000 ;
      RECT 0.085000 0.735000 1.005000 0.905000 ;
      RECT 0.085000 1.490000 1.005000 1.660000 ;
      RECT 0.085000 1.660000 0.430000 2.465000 ;
      RECT 0.655000 0.905000 1.005000 1.025000 ;
      RECT 0.655000 1.025000 1.105000 1.295000 ;
      RECT 0.655000 1.295000 1.005000 1.490000 ;
      RECT 1.175000 0.255000 1.645000 0.855000 ;
      RECT 1.195000 1.790000 1.645000 2.465000 ;
      RECT 1.470000 0.855000 1.645000 1.075000 ;
      RECT 1.470000 1.075000 2.420000 1.250000 ;
      RECT 1.470000 1.250000 1.645000 1.790000 ;
      RECT 1.815000 0.255000 2.065000 0.735000 ;
      RECT 1.815000 0.735000 2.765000 0.905000 ;
      RECT 1.815000 1.495000 2.765000 1.665000 ;
      RECT 1.815000 1.665000 2.065000 2.465000 ;
      RECT 2.595000 0.905000 2.765000 0.990000 ;
      RECT 2.595000 0.990000 3.050000 1.325000 ;
      RECT 2.595000 1.325000 2.765000 1.495000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_1
END LIBRARY

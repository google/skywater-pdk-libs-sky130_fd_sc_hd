* File: sky130_fd_sc_hd__sdfxbp_1.spice.SKY130_FD_SC_HD__SDFXBP_1.pxi
* Created: Thu Aug 27 14:47:01 2020
* 
x_PM_SKY130_FD_SC_HD__SDFXBP_1%CLK N_CLK_c_239_n N_CLK_c_243_n N_CLK_c_240_n
+ N_CLK_M1034_g N_CLK_c_244_n N_CLK_M1017_g N_CLK_c_245_n CLK
+ PM_SKY130_FD_SC_HD__SDFXBP_1%CLK
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_27_47# N_A_27_47#_M1034_s N_A_27_47#_M1017_s
+ N_A_27_47#_M1021_g N_A_27_47#_M1000_g N_A_27_47#_M1031_g N_A_27_47#_c_283_n
+ N_A_27_47#_c_284_n N_A_27_47#_M1022_g N_A_27_47#_M1006_g N_A_27_47#_c_285_n
+ N_A_27_47#_M1004_g N_A_27_47#_c_518_p N_A_27_47#_c_287_n N_A_27_47#_c_288_n
+ N_A_27_47#_c_300_n N_A_27_47#_c_289_n N_A_27_47#_c_418_p N_A_27_47#_c_301_n
+ N_A_27_47#_c_302_n N_A_27_47#_c_290_n N_A_27_47#_c_303_n N_A_27_47#_c_304_n
+ N_A_27_47#_c_305_n N_A_27_47#_c_306_n N_A_27_47#_c_307_n N_A_27_47#_c_291_n
+ N_A_27_47#_c_309_n N_A_27_47#_c_310_n N_A_27_47#_c_311_n N_A_27_47#_c_292_n
+ N_A_27_47#_c_293_n PM_SKY130_FD_SC_HD__SDFXBP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%SCE N_SCE_M1008_g N_SCE_M1026_g N_SCE_c_538_n
+ N_SCE_M1024_g N_SCE_M1029_g N_SCE_c_529_n N_SCE_c_530_n N_SCE_c_541_n
+ N_SCE_c_531_n N_SCE_c_532_n N_SCE_c_533_n N_SCE_c_534_n N_SCE_c_535_n SCE
+ PM_SKY130_FD_SC_HD__SDFXBP_1%SCE
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_299_47# N_A_299_47#_M1008_s N_A_299_47#_M1026_s
+ N_A_299_47#_M1019_g N_A_299_47#_M1018_g N_A_299_47#_c_645_n
+ N_A_299_47#_c_652_n N_A_299_47#_c_660_n N_A_299_47#_c_646_n
+ N_A_299_47#_c_662_n N_A_299_47#_c_654_n N_A_299_47#_c_647_n
+ N_A_299_47#_c_655_n N_A_299_47#_c_648_n N_A_299_47#_c_649_n
+ N_A_299_47#_c_667_n N_A_299_47#_c_656_n N_A_299_47#_c_657_n
+ PM_SKY130_FD_SC_HD__SDFXBP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%D N_D_M1027_g N_D_M1020_g D N_D_c_773_n
+ N_D_c_774_n PM_SKY130_FD_SC_HD__SDFXBP_1%D
x_PM_SKY130_FD_SC_HD__SDFXBP_1%SCD N_SCD_M1012_g N_SCD_M1014_g SCD N_SCD_c_822_n
+ PM_SKY130_FD_SC_HD__SDFXBP_1%SCD
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_193_47# N_A_193_47#_M1021_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1003_g N_A_193_47#_M1032_g N_A_193_47#_c_869_n
+ N_A_193_47#_M1002_g N_A_193_47#_M1035_g N_A_193_47#_c_870_n
+ N_A_193_47#_c_885_n N_A_193_47#_c_871_n N_A_193_47#_c_872_n
+ N_A_193_47#_c_887_n N_A_193_47#_c_888_n N_A_193_47#_c_873_n
+ N_A_193_47#_c_874_n N_A_193_47#_c_875_n N_A_193_47#_c_1005_p
+ N_A_193_47#_c_876_n N_A_193_47#_c_877_n N_A_193_47#_c_878_n
+ N_A_193_47#_c_879_n N_A_193_47#_c_880_n N_A_193_47#_c_881_n
+ PM_SKY130_FD_SC_HD__SDFXBP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_1089_183# N_A_1089_183#_M1013_d
+ N_A_1089_183#_M1025_d N_A_1089_183#_M1005_g N_A_1089_183#_M1009_g
+ N_A_1089_183#_c_1083_n N_A_1089_183#_c_1109_n N_A_1089_183#_c_1129_p
+ N_A_1089_183#_c_1110_n N_A_1089_183#_c_1084_n N_A_1089_183#_c_1085_n
+ N_A_1089_183#_c_1097_n N_A_1089_183#_c_1086_n N_A_1089_183#_c_1087_n
+ PM_SKY130_FD_SC_HD__SDFXBP_1%A_1089_183#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_930_413# N_A_930_413#_M1031_d
+ N_A_930_413#_M1003_d N_A_930_413#_c_1176_n N_A_930_413#_M1025_g
+ N_A_930_413#_c_1177_n N_A_930_413#_M1013_g N_A_930_413#_c_1178_n
+ N_A_930_413#_c_1179_n N_A_930_413#_c_1180_n N_A_930_413#_c_1194_n
+ N_A_930_413#_c_1220_n N_A_930_413#_c_1181_n N_A_930_413#_c_1186_n
+ N_A_930_413#_c_1182_n PM_SKY130_FD_SC_HD__SDFXBP_1%A_930_413#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_1517_315# N_A_1517_315#_M1011_s
+ N_A_1517_315#_M1001_s N_A_1517_315#_M1015_g N_A_1517_315#_M1016_g
+ N_A_1517_315#_c_1285_n N_A_1517_315#_M1010_g N_A_1517_315#_M1028_g
+ N_A_1517_315#_c_1286_n N_A_1517_315#_c_1287_n N_A_1517_315#_c_1288_n
+ N_A_1517_315#_M1033_g N_A_1517_315#_M1030_g N_A_1517_315#_c_1300_n
+ N_A_1517_315#_c_1301_n N_A_1517_315#_c_1302_n N_A_1517_315#_c_1303_n
+ N_A_1517_315#_c_1289_n N_A_1517_315#_c_1316_p N_A_1517_315#_c_1290_n
+ N_A_1517_315#_c_1304_n N_A_1517_315#_c_1291_n N_A_1517_315#_c_1292_n
+ N_A_1517_315#_c_1293_n N_A_1517_315#_c_1318_p N_A_1517_315#_c_1323_p
+ PM_SKY130_FD_SC_HD__SDFXBP_1%A_1517_315#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_1346_413# N_A_1346_413#_M1002_d
+ N_A_1346_413#_M1006_d N_A_1346_413#_c_1409_n N_A_1346_413#_M1011_g
+ N_A_1346_413#_M1001_g N_A_1346_413#_c_1410_n N_A_1346_413#_c_1411_n
+ N_A_1346_413#_c_1421_n N_A_1346_413#_c_1424_n N_A_1346_413#_c_1418_n
+ N_A_1346_413#_c_1412_n N_A_1346_413#_c_1413_n N_A_1346_413#_c_1414_n
+ PM_SKY130_FD_SC_HD__SDFXBP_1%A_1346_413#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_1948_47# N_A_1948_47#_M1033_s
+ N_A_1948_47#_M1030_s N_A_1948_47#_M1023_g N_A_1948_47#_M1007_g
+ N_A_1948_47#_c_1503_n N_A_1948_47#_c_1504_n N_A_1948_47#_c_1497_n
+ N_A_1948_47#_c_1498_n N_A_1948_47#_c_1499_n N_A_1948_47#_c_1500_n
+ N_A_1948_47#_c_1507_n N_A_1948_47#_c_1523_n N_A_1948_47#_c_1501_n
+ PM_SKY130_FD_SC_HD__SDFXBP_1%A_1948_47#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%VPWR N_VPWR_M1017_d N_VPWR_M1026_d N_VPWR_M1014_d
+ N_VPWR_M1005_d N_VPWR_M1015_d N_VPWR_M1001_d N_VPWR_M1030_d N_VPWR_c_1558_n
+ N_VPWR_c_1559_n N_VPWR_c_1560_n N_VPWR_c_1561_n N_VPWR_c_1562_n
+ N_VPWR_c_1563_n N_VPWR_c_1564_n N_VPWR_c_1565_n N_VPWR_c_1566_n
+ N_VPWR_c_1567_n N_VPWR_c_1568_n N_VPWR_c_1569_n N_VPWR_c_1570_n VPWR
+ N_VPWR_c_1571_n N_VPWR_c_1572_n N_VPWR_c_1573_n N_VPWR_c_1574_n
+ N_VPWR_c_1575_n N_VPWR_c_1557_n N_VPWR_c_1577_n N_VPWR_c_1578_n
+ N_VPWR_c_1579_n N_VPWR_c_1580_n PM_SKY130_FD_SC_HD__SDFXBP_1%VPWR
x_PM_SKY130_FD_SC_HD__SDFXBP_1%A_556_369# N_A_556_369#_M1020_d
+ N_A_556_369#_M1031_s N_A_556_369#_M1027_d N_A_556_369#_M1003_s
+ N_A_556_369#_c_1739_n N_A_556_369#_c_1751_n N_A_556_369#_c_1763_n
+ N_A_556_369#_c_1728_n N_A_556_369#_c_1735_n N_A_556_369#_c_1736_n
+ N_A_556_369#_c_1729_n N_A_556_369#_c_1730_n N_A_556_369#_c_1731_n
+ N_A_556_369#_c_1732_n N_A_556_369#_c_1733_n N_A_556_369#_c_1734_n
+ N_A_556_369#_c_1738_n PM_SKY130_FD_SC_HD__SDFXBP_1%A_556_369#
x_PM_SKY130_FD_SC_HD__SDFXBP_1%Q N_Q_M1010_d N_Q_M1028_d N_Q_c_1854_n
+ N_Q_c_1851_n N_Q_c_1852_n Q N_Q_c_1853_n PM_SKY130_FD_SC_HD__SDFXBP_1%Q
x_PM_SKY130_FD_SC_HD__SDFXBP_1%Q_N N_Q_N_M1023_d N_Q_N_M1007_d N_Q_N_c_1894_n
+ N_Q_N_c_1895_n Q_N Q_N PM_SKY130_FD_SC_HD__SDFXBP_1%Q_N
x_PM_SKY130_FD_SC_HD__SDFXBP_1%VGND N_VGND_M1034_d N_VGND_M1008_d N_VGND_M1012_d
+ N_VGND_M1009_d N_VGND_M1016_d N_VGND_M1011_d N_VGND_M1033_d N_VGND_c_1909_n
+ N_VGND_c_1910_n N_VGND_c_1911_n N_VGND_c_1912_n N_VGND_c_1913_n
+ N_VGND_c_1914_n N_VGND_c_1915_n N_VGND_c_1916_n N_VGND_c_1917_n
+ N_VGND_c_1918_n VGND N_VGND_c_1919_n N_VGND_c_1920_n N_VGND_c_1921_n
+ N_VGND_c_1922_n N_VGND_c_1923_n N_VGND_c_1924_n N_VGND_c_1925_n
+ N_VGND_c_1926_n N_VGND_c_1927_n N_VGND_c_1928_n N_VGND_c_1929_n
+ N_VGND_c_1930_n N_VGND_c_1931_n PM_SKY130_FD_SC_HD__SDFXBP_1%VGND
cc_1 VNB N_CLK_c_239_n 0.0573151f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_240_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0185843f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1021_g 0.0410581f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1031_g 0.0525494f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_6 VNB N_A_27_47#_c_283_n 0.0136466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_284_n 0.00284024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_285_n 0.0158261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1004_g 0.043789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_287_n 0.00318197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_288_n 0.00642096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_289_n 8.11193e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_290_n 0.00236945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_291_n 0.0224414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_292_n 0.00980165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_293_n 0.00148891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_SCE_M1008_g 0.0506763f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_18 VNB N_SCE_M1029_g 0.016865f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_19 VNB N_SCE_c_529_n 0.00224546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_SCE_c_530_n 0.00335978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_531_n 0.00187885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_532_n 0.00348269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_533_n 0.00118673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_534_n 0.0272701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_SCE_c_535_n 0.00148358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_299_47#_M1019_g 0.0216917f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_27 VNB N_A_299_47#_c_645_n 0.0128083f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_28 VNB N_A_299_47#_c_646_n 0.00262794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_299_47#_c_647_n 0.00450023f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_299_47#_c_648_n 0.00285099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_299_47#_c_649_n 0.0296746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_D_M1020_g 0.0443734f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_33 VNB N_SCD_M1012_g 0.0446303f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_34 VNB SCD 0.0123904f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_35 VNB N_SCD_c_822_n 0.0122397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_869_n 0.0180432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_870_n 0.00330484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_871_n 0.00369255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_193_47#_c_872_n 0.00632811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_873_n 0.0497048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_193_47#_c_874_n 0.00617885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_193_47#_c_875_n 0.0101801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_193_47#_c_876_n 0.00567379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_193_47#_c_877_n 9.18319e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_193_47#_c_878_n 0.0266741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_193_47#_c_879_n 0.0176138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_193_47#_c_880_n 0.0285203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_193_47#_c_881_n 0.0117653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1089_183#_M1005_g 0.0146965f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_50 VNB N_A_1089_183#_M1009_g 0.0210316f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_51 VNB N_A_1089_183#_c_1083_n 0.00354578f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_52 VNB N_A_1089_183#_c_1084_n 0.00364457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1089_183#_c_1085_n 0.00130441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1089_183#_c_1086_n 0.00302393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1089_183#_c_1087_n 0.0338642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_930_413#_c_1176_n 0.0118275f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_57 VNB N_A_930_413#_c_1177_n 0.0158415f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_58 VNB N_A_930_413#_c_1178_n 0.0152351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_930_413#_c_1179_n 0.00913873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_930_413#_c_1180_n 8.51874e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_930_413#_c_1181_n 0.0118177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_930_413#_c_1182_n 0.00180949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1517_315#_M1016_g 0.0476879f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_64 VNB N_A_1517_315#_c_1285_n 0.0195286f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_65 VNB N_A_1517_315#_c_1286_n 0.0415081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1517_315#_c_1287_n 0.0304242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1517_315#_c_1288_n 0.0178307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1517_315#_c_1289_n 0.00408987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1517_315#_c_1290_n 0.00158679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1517_315#_c_1291_n 0.00373683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1517_315#_c_1292_n 0.0128859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1517_315#_c_1293_n 0.00292904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1346_413#_c_1409_n 0.0201807f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_74 VNB N_A_1346_413#_c_1410_n 0.0419509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1346_413#_c_1411_n 0.00807206f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_76 VNB N_A_1346_413#_c_1412_n 0.00867958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1346_413#_c_1413_n 0.00584041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1346_413#_c_1414_n 0.00344545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1948_47#_c_1497_n 0.00309662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1948_47#_c_1498_n 0.00338009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1948_47#_c_1499_n 0.0240537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1948_47#_c_1500_n 0.00317036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1948_47#_c_1501_n 0.0199524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VPWR_c_1557_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_556_369#_c_1728_n 3.46824e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_556_369#_c_1729_n 0.0111787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_556_369#_c_1730_n 0.00215513f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_556_369#_c_1731_n 0.0038877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_556_369#_c_1732_n 0.00876794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_556_369#_c_1733_n 0.00235887f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_556_369#_c_1734_n 0.00172885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_Q_c_1851_n 0.00221068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_Q_c_1852_n 0.00248461f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_94 VNB N_Q_c_1853_n 0.00467334f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_95 VNB N_Q_N_c_1894_n 0.0154962f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_96 VNB N_Q_N_c_1895_n 0.00479254f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_97 VNB Q_N 0.0240401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1909_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1910_n 0.00286037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1911_n 0.00486519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1912_n 0.0452421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1913_n 0.0058544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1914_n 0.00237946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1915_n 0.0046493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1916_n 0.00436529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1917_n 0.0430904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1918_n 0.00513917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1919_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1920_n 0.029404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1921_n 0.0346399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1922_n 0.0216134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1923_n 0.0322774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1924_n 0.0154689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1925_n 0.527847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1926_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1927_n 0.00512961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1928_n 0.0038195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1929_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1930_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1931_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VPB N_CLK_c_239_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_122 VPB N_CLK_c_243_n 0.0162092f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_123 VPB N_CLK_c_244_n 0.01861f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_124 VPB N_CLK_c_245_n 0.0230979f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_125 VPB CLK 0.017656f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_126 VPB N_A_27_47#_M1000_g 0.038975f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_127 VPB N_A_27_47#_c_283_n 0.0143056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_284_n 0.0057729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_M1022_g 0.0191311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_M1006_g 0.033754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_285_n 0.0211417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_300_n 0.00202859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_301_n 0.00333071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_302_n 0.00357396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_303_n 0.0580659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_304_n 0.00130312f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_305_n 0.00111253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_27_47#_c_306_n 9.17012e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_27_47#_c_307_n 0.00543917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_291_n 0.0114072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_309_n 0.0266783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_310_n 0.00853708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_311_n 0.0106236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_292_n 0.0208929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_293_n 0.00437972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_SCE_M1008_g 0.00509208f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_147 VPB N_SCE_M1026_g 0.0236415f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_148 VPB N_SCE_c_538_n 0.0166224f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_149 VPB N_SCE_M1024_g 0.0194307f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_150 VPB N_SCE_c_530_n 0.0010494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_SCE_c_541_n 0.0293624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_299_47#_M1018_g 0.0184813f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_153 VPB N_A_299_47#_c_645_n 0.0107801f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_154 VPB N_A_299_47#_c_652_n 0.00446885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_299_47#_c_646_n 0.00415603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_299_47#_c_654_n 0.00158406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_299_47#_c_655_n 0.00201239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_299_47#_c_656_n 0.0014433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_299_47#_c_657_n 0.027856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_D_M1027_g 0.0190456f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_161 VPB N_D_M1020_g 0.00360779f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_162 VPB N_D_c_773_n 0.0269869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_D_c_774_n 0.0044856f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_164 VPB N_SCD_M1014_g 0.0328228f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_165 VPB SCD 0.00992144f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_166 VPB N_SCD_c_822_n 0.0182053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_193_47#_M1003_g 0.024991f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_168 VPB N_A_193_47#_M1035_g 0.0221869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_193_47#_c_870_n 0.00462988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_193_47#_c_885_n 0.0328226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_193_47#_c_871_n 0.00311128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_193_47#_c_887_n 0.00568481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_193_47#_c_888_n 0.0266658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_193_47#_c_881_n 0.0113861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1089_183#_M1005_g 0.049805f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_176 VPB N_A_1089_183#_c_1086_n 0.00255179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_930_413#_M1025_g 0.0226707f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_178 VPB N_A_930_413#_c_1179_n 0.0189969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_930_413#_c_1180_n 0.00681499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_930_413#_c_1186_n 0.00161138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_930_413#_c_1182_n 0.00887906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1517_315#_M1015_g 0.0252633f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_183 VPB N_A_1517_315#_M1016_g 0.0178079f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_184 VPB N_A_1517_315#_M1028_g 0.0223568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1517_315#_c_1286_n 0.0189622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1517_315#_c_1287_n 5.42563e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1517_315#_M1030_g 0.0252559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1517_315#_c_1300_n 0.0126982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1517_315#_c_1301_n 0.0137898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1517_315#_c_1302_n 0.0129003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_1517_315#_c_1303_n 0.040764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1517_315#_c_1304_n 0.00231467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1517_315#_c_1291_n 0.00373683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1517_315#_c_1292_n 0.00347878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_1346_413#_M1001_g 0.0233466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_1346_413#_c_1410_n 0.0157032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1346_413#_c_1411_n 5.11281e-19 $X=-0.19 $Y=1.305 $X2=0.33
+ $Y2=1.16
cc_198 VPB N_A_1346_413#_c_1418_n 0.0126839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1346_413#_c_1412_n 0.00349335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1346_413#_c_1413_n 0.0050339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1948_47#_M1007_g 0.0229554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_1948_47#_c_1503_n 0.0026305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1948_47#_c_1504_n 0.00527279f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_204 VPB N_A_1948_47#_c_1498_n 0.00405051f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1948_47#_c_1499_n 0.00481435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_1948_47#_c_1507_n 0.00281561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1558_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1559_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1560_n 0.00470486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1561_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1562_n 0.00548955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1563_n 0.00467156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1564_n 0.00507267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1565_n 0.0374334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1566_n 0.00324297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1567_n 0.0511015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1568_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1569_n 0.0449606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1570_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1571_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1572_n 0.0259272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1573_n 0.0217823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1574_n 0.0320609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1575_n 0.0159936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1557_n 0.0701627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1577_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1578_n 0.00436214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1579_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1580_n 0.00459796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_A_556_369#_c_1735_n 0.00775461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_556_369#_c_1736_n 0.00155557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_556_369#_c_1732_n 0.0110086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_556_369#_c_1738_n 0.00883626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_Q_c_1854_n 0.00941153f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_235 VPB N_Q_c_1851_n 0.00672426f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB Q_N 0.0420025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 N_CLK_c_239_n N_A_27_47#_M1021_g 0.0049062f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_238 N_CLK_c_240_n N_A_27_47#_M1021_g 0.0187731f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_239 CLK N_A_27_47#_M1021_g 3.14819e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_240 N_CLK_c_243_n N_A_27_47#_M1000_g 0.00541775f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_241 N_CLK_c_245_n N_A_27_47#_M1000_g 0.0276441f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_242 CLK N_A_27_47#_M1000_g 5.77812e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_243 N_CLK_c_239_n N_A_27_47#_c_287_n 0.00761961f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_244 N_CLK_c_240_n N_A_27_47#_c_287_n 0.00668648f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_245 CLK N_A_27_47#_c_287_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_246 N_CLK_c_239_n N_A_27_47#_c_288_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_247 CLK N_A_27_47#_c_288_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_248 N_CLK_c_244_n N_A_27_47#_c_300_n 0.0126874f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_249 N_CLK_c_245_n N_A_27_47#_c_300_n 0.00142281f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_250 CLK N_A_27_47#_c_300_n 0.00766156f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_251 N_CLK_c_239_n N_A_27_47#_c_289_n 3.98708e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_252 CLK N_A_27_47#_c_289_n 0.0516739f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_253 N_CLK_c_239_n N_A_27_47#_c_301_n 2.90926e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_254 N_CLK_c_243_n N_A_27_47#_c_301_n 7.07325e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_255 N_CLK_c_245_n N_A_27_47#_c_301_n 0.00436768f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_256 N_CLK_c_239_n N_A_27_47#_c_302_n 2.46885e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_257 N_CLK_c_244_n N_A_27_47#_c_302_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_258 N_CLK_c_245_n N_A_27_47#_c_302_n 0.00343236f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_259 CLK N_A_27_47#_c_302_n 0.0153591f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_260 N_CLK_c_239_n N_A_27_47#_c_290_n 0.00381855f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_261 N_CLK_c_244_n N_A_27_47#_c_304_n 0.00100532f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_262 N_CLK_c_239_n N_A_27_47#_c_291_n 0.0169118f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_263 CLK N_A_27_47#_c_291_n 0.00161603f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_264 N_CLK_c_244_n N_VPWR_c_1558_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_265 N_CLK_c_244_n N_VPWR_c_1571_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_266 N_CLK_c_244_n N_VPWR_c_1557_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_267 N_CLK_c_240_n N_VGND_c_1909_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_268 N_CLK_c_239_n N_VGND_c_1919_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_269 N_CLK_c_240_n N_VGND_c_1919_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_270 N_CLK_c_240_n N_VGND_c_1925_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_303_n N_SCE_M1026_g 0.002769f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_303_n N_SCE_M1024_g 0.00141925f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_303_n N_SCE_c_530_n 0.00408513f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_274 N_A_27_47#_M1000_g N_SCE_c_541_n 0.0023159f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_303_n N_SCE_c_541_n 0.00373131f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_303_n N_A_299_47#_M1018_g 7.69535e-19 $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_303_n N_A_299_47#_c_645_n 0.0121775f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_303_n N_A_299_47#_c_660_n 0.0158079f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_303_n N_A_299_47#_c_646_n 0.00932251f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_303_n N_A_299_47#_c_662_n 0.0368525f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_303_n N_A_299_47#_c_654_n 0.0113096f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1021_g N_A_299_47#_c_647_n 0.00159333f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_303_n N_A_299_47#_c_655_n 0.0137968f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_303_n N_A_299_47#_c_649_n 0.00262198f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_303_n N_A_299_47#_c_667_n 0.0046091f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_303_n N_A_299_47#_c_656_n 7.81108e-19 $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_303_n N_A_299_47#_c_657_n 0.0016565f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_303_n N_D_M1027_g 0.00217769f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_303_n N_D_c_773_n 0.00308822f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_303_n N_D_c_774_n 0.0085184f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_303_n N_SCD_M1014_g 0.00188492f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_303_n SCD 0.0122303f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_293 N_A_27_47#_M1031_g N_SCD_c_822_n 0.00189664f $X=4.58 $Y=0.415 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_303_n N_A_193_47#_M1000_d 0.00126326f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_303_n N_A_193_47#_M1003_g 0.00371812f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_309_n N_A_193_47#_M1003_g 0.0144149f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_310_n N_A_193_47#_M1003_g 9.60176e-19 $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1004_g N_A_193_47#_c_869_n 0.0144677f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1006_g N_A_193_47#_M1035_g 0.0175056f $X=6.655 $Y=2.275 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_307_n N_A_193_47#_M1035_g 0.00135837f $X=6.66 $Y=1.87 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_293_n N_A_193_47#_M1035_g 5.16255e-19 $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1031_g N_A_193_47#_c_870_n 0.00772854f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_283_n N_A_193_47#_c_870_n 0.00687115f $X=4.965 $Y=1.32 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_284_n N_A_193_47#_c_870_n 0.00418731f $X=4.655 $Y=1.32 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_303_n N_A_193_47#_c_870_n 0.0139192f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_306_n N_A_193_47#_c_870_n 2.15174e-19 $X=5.395 $Y=1.87 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_309_n N_A_193_47#_c_870_n 7.29366e-19 $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_310_n N_A_193_47#_c_870_n 0.0168988f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_311_n N_A_193_47#_c_870_n 0.00604391f $X=5.1 $Y=1.575 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_284_n N_A_193_47#_c_885_n 0.0162569f $X=4.655 $Y=1.32 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_303_n N_A_193_47#_c_885_n 0.00545515f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_309_n N_A_193_47#_c_885_n 0.0174998f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_310_n N_A_193_47#_c_885_n 0.00118389f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_285_n N_A_193_47#_c_871_n 0.0117161f $X=7.225 $Y=1.32 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_M1004_g N_A_193_47#_c_871_n 0.00430042f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_292_n N_A_193_47#_c_871_n 0.00402309f $X=6.65 $Y=1.32 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_293_n N_A_193_47#_c_871_n 0.0234373f $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_M1004_g N_A_193_47#_c_872_n 0.0020279f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_292_n N_A_193_47#_c_872_n 0.00222109f $X=6.65 $Y=1.32 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_293_n N_A_193_47#_c_872_n 0.0119224f $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_M1006_g N_A_193_47#_c_887_n 0.00117691f $X=6.655 $Y=2.275
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_c_285_n N_A_193_47#_c_887_n 0.00338756f $X=7.225 $Y=1.32 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_307_n N_A_193_47#_c_887_n 0.00508223f $X=6.66 $Y=1.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_293_n N_A_193_47#_c_887_n 0.0245744f $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1006_g N_A_193_47#_c_888_n 0.0130792f $X=6.655 $Y=2.275 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_285_n N_A_193_47#_c_888_n 0.0212127f $X=7.225 $Y=1.32 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_293_n N_A_193_47#_c_888_n 6.54911e-19 $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_M1031_g N_A_193_47#_c_873_n 0.00225641f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_M1021_g N_A_193_47#_c_874_n 0.00586129f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_287_n N_A_193_47#_c_874_n 0.002018f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_290_n N_A_193_47#_c_874_n 0.00471471f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_292_n N_A_193_47#_c_875_n 2.10748e-19 $X=6.65 $Y=1.32 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_M1031_g N_A_193_47#_c_876_n 0.0116466f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_283_n N_A_193_47#_c_876_n 0.00587088f $X=4.965 $Y=1.32 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_310_n N_A_193_47#_c_876_n 0.00398178f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_292_n N_A_193_47#_c_877_n 9.82747e-19 $X=6.65 $Y=1.32 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_293_n N_A_193_47#_c_877_n 0.00125233f $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_M1031_g N_A_193_47#_c_878_n 0.0213105f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_283_n N_A_193_47#_c_878_n 0.0174066f $X=4.965 $Y=1.32 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_309_n N_A_193_47#_c_878_n 5.43883e-19 $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_310_n N_A_193_47#_c_878_n 4.76262e-19 $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_M1031_g N_A_193_47#_c_879_n 0.0102605f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_M1004_g N_A_193_47#_c_880_n 0.0193601f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_292_n N_A_193_47#_c_880_n 0.020308f $X=6.65 $Y=1.32 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_M1021_g N_A_193_47#_c_881_n 0.0237597f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_287_n N_A_193_47#_c_881_n 0.00996571f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_289_n N_A_193_47#_c_881_n 0.0597702f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_418_p N_A_193_47#_c_881_n 0.00849955f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_290_n N_A_193_47#_c_881_n 0.00895075f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_303_n N_A_193_47#_c_881_n 0.0195358f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_304_n N_A_193_47#_c_881_n 0.00244986f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_305_n N_A_1089_183#_M1025_d 0.00523078f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_283_n N_A_1089_183#_M1005_g 0.0113457f $X=4.965 $Y=1.32
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_M1022_g N_A_1089_183#_M1005_g 0.0276008f $X=5.04 $Y=2.275
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_305_n N_A_1089_183#_M1005_g 0.00281129f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_306_n N_A_1089_183#_M1005_g 0.00148824f $X=5.395 $Y=1.87
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_c_309_n N_A_1089_183#_M1005_g 0.0206011f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_310_n N_A_1089_183#_M1005_g 0.0022f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_305_n N_A_1089_183#_c_1097_n 0.00261642f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_M1006_g N_A_1089_183#_c_1086_n 0.00455971f $X=6.655 $Y=2.275
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_305_n N_A_1089_183#_c_1086_n 0.0193938f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_307_n N_A_1089_183#_c_1086_n 0.00314501f $X=6.66 $Y=1.87
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_292_n N_A_1089_183#_c_1086_n 0.00225153f $X=6.65 $Y=1.32
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_293_n N_A_1089_183#_c_1086_n 0.0517078f $X=6.65 $Y=1.41
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_292_n N_A_930_413#_c_1176_n 0.0158005f $X=6.65 $Y=1.32 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_293_n N_A_930_413#_c_1176_n 3.03019e-19 $X=6.65 $Y=1.41
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_M1006_g N_A_930_413#_M1025_g 0.0247799f $X=6.655 $Y=2.275
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_c_305_n N_A_930_413#_M1025_g 0.00700233f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_293_n N_A_930_413#_M1025_g 8.29633e-19 $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_305_n N_A_930_413#_c_1179_n 0.00109659f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_M1022_g N_A_930_413#_c_1194_n 0.00859863f $X=5.04 $Y=2.275
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_303_n N_A_930_413#_c_1194_n 0.00699281f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_305_n N_A_930_413#_c_1194_n 0.00369623f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_306_n N_A_930_413#_c_1194_n 0.00172439f $X=5.395 $Y=1.87
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_309_n N_A_930_413#_c_1194_n 5.38487e-19 $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_310_n N_A_930_413#_c_1194_n 0.0252832f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_M1031_g N_A_930_413#_c_1181_n 9.86268e-19 $X=4.58 $Y=0.415
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_283_n N_A_930_413#_c_1181_n 8.14452e-19 $X=4.965 $Y=1.32
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_M1022_g N_A_930_413#_c_1186_n 9.97608e-19 $X=5.04 $Y=2.275
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_305_n N_A_930_413#_c_1186_n 0.0183205f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_306_n N_A_930_413#_c_1186_n 0.00258875f $X=5.395 $Y=1.87
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_c_309_n N_A_930_413#_c_1186_n 7.00613e-19 $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_310_n N_A_930_413#_c_1186_n 0.0250097f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_283_n N_A_930_413#_c_1182_n 0.00225879f $X=4.965 $Y=1.32
+ $X2=0 $Y2=0
cc_385 N_A_27_47#_c_305_n N_A_930_413#_c_1182_n 0.0173913f $X=6.515 $Y=1.87
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_306_n N_A_930_413#_c_1182_n 0.00179088f $X=5.395 $Y=1.87
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_310_n N_A_930_413#_c_1182_n 0.00980238f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_311_n N_A_930_413#_c_1182_n 4.44848e-19 $X=5.1 $Y=1.575
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_M1004_g N_A_1517_315#_M1016_g 0.0463015f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_M1006_g N_A_1346_413#_c_1421_n 0.00281529f $X=6.655 $Y=2.275
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_307_n N_A_1346_413#_c_1421_n 0.00210372f $X=6.66 $Y=1.87
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_293_n N_A_1346_413#_c_1421_n 0.0022468f $X=6.65 $Y=1.41
+ $X2=0 $Y2=0
cc_393 N_A_27_47#_M1004_g N_A_1346_413#_c_1424_n 0.00800808f $X=7.3 $Y=0.415
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_307_n N_A_1346_413#_c_1418_n 0.00228172f $X=6.66 $Y=1.87
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_293_n N_A_1346_413#_c_1418_n 9.63849e-19 $X=6.65 $Y=1.41
+ $X2=0 $Y2=0
cc_396 N_A_27_47#_M1004_g N_A_1346_413#_c_1412_n 3.1587e-19 $X=7.3 $Y=0.415
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_285_n N_A_1346_413#_c_1413_n 0.00557118f $X=7.225 $Y=1.32
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_M1004_g N_A_1346_413#_c_1413_n 0.0061466f $X=7.3 $Y=0.415
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_M1004_g N_A_1346_413#_c_1414_n 0.0110517f $X=7.3 $Y=0.415
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_418_p N_VPWR_M1017_d 6.67509e-19 $X=0.73 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_401 N_A_27_47#_c_304_n N_VPWR_M1017_d 0.00172249f $X=0.875 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_402 N_A_27_47#_c_305_n N_VPWR_M1005_d 0.00678497f $X=6.515 $Y=1.87 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_M1000_g N_VPWR_c_1558_n 0.00944765f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_300_n N_VPWR_c_1558_n 0.00328537f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_c_418_p N_VPWR_c_1558_n 0.013292f $X=0.73 $Y=1.795 $X2=0 $Y2=0
cc_406 N_A_27_47#_c_302_n N_VPWR_c_1558_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_407 N_A_27_47#_c_304_n N_VPWR_c_1558_n 0.00309407f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_c_303_n N_VPWR_c_1559_n 0.00124161f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_303_n N_VPWR_c_1560_n 8.00522e-19 $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_c_305_n N_VPWR_c_1561_n 0.00950843f $X=6.515 $Y=1.87 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_M1022_g N_VPWR_c_1567_n 0.0037886f $X=5.04 $Y=2.275 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_M1006_g N_VPWR_c_1569_n 0.00430107f $X=6.655 $Y=2.275 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_293_n N_VPWR_c_1569_n 0.00157744f $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_300_n N_VPWR_c_1571_n 0.0018545f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_302_n N_VPWR_c_1571_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_416 N_A_27_47#_M1000_g N_VPWR_c_1572_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_M1000_g N_VPWR_c_1557_n 0.00533769f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_M1022_g N_VPWR_c_1557_n 0.00557377f $X=5.04 $Y=2.275 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_M1006_g N_VPWR_c_1557_n 0.0057371f $X=6.655 $Y=2.275 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_300_n N_VPWR_c_1557_n 0.0040694f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_302_n N_VPWR_c_1557_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_303_n N_VPWR_c_1557_n 0.197356f $X=5.105 $Y=1.87 $X2=0 $Y2=0
cc_423 N_A_27_47#_c_304_n N_VPWR_c_1557_n 0.0146019f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_305_n N_VPWR_c_1557_n 0.053022f $X=6.515 $Y=1.87 $X2=0 $Y2=0
cc_425 N_A_27_47#_c_306_n N_VPWR_c_1557_n 0.0147031f $X=5.395 $Y=1.87 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_c_307_n N_VPWR_c_1557_n 0.0159329f $X=6.66 $Y=1.87 $X2=0 $Y2=0
cc_427 N_A_27_47#_c_293_n N_VPWR_c_1557_n 0.00100625f $X=6.65 $Y=1.41 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_303_n N_A_556_369#_c_1739_n 0.00584375f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_303_n N_A_556_369#_c_1735_n 0.0216422f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_303_n N_A_556_369#_c_1736_n 0.0102354f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_M1031_g N_A_556_369#_c_1731_n 0.00490278f $X=4.58 $Y=0.415
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_M1031_g N_A_556_369#_c_1732_n 0.00639354f $X=4.58 $Y=0.415
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_303_n N_A_556_369#_c_1732_n 0.0104876f $X=5.105 $Y=1.87
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_M1031_g N_A_556_369#_c_1733_n 0.00178202f $X=4.58 $Y=0.415
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_M1031_g N_A_556_369#_c_1734_n 0.00125885f $X=4.58 $Y=0.415
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_303_n N_A_556_369#_c_1738_n 0.01281f $X=5.105 $Y=1.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_310_n N_A_556_369#_c_1738_n 0.00314032f $X=5.1 $Y=1.74 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_303_n A_640_369# 0.00134881f $X=5.105 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_439 N_A_27_47#_c_287_n N_VGND_M1034_d 0.00166329f $X=0.615 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_440 N_A_27_47#_M1021_g N_VGND_c_1909_n 0.00954815f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_c_287_n N_VGND_c_1909_n 0.0150403f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_289_n N_VGND_c_1909_n 0.00108069f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_291_n N_VGND_c_1909_n 5.70216e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_M1031_g N_VGND_c_1911_n 0.00353857f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_M1031_g N_VGND_c_1912_n 0.00431421f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_M1004_g N_VGND_c_1914_n 0.00230753f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_M1004_g N_VGND_c_1917_n 0.00379696f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_518_p N_VGND_c_1919_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_287_n N_VGND_c_1919_n 0.00243651f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_M1021_g N_VGND_c_1920_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_M1034_s N_VGND_c_1925_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_M1021_g N_VGND_c_1925_n 0.00904511f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_M1031_g N_VGND_c_1925_n 0.00721977f $X=4.58 $Y=0.415 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_M1004_g N_VGND_c_1925_n 0.00575728f $X=7.3 $Y=0.415 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_518_p N_VGND_c_1925_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_287_n N_VGND_c_1925_n 0.00564532f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_457 N_SCE_M1008_g N_A_299_47#_M1019_g 0.0204149f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_458 N_SCE_c_529_n N_A_299_47#_M1019_g 0.00132188f $X=1.845 $Y=0.88 $X2=0
+ $Y2=0
cc_459 N_SCE_c_530_n N_A_299_47#_M1019_g 2.97105e-19 $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_460 N_SCE_c_531_n N_A_299_47#_M1019_g 0.0107276f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_461 N_SCE_M1008_g N_A_299_47#_c_645_n 0.0148807f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_462 N_SCE_M1026_g N_A_299_47#_c_645_n 0.00426482f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_463 N_SCE_c_529_n N_A_299_47#_c_645_n 0.0170444f $X=1.845 $Y=0.88 $X2=0 $Y2=0
cc_464 N_SCE_c_530_n N_A_299_47#_c_645_n 0.0572202f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_465 N_SCE_c_541_n N_A_299_47#_c_645_n 0.00366738f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_466 N_SCE_M1026_g N_A_299_47#_c_660_n 0.0123328f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_467 N_SCE_c_530_n N_A_299_47#_c_660_n 0.0104864f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_468 N_SCE_c_541_n N_A_299_47#_c_660_n 0.0039259f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_469 N_SCE_M1008_g N_A_299_47#_c_646_n 0.00145274f $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_470 N_SCE_M1026_g N_A_299_47#_c_646_n 0.00146747f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_471 N_SCE_c_538_n N_A_299_47#_c_646_n 0.00768679f $X=2.175 $Y=1.58 $X2=0
+ $Y2=0
cc_472 N_SCE_M1024_g N_A_299_47#_c_646_n 0.00565974f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_473 N_SCE_c_530_n N_A_299_47#_c_646_n 0.0405813f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_474 N_SCE_c_541_n N_A_299_47#_c_646_n 0.00129443f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_475 N_SCE_M1024_g N_A_299_47#_c_662_n 0.00619128f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_476 N_SCE_c_541_n N_A_299_47#_c_655_n 7.87955e-19 $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_477 N_SCE_M1008_g N_A_299_47#_c_648_n 5.26825e-19 $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_478 N_SCE_c_538_n N_A_299_47#_c_648_n 4.94909e-19 $X=2.175 $Y=1.58 $X2=0
+ $Y2=0
cc_479 N_SCE_c_530_n N_A_299_47#_c_648_n 0.0134242f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_480 N_SCE_c_531_n N_A_299_47#_c_648_n 0.0208599f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_481 N_SCE_c_533_n N_A_299_47#_c_648_n 0.00389077f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_482 N_SCE_M1008_g N_A_299_47#_c_649_n 0.0174183f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_483 N_SCE_c_538_n N_A_299_47#_c_649_n 0.00808785f $X=2.175 $Y=1.58 $X2=0
+ $Y2=0
cc_484 N_SCE_c_530_n N_A_299_47#_c_649_n 0.00156762f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_485 N_SCE_c_531_n N_A_299_47#_c_649_n 0.00319888f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_486 N_SCE_M1024_g N_A_299_47#_c_667_n 0.00630723f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_487 N_SCE_c_533_n N_A_299_47#_c_656_n 0.00959271f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_488 N_SCE_c_534_n N_A_299_47#_c_656_n 3.983e-19 $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_489 N_SCE_c_533_n N_A_299_47#_c_657_n 2.12418e-19 $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_490 N_SCE_c_534_n N_A_299_47#_c_657_n 0.0144723f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_491 N_SCE_M1024_g N_D_M1027_g 0.0391224f $X=2.25 $Y=2.165 $X2=0 $Y2=0
cc_492 N_SCE_M1029_g N_D_M1020_g 0.0137065f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_493 N_SCE_c_532_n N_D_M1020_g 0.0126031f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_494 N_SCE_c_533_n N_D_M1020_g 0.00203037f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_495 N_SCE_c_534_n N_D_M1020_g 0.0213831f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_496 N_SCE_M1008_g N_D_c_773_n 3.44894e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_497 N_SCE_c_538_n N_D_c_773_n 0.0102458f $X=2.175 $Y=1.58 $X2=0 $Y2=0
cc_498 N_SCE_c_541_n N_D_c_773_n 0.00183935f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_499 N_SCE_c_532_n N_D_c_773_n 8.44684e-19 $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_500 N_SCE_c_535_n N_D_c_773_n 0.0011605f $X=2.542 $Y=0.7 $X2=0 $Y2=0
cc_501 N_SCE_c_538_n N_D_c_774_n 0.00125385f $X=2.175 $Y=1.58 $X2=0 $Y2=0
cc_502 N_SCE_c_532_n N_D_c_774_n 0.00197762f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_503 N_SCE_c_535_n N_D_c_774_n 0.00315365f $X=2.542 $Y=0.7 $X2=0 $Y2=0
cc_504 N_SCE_M1029_g N_SCD_M1012_g 0.057299f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_505 N_SCE_c_533_n N_SCD_M1012_g 0.00132819f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_506 N_SCE_c_533_n SCD 0.00292467f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_507 N_SCE_c_534_n SCD 2.12952e-19 $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_508 N_SCE_M1008_g N_A_193_47#_c_873_n 0.0025855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_509 N_SCE_c_538_n N_A_193_47#_c_873_n 0.00157934f $X=2.175 $Y=1.58 $X2=0
+ $Y2=0
cc_510 N_SCE_M1029_g N_A_193_47#_c_873_n 5.27825e-19 $X=3.21 $Y=0.445 $X2=0
+ $Y2=0
cc_511 N_SCE_c_529_n N_A_193_47#_c_873_n 0.0131123f $X=1.845 $Y=0.88 $X2=0 $Y2=0
cc_512 N_SCE_c_530_n N_A_193_47#_c_873_n 0.0107908f $X=1.845 $Y=1.52 $X2=0 $Y2=0
cc_513 N_SCE_c_541_n N_A_193_47#_c_873_n 0.00331116f $X=1.845 $Y=1.52 $X2=0
+ $Y2=0
cc_514 N_SCE_c_531_n N_A_193_47#_c_873_n 0.0130577f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_515 N_SCE_c_532_n N_A_193_47#_c_873_n 0.0205248f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_516 N_SCE_c_533_n N_A_193_47#_c_873_n 0.0105367f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_517 N_SCE_c_534_n N_A_193_47#_c_873_n 0.0037338f $X=3.15 $Y=0.95 $X2=0 $Y2=0
cc_518 N_SCE_c_535_n N_A_193_47#_c_873_n 0.00735012f $X=2.542 $Y=0.7 $X2=0 $Y2=0
cc_519 N_SCE_M1026_g N_A_193_47#_c_881_n 0.00175323f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_520 N_SCE_M1026_g N_VPWR_c_1559_n 0.00910475f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_521 N_SCE_M1024_g N_VPWR_c_1559_n 0.00946067f $X=2.25 $Y=2.165 $X2=0 $Y2=0
cc_522 N_SCE_M1024_g N_VPWR_c_1565_n 0.00340471f $X=2.25 $Y=2.165 $X2=0 $Y2=0
cc_523 N_SCE_M1026_g N_VPWR_c_1572_n 0.00340533f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_524 N_SCE_M1026_g N_VPWR_c_1557_n 0.00515557f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_525 N_SCE_M1024_g N_VPWR_c_1557_n 0.00389325f $X=2.25 $Y=2.165 $X2=0 $Y2=0
cc_526 N_SCE_c_532_n N_A_556_369#_M1020_d 0.00218892f $X=3.065 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_527 N_SCE_M1024_g N_A_556_369#_c_1739_n 5.68908e-19 $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_528 N_SCE_M1029_g N_A_556_369#_c_1751_n 0.00763758f $X=3.21 $Y=0.445 $X2=0
+ $Y2=0
cc_529 N_SCE_c_532_n N_A_556_369#_c_1751_n 0.0207306f $X=3.065 $Y=0.7 $X2=0
+ $Y2=0
cc_530 N_SCE_c_534_n N_A_556_369#_c_1751_n 2.32966e-19 $X=3.15 $Y=0.95 $X2=0
+ $Y2=0
cc_531 N_SCE_M1029_g N_A_556_369#_c_1728_n 0.0041669f $X=3.21 $Y=0.445 $X2=0
+ $Y2=0
cc_532 N_SCE_c_532_n N_A_556_369#_c_1728_n 0.00790081f $X=3.065 $Y=0.7 $X2=0
+ $Y2=0
cc_533 N_SCE_M1029_g N_A_556_369#_c_1730_n 9.50994e-19 $X=3.21 $Y=0.445 $X2=0
+ $Y2=0
cc_534 N_SCE_c_532_n N_A_556_369#_c_1730_n 0.0061514f $X=3.065 $Y=0.7 $X2=0
+ $Y2=0
cc_535 N_SCE_c_533_n N_A_556_369#_c_1730_n 0.00693983f $X=3.15 $Y=0.95 $X2=0
+ $Y2=0
cc_536 N_SCE_c_529_n N_VGND_M1008_d 4.59986e-19 $X=1.845 $Y=0.88 $X2=0 $Y2=0
cc_537 N_SCE_c_531_n N_VGND_M1008_d 0.00200685f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_538 N_SCE_M1008_g N_VGND_c_1910_n 0.00411511f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_539 N_SCE_c_529_n N_VGND_c_1910_n 0.00345278f $X=1.845 $Y=0.88 $X2=0 $Y2=0
cc_540 N_SCE_c_531_n N_VGND_c_1910_n 0.0151465f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_541 N_SCE_M1008_g N_VGND_c_1920_n 0.00438392f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_542 N_SCE_c_529_n N_VGND_c_1920_n 0.00280973f $X=1.845 $Y=0.88 $X2=0 $Y2=0
cc_543 N_SCE_M1029_g N_VGND_c_1921_n 0.00362032f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_544 N_SCE_c_531_n N_VGND_c_1921_n 0.00263191f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_545 N_SCE_c_532_n N_VGND_c_1921_n 0.00274476f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_546 SCE N_VGND_c_1921_n 0.00782706f $X=2.455 $Y=0.425 $X2=0 $Y2=0
cc_547 N_SCE_M1008_g N_VGND_c_1925_n 0.00703621f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_548 N_SCE_M1029_g N_VGND_c_1925_n 0.00526606f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_549 N_SCE_c_529_n N_VGND_c_1925_n 0.00244209f $X=1.845 $Y=0.88 $X2=0 $Y2=0
cc_550 N_SCE_c_531_n N_VGND_c_1925_n 0.00260067f $X=2.455 $Y=0.7 $X2=0 $Y2=0
cc_551 N_SCE_c_532_n N_VGND_c_1925_n 0.00232388f $X=3.065 $Y=0.7 $X2=0 $Y2=0
cc_552 SCE N_VGND_c_1925_n 0.00302552f $X=2.455 $Y=0.425 $X2=0 $Y2=0
cc_553 SCE A_483_47# 0.00226988f $X=2.455 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_554 N_A_299_47#_M1018_g N_D_M1027_g 0.028319f $X=3.125 $Y=2.165 $X2=0 $Y2=0
cc_555 N_A_299_47#_c_646_n N_D_M1027_g 0.00111909f $X=2.185 $Y=1.86 $X2=0 $Y2=0
cc_556 N_A_299_47#_c_662_n N_D_M1027_g 0.0118122f $X=3.06 $Y=1.967 $X2=0 $Y2=0
cc_557 N_A_299_47#_c_654_n N_D_M1027_g 0.00126571f $X=3.145 $Y=1.86 $X2=0 $Y2=0
cc_558 N_A_299_47#_M1019_g N_D_M1020_g 0.0412183f $X=2.34 $Y=0.445 $X2=0 $Y2=0
cc_559 N_A_299_47#_c_646_n N_D_M1020_g 0.00512253f $X=2.185 $Y=1.86 $X2=0 $Y2=0
cc_560 N_A_299_47#_c_648_n N_D_M1020_g 6.95345e-19 $X=2.28 $Y=1.04 $X2=0 $Y2=0
cc_561 N_A_299_47#_c_649_n N_D_M1020_g 0.0168474f $X=2.28 $Y=1.04 $X2=0 $Y2=0
cc_562 N_A_299_47#_c_646_n N_D_c_773_n 6.00877e-19 $X=2.185 $Y=1.86 $X2=0 $Y2=0
cc_563 N_A_299_47#_c_662_n N_D_c_773_n 0.00290918f $X=3.06 $Y=1.967 $X2=0 $Y2=0
cc_564 N_A_299_47#_c_656_n N_D_c_773_n 0.0011165f $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_565 N_A_299_47#_c_657_n N_D_c_773_n 0.0197807f $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_566 N_A_299_47#_c_646_n N_D_c_774_n 0.0254459f $X=2.185 $Y=1.86 $X2=0 $Y2=0
cc_567 N_A_299_47#_c_662_n N_D_c_774_n 0.0199968f $X=3.06 $Y=1.967 $X2=0 $Y2=0
cc_568 N_A_299_47#_c_648_n N_D_c_774_n 2.73452e-19 $X=2.28 $Y=1.04 $X2=0 $Y2=0
cc_569 N_A_299_47#_c_656_n N_D_c_774_n 0.0157256f $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_570 N_A_299_47#_c_657_n N_D_c_774_n 0.00104184f $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_571 N_A_299_47#_M1018_g N_SCD_M1014_g 0.0359024f $X=3.125 $Y=2.165 $X2=0
+ $Y2=0
cc_572 N_A_299_47#_c_662_n N_SCD_M1014_g 2.17192e-19 $X=3.06 $Y=1.967 $X2=0
+ $Y2=0
cc_573 N_A_299_47#_c_654_n N_SCD_M1014_g 0.002483f $X=3.145 $Y=1.86 $X2=0 $Y2=0
cc_574 N_A_299_47#_c_656_n SCD 0.015857f $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_575 N_A_299_47#_c_657_n SCD 0.00104256f $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_576 N_A_299_47#_c_656_n N_SCD_c_822_n 3.53677e-19 $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_577 N_A_299_47#_c_657_n N_SCD_c_822_n 0.0204284f $X=3.17 $Y=1.52 $X2=0 $Y2=0
cc_578 N_A_299_47#_M1019_g N_A_193_47#_c_873_n 0.00170787f $X=2.34 $Y=0.445
+ $X2=0 $Y2=0
cc_579 N_A_299_47#_c_645_n N_A_193_47#_c_873_n 0.0177002f $X=1.505 $Y=1.86 $X2=0
+ $Y2=0
cc_580 N_A_299_47#_c_647_n N_A_193_47#_c_873_n 0.00409336f $X=1.62 $Y=0.42 $X2=0
+ $Y2=0
cc_581 N_A_299_47#_c_648_n N_A_193_47#_c_873_n 0.00873594f $X=2.28 $Y=1.04 $X2=0
+ $Y2=0
cc_582 N_A_299_47#_c_649_n N_A_193_47#_c_873_n 0.00457609f $X=2.28 $Y=1.04 $X2=0
+ $Y2=0
cc_583 N_A_299_47#_c_656_n N_A_193_47#_c_873_n 0.00166362f $X=3.17 $Y=1.52 $X2=0
+ $Y2=0
cc_584 N_A_299_47#_c_657_n N_A_193_47#_c_873_n 6.70678e-19 $X=3.17 $Y=1.52 $X2=0
+ $Y2=0
cc_585 N_A_299_47#_c_645_n N_A_193_47#_c_874_n 0.00265152f $X=1.505 $Y=1.86
+ $X2=0 $Y2=0
cc_586 N_A_299_47#_c_645_n N_A_193_47#_c_881_n 0.0733023f $X=1.505 $Y=1.86 $X2=0
+ $Y2=0
cc_587 N_A_299_47#_c_652_n N_A_193_47#_c_881_n 0.0225669f $X=1.62 $Y=2.175 $X2=0
+ $Y2=0
cc_588 N_A_299_47#_c_647_n N_A_193_47#_c_881_n 0.0146505f $X=1.62 $Y=0.42 $X2=0
+ $Y2=0
cc_589 N_A_299_47#_c_655_n N_A_193_47#_c_881_n 0.0128115f $X=1.562 $Y=1.967
+ $X2=0 $Y2=0
cc_590 N_A_299_47#_c_660_n N_VPWR_M1026_d 0.00374995f $X=2.1 $Y=1.967 $X2=0
+ $Y2=0
cc_591 N_A_299_47#_c_660_n N_VPWR_c_1559_n 0.0117994f $X=2.1 $Y=1.967 $X2=0
+ $Y2=0
cc_592 N_A_299_47#_c_667_n N_VPWR_c_1559_n 0.00348388f $X=2.185 $Y=1.967 $X2=0
+ $Y2=0
cc_593 N_A_299_47#_M1018_g N_VPWR_c_1565_n 0.00368123f $X=3.125 $Y=2.165 $X2=0
+ $Y2=0
cc_594 N_A_299_47#_c_662_n N_VPWR_c_1565_n 0.00602507f $X=3.06 $Y=1.967 $X2=0
+ $Y2=0
cc_595 N_A_299_47#_c_667_n N_VPWR_c_1565_n 0.00112385f $X=2.185 $Y=1.967 $X2=0
+ $Y2=0
cc_596 N_A_299_47#_c_652_n N_VPWR_c_1572_n 0.0174764f $X=1.62 $Y=2.175 $X2=0
+ $Y2=0
cc_597 N_A_299_47#_c_660_n N_VPWR_c_1572_n 0.00240758f $X=2.1 $Y=1.967 $X2=0
+ $Y2=0
cc_598 N_A_299_47#_M1026_s N_VPWR_c_1557_n 0.00184114f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_599 N_A_299_47#_M1018_g N_VPWR_c_1557_n 0.00535446f $X=3.125 $Y=2.165 $X2=0
+ $Y2=0
cc_600 N_A_299_47#_c_652_n N_VPWR_c_1557_n 0.00512382f $X=1.62 $Y=2.175 $X2=0
+ $Y2=0
cc_601 N_A_299_47#_c_660_n N_VPWR_c_1557_n 0.00243889f $X=2.1 $Y=1.967 $X2=0
+ $Y2=0
cc_602 N_A_299_47#_c_662_n N_VPWR_c_1557_n 0.00552167f $X=3.06 $Y=1.967 $X2=0
+ $Y2=0
cc_603 N_A_299_47#_c_667_n N_VPWR_c_1557_n 0.00108805f $X=2.185 $Y=1.967 $X2=0
+ $Y2=0
cc_604 N_A_299_47#_c_662_n A_465_369# 0.005036f $X=3.06 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_605 N_A_299_47#_c_662_n N_A_556_369#_M1027_d 0.00427378f $X=3.06 $Y=1.967
+ $X2=0 $Y2=0
cc_606 N_A_299_47#_M1018_g N_A_556_369#_c_1739_n 0.00811134f $X=3.125 $Y=2.165
+ $X2=0 $Y2=0
cc_607 N_A_299_47#_c_662_n N_A_556_369#_c_1739_n 0.0265702f $X=3.06 $Y=1.967
+ $X2=0 $Y2=0
cc_608 N_A_299_47#_c_657_n N_A_556_369#_c_1739_n 0.0012413f $X=3.17 $Y=1.52
+ $X2=0 $Y2=0
cc_609 N_A_299_47#_M1018_g N_A_556_369#_c_1763_n 0.00367162f $X=3.125 $Y=2.165
+ $X2=0 $Y2=0
cc_610 N_A_299_47#_M1018_g N_A_556_369#_c_1736_n 5.41855e-19 $X=3.125 $Y=2.165
+ $X2=0 $Y2=0
cc_611 N_A_299_47#_c_662_n N_A_556_369#_c_1736_n 0.00683183f $X=3.06 $Y=1.967
+ $X2=0 $Y2=0
cc_612 N_A_299_47#_c_654_n N_A_556_369#_c_1736_n 0.00221463f $X=3.145 $Y=1.86
+ $X2=0 $Y2=0
cc_613 N_A_299_47#_c_647_n N_VGND_c_1909_n 0.00278086f $X=1.62 $Y=0.42 $X2=0
+ $Y2=0
cc_614 N_A_299_47#_M1019_g N_VGND_c_1910_n 0.00745268f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_615 N_A_299_47#_c_647_n N_VGND_c_1920_n 0.0187745f $X=1.62 $Y=0.42 $X2=0
+ $Y2=0
cc_616 N_A_299_47#_M1019_g N_VGND_c_1921_n 0.00365142f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_617 N_A_299_47#_M1008_s N_VGND_c_1925_n 0.00210555f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_618 N_A_299_47#_M1019_g N_VGND_c_1925_n 0.00396023f $X=2.34 $Y=0.445 $X2=0
+ $Y2=0
cc_619 N_A_299_47#_c_647_n N_VGND_c_1925_n 0.00502839f $X=1.62 $Y=0.42 $X2=0
+ $Y2=0
cc_620 N_D_M1020_g N_SCD_M1012_g 0.00367381f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_621 N_D_M1020_g N_A_193_47#_c_873_n 0.00435261f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_622 N_D_c_773_n N_A_193_47#_c_873_n 0.00255857f $X=2.69 $Y=1.52 $X2=0 $Y2=0
cc_623 N_D_c_774_n N_A_193_47#_c_873_n 0.00706402f $X=2.69 $Y=1.52 $X2=0 $Y2=0
cc_624 N_D_M1027_g N_VPWR_c_1559_n 0.0018346f $X=2.705 $Y=2.165 $X2=0 $Y2=0
cc_625 N_D_M1027_g N_VPWR_c_1565_n 0.00385655f $X=2.705 $Y=2.165 $X2=0 $Y2=0
cc_626 N_D_M1027_g N_VPWR_c_1557_n 0.00544811f $X=2.705 $Y=2.165 $X2=0 $Y2=0
cc_627 N_D_M1027_g N_A_556_369#_c_1739_n 0.00614015f $X=2.705 $Y=2.165 $X2=0
+ $Y2=0
cc_628 N_D_M1020_g N_A_556_369#_c_1751_n 0.00166377f $X=2.73 $Y=0.445 $X2=0
+ $Y2=0
cc_629 N_D_M1020_g N_VGND_c_1910_n 0.00138865f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_630 N_D_M1020_g N_VGND_c_1921_n 0.0042011f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_631 N_D_M1020_g N_VGND_c_1925_n 0.00560912f $X=2.73 $Y=0.445 $X2=0 $Y2=0
cc_632 N_SCD_M1012_g N_A_193_47#_c_873_n 0.00204716f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_633 SCD N_A_193_47#_c_873_n 0.0123778f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_634 N_SCD_M1014_g N_VPWR_c_1560_n 0.00615911f $X=3.59 $Y=2.165 $X2=0 $Y2=0
cc_635 N_SCD_M1014_g N_VPWR_c_1565_n 0.00412211f $X=3.59 $Y=2.165 $X2=0 $Y2=0
cc_636 N_SCD_M1014_g N_VPWR_c_1557_n 0.00690372f $X=3.59 $Y=2.165 $X2=0 $Y2=0
cc_637 N_SCD_M1014_g N_A_556_369#_c_1739_n 0.00495708f $X=3.59 $Y=2.165 $X2=0
+ $Y2=0
cc_638 N_SCD_M1012_g N_A_556_369#_c_1751_n 0.00446703f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_639 N_SCD_M1014_g N_A_556_369#_c_1763_n 0.00670328f $X=3.59 $Y=2.165 $X2=0
+ $Y2=0
cc_640 N_SCD_M1012_g N_A_556_369#_c_1728_n 0.00659625f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_641 N_SCD_M1014_g N_A_556_369#_c_1735_n 0.0085544f $X=3.59 $Y=2.165 $X2=0
+ $Y2=0
cc_642 SCD N_A_556_369#_c_1735_n 0.0298783f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_643 N_SCD_c_822_n N_A_556_369#_c_1735_n 5.47858e-19 $X=3.65 $Y=1.355 $X2=0
+ $Y2=0
cc_644 N_SCD_M1014_g N_A_556_369#_c_1736_n 0.00253324f $X=3.59 $Y=2.165 $X2=0
+ $Y2=0
cc_645 SCD N_A_556_369#_c_1736_n 0.00364089f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_646 N_SCD_M1012_g N_A_556_369#_c_1729_n 0.00828793f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_647 SCD N_A_556_369#_c_1729_n 0.0294885f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_648 N_SCD_c_822_n N_A_556_369#_c_1729_n 5.47858e-19 $X=3.65 $Y=1.355 $X2=0
+ $Y2=0
cc_649 N_SCD_M1012_g N_A_556_369#_c_1730_n 0.00228445f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_650 SCD N_A_556_369#_c_1730_n 0.00396416f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_651 N_SCD_M1012_g N_A_556_369#_c_1731_n 0.00230408f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_652 N_SCD_M1012_g N_A_556_369#_c_1732_n 0.00428501f $X=3.59 $Y=0.445 $X2=0
+ $Y2=0
cc_653 N_SCD_M1014_g N_A_556_369#_c_1732_n 0.00437572f $X=3.59 $Y=2.165 $X2=0
+ $Y2=0
cc_654 SCD N_A_556_369#_c_1732_n 0.0490827f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_655 N_SCD_c_822_n N_A_556_369#_c_1732_n 0.00106245f $X=3.65 $Y=1.355 $X2=0
+ $Y2=0
cc_656 N_SCD_M1014_g N_A_556_369#_c_1738_n 0.00288252f $X=3.59 $Y=2.165 $X2=0
+ $Y2=0
cc_657 N_SCD_M1012_g N_VGND_c_1911_n 0.00568381f $X=3.59 $Y=0.445 $X2=0 $Y2=0
cc_658 N_SCD_M1012_g N_VGND_c_1921_n 0.00406622f $X=3.59 $Y=0.445 $X2=0 $Y2=0
cc_659 N_SCD_M1012_g N_VGND_c_1925_n 0.00667021f $X=3.59 $Y=0.445 $X2=0 $Y2=0
cc_660 N_A_193_47#_c_872_n N_A_1089_183#_M1013_d 0.00133652f $X=6.925 $Y=0.87
+ $X2=-0.19 $Y2=-0.24
cc_661 N_A_193_47#_c_875_n N_A_1089_183#_M1013_d 9.65449e-19 $X=6.525 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_662 N_A_193_47#_c_877_n N_A_1089_183#_M1013_d 6.4695e-19 $X=6.67 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_663 N_A_193_47#_c_875_n N_A_1089_183#_M1009_g 0.00208483f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_664 N_A_193_47#_c_879_n N_A_1089_183#_M1009_g 0.013781f $X=5 $Y=0.705 $X2=0
+ $Y2=0
cc_665 N_A_193_47#_c_875_n N_A_1089_183#_c_1083_n 0.0221014f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_666 N_A_193_47#_c_877_n N_A_1089_183#_c_1109_n 8.93965e-19 $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_667 N_A_193_47#_c_872_n N_A_1089_183#_c_1110_n 0.00716698f $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_668 N_A_193_47#_c_875_n N_A_1089_183#_c_1110_n 0.00363224f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_669 N_A_193_47#_c_877_n N_A_1089_183#_c_1110_n 0.00168986f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_670 N_A_193_47#_c_875_n N_A_1089_183#_c_1084_n 0.00899288f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_671 N_A_193_47#_c_871_n N_A_1089_183#_c_1085_n 0.00114045f $X=7.02 $Y=1.575
+ $X2=0 $Y2=0
cc_672 N_A_193_47#_c_872_n N_A_1089_183#_c_1085_n 0.018732f $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_673 N_A_193_47#_c_875_n N_A_1089_183#_c_1085_n 0.0176435f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_674 N_A_193_47#_c_877_n N_A_1089_183#_c_1085_n 0.00185392f $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_675 N_A_193_47#_c_880_n N_A_1089_183#_c_1085_n 5.82389e-19 $X=6.88 $Y=0.87
+ $X2=0 $Y2=0
cc_676 N_A_193_47#_c_871_n N_A_1089_183#_c_1086_n 0.00620052f $X=7.02 $Y=1.575
+ $X2=0 $Y2=0
cc_677 N_A_193_47#_c_875_n N_A_1089_183#_c_1087_n 0.00299829f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_678 N_A_193_47#_c_878_n N_A_1089_183#_c_1087_n 0.0179412f $X=5 $Y=0.87 $X2=0
+ $Y2=0
cc_679 N_A_193_47#_c_871_n N_A_930_413#_c_1176_n 6.31337e-19 $X=7.02 $Y=1.575
+ $X2=0 $Y2=0
cc_680 N_A_193_47#_c_869_n N_A_930_413#_c_1177_n 0.00957285f $X=6.785 $Y=0.705
+ $X2=0 $Y2=0
cc_681 N_A_193_47#_c_872_n N_A_930_413#_c_1177_n 0.00100831f $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_682 N_A_193_47#_c_871_n N_A_930_413#_c_1178_n 3.37852e-19 $X=7.02 $Y=1.575
+ $X2=0 $Y2=0
cc_683 N_A_193_47#_c_880_n N_A_930_413#_c_1178_n 0.00957285f $X=6.88 $Y=0.87
+ $X2=0 $Y2=0
cc_684 N_A_193_47#_M1003_g N_A_930_413#_c_1194_n 0.00166902f $X=4.575 $Y=2.275
+ $X2=0 $Y2=0
cc_685 N_A_193_47#_c_870_n N_A_930_413#_c_1194_n 0.00286257f $X=4.59 $Y=1.74
+ $X2=0 $Y2=0
cc_686 N_A_193_47#_c_885_n N_A_930_413#_c_1194_n 6.94615e-19 $X=4.59 $Y=1.74
+ $X2=0 $Y2=0
cc_687 N_A_193_47#_c_875_n N_A_930_413#_c_1220_n 0.00489874f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_688 N_A_193_47#_c_1005_p N_A_930_413#_c_1220_n 0.00119052f $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_689 N_A_193_47#_c_876_n N_A_930_413#_c_1220_n 0.0237558f $X=4.83 $Y=0.85
+ $X2=0 $Y2=0
cc_690 N_A_193_47#_c_878_n N_A_930_413#_c_1220_n 0.00256542f $X=5 $Y=0.87 $X2=0
+ $Y2=0
cc_691 N_A_193_47#_c_879_n N_A_930_413#_c_1220_n 0.00840911f $X=5 $Y=0.705 $X2=0
+ $Y2=0
cc_692 N_A_193_47#_c_870_n N_A_930_413#_c_1181_n 0.00981359f $X=4.59 $Y=1.74
+ $X2=0 $Y2=0
cc_693 N_A_193_47#_c_875_n N_A_930_413#_c_1181_n 0.0188221f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_694 N_A_193_47#_c_1005_p N_A_930_413#_c_1181_n 5.13248e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_695 N_A_193_47#_c_876_n N_A_930_413#_c_1181_n 0.0239322f $X=4.83 $Y=0.85
+ $X2=0 $Y2=0
cc_696 N_A_193_47#_c_879_n N_A_930_413#_c_1181_n 0.00604394f $X=5 $Y=0.705 $X2=0
+ $Y2=0
cc_697 N_A_193_47#_c_870_n N_A_930_413#_c_1182_n 0.00649323f $X=4.59 $Y=1.74
+ $X2=0 $Y2=0
cc_698 N_A_193_47#_c_875_n N_A_930_413#_c_1182_n 0.00803733f $X=6.525 $Y=0.85
+ $X2=0 $Y2=0
cc_699 N_A_193_47#_M1035_g N_A_1517_315#_c_1303_n 0.018025f $X=7.075 $Y=2.275
+ $X2=0 $Y2=0
cc_700 N_A_193_47#_c_888_n N_A_1517_315#_c_1303_n 0.0119764f $X=7.16 $Y=1.74
+ $X2=0 $Y2=0
cc_701 N_A_193_47#_M1035_g N_A_1346_413#_c_1421_n 0.00974744f $X=7.075 $Y=2.275
+ $X2=0 $Y2=0
cc_702 N_A_193_47#_c_887_n N_A_1346_413#_c_1421_n 0.012999f $X=7.16 $Y=1.74
+ $X2=0 $Y2=0
cc_703 N_A_193_47#_c_888_n N_A_1346_413#_c_1421_n 0.00300896f $X=7.16 $Y=1.74
+ $X2=0 $Y2=0
cc_704 N_A_193_47#_c_872_n N_A_1346_413#_c_1424_n 0.0153172f $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_705 N_A_193_47#_c_880_n N_A_1346_413#_c_1424_n 8.54271e-19 $X=6.88 $Y=0.87
+ $X2=0 $Y2=0
cc_706 N_A_193_47#_M1035_g N_A_1346_413#_c_1418_n 0.0046302f $X=7.075 $Y=2.275
+ $X2=0 $Y2=0
cc_707 N_A_193_47#_c_871_n N_A_1346_413#_c_1418_n 0.00868218f $X=7.02 $Y=1.575
+ $X2=0 $Y2=0
cc_708 N_A_193_47#_c_887_n N_A_1346_413#_c_1418_n 0.0246912f $X=7.16 $Y=1.74
+ $X2=0 $Y2=0
cc_709 N_A_193_47#_c_888_n N_A_1346_413#_c_1418_n 0.00187857f $X=7.16 $Y=1.74
+ $X2=0 $Y2=0
cc_710 N_A_193_47#_c_871_n N_A_1346_413#_c_1413_n 0.0272384f $X=7.02 $Y=1.575
+ $X2=0 $Y2=0
cc_711 N_A_193_47#_c_888_n N_A_1346_413#_c_1413_n 0.00102186f $X=7.16 $Y=1.74
+ $X2=0 $Y2=0
cc_712 N_A_193_47#_c_869_n N_A_1346_413#_c_1414_n 8.96907e-19 $X=6.785 $Y=0.705
+ $X2=0 $Y2=0
cc_713 N_A_193_47#_c_872_n N_A_1346_413#_c_1414_n 0.025625f $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_714 N_A_193_47#_c_877_n N_A_1346_413#_c_1414_n 8.16973e-19 $X=6.67 $Y=0.85
+ $X2=0 $Y2=0
cc_715 N_A_193_47#_c_880_n N_A_1346_413#_c_1414_n 3.08898e-19 $X=6.88 $Y=0.87
+ $X2=0 $Y2=0
cc_716 N_A_193_47#_c_881_n N_VPWR_c_1558_n 0.012721f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_717 N_A_193_47#_M1003_g N_VPWR_c_1560_n 0.00271302f $X=4.575 $Y=2.275 $X2=0
+ $Y2=0
cc_718 N_A_193_47#_M1003_g N_VPWR_c_1567_n 0.005785f $X=4.575 $Y=2.275 $X2=0
+ $Y2=0
cc_719 N_A_193_47#_M1035_g N_VPWR_c_1569_n 0.00383564f $X=7.075 $Y=2.275 $X2=0
+ $Y2=0
cc_720 N_A_193_47#_c_881_n N_VPWR_c_1572_n 0.0120448f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_721 N_A_193_47#_M1003_g N_VPWR_c_1557_n 0.00734982f $X=4.575 $Y=2.275 $X2=0
+ $Y2=0
cc_722 N_A_193_47#_M1035_g N_VPWR_c_1557_n 0.00579176f $X=7.075 $Y=2.275 $X2=0
+ $Y2=0
cc_723 N_A_193_47#_c_870_n N_VPWR_c_1557_n 0.00189161f $X=4.59 $Y=1.74 $X2=0
+ $Y2=0
cc_724 N_A_193_47#_c_885_n N_VPWR_c_1557_n 2.76897e-19 $X=4.59 $Y=1.74 $X2=0
+ $Y2=0
cc_725 N_A_193_47#_c_881_n N_VPWR_c_1557_n 0.00308197f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_726 N_A_193_47#_c_873_n N_A_556_369#_c_1751_n 0.00537221f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_727 N_A_193_47#_c_873_n N_A_556_369#_c_1729_n 0.0211891f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_728 N_A_193_47#_c_873_n N_A_556_369#_c_1730_n 0.0100881f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_729 N_A_193_47#_c_876_n N_A_556_369#_c_1731_n 6.72385e-19 $X=4.83 $Y=0.85
+ $X2=0 $Y2=0
cc_730 N_A_193_47#_c_870_n N_A_556_369#_c_1732_n 0.058581f $X=4.59 $Y=1.74 $X2=0
+ $Y2=0
cc_731 N_A_193_47#_c_885_n N_A_556_369#_c_1732_n 0.0052844f $X=4.59 $Y=1.74
+ $X2=0 $Y2=0
cc_732 N_A_193_47#_c_873_n N_A_556_369#_c_1732_n 0.011116f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_733 N_A_193_47#_c_1005_p N_A_556_369#_c_1732_n 2.21941e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_734 N_A_193_47#_c_876_n N_A_556_369#_c_1732_n 0.0111587f $X=4.83 $Y=0.85
+ $X2=0 $Y2=0
cc_735 N_A_193_47#_c_873_n N_A_556_369#_c_1733_n 0.00506513f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_736 N_A_193_47#_c_876_n N_A_556_369#_c_1733_n 6.01474e-19 $X=4.83 $Y=0.85
+ $X2=0 $Y2=0
cc_737 N_A_193_47#_c_873_n N_A_556_369#_c_1734_n 0.00620857f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_738 N_A_193_47#_c_1005_p N_A_556_369#_c_1734_n 2.5118e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_739 N_A_193_47#_c_876_n N_A_556_369#_c_1734_n 0.0128887f $X=4.83 $Y=0.85
+ $X2=0 $Y2=0
cc_740 N_A_193_47#_M1003_g N_A_556_369#_c_1738_n 0.00502759f $X=4.575 $Y=2.275
+ $X2=0 $Y2=0
cc_741 N_A_193_47#_c_870_n N_A_556_369#_c_1738_n 0.00558861f $X=4.59 $Y=1.74
+ $X2=0 $Y2=0
cc_742 N_A_193_47#_c_885_n N_A_556_369#_c_1738_n 0.00169363f $X=4.59 $Y=1.74
+ $X2=0 $Y2=0
cc_743 N_A_193_47#_c_873_n N_VGND_c_1910_n 0.00117884f $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_744 N_A_193_47#_c_873_n N_VGND_c_1911_n 9.19202e-19 $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_745 N_A_193_47#_c_876_n N_VGND_c_1912_n 0.00254426f $X=4.83 $Y=0.85 $X2=0
+ $Y2=0
cc_746 N_A_193_47#_c_879_n N_VGND_c_1912_n 0.0037981f $X=5 $Y=0.705 $X2=0 $Y2=0
cc_747 N_A_193_47#_c_875_n N_VGND_c_1913_n 0.00197288f $X=6.525 $Y=0.85 $X2=0
+ $Y2=0
cc_748 N_A_193_47#_c_869_n N_VGND_c_1917_n 0.00435108f $X=6.785 $Y=0.705 $X2=0
+ $Y2=0
cc_749 N_A_193_47#_c_872_n N_VGND_c_1917_n 0.00341023f $X=6.925 $Y=0.87 $X2=0
+ $Y2=0
cc_750 N_A_193_47#_c_880_n N_VGND_c_1917_n 8.04624e-19 $X=6.88 $Y=0.87 $X2=0
+ $Y2=0
cc_751 N_A_193_47#_c_881_n N_VGND_c_1920_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_752 N_A_193_47#_M1021_d N_VGND_c_1925_n 0.00238313f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_753 N_A_193_47#_c_869_n N_VGND_c_1925_n 0.00623562f $X=6.785 $Y=0.705 $X2=0
+ $Y2=0
cc_754 N_A_193_47#_c_872_n N_VGND_c_1925_n 0.00402561f $X=6.925 $Y=0.87 $X2=0
+ $Y2=0
cc_755 N_A_193_47#_c_873_n N_VGND_c_1925_n 0.158662f $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_756 N_A_193_47#_c_874_n N_VGND_c_1925_n 0.0154435f $X=1.245 $Y=0.85 $X2=0
+ $Y2=0
cc_757 N_A_193_47#_c_875_n N_VGND_c_1925_n 0.0711725f $X=6.525 $Y=0.85 $X2=0
+ $Y2=0
cc_758 N_A_193_47#_c_1005_p N_VGND_c_1925_n 0.0146104f $X=4.975 $Y=0.85 $X2=0
+ $Y2=0
cc_759 N_A_193_47#_c_876_n N_VGND_c_1925_n 0.00248905f $X=4.83 $Y=0.85 $X2=0
+ $Y2=0
cc_760 N_A_193_47#_c_877_n N_VGND_c_1925_n 0.0147739f $X=6.67 $Y=0.85 $X2=0
+ $Y2=0
cc_761 N_A_193_47#_c_879_n N_VGND_c_1925_n 0.00563926f $X=5 $Y=0.705 $X2=0 $Y2=0
cc_762 N_A_193_47#_c_880_n N_VGND_c_1925_n 0.00134095f $X=6.88 $Y=0.87 $X2=0
+ $Y2=0
cc_763 N_A_193_47#_c_881_n N_VGND_c_1925_n 0.00280714f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_764 N_A_1089_183#_c_1086_n N_A_930_413#_c_1176_n 0.00595764f $X=6.35 $Y=2.135
+ $X2=0 $Y2=0
cc_765 N_A_1089_183#_M1005_g N_A_930_413#_M1025_g 0.0139082f $X=5.52 $Y=2.275
+ $X2=0 $Y2=0
cc_766 N_A_1089_183#_c_1097_n N_A_930_413#_M1025_g 0.00378805f $X=6.39 $Y=2.3
+ $X2=0 $Y2=0
cc_767 N_A_1089_183#_c_1086_n N_A_930_413#_M1025_g 0.0122998f $X=6.35 $Y=2.135
+ $X2=0 $Y2=0
cc_768 N_A_1089_183#_M1009_g N_A_930_413#_c_1177_n 0.0109128f $X=5.55 $Y=0.445
+ $X2=0 $Y2=0
cc_769 N_A_1089_183#_c_1083_n N_A_930_413#_c_1177_n 0.00351053f $X=6.225
+ $Y=0.915 $X2=0 $Y2=0
cc_770 N_A_1089_183#_c_1109_n N_A_930_413#_c_1177_n 0.00675936f $X=6.31 $Y=0.765
+ $X2=0 $Y2=0
cc_771 N_A_1089_183#_c_1129_p N_A_930_413#_c_1177_n 0.004701f $X=6.395 $Y=0.45
+ $X2=0 $Y2=0
cc_772 N_A_1089_183#_c_1085_n N_A_930_413#_c_1177_n 0.00333126f $X=6.31 $Y=0.915
+ $X2=0 $Y2=0
cc_773 N_A_1089_183#_c_1087_n N_A_930_413#_c_1177_n 0.00500517f $X=5.55 $Y=0.93
+ $X2=0 $Y2=0
cc_774 N_A_1089_183#_M1005_g N_A_930_413#_c_1178_n 0.00398999f $X=5.52 $Y=2.275
+ $X2=0 $Y2=0
cc_775 N_A_1089_183#_c_1083_n N_A_930_413#_c_1178_n 0.00996228f $X=6.225
+ $Y=0.915 $X2=0 $Y2=0
cc_776 N_A_1089_183#_c_1084_n N_A_930_413#_c_1178_n 2.46578e-19 $X=5.765 $Y=0.93
+ $X2=0 $Y2=0
cc_777 N_A_1089_183#_c_1085_n N_A_930_413#_c_1178_n 0.00234347f $X=6.31 $Y=0.915
+ $X2=0 $Y2=0
cc_778 N_A_1089_183#_c_1086_n N_A_930_413#_c_1178_n 0.00394884f $X=6.35 $Y=2.135
+ $X2=0 $Y2=0
cc_779 N_A_1089_183#_c_1087_n N_A_930_413#_c_1178_n 0.00573363f $X=5.55 $Y=0.93
+ $X2=0 $Y2=0
cc_780 N_A_1089_183#_M1005_g N_A_930_413#_c_1179_n 0.0173592f $X=5.52 $Y=2.275
+ $X2=0 $Y2=0
cc_781 N_A_1089_183#_c_1083_n N_A_930_413#_c_1179_n 0.00400764f $X=6.225
+ $Y=0.915 $X2=0 $Y2=0
cc_782 N_A_1089_183#_c_1087_n N_A_930_413#_c_1179_n 0.00238133f $X=5.55 $Y=0.93
+ $X2=0 $Y2=0
cc_783 N_A_1089_183#_c_1086_n N_A_930_413#_c_1180_n 0.00611615f $X=6.35 $Y=2.135
+ $X2=0 $Y2=0
cc_784 N_A_1089_183#_M1005_g N_A_930_413#_c_1194_n 0.0101048f $X=5.52 $Y=2.275
+ $X2=0 $Y2=0
cc_785 N_A_1089_183#_M1009_g N_A_930_413#_c_1181_n 0.00441151f $X=5.55 $Y=0.445
+ $X2=0 $Y2=0
cc_786 N_A_1089_183#_c_1084_n N_A_930_413#_c_1181_n 0.0242417f $X=5.765 $Y=0.93
+ $X2=0 $Y2=0
cc_787 N_A_1089_183#_c_1087_n N_A_930_413#_c_1181_n 0.0095167f $X=5.55 $Y=0.93
+ $X2=0 $Y2=0
cc_788 N_A_1089_183#_M1005_g N_A_930_413#_c_1186_n 0.0153783f $X=5.52 $Y=2.275
+ $X2=0 $Y2=0
cc_789 N_A_1089_183#_c_1086_n N_A_930_413#_c_1186_n 0.00754007f $X=6.35 $Y=2.135
+ $X2=0 $Y2=0
cc_790 N_A_1089_183#_M1005_g N_A_930_413#_c_1182_n 0.0138593f $X=5.52 $Y=2.275
+ $X2=0 $Y2=0
cc_791 N_A_1089_183#_c_1083_n N_A_930_413#_c_1182_n 0.0186614f $X=6.225 $Y=0.915
+ $X2=0 $Y2=0
cc_792 N_A_1089_183#_c_1084_n N_A_930_413#_c_1182_n 0.0112018f $X=5.765 $Y=0.93
+ $X2=0 $Y2=0
cc_793 N_A_1089_183#_c_1086_n N_A_930_413#_c_1182_n 0.0245884f $X=6.35 $Y=2.135
+ $X2=0 $Y2=0
cc_794 N_A_1089_183#_c_1087_n N_A_930_413#_c_1182_n 0.00213749f $X=5.55 $Y=0.93
+ $X2=0 $Y2=0
cc_795 N_A_1089_183#_c_1097_n N_A_1346_413#_c_1421_n 0.0109209f $X=6.39 $Y=2.3
+ $X2=0 $Y2=0
cc_796 N_A_1089_183#_M1005_g N_VPWR_c_1561_n 0.0057281f $X=5.52 $Y=2.275 $X2=0
+ $Y2=0
cc_797 N_A_1089_183#_c_1086_n N_VPWR_c_1561_n 0.0237f $X=6.35 $Y=2.135 $X2=0
+ $Y2=0
cc_798 N_A_1089_183#_M1005_g N_VPWR_c_1567_n 0.00378797f $X=5.52 $Y=2.275 $X2=0
+ $Y2=0
cc_799 N_A_1089_183#_c_1097_n N_VPWR_c_1569_n 0.015079f $X=6.39 $Y=2.3 $X2=0
+ $Y2=0
cc_800 N_A_1089_183#_M1025_d N_VPWR_c_1557_n 0.00285154f $X=6.255 $Y=1.735 $X2=0
+ $Y2=0
cc_801 N_A_1089_183#_M1005_g N_VPWR_c_1557_n 0.00596544f $X=5.52 $Y=2.275 $X2=0
+ $Y2=0
cc_802 N_A_1089_183#_c_1097_n N_VPWR_c_1557_n 0.00439826f $X=6.39 $Y=2.3 $X2=0
+ $Y2=0
cc_803 N_A_1089_183#_c_1083_n N_VGND_M1009_d 0.00306998f $X=6.225 $Y=0.915 $X2=0
+ $Y2=0
cc_804 N_A_1089_183#_M1009_g N_VGND_c_1912_n 0.00585385f $X=5.55 $Y=0.445 $X2=0
+ $Y2=0
cc_805 N_A_1089_183#_M1009_g N_VGND_c_1913_n 0.00603751f $X=5.55 $Y=0.445 $X2=0
+ $Y2=0
cc_806 N_A_1089_183#_c_1109_n N_VGND_c_1913_n 0.00354103f $X=6.31 $Y=0.765 $X2=0
+ $Y2=0
cc_807 N_A_1089_183#_c_1129_p N_VGND_c_1913_n 0.013122f $X=6.395 $Y=0.45 $X2=0
+ $Y2=0
cc_808 N_A_1089_183#_c_1084_n N_VGND_c_1913_n 0.0258565f $X=5.765 $Y=0.93 $X2=0
+ $Y2=0
cc_809 N_A_1089_183#_c_1087_n N_VGND_c_1913_n 0.00122075f $X=5.55 $Y=0.93 $X2=0
+ $Y2=0
cc_810 N_A_1089_183#_c_1129_p N_VGND_c_1917_n 0.00594819f $X=6.395 $Y=0.45 $X2=0
+ $Y2=0
cc_811 N_A_1089_183#_c_1110_n N_VGND_c_1917_n 0.0100275f $X=6.52 $Y=0.45 $X2=0
+ $Y2=0
cc_812 N_A_1089_183#_M1013_d N_VGND_c_1925_n 0.00246577f $X=6.355 $Y=0.235 $X2=0
+ $Y2=0
cc_813 N_A_1089_183#_M1009_g N_VGND_c_1925_n 0.0070154f $X=5.55 $Y=0.445 $X2=0
+ $Y2=0
cc_814 N_A_1089_183#_c_1083_n N_VGND_c_1925_n 0.0042145f $X=6.225 $Y=0.915 $X2=0
+ $Y2=0
cc_815 N_A_1089_183#_c_1129_p N_VGND_c_1925_n 0.00261981f $X=6.395 $Y=0.45 $X2=0
+ $Y2=0
cc_816 N_A_1089_183#_c_1110_n N_VGND_c_1925_n 0.00441842f $X=6.52 $Y=0.45 $X2=0
+ $Y2=0
cc_817 N_A_1089_183#_c_1084_n N_VGND_c_1925_n 0.00269026f $X=5.765 $Y=0.93 $X2=0
+ $Y2=0
cc_818 N_A_930_413#_c_1194_n N_VPWR_M1005_d 0.00236303f $X=5.545 $Y=2.275 $X2=0
+ $Y2=0
cc_819 N_A_930_413#_c_1186_n N_VPWR_M1005_d 0.00412006f $X=5.63 $Y=2.19 $X2=0
+ $Y2=0
cc_820 N_A_930_413#_M1025_g N_VPWR_c_1561_n 0.00314007f $X=6.18 $Y=2.11 $X2=0
+ $Y2=0
cc_821 N_A_930_413#_c_1179_n N_VPWR_c_1561_n 9.53331e-19 $X=6.105 $Y=1.41 $X2=0
+ $Y2=0
cc_822 N_A_930_413#_c_1194_n N_VPWR_c_1561_n 0.0138309f $X=5.545 $Y=2.275 $X2=0
+ $Y2=0
cc_823 N_A_930_413#_c_1186_n N_VPWR_c_1561_n 0.0252361f $X=5.63 $Y=2.19 $X2=0
+ $Y2=0
cc_824 N_A_930_413#_c_1182_n N_VPWR_c_1561_n 0.00741701f $X=5.63 $Y=1.41 $X2=0
+ $Y2=0
cc_825 N_A_930_413#_c_1194_n N_VPWR_c_1567_n 0.0359536f $X=5.545 $Y=2.275 $X2=0
+ $Y2=0
cc_826 N_A_930_413#_M1025_g N_VPWR_c_1569_n 0.00541359f $X=6.18 $Y=2.11 $X2=0
+ $Y2=0
cc_827 N_A_930_413#_M1003_d N_VPWR_c_1557_n 0.00217001f $X=4.65 $Y=2.065 $X2=0
+ $Y2=0
cc_828 N_A_930_413#_M1025_g N_VPWR_c_1557_n 0.00665748f $X=6.18 $Y=2.11 $X2=0
+ $Y2=0
cc_829 N_A_930_413#_c_1194_n N_VPWR_c_1557_n 0.0161661f $X=5.545 $Y=2.275 $X2=0
+ $Y2=0
cc_830 N_A_930_413#_c_1194_n A_1023_413# 0.0045944f $X=5.545 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_831 N_A_930_413#_c_1220_n N_VGND_c_1912_n 0.0255873f $X=5.255 $Y=0.45 $X2=0
+ $Y2=0
cc_832 N_A_930_413#_c_1177_n N_VGND_c_1913_n 0.00816054f $X=6.28 $Y=0.95 $X2=0
+ $Y2=0
cc_833 N_A_930_413#_c_1177_n N_VGND_c_1917_n 0.00407056f $X=6.28 $Y=0.95 $X2=0
+ $Y2=0
cc_834 N_A_930_413#_M1031_d N_VGND_c_1925_n 0.00228204f $X=4.655 $Y=0.235 $X2=0
+ $Y2=0
cc_835 N_A_930_413#_c_1177_n N_VGND_c_1925_n 0.00620172f $X=6.28 $Y=0.95 $X2=0
+ $Y2=0
cc_836 N_A_930_413#_c_1220_n N_VGND_c_1925_n 0.0112934f $X=5.255 $Y=0.45 $X2=0
+ $Y2=0
cc_837 N_A_930_413#_c_1220_n A_1027_47# 0.00455507f $X=5.255 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_838 N_A_930_413#_c_1181_n A_1027_47# 0.00200718f $X=5.34 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_839 N_A_1517_315#_c_1285_n N_A_1346_413#_c_1409_n 0.0222022f $X=9.135
+ $Y=0.995 $X2=0 $Y2=0
cc_840 N_A_1517_315#_c_1289_n N_A_1346_413#_c_1409_n 0.00404044f $X=8.505
+ $Y=0.385 $X2=0 $Y2=0
cc_841 N_A_1517_315#_c_1290_n N_A_1346_413#_c_1409_n 0.00482817f $X=8.577
+ $Y=0.995 $X2=0 $Y2=0
cc_842 N_A_1517_315#_c_1293_n N_A_1346_413#_c_1409_n 0.0026257f $X=8.505
+ $Y=0.825 $X2=0 $Y2=0
cc_843 N_A_1517_315#_M1028_g N_A_1346_413#_M1001_g 0.0225853f $X=9.135 $Y=1.985
+ $X2=0 $Y2=0
cc_844 N_A_1517_315#_c_1303_n N_A_1346_413#_M1001_g 0.00279976f $X=7.84 $Y=1.74
+ $X2=0 $Y2=0
cc_845 N_A_1517_315#_c_1316_p N_A_1346_413#_M1001_g 0.00597831f $X=8.505 $Y=1.95
+ $X2=0 $Y2=0
cc_846 N_A_1517_315#_c_1304_n N_A_1346_413#_M1001_g 0.00869923f $X=8.577
+ $Y=1.575 $X2=0 $Y2=0
cc_847 N_A_1517_315#_c_1318_p N_A_1346_413#_M1001_g 0.00748031f $X=8.525 $Y=1.74
+ $X2=0 $Y2=0
cc_848 N_A_1517_315#_M1016_g N_A_1346_413#_c_1410_n 0.0177134f $X=7.775 $Y=0.445
+ $X2=0 $Y2=0
cc_849 N_A_1517_315#_c_1302_n N_A_1346_413#_c_1410_n 0.00716149f $X=8.38 $Y=1.74
+ $X2=0 $Y2=0
cc_850 N_A_1517_315#_c_1293_n N_A_1346_413#_c_1410_n 0.00615736f $X=8.505
+ $Y=0.825 $X2=0 $Y2=0
cc_851 N_A_1517_315#_c_1318_p N_A_1346_413#_c_1410_n 0.00428237f $X=8.525
+ $Y=1.74 $X2=0 $Y2=0
cc_852 N_A_1517_315#_c_1323_p N_A_1346_413#_c_1410_n 0.0168182f $X=8.577 $Y=1.16
+ $X2=0 $Y2=0
cc_853 N_A_1517_315#_c_1291_n N_A_1346_413#_c_1411_n 0.0180498f $X=9.135 $Y=1.16
+ $X2=0 $Y2=0
cc_854 N_A_1517_315#_c_1292_n N_A_1346_413#_c_1411_n 0.0216171f $X=9.135 $Y=1.16
+ $X2=0 $Y2=0
cc_855 N_A_1517_315#_c_1323_p N_A_1346_413#_c_1411_n 9.32228e-19 $X=8.577
+ $Y=1.16 $X2=0 $Y2=0
cc_856 N_A_1517_315#_M1015_g N_A_1346_413#_c_1421_n 0.00194535f $X=7.66 $Y=2.275
+ $X2=0 $Y2=0
cc_857 N_A_1517_315#_M1016_g N_A_1346_413#_c_1424_n 0.00114979f $X=7.775
+ $Y=0.445 $X2=0 $Y2=0
cc_858 N_A_1517_315#_c_1302_n N_A_1346_413#_c_1418_n 0.0262086f $X=8.38 $Y=1.74
+ $X2=0 $Y2=0
cc_859 N_A_1517_315#_c_1303_n N_A_1346_413#_c_1418_n 0.00865902f $X=7.84 $Y=1.74
+ $X2=0 $Y2=0
cc_860 N_A_1517_315#_M1016_g N_A_1346_413#_c_1412_n 0.017942f $X=7.775 $Y=0.445
+ $X2=0 $Y2=0
cc_861 N_A_1517_315#_c_1302_n N_A_1346_413#_c_1412_n 0.033362f $X=8.38 $Y=1.74
+ $X2=0 $Y2=0
cc_862 N_A_1517_315#_c_1303_n N_A_1346_413#_c_1412_n 0.00739167f $X=7.84 $Y=1.74
+ $X2=0 $Y2=0
cc_863 N_A_1517_315#_c_1323_p N_A_1346_413#_c_1412_n 0.0277655f $X=8.577 $Y=1.16
+ $X2=0 $Y2=0
cc_864 N_A_1517_315#_M1016_g N_A_1346_413#_c_1413_n 0.00880678f $X=7.775
+ $Y=0.445 $X2=0 $Y2=0
cc_865 N_A_1517_315#_M1016_g N_A_1346_413#_c_1414_n 0.00779225f $X=7.775
+ $Y=0.445 $X2=0 $Y2=0
cc_866 N_A_1517_315#_c_1300_n N_A_1948_47#_M1007_g 0.00474627f $X=10.047
+ $Y=1.515 $X2=0 $Y2=0
cc_867 N_A_1517_315#_c_1301_n N_A_1948_47#_M1007_g 0.0181632f $X=10.047 $Y=1.665
+ $X2=0 $Y2=0
cc_868 N_A_1517_315#_M1028_g N_A_1948_47#_c_1503_n 0.00161237f $X=9.135 $Y=1.985
+ $X2=0 $Y2=0
cc_869 N_A_1517_315#_c_1286_n N_A_1948_47#_c_1503_n 0.00286889f $X=9.945 $Y=1.16
+ $X2=0 $Y2=0
cc_870 N_A_1517_315#_M1030_g N_A_1948_47#_c_1503_n 0.00498986f $X=10.075
+ $Y=2.165 $X2=0 $Y2=0
cc_871 N_A_1517_315#_M1030_g N_A_1948_47#_c_1504_n 0.00647251f $X=10.075
+ $Y=2.165 $X2=0 $Y2=0
cc_872 N_A_1517_315#_c_1287_n N_A_1948_47#_c_1497_n 0.00880948f $X=10.02
+ $Y=1.325 $X2=0 $Y2=0
cc_873 N_A_1517_315#_c_1288_n N_A_1948_47#_c_1497_n 0.00170371f $X=10.075
+ $Y=0.73 $X2=0 $Y2=0
cc_874 N_A_1517_315#_c_1287_n N_A_1948_47#_c_1498_n 0.0133342f $X=10.02 $Y=1.325
+ $X2=0 $Y2=0
cc_875 N_A_1517_315#_c_1301_n N_A_1948_47#_c_1498_n 0.00159098f $X=10.047
+ $Y=1.665 $X2=0 $Y2=0
cc_876 N_A_1517_315#_c_1287_n N_A_1948_47#_c_1499_n 0.0177772f $X=10.02 $Y=1.325
+ $X2=0 $Y2=0
cc_877 N_A_1517_315#_c_1286_n N_A_1948_47#_c_1500_n 0.00252128f $X=9.945 $Y=1.16
+ $X2=0 $Y2=0
cc_878 N_A_1517_315#_M1030_g N_A_1948_47#_c_1507_n 5.32975e-19 $X=10.075
+ $Y=2.165 $X2=0 $Y2=0
cc_879 N_A_1517_315#_c_1300_n N_A_1948_47#_c_1507_n 0.00764243f $X=10.047
+ $Y=1.515 $X2=0 $Y2=0
cc_880 N_A_1517_315#_c_1301_n N_A_1948_47#_c_1507_n 0.00643794f $X=10.047
+ $Y=1.665 $X2=0 $Y2=0
cc_881 N_A_1517_315#_c_1286_n N_A_1948_47#_c_1523_n 0.0134399f $X=9.945 $Y=1.16
+ $X2=0 $Y2=0
cc_882 N_A_1517_315#_c_1287_n N_A_1948_47#_c_1523_n 0.00652717f $X=10.02
+ $Y=1.325 $X2=0 $Y2=0
cc_883 N_A_1517_315#_c_1287_n N_A_1948_47#_c_1501_n 0.00317818f $X=10.02
+ $Y=1.325 $X2=0 $Y2=0
cc_884 N_A_1517_315#_c_1288_n N_A_1948_47#_c_1501_n 0.0140671f $X=10.075 $Y=0.73
+ $X2=0 $Y2=0
cc_885 N_A_1517_315#_M1015_g N_VPWR_c_1562_n 0.0115962f $X=7.66 $Y=2.275 $X2=0
+ $Y2=0
cc_886 N_A_1517_315#_c_1302_n N_VPWR_c_1562_n 0.0182102f $X=8.38 $Y=1.74 $X2=0
+ $Y2=0
cc_887 N_A_1517_315#_c_1303_n N_VPWR_c_1562_n 0.0049226f $X=7.84 $Y=1.74 $X2=0
+ $Y2=0
cc_888 N_A_1517_315#_c_1316_p N_VPWR_c_1562_n 0.01625f $X=8.505 $Y=1.95 $X2=0
+ $Y2=0
cc_889 N_A_1517_315#_M1028_g N_VPWR_c_1563_n 0.00313741f $X=9.135 $Y=1.985 $X2=0
+ $Y2=0
cc_890 N_A_1517_315#_c_1291_n N_VPWR_c_1563_n 0.00929281f $X=9.135 $Y=1.16 $X2=0
+ $Y2=0
cc_891 N_A_1517_315#_c_1301_n N_VPWR_c_1564_n 0.0119616f $X=10.047 $Y=1.665
+ $X2=0 $Y2=0
cc_892 N_A_1517_315#_M1015_g N_VPWR_c_1569_n 0.00585385f $X=7.66 $Y=2.275 $X2=0
+ $Y2=0
cc_893 N_A_1517_315#_c_1316_p N_VPWR_c_1573_n 0.0170823f $X=8.505 $Y=1.95 $X2=0
+ $Y2=0
cc_894 N_A_1517_315#_M1028_g N_VPWR_c_1574_n 0.00571722f $X=9.135 $Y=1.985 $X2=0
+ $Y2=0
cc_895 N_A_1517_315#_M1030_g N_VPWR_c_1574_n 0.00542953f $X=10.075 $Y=2.165
+ $X2=0 $Y2=0
cc_896 N_A_1517_315#_M1001_s N_VPWR_c_1557_n 0.00208837f $X=8.38 $Y=1.485 $X2=0
+ $Y2=0
cc_897 N_A_1517_315#_M1015_g N_VPWR_c_1557_n 0.0124099f $X=7.66 $Y=2.275 $X2=0
+ $Y2=0
cc_898 N_A_1517_315#_M1028_g N_VPWR_c_1557_n 0.0116712f $X=9.135 $Y=1.985 $X2=0
+ $Y2=0
cc_899 N_A_1517_315#_M1030_g N_VPWR_c_1557_n 0.0111168f $X=10.075 $Y=2.165 $X2=0
+ $Y2=0
cc_900 N_A_1517_315#_c_1302_n N_VPWR_c_1557_n 0.0130411f $X=8.38 $Y=1.74 $X2=0
+ $Y2=0
cc_901 N_A_1517_315#_c_1303_n N_VPWR_c_1557_n 7.75814e-19 $X=7.84 $Y=1.74 $X2=0
+ $Y2=0
cc_902 N_A_1517_315#_c_1316_p N_VPWR_c_1557_n 0.0108334f $X=8.505 $Y=1.95 $X2=0
+ $Y2=0
cc_903 N_A_1517_315#_M1028_g N_Q_c_1854_n 0.0143565f $X=9.135 $Y=1.985 $X2=0
+ $Y2=0
cc_904 N_A_1517_315#_M1030_g N_Q_c_1854_n 0.00157346f $X=10.075 $Y=2.165 $X2=0
+ $Y2=0
cc_905 N_A_1517_315#_c_1301_n N_Q_c_1854_n 6.22549e-19 $X=10.047 $Y=1.665 $X2=0
+ $Y2=0
cc_906 N_A_1517_315#_c_1304_n N_Q_c_1854_n 9.62634e-19 $X=8.577 $Y=1.575 $X2=0
+ $Y2=0
cc_907 N_A_1517_315#_c_1318_p N_Q_c_1854_n 0.00156781f $X=8.525 $Y=1.74 $X2=0
+ $Y2=0
cc_908 N_A_1517_315#_c_1285_n N_Q_c_1851_n 0.00489844f $X=9.135 $Y=0.995 $X2=0
+ $Y2=0
cc_909 N_A_1517_315#_M1028_g N_Q_c_1851_n 0.00676807f $X=9.135 $Y=1.985 $X2=0
+ $Y2=0
cc_910 N_A_1517_315#_c_1286_n N_Q_c_1851_n 0.0281429f $X=9.945 $Y=1.16 $X2=0
+ $Y2=0
cc_911 N_A_1517_315#_c_1287_n N_Q_c_1851_n 8.4021e-19 $X=10.02 $Y=1.325 $X2=0
+ $Y2=0
cc_912 N_A_1517_315#_c_1300_n N_Q_c_1851_n 0.00105777f $X=10.047 $Y=1.515 $X2=0
+ $Y2=0
cc_913 N_A_1517_315#_c_1304_n N_Q_c_1851_n 0.00101051f $X=8.577 $Y=1.575 $X2=0
+ $Y2=0
cc_914 N_A_1517_315#_c_1291_n N_Q_c_1851_n 0.0264832f $X=9.135 $Y=1.16 $X2=0
+ $Y2=0
cc_915 N_A_1517_315#_c_1285_n N_Q_c_1852_n 0.00214656f $X=9.135 $Y=0.995 $X2=0
+ $Y2=0
cc_916 N_A_1517_315#_c_1286_n N_Q_c_1852_n 0.00263236f $X=9.945 $Y=1.16 $X2=0
+ $Y2=0
cc_917 N_A_1517_315#_c_1287_n N_Q_c_1852_n 4.86053e-19 $X=10.02 $Y=1.325 $X2=0
+ $Y2=0
cc_918 N_A_1517_315#_c_1291_n N_Q_c_1852_n 0.00264474f $X=9.135 $Y=1.16 $X2=0
+ $Y2=0
cc_919 N_A_1517_315#_c_1293_n N_Q_c_1852_n 0.00310961f $X=8.505 $Y=0.825 $X2=0
+ $Y2=0
cc_920 N_A_1517_315#_c_1285_n N_Q_c_1853_n 0.00487455f $X=9.135 $Y=0.995 $X2=0
+ $Y2=0
cc_921 N_A_1517_315#_c_1288_n N_Q_c_1853_n 9.486e-19 $X=10.075 $Y=0.73 $X2=0
+ $Y2=0
cc_922 N_A_1517_315#_c_1293_n N_Q_c_1853_n 9.0648e-19 $X=8.505 $Y=0.825 $X2=0
+ $Y2=0
cc_923 N_A_1517_315#_M1016_g N_VGND_c_1914_n 0.0215676f $X=7.775 $Y=0.445 $X2=0
+ $Y2=0
cc_924 N_A_1517_315#_c_1289_n N_VGND_c_1914_n 0.0186495f $X=8.505 $Y=0.385 $X2=0
+ $Y2=0
cc_925 N_A_1517_315#_c_1285_n N_VGND_c_1915_n 0.00309623f $X=9.135 $Y=0.995
+ $X2=0 $Y2=0
cc_926 N_A_1517_315#_c_1291_n N_VGND_c_1915_n 0.00929281f $X=9.135 $Y=1.16 $X2=0
+ $Y2=0
cc_927 N_A_1517_315#_c_1288_n N_VGND_c_1916_n 0.00667732f $X=10.075 $Y=0.73
+ $X2=0 $Y2=0
cc_928 N_A_1517_315#_c_1289_n N_VGND_c_1922_n 0.0161941f $X=8.505 $Y=0.385 $X2=0
+ $Y2=0
cc_929 N_A_1517_315#_c_1285_n N_VGND_c_1923_n 0.00543342f $X=9.135 $Y=0.995
+ $X2=0 $Y2=0
cc_930 N_A_1517_315#_c_1287_n N_VGND_c_1923_n 0.00105583f $X=10.02 $Y=1.325
+ $X2=0 $Y2=0
cc_931 N_A_1517_315#_c_1288_n N_VGND_c_1923_n 0.00585385f $X=10.075 $Y=0.73
+ $X2=0 $Y2=0
cc_932 N_A_1517_315#_M1011_s N_VGND_c_1925_n 0.00212021f $X=8.38 $Y=0.235 $X2=0
+ $Y2=0
cc_933 N_A_1517_315#_M1016_g N_VGND_c_1925_n 9.61436e-19 $X=7.775 $Y=0.445 $X2=0
+ $Y2=0
cc_934 N_A_1517_315#_c_1285_n N_VGND_c_1925_n 0.0109354f $X=9.135 $Y=0.995 $X2=0
+ $Y2=0
cc_935 N_A_1517_315#_c_1287_n N_VGND_c_1925_n 0.00138273f $X=10.02 $Y=1.325
+ $X2=0 $Y2=0
cc_936 N_A_1517_315#_c_1288_n N_VGND_c_1925_n 0.0122138f $X=10.075 $Y=0.73 $X2=0
+ $Y2=0
cc_937 N_A_1517_315#_c_1289_n N_VGND_c_1925_n 0.0121006f $X=8.505 $Y=0.385 $X2=0
+ $Y2=0
cc_938 N_A_1346_413#_M1001_g N_VPWR_c_1562_n 0.0021703f $X=8.715 $Y=1.985 $X2=0
+ $Y2=0
cc_939 N_A_1346_413#_M1001_g N_VPWR_c_1563_n 0.00313741f $X=8.715 $Y=1.985 $X2=0
+ $Y2=0
cc_940 N_A_1346_413#_c_1421_n N_VPWR_c_1569_n 0.0273845f $X=7.415 $Y=2.25 $X2=0
+ $Y2=0
cc_941 N_A_1346_413#_M1001_g N_VPWR_c_1573_n 0.00541763f $X=8.715 $Y=1.985 $X2=0
+ $Y2=0
cc_942 N_A_1346_413#_M1006_d N_VPWR_c_1557_n 0.00219484f $X=6.73 $Y=2.065 $X2=0
+ $Y2=0
cc_943 N_A_1346_413#_M1001_g N_VPWR_c_1557_n 0.0109319f $X=8.715 $Y=1.985 $X2=0
+ $Y2=0
cc_944 N_A_1346_413#_c_1421_n N_VPWR_c_1557_n 0.0276628f $X=7.415 $Y=2.25 $X2=0
+ $Y2=0
cc_945 N_A_1346_413#_c_1421_n A_1430_413# 0.0105858f $X=7.415 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_946 N_A_1346_413#_c_1418_n A_1430_413# 0.00184879f $X=7.5 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_947 N_A_1346_413#_M1001_g N_Q_c_1854_n 4.38906e-19 $X=8.715 $Y=1.985 $X2=0
+ $Y2=0
cc_948 N_A_1346_413#_c_1409_n N_Q_c_1852_n 2.93604e-19 $X=8.715 $Y=0.995 $X2=0
+ $Y2=0
cc_949 N_A_1346_413#_c_1409_n N_VGND_c_1914_n 0.00268732f $X=8.715 $Y=0.995
+ $X2=0 $Y2=0
cc_950 N_A_1346_413#_c_1424_n N_VGND_c_1914_n 0.0104892f $X=7.285 $Y=0.45 $X2=0
+ $Y2=0
cc_951 N_A_1346_413#_c_1412_n N_VGND_c_1914_n 0.0154767f $X=8.23 $Y=1.16 $X2=0
+ $Y2=0
cc_952 N_A_1346_413#_c_1414_n N_VGND_c_1914_n 0.00447237f $X=7.435 $Y=0.995
+ $X2=0 $Y2=0
cc_953 N_A_1346_413#_c_1409_n N_VGND_c_1915_n 0.00309623f $X=8.715 $Y=0.995
+ $X2=0 $Y2=0
cc_954 N_A_1346_413#_c_1424_n N_VGND_c_1917_n 0.0184388f $X=7.285 $Y=0.45 $X2=0
+ $Y2=0
cc_955 N_A_1346_413#_c_1409_n N_VGND_c_1922_n 0.00543148f $X=8.715 $Y=0.995
+ $X2=0 $Y2=0
cc_956 N_A_1346_413#_M1002_d N_VGND_c_1925_n 0.00333348f $X=6.86 $Y=0.235 $X2=0
+ $Y2=0
cc_957 N_A_1346_413#_c_1409_n N_VGND_c_1925_n 0.0109348f $X=8.715 $Y=0.995 $X2=0
+ $Y2=0
cc_958 N_A_1346_413#_c_1424_n N_VGND_c_1925_n 0.0182474f $X=7.285 $Y=0.45 $X2=0
+ $Y2=0
cc_959 N_A_1346_413#_c_1424_n A_1475_47# 0.00201232f $X=7.285 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_960 N_A_1346_413#_c_1414_n A_1475_47# 0.00127737f $X=7.435 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_961 N_A_1948_47#_M1007_g N_VPWR_c_1564_n 0.0211857f $X=10.56 $Y=1.985 $X2=0
+ $Y2=0
cc_962 N_A_1948_47#_c_1498_n N_VPWR_c_1564_n 0.0228967f $X=10.475 $Y=1.16 $X2=0
+ $Y2=0
cc_963 N_A_1948_47#_c_1499_n N_VPWR_c_1564_n 0.00320419f $X=10.475 $Y=1.16 $X2=0
+ $Y2=0
cc_964 N_A_1948_47#_c_1507_n N_VPWR_c_1564_n 0.0687607f $X=9.865 $Y=1.685 $X2=0
+ $Y2=0
cc_965 N_A_1948_47#_c_1504_n N_VPWR_c_1574_n 0.016757f $X=9.865 $Y=2 $X2=0 $Y2=0
cc_966 N_A_1948_47#_M1007_g N_VPWR_c_1575_n 0.0046653f $X=10.56 $Y=1.985 $X2=0
+ $Y2=0
cc_967 N_A_1948_47#_M1030_s N_VPWR_c_1557_n 0.00211564f $X=9.74 $Y=1.845 $X2=0
+ $Y2=0
cc_968 N_A_1948_47#_M1007_g N_VPWR_c_1557_n 0.00896841f $X=10.56 $Y=1.985 $X2=0
+ $Y2=0
cc_969 N_A_1948_47#_c_1504_n N_VPWR_c_1557_n 0.0121755f $X=9.865 $Y=2 $X2=0
+ $Y2=0
cc_970 N_A_1948_47#_c_1503_n N_Q_c_1854_n 0.0615769f $X=9.865 $Y=1.85 $X2=0
+ $Y2=0
cc_971 N_A_1948_47#_c_1507_n N_Q_c_1854_n 0.00897636f $X=9.865 $Y=1.685 $X2=0
+ $Y2=0
cc_972 N_A_1948_47#_c_1497_n N_Q_c_1851_n 0.0129793f $X=9.865 $Y=0.995 $X2=0
+ $Y2=0
cc_973 N_A_1948_47#_c_1507_n N_Q_c_1851_n 0.017165f $X=9.865 $Y=1.685 $X2=0
+ $Y2=0
cc_974 N_A_1948_47#_c_1523_n N_Q_c_1851_n 0.0255923f $X=9.905 $Y=1.16 $X2=0
+ $Y2=0
cc_975 N_A_1948_47#_c_1497_n N_Q_c_1852_n 0.00721425f $X=9.865 $Y=0.995 $X2=0
+ $Y2=0
cc_976 N_A_1948_47#_c_1497_n N_Q_c_1853_n 0.00628298f $X=9.865 $Y=0.995 $X2=0
+ $Y2=0
cc_977 N_A_1948_47#_c_1500_n N_Q_c_1853_n 0.0225298f $X=9.865 $Y=0.51 $X2=0
+ $Y2=0
cc_978 N_A_1948_47#_M1007_g Q_N 0.00384193f $X=10.56 $Y=1.985 $X2=0 $Y2=0
cc_979 N_A_1948_47#_c_1498_n Q_N 0.0266145f $X=10.475 $Y=1.16 $X2=0 $Y2=0
cc_980 N_A_1948_47#_c_1507_n Q_N 0.00118007f $X=9.865 $Y=1.685 $X2=0 $Y2=0
cc_981 N_A_1948_47#_c_1501_n Q_N 0.0193867f $X=10.487 $Y=0.995 $X2=0 $Y2=0
cc_982 N_A_1948_47#_c_1497_n N_VGND_c_1916_n 0.00912263f $X=9.865 $Y=0.995 $X2=0
+ $Y2=0
cc_983 N_A_1948_47#_c_1498_n N_VGND_c_1916_n 0.0230938f $X=10.475 $Y=1.16 $X2=0
+ $Y2=0
cc_984 N_A_1948_47#_c_1499_n N_VGND_c_1916_n 0.00315906f $X=10.475 $Y=1.16 $X2=0
+ $Y2=0
cc_985 N_A_1948_47#_c_1501_n N_VGND_c_1916_n 0.0124584f $X=10.487 $Y=0.995 $X2=0
+ $Y2=0
cc_986 N_A_1948_47#_c_1500_n N_VGND_c_1923_n 0.0107099f $X=9.865 $Y=0.51 $X2=0
+ $Y2=0
cc_987 N_A_1948_47#_c_1501_n N_VGND_c_1924_n 0.0046653f $X=10.487 $Y=0.995 $X2=0
+ $Y2=0
cc_988 N_A_1948_47#_M1033_s N_VGND_c_1925_n 0.00272276f $X=9.74 $Y=0.235 $X2=0
+ $Y2=0
cc_989 N_A_1948_47#_c_1500_n N_VGND_c_1925_n 0.00902066f $X=9.865 $Y=0.51 $X2=0
+ $Y2=0
cc_990 N_A_1948_47#_c_1501_n N_VGND_c_1925_n 0.00896841f $X=10.487 $Y=0.995
+ $X2=0 $Y2=0
cc_991 N_VPWR_c_1557_n A_465_369# 0.00270153f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_992 N_VPWR_c_1557_n N_A_556_369#_M1027_d 0.00179277f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_993 N_VPWR_c_1557_n N_A_556_369#_M1003_s 0.00201964f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_994 N_VPWR_c_1559_n N_A_556_369#_c_1739_n 0.00585291f $X=2.04 $Y=2.33 $X2=0
+ $Y2=0
cc_995 N_VPWR_c_1560_n N_A_556_369#_c_1739_n 0.0133617f $X=3.825 $Y=2.33 $X2=0
+ $Y2=0
cc_996 N_VPWR_c_1565_n N_A_556_369#_c_1739_n 0.0382569f $X=3.74 $Y=2.72 $X2=0
+ $Y2=0
cc_997 N_VPWR_c_1557_n N_A_556_369#_c_1739_n 0.0141922f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_998 N_VPWR_c_1560_n N_A_556_369#_c_1763_n 0.00558244f $X=3.825 $Y=2.33 $X2=0
+ $Y2=0
cc_999 N_VPWR_M1014_d N_A_556_369#_c_1735_n 0.00372198f $X=3.665 $Y=1.845 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1560_n N_A_556_369#_c_1735_n 0.0119067f $X=3.825 $Y=2.33 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1565_n N_A_556_369#_c_1735_n 0.00196122f $X=3.74 $Y=2.72 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1567_n N_A_556_369#_c_1735_n 0.00384075f $X=5.885 $Y=2.72 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1557_n N_A_556_369#_c_1735_n 0.00499201f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_1004 N_VPWR_c_1560_n N_A_556_369#_c_1738_n 0.0159048f $X=3.825 $Y=2.33 $X2=0
+ $Y2=0
cc_1005 N_VPWR_c_1567_n N_A_556_369#_c_1738_n 0.0168495f $X=5.885 $Y=2.72 $X2=0
+ $Y2=0
cc_1006 N_VPWR_c_1557_n N_A_556_369#_c_1738_n 0.0050874f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_1007 N_VPWR_c_1557_n A_640_369# 0.00210687f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1008 N_VPWR_c_1557_n A_1023_413# 0.00220519f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1009 N_VPWR_c_1557_n A_1430_413# 0.00377587f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1010 N_VPWR_c_1557_n N_Q_M1028_d 0.00209319f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1011 N_VPWR_c_1574_n N_Q_c_1854_n 0.0211085f $X=10.21 $Y=2.72 $X2=0 $Y2=0
cc_1012 N_VPWR_c_1557_n N_Q_c_1854_n 0.0125182f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1013 N_VPWR_c_1557_n N_Q_N_M1007_d 0.00401809f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1014 N_VPWR_c_1575_n Q_N 0.00923202f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1015 N_VPWR_c_1557_n Q_N 0.00900352f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1016 N_A_556_369#_c_1739_n A_640_369# 0.00382565f $X=3.4 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_1017 N_A_556_369#_c_1763_n A_640_369# 0.00266005f $X=3.485 $Y=2.245 $X2=-0.19
+ $Y2=-0.24
cc_1018 N_A_556_369#_c_1736_n A_640_369# 9.25434e-19 $X=3.57 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_1019 N_A_556_369#_c_1751_n N_VGND_c_1910_n 9.32728e-19 $X=3.405 $Y=0.36 $X2=0
+ $Y2=0
cc_1020 N_A_556_369#_c_1751_n N_VGND_c_1911_n 0.0135146f $X=3.405 $Y=0.36 $X2=0
+ $Y2=0
cc_1021 N_A_556_369#_c_1728_n N_VGND_c_1911_n 0.00707611f $X=3.49 $Y=0.715 $X2=0
+ $Y2=0
cc_1022 N_A_556_369#_c_1729_n N_VGND_c_1911_n 0.0142754f $X=4.165 $Y=0.8 $X2=0
+ $Y2=0
cc_1023 N_A_556_369#_c_1731_n N_VGND_c_1911_n 6.21916e-19 $X=4.25 $Y=0.715 $X2=0
+ $Y2=0
cc_1024 N_A_556_369#_c_1733_n N_VGND_c_1911_n 0.0111003f $X=4.35 $Y=0.45 $X2=0
+ $Y2=0
cc_1025 N_A_556_369#_c_1729_n N_VGND_c_1912_n 0.00340284f $X=4.165 $Y=0.8 $X2=0
+ $Y2=0
cc_1026 N_A_556_369#_c_1733_n N_VGND_c_1912_n 0.012161f $X=4.35 $Y=0.45 $X2=0
+ $Y2=0
cc_1027 N_A_556_369#_c_1751_n N_VGND_c_1921_n 0.0381445f $X=3.405 $Y=0.36 $X2=0
+ $Y2=0
cc_1028 N_A_556_369#_c_1729_n N_VGND_c_1921_n 0.00246058f $X=4.165 $Y=0.8 $X2=0
+ $Y2=0
cc_1029 N_A_556_369#_M1020_d N_VGND_c_1925_n 0.00217379f $X=2.805 $Y=0.235 $X2=0
+ $Y2=0
cc_1030 N_A_556_369#_M1031_s N_VGND_c_1925_n 0.00195217f $X=4.225 $Y=0.235 $X2=0
+ $Y2=0
cc_1031 N_A_556_369#_c_1751_n N_VGND_c_1925_n 0.012723f $X=3.405 $Y=0.36 $X2=0
+ $Y2=0
cc_1032 N_A_556_369#_c_1729_n N_VGND_c_1925_n 0.00472438f $X=4.165 $Y=0.8 $X2=0
+ $Y2=0
cc_1033 N_A_556_369#_c_1733_n N_VGND_c_1925_n 0.00544577f $X=4.35 $Y=0.45 $X2=0
+ $Y2=0
cc_1034 N_A_556_369#_c_1751_n A_657_47# 0.00210941f $X=3.405 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1035 N_A_556_369#_c_1728_n A_657_47# 0.00222412f $X=3.49 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_1036 N_Q_c_1852_n N_VGND_c_1923_n 5.10712e-19 $X=9.355 $Y=0.725 $X2=0 $Y2=0
cc_1037 N_Q_c_1853_n N_VGND_c_1923_n 0.016881f $X=9.345 $Y=0.395 $X2=0 $Y2=0
cc_1038 N_Q_M1010_d N_VGND_c_1925_n 0.00212516f $X=9.21 $Y=0.235 $X2=0 $Y2=0
cc_1039 N_Q_c_1852_n N_VGND_c_1925_n 0.00289201f $X=9.355 $Y=0.725 $X2=0 $Y2=0
cc_1040 N_Q_c_1853_n N_VGND_c_1925_n 0.0127972f $X=9.345 $Y=0.395 $X2=0 $Y2=0
cc_1041 Q_N N_VGND_c_1916_n 5.94513e-19 $X=10.715 $Y=1.445 $X2=0 $Y2=0
cc_1042 N_Q_N_c_1894_n N_VGND_c_1924_n 0.0165374f $X=10.812 $Y=0.668 $X2=0 $Y2=0
cc_1043 N_Q_N_M1023_d N_VGND_c_1925_n 0.00387432f $X=10.635 $Y=0.235 $X2=0 $Y2=0
cc_1044 N_Q_N_c_1894_n N_VGND_c_1925_n 0.00968619f $X=10.812 $Y=0.668 $X2=0
+ $Y2=0
cc_1045 N_VGND_c_1925_n A_483_47# 0.00171756f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1046 N_VGND_c_1925_n A_657_47# 0.00152414f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1047 N_VGND_c_1925_n A_1027_47# 0.00272292f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1048 N_VGND_c_1925_n A_1475_47# 0.0111093f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24

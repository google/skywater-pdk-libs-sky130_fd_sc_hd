* File: sky130_fd_sc_hd__buf_2.spice
* Created: Thu Aug 27 14:09:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__buf_2.spice.pex"
.subckt sky130_fd_sc_hd__buf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=11.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1004_d N_A_27_47#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.08775 PD=1.18458 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_27_47#_M1005_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.08775 PD=1.83 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=12.2928 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1001_d N_A_27_47#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.181707 AS=0.135 PD=1.61585 PS=1.27 NRD=0.9653 NRS=0 M=1 R=6.66667
+ SA=75000.5 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_27_47#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.135 PD=2.53 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=3.5631 P=7.65
c_38 VPB 0 1.42894e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__buf_2.spice.SKY130_FD_SC_HD__BUF_2.pxi"
*
.ends
*
*

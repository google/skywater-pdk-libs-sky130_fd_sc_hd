* File: sky130_fd_sc_hd__a311o_2.pex.spice
* Created: Thu Aug 27 14:04:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A311O_2%A_79_21# 1 2 3 10 12 15 17 19 22 27 28 29 30
+ 31 32 34 35 36 40 41 42 45 49
c116 28 0 1.86031e-19 $X=1.1 $Y=1.16
c117 27 0 1.11805e-19 $X=1.1 $Y=1.16
r118 51 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r119 47 49 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.88 $Y=1.665
+ $X2=3.88 $Y2=1.96
r120 43 45 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.88 $Y=0.655
+ $X2=3.88 $Y2=0.42
r121 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.795 $Y=0.74
+ $X2=3.88 $Y2=0.655
r122 41 42 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.795 $Y=0.74
+ $X2=2.96 $Y2=0.74
r123 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.875 $Y=0.655
+ $X2=2.96 $Y2=0.74
r124 38 40 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.655
+ $X2=2.875 $Y2=0.57
r125 37 40 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.875 $Y=0.425
+ $X2=2.875 $Y2=0.57
r126 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.79 $Y=0.34
+ $X2=2.875 $Y2=0.425
r127 35 36 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=2.79 $Y=0.34
+ $X2=1.695 $Y2=0.34
r128 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.61 $Y=0.425
+ $X2=1.695 $Y2=0.34
r129 33 34 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.61 $Y=0.425
+ $X2=1.61 $Y2=0.655
r130 31 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.795 $Y=1.58
+ $X2=3.88 $Y2=1.665
r131 31 32 170.278 $w=1.68e-07 $l=2.61e-06 $layer=LI1_cond $X=3.795 $Y=1.58
+ $X2=1.185 $Y2=1.58
r132 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=0.74
+ $X2=1.61 $Y2=0.655
r133 29 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.525 $Y=0.74
+ $X2=1.185 $Y2=0.74
r134 28 53 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.1 $Y=1.16
+ $X2=0.89 $Y2=1.16
r135 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r136 25 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.1 $Y=1.495
+ $X2=1.185 $Y2=1.58
r137 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=1.495
+ $X2=1.1 $Y2=1.16
r138 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.1 $Y=0.825
+ $X2=1.185 $Y2=0.74
r139 24 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=0.825
+ $X2=1.1 $Y2=1.16
r140 20 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r141 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r142 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r143 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r144 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r145 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r146 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r147 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r148 3 49 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=1.96
r149 2 45 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.42
r150 1 40 182 $w=1.7e-07 $l=4.50194e-07 $layer=licon1_NDIFF $count=1 $X=2.605
+ $Y=0.235 $X2=2.875 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%A3 3 6 8 11 13
r39 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.16
+ $X2=1.58 $Y2=1.325
r40 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.16
+ $X2=1.58 $Y2=0.995
r41 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.16 $X2=1.58 $Y2=1.16
r42 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.52 $Y=1.985
+ $X2=1.52 $Y2=1.325
r43 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.52 $Y=0.56 $X2=1.52
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%A2 3 6 8 11 13
r36 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.16
+ $X2=2.07 $Y2=1.325
r37 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.16
+ $X2=2.07 $Y2=0.995
r38 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.16 $X2=2.07 $Y2=1.16
r39 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.01 $Y=1.985
+ $X2=2.01 $Y2=1.325
r40 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.01 $Y=0.56 $X2=2.01
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%A1 3 6 10 13 15
r36 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.59 $Y2=1.325
r37 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.59 $Y2=0.995
r38 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.16 $X2=2.59 $Y2=1.16
r39 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.53 $Y=1.985
+ $X2=2.53 $Y2=1.325
r40 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.53 $Y=0.56 $X2=2.53
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%B1 3 6 8 11 12 13
r31 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.16
+ $X2=3.15 $Y2=1.325
r32 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.16
+ $X2=3.15 $Y2=0.995
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.16 $X2=3.15 $Y2=1.16
r34 8 12 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=3.15 $Y2=1.16
r35 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.1 $Y=1.985 $X2=3.1
+ $Y2=1.325
r36 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.09 $Y=0.56 $X2=3.09
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%C1 3 6 8 11 13
r23 11 14 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.16
+ $X2=3.755 $Y2=1.325
r24 11 13 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.16
+ $X2=3.755 $Y2=0.995
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.16 $X2=3.78 $Y2=1.16
r26 8 12 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.905 $Y=1.16
+ $X2=3.78 $Y2=1.16
r27 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.985
+ $X2=3.67 $Y2=1.325
r28 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.67 $Y=0.56 $X2=3.67
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%VPWR 1 2 3 10 12 18 22 25 26 28 29 30 43 44
c58 18 0 1.86031e-19 $X=1.245 $Y=2
c59 2 0 1.11805e-19 $X=0.965 $Y=1.485
r60 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 41 44 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 40 43 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 38 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 32 47 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r69 32 34 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 30 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 30 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 28 37 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.07 $Y2=2.72
r73 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.29 $Y2=2.72
r74 27 40 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=2.53 $Y2=2.72
r75 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=2.29 $Y2=2.72
r76 25 34 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=2.72 $X2=1.15
+ $Y2=2.72
r77 25 26 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.16 $Y=2.72 $X2=1.27
+ $Y2=2.72
r78 24 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.38 $Y=2.72 $X2=2.07
+ $Y2=2.72
r79 24 26 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.38 $Y=2.72 $X2=1.27
+ $Y2=2.72
r80 20 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.635
+ $X2=2.29 $Y2=2.72
r81 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.29 $Y=2.635
+ $X2=2.29 $Y2=2.34
r82 16 26 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.635
+ $X2=1.27 $Y2=2.72
r83 16 18 33.2637 $w=2.18e-07 $l=6.35e-07 $layer=LI1_cond $X=1.27 $Y=2.635
+ $X2=1.27 $Y2=2
r84 12 15 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r85 10 47 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r86 10 15 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r87 3 22 600 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=1.485 $X2=2.29 $Y2=2.34
r88 2 18 300 $w=1.7e-07 $l=6.39863e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.245 $Y2=2
r89 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r90 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%X 1 2 7 8 9 10 11 12 20
r15 12 37 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=2.21
+ $X2=0.68 $Y2=2.34
r16 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=2.21
r17 11 31 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=1.66
r18 10 31 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=1.53
+ $X2=0.68 $Y2=1.66
r19 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=1.19 $X2=0.68
+ $Y2=1.53
r20 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.85 $X2=0.68
+ $Y2=1.19
r21 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.51 $X2=0.68
+ $Y2=0.85
r22 7 20 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.68 $Y=0.51 $X2=0.68
+ $Y2=0.38
r23 2 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r24 2 31 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r25 1 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%A_319_297# 1 2 7 9 11 13 15
r24 13 20 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=2.005
+ $X2=2.87 $Y2=1.92
r25 13 15 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.87 $Y=2.005
+ $X2=2.87 $Y2=2.3
r26 12 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.84 $Y=1.92
+ $X2=1.715 $Y2=1.92
r27 11 20 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.715 $Y=1.92
+ $X2=2.87 $Y2=1.92
r28 11 12 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.715 $Y=1.92
+ $X2=1.84 $Y2=1.92
r29 7 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=2.005
+ $X2=1.715 $Y2=1.92
r30 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.715 $Y=2.005
+ $X2=1.715 $Y2=2.3
r31 2 20 600 $w=1.7e-07 $l=5.47859e-07 $layer=licon1_PDIFF $count=1 $X=2.605
+ $Y=1.485 $X2=2.86 $Y2=1.92
r32 2 15 600 $w=1.7e-07 $l=9.33836e-07 $layer=licon1_PDIFF $count=1 $X=2.605
+ $Y=1.485 $X2=2.86 $Y2=2.3
r33 1 18 600 $w=1.7e-07 $l=5.08748e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.485 $X2=1.755 $Y2=1.92
r34 1 9 600 $w=1.7e-07 $l=8.91417e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.485 $X2=1.755 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A311O_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r59 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r60 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 40 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r62 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r63 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.385
+ $Y2=0
r64 37 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.91
+ $Y2=0
r65 36 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r66 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r67 33 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r68 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r69 32 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r70 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r71 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.18
+ $Y2=0
r72 30 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.61
+ $Y2=0
r73 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.385
+ $Y2=0
r74 29 35 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=2.99
+ $Y2=0
r75 28 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r76 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r77 25 43 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r78 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r79 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.18
+ $Y2=0
r80 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.69
+ $Y2=0
r81 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r82 22 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r83 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=0.085
+ $X2=3.385 $Y2=0
r84 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.385 $Y=0.085
+ $X2=3.385 $Y2=0.4
r85 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0
r86 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.38
r87 10 43 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r88 10 12 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.38
r89 3 20 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.385 $Y2=0.4
r90 2 16 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.18 $Y2=0.38
r91 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


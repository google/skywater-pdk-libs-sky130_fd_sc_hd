* File: sky130_fd_sc_hd__clkdlybuf4s15_1.spice.pex
* Created: Thu Aug 27 14:11:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A 3 7 9 12 13
r31 12 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.39 $Y=1.16
+ $X2=0.39 $Y2=1.325
r32 12 14 40.7411 $w=3.2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.39 $Y=1.16
+ $X2=0.39 $Y2=1.025
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.395
+ $Y=1.16 $X2=0.395 $Y2=1.16
r34 9 13 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.395 $Y2=1.19
r35 7 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r36 3 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_27_47# 1 2 7 9 12 14 15 18 22 24
+ 25 26 27 31
r65 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.16 $X2=0.925 $Y2=1.16
r66 29 31 8.26157 $w=4.83e-07 $l=3.35e-07 $layer=LI1_cond $X=0.972 $Y=1.495
+ $X2=0.972 $Y2=1.16
r67 28 31 6.78189 $w=4.83e-07 $l=2.75e-07 $layer=LI1_cond $X=0.972 $Y=0.885
+ $X2=0.972 $Y2=1.16
r68 26 29 9.10402 $w=1.7e-07 $l=2.81308e-07 $layer=LI1_cond $X=0.73 $Y=1.58
+ $X2=0.972 $Y2=1.495
r69 26 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=1.58
+ $X2=0.425 $Y2=1.58
r70 24 28 9.10402 $w=1.7e-07 $l=2.81308e-07 $layer=LI1_cond $X=0.73 $Y=0.8
+ $X2=0.972 $Y2=0.885
r71 24 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.8
+ $X2=0.425 $Y2=0.8
r72 20 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.425 $Y2=1.58
r73 20 22 10.1686 $w=3.38e-07 $l=3e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.965
r74 16 25 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.425 $Y2=0.8
r75 16 18 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.38
r76 14 32 66.9854 $w=3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.26 $Y=1.145
+ $X2=0.925 $Y2=1.145
r77 14 15 3.90195 $w=3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.26 $Y=1.145
+ $X2=1.335 $Y2=1.145
r78 10 15 34.7346 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.335 $Y=1.295
+ $X2=1.335 $Y2=1.145
r79 10 12 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.335 $Y=1.295
+ $X2=1.335 $Y2=2.075
r80 7 15 34.7346 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=1.145
r81 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=0.56
r82 2 22 300 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.965
r83 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_282_47# 1 2 7 9 12 15 18 23 28 29
+ 31 33 34 35
c64 28 0 1.84838e-19 $X=2.52 $Y=1.16
r65 33 34 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.572 $Y=2
+ $X2=1.572 $Y2=1.835
r66 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.16 $X2=2.52 $Y2=1.16
r67 26 35 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=1.152
+ $X2=1.675 $Y2=1.152
r68 26 28 43.2261 $w=1.93e-07 $l=7.6e-07 $layer=LI1_cond $X=1.76 $Y=1.152
+ $X2=2.52 $Y2=1.152
r69 24 35 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.675 $Y=1.25
+ $X2=1.675 $Y2=1.152
r70 24 34 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.675 $Y=1.25
+ $X2=1.675 $Y2=1.835
r71 23 35 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.675 $Y=1.055
+ $X2=1.675 $Y2=1.152
r72 23 31 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.675 $Y=1.055
+ $X2=1.675 $Y2=0.825
r73 16 31 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=1.572 $Y=0.638
+ $X2=1.572 $Y2=0.825
r74 16 18 7.92881 $w=3.73e-07 $l=2.58e-07 $layer=LI1_cond $X=1.572 $Y=0.638
+ $X2=1.572 $Y2=0.38
r75 14 29 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.385 $Y=1.165
+ $X2=2.52 $Y2=1.165
r76 14 15 5.03009 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.385 $Y=1.165
+ $X2=2.2 $Y2=1.165
r77 10 15 37.0704 $w=1.5e-07 $l=2.13014e-07 $layer=POLY_cond $X=2.31 $Y=1.33
+ $X2=2.2 $Y2=1.165
r78 10 12 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.31 $Y=1.33
+ $X2=2.31 $Y2=2.075
r79 7 15 37.0704 $w=1.5e-07 $l=2.13014e-07 $layer=POLY_cond $X=2.31 $Y=1 $X2=2.2
+ $Y2=1.165
r80 7 9 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.31 $Y=1 $X2=2.31
+ $Y2=0.56
r81 2 33 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.665 $X2=1.55 $Y2=2
r82 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%A_394_47# 1 2 9 13 17 21 23 24 25 26
+ 30 31
c65 31 0 1.84838e-19 $X=3.11 $Y=1.16
r66 31 34 48.9793 $w=3e-07 $l=1.7e-07 $layer=POLY_cond $X=3.095 $Y=1.16
+ $X2=3.095 $Y2=1.33
r67 31 33 46.9797 $w=3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.095 $Y=1.16
+ $X2=3.095 $Y2=1
r68 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.16 $X2=3.11 $Y2=1.16
r69 28 30 8.8128 $w=3.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.025 $Y=1.42
+ $X2=3.025 $Y2=1.16
r70 27 30 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=3.025 $Y=0.885
+ $X2=3.025 $Y2=1.16
r71 25 28 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.855 $Y=1.505
+ $X2=3.025 $Y2=1.42
r72 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.855 $Y=1.505
+ $X2=2.41 $Y2=1.505
r73 23 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.855 $Y=0.8
+ $X2=3.025 $Y2=0.885
r74 23 24 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.855 $Y=0.8
+ $X2=2.26 $Y2=0.8
r75 19 26 9.06158 $w=1.7e-07 $l=2.79285e-07 $layer=LI1_cond $X=2.17 $Y=1.59
+ $X2=2.41 $Y2=1.505
r76 19 21 10.2165 $w=4.78e-07 $l=4.1e-07 $layer=LI1_cond $X=2.17 $Y=1.59
+ $X2=2.17 $Y2=2
r77 15 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.095 $Y=0.715
+ $X2=2.26 $Y2=0.8
r78 15 17 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.095 $Y=0.715
+ $X2=2.095 $Y2=0.38
r79 13 34 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=3.17 $Y=1.985
+ $X2=3.17 $Y2=1.33
r80 9 33 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.17 $Y=0.445
+ $X2=3.17 $Y2=1
r81 2 21 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=1.97
+ $Y=1.665 $X2=2.095 $Y2=2
r82 1 17 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.095 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
r41 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r43 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.76 $Y2=2.72
r50 25 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.76 $Y2=2.72
r52 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 16 30 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.64 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 16 17 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=2.72 $X2=2.84
+ $Y2=2.72
r57 15 33 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.04 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 15 17 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.04 $Y=2.72 $X2=2.84
+ $Y2=2.72
r59 11 17 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=2.635 $X2=2.84
+ $Y2=2.72
r60 11 13 18.295 $w=3.98e-07 $l=6.35e-07 $layer=LI1_cond $X=2.84 $Y=2.635
+ $X2=2.84 $Y2=2
r61 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.635 $X2=0.76
+ $Y2=2.72
r62 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=2
r63 2 13 300 $w=1.7e-07 $l=6.35807e-07 $layer=licon1_PDIFF $count=2 $X=2.385
+ $Y=1.665 $X2=2.875 $Y2=2
r64 1 9 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.76 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%X 1 2 7 8 9 10 11 12 41 46
r16 30 46 2.45455 $w=3.83e-07 $l=8.2e-08 $layer=LI1_cond $X=3.402 $Y=1.952
+ $X2=3.402 $Y2=1.87
r17 21 41 1.45362 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=3.48 $Y=0.545
+ $X2=3.48 $Y2=0.415
r18 11 46 0.0598672 $w=3.83e-07 $l=2e-09 $layer=LI1_cond $X=3.402 $Y=1.868
+ $X2=3.402 $Y2=1.87
r19 11 44 5.086 $w=3.83e-07 $l=1.08e-07 $layer=LI1_cond $X=3.402 $Y=1.868
+ $X2=3.402 $Y2=1.76
r20 11 12 7.69293 $w=3.83e-07 $l=2.57e-07 $layer=LI1_cond $X=3.402 $Y=1.953
+ $X2=3.402 $Y2=2.21
r21 11 30 0.0299336 $w=3.83e-07 $l=1e-09 $layer=LI1_cond $X=3.402 $Y=1.953
+ $X2=3.402 $Y2=1.952
r22 10 44 11.5244 $w=2.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.48 $Y=1.53
+ $X2=3.48 $Y2=1.76
r23 9 10 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.48 $Y=1.19 $X2=3.48
+ $Y2=1.53
r24 8 9 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.48 $Y=0.85 $X2=3.48
+ $Y2=1.19
r25 7 41 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=3.45 $Y=0.415 $X2=3.48
+ $Y2=0.415
r26 7 37 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=3.45 $Y=0.415
+ $X2=3.385 $Y2=0.415
r27 7 8 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.48 $Y=0.57 $X2=3.48
+ $Y2=0.85
r28 7 21 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.48 $Y=0.57 $X2=3.48
+ $Y2=0.545
r29 2 11 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=3.245
+ $Y=1.485 $X2=3.385 $Y2=2
r30 1 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.385 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r46 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r48 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r49 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r51 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r52 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r53 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 25 37 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.752
+ $Y2=0
r55 25 27 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.15
+ $Y2=0
r56 20 37 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.752
+ $Y2=0
r57 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r58 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r59 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r60 16 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.53
+ $Y2=0
r61 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.875
+ $Y2=0
r62 15 33 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.45
+ $Y2=0
r63 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.875
+ $Y2=0
r64 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r65 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.38
r66 7 37 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0
r67 7 9 10.7927 $w=3.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0.38
r68 2 13 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.235 $X2=2.875 $Y2=0.38
r69 1 9 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.745 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__buf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
M1000 VPWR A a_27_47# VPB phighvt w=790000u l=150000u
+  ad=2.291e+11p pd=2.16e+06u as=2.054e+11p ps=2.1e+06u
M1001 X a_27_47# VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=1.508e+11p ps=1.62e+06u
M1002 X a_27_47# VPWR VPB phighvt w=790000u l=150000u
+  ad=2.054e+11p pd=2.1e+06u as=0p ps=0u
M1003 VGND A a_27_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
.ends


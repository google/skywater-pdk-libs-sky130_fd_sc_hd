* File: sky130_fd_sc_hd__and4b_2.pxi.spice
* Created: Tue Sep  1 18:58:24 2020
* 
x_PM_SKY130_FD_SC_HD__AND4B_2%A_N N_A_N_M1011_g N_A_N_M1006_g A_N A_N A_N
+ N_A_N_c_82_n PM_SKY130_FD_SC_HD__AND4B_2%A_N
x_PM_SKY130_FD_SC_HD__AND4B_2%A_27_413# N_A_27_413#_M1011_d N_A_27_413#_M1006_s
+ N_A_27_413#_c_110_n N_A_27_413#_M1012_g N_A_27_413#_c_111_n
+ N_A_27_413#_c_112_n N_A_27_413#_M1003_g N_A_27_413#_c_117_n
+ N_A_27_413#_c_118_n N_A_27_413#_c_119_n N_A_27_413#_c_113_n
+ N_A_27_413#_c_120_n N_A_27_413#_c_156_p N_A_27_413#_c_114_n
+ PM_SKY130_FD_SC_HD__AND4B_2%A_27_413#
x_PM_SKY130_FD_SC_HD__AND4B_2%B N_B_M1009_g N_B_M1004_g N_B_c_176_n N_B_c_181_n
+ B B B B N_B_c_178_n PM_SKY130_FD_SC_HD__AND4B_2%B
x_PM_SKY130_FD_SC_HD__AND4B_2%C N_C_M1002_g N_C_M1001_g C C C C N_C_c_221_n
+ PM_SKY130_FD_SC_HD__AND4B_2%C
x_PM_SKY130_FD_SC_HD__AND4B_2%D N_D_M1008_g N_D_M1013_g D D D N_D_c_260_n
+ PM_SKY130_FD_SC_HD__AND4B_2%D
x_PM_SKY130_FD_SC_HD__AND4B_2%A_193_413# N_A_193_413#_M1003_s
+ N_A_193_413#_M1012_d N_A_193_413#_M1001_d N_A_193_413#_c_302_n
+ N_A_193_413#_M1005_g N_A_193_413#_M1000_g N_A_193_413#_c_303_n
+ N_A_193_413#_M1007_g N_A_193_413#_M1010_g N_A_193_413#_c_331_n
+ N_A_193_413#_c_309_n N_A_193_413#_c_370_p N_A_193_413#_c_310_n
+ N_A_193_413#_c_311_n N_A_193_413#_c_312_n N_A_193_413#_c_304_n
+ N_A_193_413#_c_329_n N_A_193_413#_c_314_n N_A_193_413#_c_305_n
+ N_A_193_413#_c_306_n PM_SKY130_FD_SC_HD__AND4B_2%A_193_413#
x_PM_SKY130_FD_SC_HD__AND4B_2%VPWR N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_M1013_d
+ N_VPWR_M1010_d N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_418_n
+ VPWR N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n
+ N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_414_n
+ PM_SKY130_FD_SC_HD__AND4B_2%VPWR
x_PM_SKY130_FD_SC_HD__AND4B_2%X N_X_M1005_s N_X_M1000_s X X X X X X N_X_c_490_n
+ X X PM_SKY130_FD_SC_HD__AND4B_2%X
x_PM_SKY130_FD_SC_HD__AND4B_2%VGND N_VGND_M1011_s N_VGND_M1008_d N_VGND_M1007_d
+ N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n
+ VGND N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n N_VGND_c_527_n
+ PM_SKY130_FD_SC_HD__AND4B_2%VGND
cc_1 VNB N_A_N_M1011_g 0.036913f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.0133234f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_A_N_c_82_n 0.0441123f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_413#_c_110_n 0.0437162f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_5 VNB N_A_27_413#_c_111_n 0.0362798f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_6 VNB N_A_27_413#_c_112_n 0.0169133f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_413#_c_113_n 0.00656206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_413#_c_114_n 0.00254319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_M1004_g 0.0335356f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_10 VNB N_B_c_176_n 0.00519761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB B 0.00300494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_178_n 0.022019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_C_M1002_g 0.0285467f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_14 VNB C 0.00448253f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_15 VNB N_C_c_221_n 0.021913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1008_g 0.0283603f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_17 VNB D 0.00388216f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_18 VNB N_D_c_260_n 0.0207071f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_19 VNB N_A_193_413#_c_302_n 0.0172509f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_A_193_413#_c_303_n 0.0189043f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_21 VNB N_A_193_413#_c_304_n 0.00815265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_193_413#_c_305_n 0.00262967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_193_413#_c_306_n 0.0429776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_414_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 0.00832862f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_26 VNB X 0.0225241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_519_n 0.010303f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_28 VNB N_VGND_c_520_n 0.0125358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_521_n 0.00218188f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_30 VNB N_VGND_c_522_n 0.0102396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_523_n 0.0120262f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_524_n 0.0631579f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.16
cc_33 VNB N_VGND_c_525_n 0.0152324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_526_n 0.00506835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_527_n 0.224505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A_N_M1006_g 0.0596584f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_37 VPB A_N 0.016912f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_38 VPB N_A_N_c_82_n 0.0111506f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_39 VPB N_A_27_413#_c_110_n 0.00622168f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_40 VPB N_A_27_413#_M1012_g 0.0549562f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_41 VPB N_A_27_413#_c_117_n 0.00288908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_413#_c_118_n 0.00826823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_413#_c_119_n 0.00848092f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=0.85
cc_44 VPB N_A_27_413#_c_120_n 0.00923161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_413#_c_114_n 4.75249e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_B_M1009_g 0.032991f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_47 VPB N_B_c_176_n 0.0221513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_B_c_181_n 0.0224105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB B 0.00149309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_C_M1001_g 0.0535673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_51 VPB C 0.00532326f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_52 VPB N_C_c_221_n 0.00517217f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_D_M1013_g 0.0497892f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_54 VPB D 0.00397693f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_55 VPB N_D_c_260_n 0.00451149f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_56 VPB N_A_193_413#_M1000_g 0.0186567f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_57 VPB N_A_193_413#_M1010_g 0.0218472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_193_413#_c_309_n 0.0175202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_193_413#_c_310_n 0.00454575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_193_413#_c_311_n 0.00116098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_193_413#_c_312_n 0.0139891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_193_413#_c_304_n 0.0070252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_193_413#_c_314_n 0.00424749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_193_413#_c_305_n 2.35845e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_193_413#_c_306_n 0.00864474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_415_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_67 VPB N_VPWR_c_416_n 0.00212472f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=0.85
cc_68 VPB N_VPWR_c_417_n 0.0101444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_418_n 0.0252587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_419_n 0.0152577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_420_n 0.0150966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_421_n 0.013276f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_422_n 0.00436502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_423_n 0.0171883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_424_n 0.0121855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_425_n 0.00507517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_414_n 0.0449639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB X 0.00959884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB X 0.0112983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 N_A_N_M1011_g N_A_27_413#_c_110_n 0.00780001f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_81 A_N N_A_27_413#_c_110_n 2.59894e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_82 N_A_N_c_82_n N_A_27_413#_c_110_n 0.0208351f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_N_M1006_g N_A_27_413#_M1012_g 0.0381489f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_84 N_A_N_M1006_g N_A_27_413#_c_117_n 0.00258333f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_85 N_A_N_M1006_g N_A_27_413#_c_118_n 0.017202f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_86 N_A_N_c_82_n N_A_27_413#_c_118_n 0.00130998f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_87 A_N N_A_27_413#_c_119_n 0.0132061f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_N_c_82_n N_A_27_413#_c_119_n 9.93381e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_N_M1011_g N_A_27_413#_c_113_n 0.00732262f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_90 A_N N_A_27_413#_c_113_n 0.0130789f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_91 N_A_N_M1006_g N_A_27_413#_c_120_n 0.00698621f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_92 A_N N_A_27_413#_c_120_n 0.0156434f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_93 A_N N_A_27_413#_c_114_n 0.016515f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_94 N_A_N_c_82_n N_A_27_413#_c_114_n 0.00292073f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_N_M1006_g N_VPWR_c_415_n 0.00900519f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_96 N_A_N_M1006_g N_VPWR_c_419_n 0.00348948f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_97 N_A_N_M1006_g N_VPWR_c_414_n 0.00506544f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_98 N_A_N_M1011_g N_VGND_c_520_n 0.0104655f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_99 A_N N_VGND_c_520_n 0.0114029f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A_N_c_82_n N_VGND_c_520_n 0.00256405f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_N_M1011_g N_VGND_c_524_n 0.0046653f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A_N_M1011_g N_VGND_c_527_n 0.00921786f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_103 A_N N_VGND_c_527_n 0.00107484f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A_27_413#_c_110_n N_B_M1004_g 0.00209204f $X=0.89 $Y=1.325 $X2=0 $Y2=0
cc_105 N_A_27_413#_c_112_n N_B_M1004_g 0.0481589f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_106 N_A_27_413#_M1012_g N_B_c_176_n 0.0204888f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_107 N_A_27_413#_c_112_n B 0.00255668f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_108 N_A_27_413#_c_110_n N_B_c_178_n 0.00530766f $X=0.89 $Y=1.325 $X2=0 $Y2=0
cc_109 N_A_27_413#_c_111_n N_B_c_178_n 0.0041805f $X=1.335 $Y=0.805 $X2=0 $Y2=0
cc_110 N_A_27_413#_c_110_n N_A_193_413#_c_312_n 3.57503e-19 $X=0.89 $Y=1.325
+ $X2=0 $Y2=0
cc_111 N_A_27_413#_M1012_g N_A_193_413#_c_312_n 0.00489726f $X=0.89 $Y=2.275
+ $X2=0 $Y2=0
cc_112 N_A_27_413#_c_117_n N_A_193_413#_c_312_n 0.00187617f $X=0.26 $Y=2.3 $X2=0
+ $Y2=0
cc_113 N_A_27_413#_c_118_n N_A_193_413#_c_312_n 0.0127772f $X=0.635 $Y=1.915
+ $X2=0 $Y2=0
cc_114 N_A_27_413#_c_120_n N_A_193_413#_c_312_n 0.0114902f $X=0.72 $Y=1.83 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_c_110_n N_A_193_413#_c_304_n 0.00442216f $X=0.89 $Y=1.325
+ $X2=0 $Y2=0
cc_116 N_A_27_413#_M1012_g N_A_193_413#_c_304_n 0.0030512f $X=0.89 $Y=2.275
+ $X2=0 $Y2=0
cc_117 N_A_27_413#_c_111_n N_A_193_413#_c_304_n 0.0139149f $X=1.335 $Y=0.805
+ $X2=0 $Y2=0
cc_118 N_A_27_413#_c_112_n N_A_193_413#_c_304_n 0.00253797f $X=1.41 $Y=0.73
+ $X2=0 $Y2=0
cc_119 N_A_27_413#_c_113_n N_A_193_413#_c_304_n 0.0182501f $X=0.72 $Y=0.995
+ $X2=0 $Y2=0
cc_120 N_A_27_413#_c_120_n N_A_193_413#_c_304_n 0.0155437f $X=0.72 $Y=1.83 $X2=0
+ $Y2=0
cc_121 N_A_27_413#_c_114_n N_A_193_413#_c_304_n 0.0248276f $X=0.89 $Y=1.16 $X2=0
+ $Y2=0
cc_122 N_A_27_413#_c_111_n N_A_193_413#_c_329_n 0.00187101f $X=1.335 $Y=0.805
+ $X2=0 $Y2=0
cc_123 N_A_27_413#_c_156_p N_A_193_413#_c_329_n 0.0167624f $X=0.68 $Y=0.42 $X2=0
+ $Y2=0
cc_124 N_A_27_413#_M1012_g N_VPWR_c_415_n 0.00959643f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_125 N_A_27_413#_c_118_n N_VPWR_c_415_n 0.0172745f $X=0.635 $Y=1.915 $X2=0
+ $Y2=0
cc_126 N_A_27_413#_c_117_n N_VPWR_c_419_n 0.0115478f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_127 N_A_27_413#_c_118_n N_VPWR_c_419_n 0.00237804f $X=0.635 $Y=1.915 $X2=0
+ $Y2=0
cc_128 N_A_27_413#_M1012_g N_VPWR_c_423_n 0.0046653f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_129 N_A_27_413#_M1012_g N_VPWR_c_424_n 9.4904e-19 $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_130 N_A_27_413#_M1006_s N_VPWR_c_414_n 0.00374845f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_131 N_A_27_413#_M1012_g N_VPWR_c_414_n 0.00833373f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_132 N_A_27_413#_c_117_n N_VPWR_c_414_n 0.00645836f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_133 N_A_27_413#_c_118_n N_VPWR_c_414_n 0.00516132f $X=0.635 $Y=1.915 $X2=0
+ $Y2=0
cc_134 N_A_27_413#_c_110_n N_VGND_c_524_n 0.00424743f $X=0.89 $Y=1.325 $X2=0
+ $Y2=0
cc_135 N_A_27_413#_c_111_n N_VGND_c_524_n 7.2576e-19 $X=1.335 $Y=0.805 $X2=0
+ $Y2=0
cc_136 N_A_27_413#_c_112_n N_VGND_c_524_n 0.00585385f $X=1.41 $Y=0.73 $X2=0
+ $Y2=0
cc_137 N_A_27_413#_c_156_p N_VGND_c_524_n 0.0143008f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_138 N_A_27_413#_M1011_d N_VGND_c_527_n 0.00382094f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_139 N_A_27_413#_c_110_n N_VGND_c_527_n 0.0059814f $X=0.89 $Y=1.325 $X2=0
+ $Y2=0
cc_140 N_A_27_413#_c_112_n N_VGND_c_527_n 0.0119273f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_141 N_A_27_413#_c_156_p N_VGND_c_527_n 0.00798371f $X=0.68 $Y=0.42 $X2=0
+ $Y2=0
cc_142 N_B_M1004_g N_C_M1002_g 0.0297441f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_143 B N_C_M1002_g 4.65335e-19 $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_144 N_B_M1009_g N_C_M1001_g 0.00964675f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_145 N_B_c_176_n N_C_M1001_g 0.0117015f $X=1.62 $Y=1.56 $X2=0 $Y2=0
cc_146 B N_C_M1001_g 5.77957e-19 $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_147 N_B_M1004_g C 0.00628598f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_148 N_B_c_176_n C 0.00387319f $X=1.62 $Y=1.56 $X2=0 $Y2=0
cc_149 B C 0.0814825f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_150 N_B_M1004_g N_C_c_221_n 0.0149995f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_151 N_B_c_176_n N_C_c_221_n 0.00424512f $X=1.62 $Y=1.56 $X2=0 $Y2=0
cc_152 B N_C_c_221_n 3.08294e-19 $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_153 N_B_M1009_g N_A_193_413#_c_331_n 0.00520411f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_154 N_B_M1009_g N_A_193_413#_c_309_n 0.015361f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_155 N_B_c_181_n N_A_193_413#_c_309_n 0.00363902f $X=1.62 $Y=1.745 $X2=0 $Y2=0
cc_156 B N_A_193_413#_c_309_n 0.017201f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_157 N_B_c_178_n N_A_193_413#_c_309_n 9.86952e-19 $X=1.66 $Y=1.24 $X2=0 $Y2=0
cc_158 N_B_M1009_g N_A_193_413#_c_312_n 3.29239e-19 $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_159 N_B_c_181_n N_A_193_413#_c_312_n 0.00547938f $X=1.62 $Y=1.745 $X2=0 $Y2=0
cc_160 N_B_M1004_g N_A_193_413#_c_304_n 7.04111e-19 $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_161 B N_A_193_413#_c_304_n 0.0690634f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_162 N_B_c_178_n N_A_193_413#_c_304_n 0.00547938f $X=1.66 $Y=1.24 $X2=0 $Y2=0
cc_163 N_B_M1009_g N_VPWR_c_415_n 9.24705e-19 $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_164 N_B_M1009_g N_VPWR_c_423_n 0.00339367f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_165 N_B_M1009_g N_VPWR_c_424_n 0.0100242f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_166 N_B_M1009_g N_VPWR_c_414_n 0.00443034f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_167 N_B_M1004_g N_VGND_c_524_n 0.0052149f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_168 B N_VGND_c_524_n 0.00613012f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_169 N_B_M1004_g N_VGND_c_527_n 0.00913542f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_170 B N_VGND_c_527_n 0.00739098f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_171 B A_297_47# 0.00129203f $X=1.53 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_172 N_C_M1002_g N_D_M1008_g 0.0366266f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_173 C N_D_M1008_g 0.00140998f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_174 N_C_M1001_g N_D_M1013_g 0.0334585f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_175 C N_D_M1013_g 6.66164e-19 $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_176 N_C_M1002_g D 0.00662674f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_177 C D 0.07641f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_178 C N_D_c_260_n 2.98688e-19 $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_179 N_C_c_221_n N_D_c_260_n 0.0202358f $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_180 N_C_M1001_g N_A_193_413#_c_309_n 0.0143045f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_181 C N_A_193_413#_c_309_n 0.0213768f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_182 N_C_c_221_n N_A_193_413#_c_309_n 4.56204e-19 $X=2.19 $Y=1.16 $X2=0 $Y2=0
cc_183 N_C_M1001_g N_A_193_413#_c_314_n 0.00703405f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_184 N_C_M1001_g N_VPWR_c_420_n 0.00339367f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_185 N_C_M1001_g N_VPWR_c_424_n 0.00818188f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_186 N_C_M1001_g N_VPWR_c_414_n 0.00406251f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_187 N_C_M1002_g N_VGND_c_521_n 0.0020428f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_188 C N_VGND_c_521_n 0.00143341f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_189 N_C_M1002_g N_VGND_c_524_n 0.00482371f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_190 C N_VGND_c_524_n 0.00953851f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_191 N_C_M1002_g N_VGND_c_527_n 0.00828276f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_192 C N_VGND_c_527_n 0.0105691f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_193 C A_369_47# 0.00524479f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_194 N_D_M1008_g N_A_193_413#_c_302_n 0.0231915f $X=2.715 $Y=0.445 $X2=0 $Y2=0
cc_195 D N_A_193_413#_c_302_n 0.00130937f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_196 N_D_M1013_g N_A_193_413#_M1000_g 0.0327523f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_197 D N_A_193_413#_M1000_g 2.85909e-19 $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_198 N_D_M1013_g N_A_193_413#_c_310_n 0.0126199f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_199 D N_A_193_413#_c_310_n 0.0123479f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_200 N_D_c_260_n N_A_193_413#_c_310_n 5.96205e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_201 N_D_M1013_g N_A_193_413#_c_311_n 0.00559596f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_202 D N_A_193_413#_c_311_n 0.0177517f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_203 N_D_M1013_g N_A_193_413#_c_314_n 0.00302849f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_204 D N_A_193_413#_c_314_n 0.0146459f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_205 N_D_c_260_n N_A_193_413#_c_314_n 2.273e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_206 D N_A_193_413#_c_305_n 0.0210882f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_207 N_D_c_260_n N_A_193_413#_c_305_n 0.00197118f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_208 D N_A_193_413#_c_306_n 3.50639e-19 $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_209 N_D_c_260_n N_A_193_413#_c_306_n 0.0204413f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_210 N_D_M1013_g N_VPWR_c_416_n 0.00165619f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_211 N_D_M1013_g N_VPWR_c_420_n 0.00441875f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_212 N_D_M1013_g N_VPWR_c_424_n 5.48685e-19 $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_213 N_D_M1013_g N_VPWR_c_414_n 0.00621224f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_214 D X 0.00609194f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_215 N_D_M1008_g N_X_c_490_n 0.00113119f $X=2.715 $Y=0.445 $X2=0 $Y2=0
cc_216 D X 0.00501139f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_217 N_D_M1008_g N_VGND_c_521_n 0.0101411f $X=2.715 $Y=0.445 $X2=0 $Y2=0
cc_218 D N_VGND_c_521_n 9.76265e-19 $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_219 N_D_M1008_g N_VGND_c_524_n 0.00340417f $X=2.715 $Y=0.445 $X2=0 $Y2=0
cc_220 D N_VGND_c_524_n 0.00523343f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_221 N_D_M1008_g N_VGND_c_527_n 0.00409563f $X=2.715 $Y=0.445 $X2=0 $Y2=0
cc_222 D N_VGND_c_527_n 0.00886174f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_223 D A_469_47# 0.00261754f $X=2.45 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_224 N_A_193_413#_c_309_n N_VPWR_M1009_d 0.00534726f $X=2.44 $Y=2 $X2=0 $Y2=0
cc_225 N_A_193_413#_c_310_n N_VPWR_M1013_d 0.00652168f $X=2.995 $Y=1.88 $X2=0
+ $Y2=0
cc_226 N_A_193_413#_c_311_n N_VPWR_M1013_d 0.00330702f $X=3.08 $Y=1.795 $X2=0
+ $Y2=0
cc_227 N_A_193_413#_M1000_g N_VPWR_c_416_n 0.00735045f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_193_413#_M1010_g N_VPWR_c_416_n 5.16112e-19 $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_193_413#_c_310_n N_VPWR_c_416_n 0.0157062f $X=2.995 $Y=1.88 $X2=0
+ $Y2=0
cc_230 N_A_193_413#_M1000_g N_VPWR_c_418_n 5.91467e-19 $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_193_413#_M1010_g N_VPWR_c_418_n 0.0114227f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_193_413#_c_309_n N_VPWR_c_420_n 0.00317671f $X=2.44 $Y=2 $X2=0 $Y2=0
cc_233 N_A_193_413#_c_370_p N_VPWR_c_420_n 0.0115924f $X=2.525 $Y=2.3 $X2=0
+ $Y2=0
cc_234 N_A_193_413#_c_310_n N_VPWR_c_420_n 0.00302941f $X=2.995 $Y=1.88 $X2=0
+ $Y2=0
cc_235 N_A_193_413#_M1000_g N_VPWR_c_421_n 0.0046653f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_193_413#_M1010_g N_VPWR_c_421_n 0.0046653f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_193_413#_c_331_n N_VPWR_c_423_n 0.0116048f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_238 N_A_193_413#_c_309_n N_VPWR_c_423_n 0.0036143f $X=2.44 $Y=2 $X2=0 $Y2=0
cc_239 N_A_193_413#_c_312_n N_VPWR_c_423_n 0.00249276f $X=1.165 $Y=2 $X2=0 $Y2=0
cc_240 N_A_193_413#_c_331_n N_VPWR_c_424_n 0.00898144f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_241 N_A_193_413#_c_309_n N_VPWR_c_424_n 0.0418204f $X=2.44 $Y=2 $X2=0 $Y2=0
cc_242 N_A_193_413#_c_370_p N_VPWR_c_424_n 0.0136736f $X=2.525 $Y=2.3 $X2=0
+ $Y2=0
cc_243 N_A_193_413#_M1012_d N_VPWR_c_414_n 0.00641078f $X=0.965 $Y=2.065 $X2=0
+ $Y2=0
cc_244 N_A_193_413#_M1001_d N_VPWR_c_414_n 0.00310578f $X=2.345 $Y=2.065 $X2=0
+ $Y2=0
cc_245 N_A_193_413#_M1000_g N_VPWR_c_414_n 0.00798194f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_246 N_A_193_413#_M1010_g N_VPWR_c_414_n 0.00798194f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_193_413#_c_331_n N_VPWR_c_414_n 0.00646998f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_248 N_A_193_413#_c_309_n N_VPWR_c_414_n 0.0146105f $X=2.44 $Y=2 $X2=0 $Y2=0
cc_249 N_A_193_413#_c_370_p N_VPWR_c_414_n 0.00646745f $X=2.525 $Y=2.3 $X2=0
+ $Y2=0
cc_250 N_A_193_413#_c_310_n N_VPWR_c_414_n 0.00654502f $X=2.995 $Y=1.88 $X2=0
+ $Y2=0
cc_251 N_A_193_413#_c_312_n N_VPWR_c_414_n 0.00388138f $X=1.165 $Y=2 $X2=0 $Y2=0
cc_252 N_A_193_413#_c_302_n X 0.00709144f $X=3.215 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_193_413#_c_303_n X 0.0119163f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_193_413#_c_306_n X 0.00194336f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_193_413#_M1010_g X 0.0160638f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A_193_413#_c_306_n X 0.00191553f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_193_413#_c_302_n N_X_c_490_n 0.00607657f $X=3.215 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A_193_413#_c_302_n X 0.00234616f $X=3.215 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_193_413#_M1000_g X 0.00178368f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_193_413#_c_303_n X 0.00719617f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_193_413#_M1010_g X 0.00890955f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A_193_413#_c_311_n X 0.0120832f $X=3.08 $Y=1.795 $X2=0 $Y2=0
cc_263 N_A_193_413#_c_305_n X 0.0255867f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_193_413#_c_306_n X 0.0250729f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_193_413#_c_302_n N_VGND_c_521_n 0.00279623f $X=3.215 $Y=0.995 $X2=0
+ $Y2=0
cc_266 N_A_193_413#_c_305_n N_VGND_c_521_n 0.00319889f $X=3.17 $Y=1.16 $X2=0
+ $Y2=0
cc_267 N_A_193_413#_c_306_n N_VGND_c_521_n 9.49739e-19 $X=3.67 $Y=1.16 $X2=0
+ $Y2=0
cc_268 N_A_193_413#_c_302_n N_VGND_c_523_n 4.73778e-19 $X=3.215 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A_193_413#_c_303_n N_VGND_c_523_n 0.0080377f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A_193_413#_c_329_n N_VGND_c_524_n 0.0139021f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_271 N_A_193_413#_c_302_n N_VGND_c_525_n 0.00541359f $X=3.215 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A_193_413#_c_303_n N_VGND_c_525_n 0.00339835f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_273 N_A_193_413#_M1003_s N_VGND_c_527_n 0.00256467f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_274 N_A_193_413#_c_302_n N_VGND_c_527_n 0.00988683f $X=3.215 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A_193_413#_c_303_n N_VGND_c_527_n 0.00404195f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_A_193_413#_c_329_n N_VGND_c_527_n 0.00836197f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_414_n N_X_M1000_s 0.00590463f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_421_n X 0.013857f $X=3.715 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_414_n X 0.00781789f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_M1010_d X 0.00317633f $X=3.745 $Y=1.485 $X2=0 $Y2=0
cc_281 N_VPWR_c_418_n X 0.0248381f $X=3.88 $Y=2 $X2=0 $Y2=0
cc_282 N_VPWR_M1010_d X 2.16973e-19 $X=3.745 $Y=1.485 $X2=0 $Y2=0
cc_283 X N_VGND_M1007_d 0.00300766f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_284 X N_VGND_M1007_d 2.61253e-19 $X=3.905 $Y=0.85 $X2=0 $Y2=0
cc_285 X N_VGND_c_523_n 0.0226502f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_286 X N_VGND_c_525_n 0.00260571f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_287 N_X_c_490_n N_VGND_c_525_n 0.0175166f $X=3.46 $Y=0.42 $X2=0 $Y2=0
cc_288 N_X_M1005_s N_VGND_c_527_n 0.00260662f $X=3.29 $Y=0.235 $X2=0 $Y2=0
cc_289 X N_VGND_c_527_n 0.00638723f $X=3.82 $Y=0.765 $X2=0 $Y2=0
cc_290 N_X_c_490_n N_VGND_c_527_n 0.0106652f $X=3.46 $Y=0.42 $X2=0 $Y2=0
cc_291 N_VGND_c_527_n A_297_47# 0.00326666f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_292 N_VGND_c_527_n A_369_47# 0.00705492f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_293 N_VGND_c_527_n A_469_47# 0.00660809f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a31o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 1.705000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725000 1.075000 1.055000 1.245000 ;
        RECT 0.805000 0.735000 2.170000 0.905000 ;
        RECT 0.805000 0.905000 0.975000 1.075000 ;
        RECT 1.985000 0.905000 2.170000 1.075000 ;
        RECT 1.985000 1.075000 2.315000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.525000 1.445000 ;
        RECT 0.150000 1.445000 2.855000 1.615000 ;
        RECT 2.525000 1.075000 2.855000 1.445000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.575000 1.075000 4.030000 1.285000 ;
        RECT 3.815000 0.745000 4.030000 1.075000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505000 0.655000 6.295000 0.825000 ;
        RECT 4.535000 1.785000 6.295000 1.955000 ;
        RECT 4.595000 1.955000 4.765000 2.465000 ;
        RECT 5.435000 1.955000 5.605000 2.465000 ;
        RECT 6.125000 0.825000 6.295000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.175000  0.085000 0.345000 0.905000 ;
        RECT 2.700000  0.085000 2.985000 0.530000 ;
        RECT 3.735000  0.085000 4.265000 0.565000 ;
        RECT 4.935000  0.085000 5.265000 0.485000 ;
        RECT 5.775000  0.085000 6.105000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.515000 2.125000 0.845000 2.635000 ;
        RECT 1.355000 2.125000 1.685000 2.635000 ;
        RECT 2.195000 2.125000 2.525000 2.635000 ;
        RECT 4.095000 2.125000 4.425000 2.635000 ;
        RECT 4.935000 2.125000 5.265000 2.635000 ;
        RECT 5.775000 2.125000 6.105000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 1.785000 2.985000 1.955000 ;
      RECT 0.175000 1.955000 0.345000 2.465000 ;
      RECT 1.015000 1.955000 1.185000 2.465000 ;
      RECT 1.355000 0.395000 2.520000 0.565000 ;
      RECT 1.855000 1.955000 2.025000 2.465000 ;
      RECT 2.350000 0.565000 2.520000 0.700000 ;
      RECT 2.350000 0.700000 3.485000 0.805000 ;
      RECT 2.350000 0.805000 3.345000 0.870000 ;
      RECT 2.815000 1.955000 2.985000 2.295000 ;
      RECT 2.815000 2.295000 3.825000 2.465000 ;
      RECT 3.155000 0.295000 3.485000 0.700000 ;
      RECT 3.155000 0.870000 3.345000 1.455000 ;
      RECT 3.155000 1.455000 4.395000 1.625000 ;
      RECT 3.155000 1.625000 3.485000 2.115000 ;
      RECT 3.655000 1.795000 3.825000 2.295000 ;
      RECT 4.225000 0.995000 5.935000 1.325000 ;
      RECT 4.225000 1.325000 4.395000 1.455000 ;
  END
END sky130_fd_sc_hd__a31o_4

* NGSPICE file created from sky130_fd_sc_hd__o22a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=8.775e+11p ps=9.2e+06u
M1001 a_96_21# B2 a_484_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=9.165e+11p ps=9.32e+06u
M1002 a_918_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=1.975e+12p ps=1.395e+07u
M1003 VPWR a_96_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.4e+11p ps=5.08e+06u
M1004 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_96_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_96_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_96_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_918_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_566_297# B2 a_96_21# VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=5.4e+11p ps=5.08e+06u
M1010 a_96_21# B2 a_566_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_918_297# A2 a_96_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_484_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_566_297# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_484_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_484_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_484_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_96_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_484_47# B2 a_96_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_96_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_96_21# A2 a_918_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR B1 a_566_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_96_21# B1 a_484_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_484_47# B1 a_96_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


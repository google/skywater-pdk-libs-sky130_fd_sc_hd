* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_226_47# A2_N a_226_297# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_76_199# a_226_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=6.266e+11p ps=5.69e+06u
M1002 a_489_413# a_226_47# a_76_199# VPB phighvt w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=1.092e+11p ps=1.36e+06u
M1003 VGND B1 a_556_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1004 a_556_47# B2 a_76_199# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_76_199# X VPB phighvt w=1e+06u l=150000u
+  ad=4.469e+11p pd=4.25e+06u as=2.6e+11p ps=2.52e+06u
M1006 a_489_413# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2_N a_226_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1008 VPWR B2 a_489_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_226_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_226_297# A1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_76_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
.ends


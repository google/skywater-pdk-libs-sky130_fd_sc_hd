* File: sky130_fd_sc_hd__nand4_4.spice.pex
* Created: Thu Aug 27 14:30:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4_4%D 3 7 11 15 19 23 25 27 31 33 34 35 36
c80 36 0 1.88146e-19 $X=1.615 $Y=1.19
c81 27 0 1.09605e-19 $X=1.73 $Y=0.56
r82 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r83 42 44 34.1782 $w=2.75e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r84 36 49 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.52 $Y2=1.175
r85 35 49 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.52 $Y2=1.175
r86 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.155 $Y2=1.175
r87 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r88 33 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r89 25 48 36.8073 $w=2.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.52 $Y2=1.16
r90 25 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r91 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r92 17 48 36.8073 $w=2.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r93 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r94 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r95 9 17 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r96 9 44 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.47 $Y2=1.16
r97 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r98 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r99 5 44 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r100 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.985
r101 1 44 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r102 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%C 3 7 11 15 19 23 27 31 33 34 35 36 51
c80 51 0 1.88146e-19 $X=3.41 $Y=1.16
r81 49 51 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=3.2 $Y=1.16 $X2=3.41
+ $Y2=1.16
r82 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.16 $X2=3.2 $Y2=1.16
r83 47 49 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.99 $Y=1.16 $X2=3.2
+ $Y2=1.16
r84 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16 $X2=2.99
+ $Y2=1.16
r85 44 46 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=2.355 $Y=1.16
+ $X2=2.57 $Y2=1.16
r86 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.355
+ $Y=1.16 $X2=2.355 $Y2=1.16
r87 41 44 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.355 $Y2=1.16
r88 36 50 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=3.455 $Y=1.175
+ $X2=3.2 $Y2=1.175
r89 35 50 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=3.2 $Y2=1.175
r90 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.995 $Y2=1.175
r91 34 45 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.355 $Y2=1.175
r92 33 45 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=2.355 $Y2=1.175
r93 29 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r94 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r95 25 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r96 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r97 21 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r98 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r99 17 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r100 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r101 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r102 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r103 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r104 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r105 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r106 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r107 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r108 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%B 3 7 11 15 19 23 27 31 33 34 35 36 41 52
r80 50 52 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=5.4 $Y=1.16 $X2=5.61
+ $Y2=1.16
r81 48 50 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=5.19 $Y=1.16 $X2=5.4
+ $Y2=1.16
r82 47 48 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.16 $X2=5.19
+ $Y2=1.16
r83 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.35 $Y=1.16 $X2=4.77
+ $Y2=1.16
r84 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.11
+ $Y=1.16 $X2=4.11 $Y2=1.16
r85 41 46 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.275 $Y=1.16
+ $X2=4.35 $Y2=1.16
r86 41 43 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.275 $Y=1.16
+ $X2=4.11 $Y2=1.16
r87 36 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.4 $Y=1.16
+ $X2=5.4 $Y2=1.16
r88 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.855 $Y=1.175
+ $X2=5.315 $Y2=1.175
r89 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.855 $Y2=1.175
r90 34 44 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.11 $Y2=1.175
r91 33 44 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=4.11 $Y2=1.175
r92 29 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.16
r93 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.985
r94 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=1.16
r95 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=0.56
r96 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.16
r97 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.985
r98 17 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=1.16
r99 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=0.56
r100 13 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.16
r101 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.985
r102 9 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=1.16
r103 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=0.56
r104 5 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.16
r105 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.985
r106 1 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=1.16
r107 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%A 3 7 11 15 19 23 27 31 33 34 35 45
c80 45 0 1.93124e-19 $X=7.35 $Y=1.16
r81 45 47 34.1782 $w=2.75e-07 $l=1.95e-07 $layer=POLY_cond $X=7.35 $Y=1.16
+ $X2=7.545 $Y2=1.16
r82 35 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.545
+ $Y=1.16 $X2=7.545 $Y2=1.16
r83 34 35 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=7.125 $Y=1.175
+ $X2=7.545 $Y2=1.175
r84 33 34 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=6.63 $Y=1.175
+ $X2=7.125 $Y2=1.175
r85 33 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.63
+ $Y=1.16 $X2=6.63 $Y2=1.16
r86 29 45 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.35 $Y=1.305
+ $X2=7.35 $Y2=1.16
r87 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.35 $Y=1.305
+ $X2=7.35 $Y2=1.985
r88 25 45 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.35 $Y=1.015
+ $X2=7.35 $Y2=1.16
r89 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.35 $Y=1.015
+ $X2=7.35 $Y2=0.56
r90 17 45 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=6.93 $Y=1.16
+ $X2=7.35 $Y2=1.16
r91 17 42 52.5818 $w=2.75e-07 $l=3e-07 $layer=POLY_cond $X=6.93 $Y=1.16 $X2=6.63
+ $Y2=1.16
r92 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.93 $Y=1.295
+ $X2=6.93 $Y2=1.985
r93 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.93 $Y=1.025
+ $X2=6.93 $Y2=0.56
r94 9 42 21.0327 $w=2.75e-07 $l=1.2e-07 $layer=POLY_cond $X=6.51 $Y=1.16
+ $X2=6.63 $Y2=1.16
r95 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.51 $Y=1.295
+ $X2=6.51 $Y2=1.985
r96 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.51 $Y=1.025
+ $X2=6.51 $Y2=0.56
r97 1 9 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=6.09 $Y=1.16 $X2=6.51
+ $Y2=1.16
r98 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.09 $Y=1.295 $X2=6.09
+ $Y2=1.985
r99 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.09 $Y=1.025
+ $X2=6.09 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 40 44 48 52
+ 56 58 62 64 66 71 72 74 75 77 78 80 81 82 83 84 96 107 116 119 123
r124 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r125 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r126 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r127 111 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r128 111 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r129 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r130 108 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=6.72 $Y2=2.72
r131 108 110 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=7.13 $Y2=2.72
r132 107 122 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=7.475 $Y=2.72
+ $X2=7.647 $Y2=2.72
r133 107 110 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.475 $Y=2.72
+ $X2=7.13 $Y2=2.72
r134 106 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r135 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r136 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r137 103 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r138 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r139 100 116 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=3.88 $Y2=2.72
r140 100 102 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.83 $Y2=2.72
r141 99 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r142 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r143 96 116 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.88 $Y2=2.72
r144 96 98 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.72
+ $X2=3.45 $Y2=2.72
r145 95 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r146 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r147 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r148 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r149 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r150 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 86 113 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r152 86 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r153 84 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 84 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 82 105 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=5.77 $Y=2.72
+ $X2=5.75 $Y2=2.72
r156 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.77 $Y=2.72
+ $X2=5.855 $Y2=2.72
r157 80 102 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.83 $Y2=2.72
r158 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.98 $Y2=2.72
r159 79 105 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=5.75 $Y2=2.72
r160 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=4.98 $Y2=2.72
r161 77 94 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.53 $Y2=2.72
r162 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.78 $Y2=2.72
r163 76 98 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.45 $Y2=2.72
r164 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.78 $Y2=2.72
r165 74 91 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r166 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.94 $Y2=2.72
r167 73 94 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.53 $Y2=2.72
r168 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.94 $Y2=2.72
r169 71 88 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r170 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r171 70 91 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r172 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r173 66 69 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=7.605 $Y=1.66
+ $X2=7.605 $Y2=2.34
r174 64 122 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=7.605 $Y=2.635
+ $X2=7.647 $Y2=2.72
r175 64 69 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=7.605 $Y=2.635
+ $X2=7.605 $Y2=2.34
r176 60 119 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.72 $Y=2.635
+ $X2=6.72 $Y2=2.72
r177 60 62 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.72 $Y=2.635
+ $X2=6.72 $Y2=2
r178 59 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.72
+ $X2=5.855 $Y2=2.72
r179 58 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.635 $Y=2.72
+ $X2=6.72 $Y2=2.72
r180 58 59 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.635 $Y=2.72
+ $X2=5.94 $Y2=2.72
r181 54 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.855 $Y=2.635
+ $X2=5.855 $Y2=2.72
r182 54 56 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.855 $Y=2.635
+ $X2=5.855 $Y2=2
r183 50 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r184 50 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2
r185 46 116 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.72
r186 46 48 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2
r187 42 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r188 42 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r189 38 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r190 38 40 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r191 34 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r192 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r193 30 33 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r194 28 113 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r195 28 33 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r196 9 69 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.425
+ $Y=1.485 $X2=7.56 $Y2=2.34
r197 9 66 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.425
+ $Y=1.485 $X2=7.56 $Y2=1.66
r198 8 62 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.585
+ $Y=1.485 $X2=6.72 $Y2=2
r199 7 56 300 $w=1.7e-07 $l=5.93949e-07 $layer=licon1_PDIFF $count=2 $X=5.685
+ $Y=1.485 $X2=5.855 $Y2=2
r200 6 52 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2
r201 5 48 150 $w=1.7e-07 $l=8.75414e-07 $layer=licon1_PDIFF $count=4 $X=3.485
+ $Y=1.485 $X2=4.14 $Y2=2
r202 4 44 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r203 3 40 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r204 2 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r205 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r206 1 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%Y 1 2 3 4 5 6 7 8 9 10 31 33 35 39 41 45 47
+ 51 53 57 59 63 65 69 71 75 77 79 81 86 88 90 92 94 98 101
r172 96 101 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=6.2 $Y=1.445
+ $X2=6.2 $Y2=1.19
r173 96 98 2.61222 $w=1.8e-07 $l=1.47207e-07 $layer=LI1_cond $X=6.2 $Y=1.445
+ $X2=6.287 $Y2=1.555
r174 95 101 17.5606 $w=1.78e-07 $l=2.85e-07 $layer=LI1_cond $X=6.2 $Y=0.905
+ $X2=6.2 $Y2=1.19
r175 79 100 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=7.14 $Y=1.665
+ $X2=7.14 $Y2=1.555
r176 79 81 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.14 $Y=1.665
+ $X2=7.14 $Y2=2.34
r177 78 98 3.51191 $w=2.2e-07 $l=1.78e-07 $layer=LI1_cond $X=6.465 $Y=1.555
+ $X2=6.287 $Y2=1.555
r178 77 100 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=1.555
+ $X2=7.14 $Y2=1.555
r179 77 78 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=6.975 $Y=1.555
+ $X2=6.465 $Y2=1.555
r180 73 75 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=6.3 $Y=0.78
+ $X2=7.14 $Y2=0.78
r181 71 95 7.0541 $w=2.5e-07 $l=1.63936e-07 $layer=LI1_cond $X=6.29 $Y=0.78
+ $X2=6.2 $Y2=0.905
r182 71 73 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=6.29 $Y=0.78 $X2=6.3
+ $Y2=0.78
r183 67 98 2.61222 $w=3.3e-07 $l=1.16319e-07 $layer=LI1_cond $X=6.3 $Y=1.665
+ $X2=6.287 $Y2=1.555
r184 67 69 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.3 $Y=1.665
+ $X2=6.3 $Y2=2.34
r185 66 94 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=1.555
+ $X2=5.4 $Y2=1.555
r186 65 98 3.51191 $w=2.2e-07 $l=1.77e-07 $layer=LI1_cond $X=6.11 $Y=1.555
+ $X2=6.287 $Y2=1.555
r187 65 66 28.5492 $w=2.18e-07 $l=5.45e-07 $layer=LI1_cond $X=6.11 $Y=1.555
+ $X2=5.565 $Y2=1.555
r188 61 94 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=5.4 $Y=1.665
+ $X2=5.4 $Y2=1.555
r189 61 63 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.4 $Y=1.665
+ $X2=5.4 $Y2=2.34
r190 60 92 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=1.555
+ $X2=4.56 $Y2=1.555
r191 59 94 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=1.555
+ $X2=5.4 $Y2=1.555
r192 59 60 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=5.235 $Y=1.555
+ $X2=4.725 $Y2=1.555
r193 55 92 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.555
r194 55 57 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=2.34
r195 54 90 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=1.555
+ $X2=3.2 $Y2=1.555
r196 53 92 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.555
+ $X2=4.56 $Y2=1.555
r197 53 54 53.9553 $w=2.18e-07 $l=1.03e-06 $layer=LI1_cond $X=4.395 $Y=1.555
+ $X2=3.365 $Y2=1.555
r198 49 90 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.2 $Y=1.665
+ $X2=3.2 $Y2=1.555
r199 49 51 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.2 $Y=1.665
+ $X2=3.2 $Y2=2.34
r200 48 88 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=1.555
+ $X2=2.36 $Y2=1.555
r201 47 90 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=1.555
+ $X2=3.2 $Y2=1.555
r202 47 48 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=3.035 $Y=1.555
+ $X2=2.525 $Y2=1.555
r203 43 88 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=1.555
r204 43 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.36 $Y=1.665
+ $X2=2.36 $Y2=2.34
r205 42 86 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.555
+ $X2=1.52 $Y2=1.555
r206 41 88 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=2.36 $Y2=1.555
r207 41 42 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=2.195 $Y=1.555
+ $X2=1.685 $Y2=1.555
r208 37 86 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.555
r209 37 39 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r210 36 84 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.555
+ $X2=0.68 $Y2=1.555
r211 35 86 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=1.52 $Y2=1.555
r212 35 36 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.555
+ $X2=0.845 $Y2=1.555
r213 31 84 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.555
r214 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r215 10 100 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.005
+ $Y=1.485 $X2=7.14 $Y2=1.66
r216 10 81 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.005
+ $Y=1.485 $X2=7.14 $Y2=2.34
r217 9 98 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.165
+ $Y=1.485 $X2=6.3 $Y2=1.66
r218 9 69 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.165
+ $Y=1.485 $X2=6.3 $Y2=2.34
r219 8 94 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.66
r220 8 63 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=2.34
r221 7 92 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.66
r222 7 57 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2.34
r223 6 90 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.66
r224 6 51 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.34
r225 5 88 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.66
r226 5 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.34
r227 4 86 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r228 4 39 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r229 3 84 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r230 3 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r231 2 75 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=7.005
+ $Y=0.235 $X2=7.14 $Y2=0.74
r232 1 73 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=6.165
+ $Y=0.235 $X2=6.3 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%A_27_47# 1 2 3 4 5 16 19 20 21 24 30 34 36
r57 32 34 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=0.37
+ $X2=3.62 $Y2=0.37
r58 30 32 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.37
+ $X2=2.78 $Y2=0.37
r59 27 29 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.94 $Y=0.655 $X2=1.94
+ $Y2=0.625
r60 26 30 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.94 $Y=0.485
+ $X2=2.025 $Y2=0.37
r61 26 29 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.94 $Y=0.485
+ $X2=1.94 $Y2=0.625
r62 25 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.78 $X2=1.1
+ $Y2=0.78
r63 24 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.855 $Y=0.78
+ $X2=1.94 $Y2=0.655
r64 24 25 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=0.78
+ $X2=1.185 $Y2=0.78
r65 21 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.1 $Y=0.655 $X2=1.1
+ $Y2=0.78
r66 21 23 2.15294 $w=1.7e-07 $l=3e-08 $layer=LI1_cond $X=1.1 $Y=0.655 $X2=1.1
+ $Y2=0.625
r67 19 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.78 $X2=1.1
+ $Y2=0.78
r68 19 20 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.78
+ $X2=0.345 $Y2=0.78
r69 16 20 6.81736 $w=2.5e-07 $l=1.79956e-07 $layer=LI1_cond $X=0.217 $Y=0.655
+ $X2=0.345 $Y2=0.78
r70 16 18 1.43529 $w=2.55e-07 $l=3e-08 $layer=LI1_cond $X=0.217 $Y=0.655
+ $X2=0.217 $Y2=0.625
r71 5 34 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.4
r72 4 32 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.4
r73 3 29 182 $w=1.7e-07 $l=4.52493e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.625
r74 2 23 182 $w=1.7e-07 $l=4.52493e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.625
r75 1 18 182 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%VGND 1 2 9 13 15 17 22 29 30 33 36
r91 36 37 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r92 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r93 30 37 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=7.59 $Y=0 $X2=1.61
+ $Y2=0
r94 29 30 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r95 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.52
+ $Y2=0
r96 27 29 385.246 $w=1.68e-07 $l=5.905e-06 $layer=LI1_cond $X=1.685 $Y=0
+ $X2=7.59 $Y2=0
r97 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r98 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r99 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r100 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r101 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r102 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.52
+ $Y2=0
r103 22 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.15 $Y2=0
r104 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r105 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r106 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r107 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r108 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r109 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.4
r110 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r111 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r112 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r113 1 9 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%A_445_47# 1 2 3 4 21
c33 21 0 1.09605e-19 $X=5.4 $Y=0.74
r34 19 21 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=0.78 $X2=5.4
+ $Y2=0.78
r35 17 19 62.6929 $w=2.48e-07 $l=1.36e-06 $layer=LI1_cond $X=3.2 $Y=0.78
+ $X2=4.56 $Y2=0.78
r36 14 17 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.78 $X2=3.2
+ $Y2=0.78
r37 4 21 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.74
r38 3 19 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.74
r39 2 17 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.74
r40 1 14 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4_4%A_803_47# 1 2 3 4 5 16 24 26 30 32 35
c47 26 0 1.93124e-19 $X=7.475 $Y=0.37
r48 30 37 3.25045 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=7.602 $Y=0.485
+ $X2=7.602 $Y2=0.37
r49 30 32 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=7.602 $Y=0.485
+ $X2=7.602 $Y2=0.74
r50 27 35 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=0.37
+ $X2=5.855 $Y2=0.37
r51 27 29 39.0829 $w=2.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.94 $Y=0.37
+ $X2=6.72 $Y2=0.37
r52 26 37 3.58963 $w=2.3e-07 $l=1.27e-07 $layer=LI1_cond $X=7.475 $Y=0.37
+ $X2=7.602 $Y2=0.37
r53 26 29 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=7.475 $Y=0.37
+ $X2=6.72 $Y2=0.37
r54 22 35 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.855 $Y=0.485
+ $X2=5.855 $Y2=0.37
r55 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.855 $Y=0.485
+ $X2=5.855 $Y2=0.74
r56 18 21 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.37
+ $X2=4.98 $Y2=0.37
r57 16 35 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.77 $Y=0.37
+ $X2=5.855 $Y2=0.37
r58 16 21 39.5839 $w=2.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.77 $Y=0.37
+ $X2=4.98 $Y2=0.37
r59 5 37 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.56 $Y2=0.4
r60 5 32 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.56 $Y2=0.74
r61 4 29 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.585
+ $Y=0.235 $X2=6.72 $Y2=0.4
r62 3 35 182 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.855 $Y2=0.4
r63 3 24 182 $w=1.7e-07 $l=5.83845e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.855 $Y2=0.74
r64 2 21 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.4
r65 1 18 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.4
.ends


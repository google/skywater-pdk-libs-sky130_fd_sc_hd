* File: sky130_fd_sc_hd__ebufn_8.spice
* Created: Thu Aug 27 14:19:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__ebufn_8.pex.spice"
.subckt sky130_fd_sc_hd__ebufn_8  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_116_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.19175 AS=0.08775 PD=1.89 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A_M1020_g N_A_116_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.08775 PD=1.005 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1031 N_A_301_47#_M1031_d N_TE_B_M1031_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.115375 PD=1.82 PS=1.005 NRD=0 NRS=14.76 M=1 R=4.33333
+ SA=75001.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_455_47#_M1000_d N_A_301_47#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_455_47#_M1005_d N_A_301_47#_M1005_g N_VGND_M1000_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75006.3 A=0.0975 P=1.6 MULT=1
MM1007 N_A_455_47#_M1005_d N_A_301_47#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1010 N_A_455_47#_M1010_d N_A_301_47#_M1010_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1012 N_A_455_47#_M1010_d N_A_301_47#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75005.1 A=0.0975 P=1.6 MULT=1
MM1014 N_A_455_47#_M1014_d N_A_301_47#_M1014_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75004.7 A=0.0975 P=1.6 MULT=1
MM1015 N_A_455_47#_M1014_d N_A_301_47#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75004.2 A=0.0975 P=1.6 MULT=1
MM1021 N_A_455_47#_M1021_d N_A_301_47#_M1021_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.17225 AS=0.08775 PD=1.18 PS=0.92 NRD=23.988 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1001 N_Z_M1001_d N_A_116_47#_M1001_g N_A_455_47#_M1021_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.17225 PD=0.92 PS=1.18 NRD=0 NRS=22.152 M=1 R=4.33333
+ SA=75003.8 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1006 N_Z_M1001_d N_A_116_47#_M1006_g N_A_455_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75004.2 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1026 N_Z_M1026_d N_A_116_47#_M1026_g N_A_455_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75004.6 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1027 N_Z_M1026_d N_A_116_47#_M1027_g N_A_455_47#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75005.1 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1029 N_Z_M1029_d N_A_116_47#_M1029_g N_A_455_47#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75005.5 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1032 N_Z_M1029_d N_A_116_47#_M1032_g N_A_455_47#_M1032_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75005.9 SB=75001 A=0.0975 P=1.6 MULT=1
MM1033 N_Z_M1033_d N_A_116_47#_M1033_g N_A_455_47#_M1032_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75006.3 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1034 N_Z_M1033_d N_A_116_47#_M1034_g N_A_455_47#_M1034_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75006.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1019 N_VPWR_M1019_d N_A_M1019_g N_A_116_47#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1036 N_VPWR_M1036_d N_A_M1036_g N_A_116_47#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1775 AS=0.135 PD=1.355 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1025 N_A_301_47#_M1025_d N_TE_B_M1025_g N_VPWR_M1036_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1775 PD=2.52 PS=1.355 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_407_309#_M1002_d N_TE_B_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.2444 AS=0.1269 PD=2.4 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667 SA=75000.2
+ SB=75007 A=0.141 P=2.18 MULT=1
MM1008 N_A_407_309#_M1008_d N_TE_B_M1008_g N_VPWR_M1002_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75000.6 SB=75006.6 A=0.141 P=2.18 MULT=1
MM1011 N_A_407_309#_M1008_d N_TE_B_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667 SA=75001
+ SB=75006.2 A=0.141 P=2.18 MULT=1
MM1016 N_A_407_309#_M1016_d N_TE_B_M1016_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75001.4 SB=75005.7 A=0.141 P=2.18 MULT=1
MM1017 N_A_407_309#_M1016_d N_TE_B_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75001.9 SB=75005.3 A=0.141 P=2.18 MULT=1
MM1022 N_A_407_309#_M1022_d N_TE_B_M1022_g N_VPWR_M1017_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75002.3 SB=75004.9 A=0.141 P=2.18 MULT=1
MM1028 N_A_407_309#_M1022_d N_TE_B_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75002.7 SB=75004.5 A=0.141 P=2.18 MULT=1
MM1037 N_A_407_309#_M1037_d N_TE_B_M1037_g N_VPWR_M1028_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.370912 AS=0.1269 PD=1.71526 PS=1.21 NRD=16.7647 NRS=0 M=1
+ R=6.26667 SA=75003.1 SB=75004.1 A=0.141 P=2.18 MULT=1
MM1003 N_A_407_309#_M1037_d N_A_116_47#_M1003_g N_Z_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.394588 AS=0.135 PD=1.82474 PS=1.27 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75003.8 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1009 N_A_407_309#_M1009_d N_A_116_47#_M1009_g N_Z_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.3
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1013 N_A_407_309#_M1009_d N_A_116_47#_M1013_g N_Z_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.7
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1018 N_A_407_309#_M1018_d N_A_116_47#_M1018_g N_Z_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.1
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1023 N_A_407_309#_M1018_d N_A_116_47#_M1023_g N_Z_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.5
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1024 N_A_407_309#_M1024_d N_A_116_47#_M1024_g N_Z_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.9
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1030 N_A_407_309#_M1024_d N_A_116_47#_M1030_g N_Z_M1030_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1035 N_A_407_309#_M1035_d N_A_116_47#_M1035_g N_Z_M1030_s VPB PHIGHVT L=0.15
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX38_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_83 VNB 0 1.39443e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__ebufn_8.pxi.spice"
*
.ends
*
*

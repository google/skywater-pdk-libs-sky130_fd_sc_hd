* File: sky130_fd_sc_hd__or3b_2.spice
* Created: Thu Aug 27 14:43:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or3b_2.spice.pex"
.subckt sky130_fd_sc_hd__or3b_2  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_C_N_M1009_g N_A_27_47#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1009_d N_A_176_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=11.076 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_176_21#_M1004_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.123773 AS=0.08775 PD=1.2028 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_A_176_21#_M1005_d N_A_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0799766 PD=0.69 PS=0.777196 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_A_176_21#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_176_21#_M1006_d N_A_27_47#_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_C_N_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.1092 PD=0.789718 PS=1.36 NRD=70.4866 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1010_d N_A_176_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.205282 AS=0.135 PD=1.88028 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.4
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_176_21#_M1011_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.208803 AS=0.135 PD=1.88732 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 A_388_297# N_A_M1001_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0567
+ AS=0.0876972 PD=0.69 PS=0.792676 NRD=37.5088 NRS=72.1217 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_472_297# N_B_M1000_g A_388_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.0567
+ AS=0.0567 PD=0.69 PS=0.69 NRD=37.5088 NRS=37.5088 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_176_21#_M1008_d N_A_27_47#_M1008_g A_472_297# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=37.5088 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__or3b_2.spice.SKY130_FD_SC_HD__OR3B_2.pxi"
*
.ends
*
*

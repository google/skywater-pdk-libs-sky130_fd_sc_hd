# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__xnor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175000 1.075000 5.390000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.075000 1.855000 1.275000 ;
        RECT 1.685000 1.275000 1.855000 1.445000 ;
        RECT 1.685000 1.445000 5.730000 1.615000 ;
        RECT 5.560000 1.075000 7.430000 1.275000 ;
        RECT 5.560000 1.275000 5.730000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.721000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.160000 1.785000  8.250000 2.045000 ;
        RECT 7.960000 1.445000 10.035000 1.665000 ;
        RECT 7.960000 1.665000  8.250000 1.785000 ;
        RECT 7.960000 2.045000  8.250000 2.465000 ;
        RECT 8.380000 0.645000 10.035000 0.905000 ;
        RECT 8.840000 1.665000  9.090000 2.465000 ;
        RECT 9.680000 1.665000 10.035000 2.465000 ;
        RECT 9.815000 0.905000 10.035000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 2.350000  0.085000  2.520000 0.555000 ;
        RECT 3.190000  0.085000  3.360000 0.555000 ;
        RECT 4.035000  0.085000  4.310000 0.905000 ;
        RECT 4.980000  0.085000  5.150000 0.555000 ;
        RECT 5.820000  0.085000  5.990000 0.555000 ;
        RECT 6.660000  0.085000  6.830000 0.555000 ;
        RECT 7.500000  0.085000  7.770000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.630000 1.835000  0.880000 2.635000 ;
        RECT 1.470000 2.175000  1.720000 2.635000 ;
        RECT 2.310000 2.175000  2.560000 2.635000 ;
        RECT 3.150000 2.175000  3.400000 2.635000 ;
        RECT 4.520000 2.175000  4.770000 2.635000 ;
        RECT 5.360000 2.175000  5.610000 2.635000 ;
        RECT 8.420000 1.835000  8.670000 2.635000 ;
        RECT 9.260000 1.835000  9.510000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.645000 1.760000 0.905000 ;
      RECT 0.085000 0.905000 0.320000 1.445000 ;
      RECT 0.085000 1.445000 1.300000 1.615000 ;
      RECT 0.085000 1.615000 0.460000 2.465000 ;
      RECT 0.170000 0.255000 2.180000 0.475000 ;
      RECT 1.050000 1.615000 1.300000 1.785000 ;
      RECT 1.050000 1.785000 3.820000 2.005000 ;
      RECT 1.050000 2.005000 1.300000 2.465000 ;
      RECT 1.890000 2.005000 2.140000 2.465000 ;
      RECT 1.930000 0.475000 2.180000 0.725000 ;
      RECT 1.930000 0.725000 3.860000 0.905000 ;
      RECT 2.690000 0.255000 3.020000 0.725000 ;
      RECT 2.730000 2.005000 2.980000 2.465000 ;
      RECT 3.530000 0.255000 3.860000 0.725000 ;
      RECT 3.570000 2.005000 3.820000 2.465000 ;
      RECT 4.035000 1.785000 5.990000 2.005000 ;
      RECT 4.035000 2.005000 4.350000 2.465000 ;
      RECT 4.480000 0.255000 4.810000 0.725000 ;
      RECT 4.480000 0.725000 7.430000 0.735000 ;
      RECT 4.480000 0.735000 8.210000 0.905000 ;
      RECT 4.940000 2.005000 5.190000 2.465000 ;
      RECT 5.320000 0.255000 5.650000 0.725000 ;
      RECT 5.780000 2.005000 5.990000 2.215000 ;
      RECT 5.780000 2.215000 7.750000 2.465000 ;
      RECT 5.900000 1.445000 7.770000 1.615000 ;
      RECT 6.160000 0.255000 6.490000 0.725000 ;
      RECT 7.000000 0.255000 7.330000 0.725000 ;
      RECT 7.600000 1.075000 9.645000 1.275000 ;
      RECT 7.600000 1.275000 7.770000 1.445000 ;
      RECT 7.960000 0.305000 9.970000 0.475000 ;
      RECT 7.960000 0.475000 8.210000 0.735000 ;
    LAYER mcon ;
      RECT 1.065000 1.445000 1.235000 1.615000 ;
      RECT 6.125000 1.445000 6.295000 1.615000 ;
    LAYER met1 ;
      RECT 1.005000 1.415000 1.295000 1.460000 ;
      RECT 1.005000 1.460000 6.355000 1.600000 ;
      RECT 1.005000 1.600000 1.295000 1.645000 ;
      RECT 6.065000 1.415000 6.355000 1.460000 ;
      RECT 6.065000 1.600000 6.355000 1.645000 ;
  END
END sky130_fd_sc_hd__xnor2_4

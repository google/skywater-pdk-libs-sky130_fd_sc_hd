* File: sky130_fd_sc_hd__nand3b_2.pxi.spice
* Created: Thu Aug 27 14:29:53 2020
* 
x_PM_SKY130_FD_SC_HD__NAND3B_2%A_N N_A_N_M1013_g N_A_N_M1004_g A_N N_A_N_c_77_n
+ PM_SKY130_FD_SC_HD__NAND3B_2%A_N
x_PM_SKY130_FD_SC_HD__NAND3B_2%C N_C_M1005_g N_C_M1007_g N_C_M1008_g N_C_M1011_g
+ C C N_C_c_107_n PM_SKY130_FD_SC_HD__NAND3B_2%C
x_PM_SKY130_FD_SC_HD__NAND3B_2%B N_B_M1001_g N_B_M1003_g N_B_M1000_g N_B_M1002_g
+ B B B N_B_c_153_n PM_SKY130_FD_SC_HD__NAND3B_2%B
x_PM_SKY130_FD_SC_HD__NAND3B_2%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1004_s
+ N_A_27_47#_M1006_g N_A_27_47#_M1010_g N_A_27_47#_M1009_g N_A_27_47#_M1012_g
+ N_A_27_47#_c_198_n N_A_27_47#_c_204_n N_A_27_47#_c_205_n N_A_27_47#_c_199_n
+ N_A_27_47#_c_206_n N_A_27_47#_c_207_n N_A_27_47#_c_208_n N_A_27_47#_c_200_n
+ PM_SKY130_FD_SC_HD__NAND3B_2%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND3B_2%VPWR N_VPWR_M1004_d N_VPWR_M1011_d N_VPWR_M1003_d
+ N_VPWR_M1010_d N_VPWR_M1012_d N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n
+ N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n
+ VPWR N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n
+ N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_278_n
+ PM_SKY130_FD_SC_HD__NAND3B_2%VPWR
x_PM_SKY130_FD_SC_HD__NAND3B_2%Y N_Y_M1006_s N_Y_M1007_s N_Y_M1001_s N_Y_M1010_s
+ N_Y_c_355_n N_Y_c_351_n N_Y_c_349_n N_Y_c_352_n N_Y_c_354_n N_Y_c_358_n
+ N_Y_c_379_n Y Y PM_SKY130_FD_SC_HD__NAND3B_2%Y
x_PM_SKY130_FD_SC_HD__NAND3B_2%VGND N_VGND_M1013_d N_VGND_M1008_d N_VGND_c_414_n
+ N_VGND_c_415_n N_VGND_c_416_n VGND N_VGND_c_417_n N_VGND_c_418_n
+ N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n PM_SKY130_FD_SC_HD__NAND3B_2%VGND
x_PM_SKY130_FD_SC_HD__NAND3B_2%A_218_47# N_A_218_47#_M1005_s N_A_218_47#_M1000_d
+ N_A_218_47#_c_472_n N_A_218_47#_c_468_n N_A_218_47#_c_469_n
+ N_A_218_47#_c_470_n N_A_218_47#_c_471_n PM_SKY130_FD_SC_HD__NAND3B_2%A_218_47#
x_PM_SKY130_FD_SC_HD__NAND3B_2%A_408_47# N_A_408_47#_M1000_s N_A_408_47#_M1002_s
+ N_A_408_47#_M1009_d N_A_408_47#_c_502_n N_A_408_47#_c_503_n
+ N_A_408_47#_c_504_n N_A_408_47#_c_523_n PM_SKY130_FD_SC_HD__NAND3B_2%A_408_47#
cc_1 VNB N_A_N_M1013_g 0.0343996f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.00233138f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_3 VNB N_A_N_c_77_n 0.0275829f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_4 VNB N_C_M1005_g 0.0186937f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB N_C_M1007_g 4.43991e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_6 VNB N_C_M1008_g 0.0238914f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.16
cc_7 VNB N_C_M1011_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_8 VNB C 0.00583613f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_9 VNB N_C_c_107_n 0.0290308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_M1001_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_11 VNB N_B_M1003_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_12 VNB N_B_M1000_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.16
cc_13 VNB N_B_M1002_g 0.0176813f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_14 VNB B 0.00625415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B_c_153_n 0.0709095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_M1006_g 0.0176616f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_17 VNB N_A_27_47#_M1010_g 7.17814e-19 $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_18 VNB N_A_27_47#_M1009_g 0.0208563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_M1012_g 4.56514e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_198_n 0.0307423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_199_n 0.0188007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_200_n 0.0317334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_278_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_349_n 0.0199508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB Y 0.0197113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_414_n 0.0102463f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_27 VNB N_VGND_c_415_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.16
cc_28 VNB N_VGND_c_416_n 0.00826368f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_29 VNB N_VGND_c_417_n 0.0174876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_418_n 0.0557983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_419_n 0.221826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_420_n 0.00595612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_421_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_218_47#_c_468_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_35 VNB N_A_218_47#_c_469_n 0.00236711f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_36 VNB N_A_218_47#_c_470_n 0.00317456f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_37 VNB N_A_218_47#_c_471_n 0.00912193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_408_47#_c_502_n 0.00245946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_408_47#_c_503_n 0.00185524f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.175
cc_40 VNB N_A_408_47#_c_504_n 0.0103948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VPB N_A_N_M1004_g 0.0589469f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_42 VPB N_A_N_c_77_n 0.00588003f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_43 VPB N_C_M1007_g 0.020714f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_44 VPB N_C_M1011_g 0.0194911f $X=-0.19 $Y=1.305 $X2=0.562 $Y2=1.325
cc_45 VPB N_B_M1001_g 0.0194911f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_46 VPB N_B_M1003_g 0.0267252f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_47 VPB N_A_27_47#_M1010_g 0.026666f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_48 VPB N_A_27_47#_M1012_g 0.0223499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_198_n 0.00671796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_204_n 0.0302764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_205_n 0.00136269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_206_n 0.00770964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_207_n 0.0167397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_208_n 0.021328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_279_n 0.00713256f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_56 VPB N_VPWR_c_280_n 0.017296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_281_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_282_n 0.00573435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_283_n 0.00598254f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_284_n 0.00573435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_285_n 0.0106218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_286_n 0.0177765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_287_n 0.0174876f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_288_n 0.017296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_289_n 0.0178421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_290_n 0.00593022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_291_n 0.00323604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_292_n 0.00477752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_293_n 0.00477752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_278_n 0.045637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_Y_c_351_n 0.00745667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_Y_c_352_n 0.0102944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB Y 0.0200987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 N_A_N_M1013_g N_C_M1005_g 0.0146134f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_N_c_77_n N_C_M1005_g 0.0223343f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_N_M1004_g N_C_M1007_g 0.0266063f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_77 A_N C 0.0115096f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_78 A_N N_C_c_107_n 0.00152567f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_N_M1013_g N_A_27_47#_c_198_n 0.0226339f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_80 A_N N_A_27_47#_c_198_n 0.0150209f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A_N_M1004_g N_A_27_47#_c_204_n 0.0177669f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_82 A_N N_A_27_47#_c_204_n 0.0250954f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_N_c_77_n N_A_27_47#_c_204_n 0.00439952f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_N_M1013_g N_A_27_47#_c_199_n 0.00544454f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_N_M1004_g N_A_27_47#_c_207_n 0.00507425f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_86 N_A_N_M1004_g N_A_27_47#_c_208_n 0.0127931f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_87 N_A_N_M1004_g N_VPWR_c_279_n 0.00829144f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_88 N_A_N_M1004_g N_VPWR_c_287_n 0.00564131f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_89 N_A_N_M1004_g N_VPWR_c_278_n 0.011364f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_90 N_A_N_M1004_g N_Y_c_354_n 2.66813e-19 $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_91 N_A_N_M1013_g N_VGND_c_414_n 0.00852603f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_92 A_N N_VGND_c_414_n 0.0164192f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A_N_c_77_n N_VGND_c_414_n 0.00382571f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_N_M1013_g N_VGND_c_417_n 0.00564131f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_N_M1013_g N_VGND_c_419_n 0.011364f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_96 N_C_M1011_g N_B_M1001_g 0.0309508f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_97 C B 0.0150406f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_98 C N_B_c_153_n 0.00213358f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_99 N_C_c_107_n N_B_c_153_n 0.0309508f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_100 N_C_M1007_g N_A_27_47#_c_204_n 0.0183009f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_101 N_C_M1011_g N_A_27_47#_c_204_n 0.0103223f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_102 C N_A_27_47#_c_204_n 0.0494367f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_103 N_C_c_107_n N_A_27_47#_c_204_n 0.00198252f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_104 N_C_M1007_g N_VPWR_c_279_n 0.00172108f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_105 N_C_M1007_g N_VPWR_c_280_n 0.00541359f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_106 N_C_M1011_g N_VPWR_c_280_n 0.00422241f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_107 N_C_M1011_g N_VPWR_c_281_n 0.00146448f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_108 N_C_M1007_g N_VPWR_c_278_n 0.00980531f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_109 N_C_M1011_g N_VPWR_c_278_n 0.00572376f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_110 N_C_M1011_g N_Y_c_355_n 0.00954125f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_111 N_C_M1007_g N_Y_c_354_n 0.00868254f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_112 N_C_M1011_g N_Y_c_354_n 0.00745991f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_113 N_C_M1011_g N_Y_c_358_n 5.19281e-19 $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_114 N_C_M1005_g N_VGND_c_414_n 0.0018963f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_115 N_C_M1005_g N_VGND_c_415_n 0.00541359f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_116 N_C_M1008_g N_VGND_c_415_n 0.00422241f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_117 N_C_M1008_g N_VGND_c_416_n 0.00321269f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_118 N_C_M1005_g N_VGND_c_419_n 0.00980531f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_119 N_C_M1008_g N_VGND_c_419_n 0.00702263f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_120 N_C_M1005_g N_A_218_47#_c_472_n 0.00511586f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_121 N_C_M1008_g N_A_218_47#_c_472_n 0.00907724f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_122 N_C_M1005_g N_A_218_47#_c_468_n 0.00266814f $X=1.015 $Y=0.56 $X2=0 $Y2=0
cc_123 N_C_M1008_g N_A_218_47#_c_468_n 0.00116017f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_124 C N_A_218_47#_c_468_n 0.0265408f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_125 N_C_c_107_n N_A_218_47#_c_468_n 0.00213429f $X=1.435 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C_M1008_g N_A_218_47#_c_469_n 0.00137399f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_127 N_C_M1008_g N_A_218_47#_c_471_n 0.0112581f $X=1.435 $Y=0.56 $X2=0 $Y2=0
cc_128 C N_A_218_47#_c_471_n 0.0259558f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B_M1002_g N_A_27_47#_M1006_g 0.0139248f $X=2.795 $Y=0.56 $X2=0 $Y2=0
cc_130 N_B_M1001_g N_A_27_47#_c_204_n 0.0116623f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_131 N_B_M1003_g N_A_27_47#_c_204_n 0.0124694f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_132 B N_A_27_47#_c_204_n 0.0866172f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B_c_153_n N_A_27_47#_c_204_n 0.015566f $X=2.795 $Y=1.16 $X2=0 $Y2=0
cc_134 B N_A_27_47#_c_205_n 0.0150931f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_135 N_B_c_153_n N_A_27_47#_c_205_n 2.36933e-19 $X=2.795 $Y=1.16 $X2=0 $Y2=0
cc_136 B N_A_27_47#_c_200_n 0.0021379f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_137 N_B_c_153_n N_A_27_47#_c_200_n 0.0139248f $X=2.795 $Y=1.16 $X2=0 $Y2=0
cc_138 N_B_M1001_g N_VPWR_c_281_n 0.00146448f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_139 N_B_M1003_g N_VPWR_c_282_n 0.00321269f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B_M1001_g N_VPWR_c_288_n 0.00422241f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B_M1003_g N_VPWR_c_288_n 0.00541359f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B_M1001_g N_VPWR_c_278_n 0.00572376f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B_M1003_g N_VPWR_c_278_n 0.00712156f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B_M1001_g N_Y_c_355_n 0.00954125f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B_M1003_g N_Y_c_351_n 0.0101664f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_146 N_B_M1001_g N_Y_c_354_n 5.19281e-19 $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_147 N_B_M1001_g N_Y_c_358_n 0.00745991f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B_M1003_g N_Y_c_358_n 0.0143133f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B_M1000_g N_VGND_c_416_n 0.00231165f $X=2.375 $Y=0.56 $X2=0 $Y2=0
cc_150 N_B_M1000_g N_VGND_c_418_n 0.00357877f $X=2.375 $Y=0.56 $X2=0 $Y2=0
cc_151 N_B_M1002_g N_VGND_c_418_n 0.00357877f $X=2.795 $Y=0.56 $X2=0 $Y2=0
cc_152 N_B_M1000_g N_VGND_c_419_n 0.00655123f $X=2.375 $Y=0.56 $X2=0 $Y2=0
cc_153 N_B_M1002_g N_VGND_c_419_n 0.00525237f $X=2.795 $Y=0.56 $X2=0 $Y2=0
cc_154 N_B_M1000_g N_A_218_47#_c_470_n 0.0142655f $X=2.375 $Y=0.56 $X2=0 $Y2=0
cc_155 N_B_M1002_g N_A_218_47#_c_470_n 0.00383673f $X=2.795 $Y=0.56 $X2=0 $Y2=0
cc_156 N_B_c_153_n N_A_218_47#_c_470_n 0.00207887f $X=2.795 $Y=1.16 $X2=0 $Y2=0
cc_157 B N_A_218_47#_c_471_n 0.0591961f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_158 N_B_c_153_n N_A_218_47#_c_471_n 0.0148894f $X=2.795 $Y=1.16 $X2=0 $Y2=0
cc_159 N_B_M1000_g N_A_408_47#_c_502_n 0.00866705f $X=2.375 $Y=0.56 $X2=0 $Y2=0
cc_160 N_B_M1002_g N_A_408_47#_c_502_n 0.0103313f $X=2.795 $Y=0.56 $X2=0 $Y2=0
cc_161 B N_A_408_47#_c_502_n 0.00368637f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_162 B N_A_408_47#_c_503_n 0.0142952f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_204_n N_VPWR_M1004_d 0.00337911f $X=3.32 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_164 N_A_27_47#_c_204_n N_VPWR_M1011_d 0.00166235f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_204_n N_VPWR_M1003_d 0.0027344f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_204_n N_VPWR_M1010_d 0.0027344f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_204_n N_VPWR_c_279_n 0.0204137f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_208_n N_VPWR_c_279_n 0.0116244f $X=0.25 $Y=2.065 $X2=0 $Y2=0
cc_169 N_A_27_47#_M1010_g N_VPWR_c_284_n 0.00321269f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_M1012_g N_VPWR_c_286_n 0.0032322f $X=3.635 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_207_n N_VPWR_c_287_n 0.0201353f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1010_g N_VPWR_c_289_n 0.00541359f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1012_g N_VPWR_c_289_n 0.00436487f $X=3.635 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_M1004_s N_VPWR_c_278_n 0.00209319f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_M1010_g N_VPWR_c_278_n 0.00712156f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1012_g N_VPWR_c_278_n 0.00684832f $X=3.635 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_207_n N_VPWR_c_278_n 0.012035f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_204_n N_Y_M1007_s 0.00165831f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_204_n N_Y_M1001_s 0.00165831f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_204_n N_Y_M1010_s 0.00171424f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_204_n N_Y_c_355_n 0.0280797f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1010_g N_Y_c_351_n 0.0101664f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_204_n N_Y_c_351_n 0.0660197f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1006_g N_Y_c_349_n 0.00420883f $X=3.215 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1009_g N_Y_c_349_n 0.015665f $X=3.635 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_204_n N_Y_c_349_n 0.00185145f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_205_n N_Y_c_349_n 0.0262855f $X=3.485 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_200_n N_Y_c_349_n 0.00207755f $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_27_47#_M1012_g N_Y_c_352_n 0.0152618f $X=3.635 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_204_n N_Y_c_352_n 0.00677293f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_204_n N_Y_c_354_n 0.0172624f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_204_n N_Y_c_358_n 0.0172624f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_193 N_A_27_47#_M1010_g N_Y_c_379_n 0.0138434f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_204_n N_Y_c_379_n 0.016072f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_200_n N_Y_c_379_n 3.59001e-19 $X=3.635 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_27_47#_M1009_g Y 0.024803f $X=3.635 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_204_n Y 0.0119682f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_205_n Y 0.0248539f $X=3.485 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_198_n N_VGND_c_414_n 0.0126396f $X=0.175 $Y=1.445 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_204_n N_VGND_c_414_n 0.00412107f $X=3.32 $Y=1.53 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_199_n N_VGND_c_417_n 0.0201353f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1006_g N_VGND_c_418_n 0.00357877f $X=3.215 $Y=0.56 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1009_g N_VGND_c_418_n 0.00357877f $X=3.635 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_M1013_s N_VGND_c_419_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_M1006_g N_VGND_c_419_n 0.00525237f $X=3.215 $Y=0.56 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_M1009_g N_VGND_c_419_n 0.00621133f $X=3.635 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_199_n N_VGND_c_419_n 0.012035f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_204_n N_A_218_47#_c_471_n 0.00656263f $X=3.32 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_M1006_g N_A_408_47#_c_504_n 0.0124168f $X=3.215 $Y=0.56 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_M1009_g N_A_408_47#_c_504_n 0.00866705f $X=3.635 $Y=0.56 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_278_n N_Y_M1007_s 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_212 N_VPWR_c_278_n N_Y_M1001_s 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_278_n N_Y_M1010_s 0.00238028f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_M1011_d N_Y_c_355_n 0.00330444f $X=1.51 $Y=1.485 $X2=0 $Y2=0
cc_215 N_VPWR_c_280_n N_Y_c_355_n 0.00205325f $X=1.56 $Y=2.72 $X2=0 $Y2=0
cc_216 N_VPWR_c_281_n N_Y_c_355_n 0.0123861f $X=1.645 $Y=2.34 $X2=0 $Y2=0
cc_217 N_VPWR_c_288_n N_Y_c_355_n 0.00205325f $X=2.4 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_278_n N_Y_c_355_n 0.00852004f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_219 N_VPWR_M1003_d N_Y_c_351_n 0.00502005f $X=2.35 $Y=1.485 $X2=0 $Y2=0
cc_220 N_VPWR_M1010_d N_Y_c_351_n 0.00526687f $X=2.88 $Y=1.485 $X2=0 $Y2=0
cc_221 N_VPWR_c_282_n N_Y_c_351_n 0.0154104f $X=2.485 $Y=2.34 $X2=0 $Y2=0
cc_222 N_VPWR_c_284_n N_Y_c_351_n 0.0154104f $X=3.005 $Y=2.34 $X2=0 $Y2=0
cc_223 N_VPWR_c_278_n N_Y_c_351_n 0.0196453f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_M1012_d N_Y_c_352_n 0.00634141f $X=3.71 $Y=1.485 $X2=0 $Y2=0
cc_225 N_VPWR_c_286_n N_Y_c_352_n 0.0239447f $X=3.845 $Y=2.34 $X2=0 $Y2=0
cc_226 N_VPWR_c_289_n N_Y_c_352_n 0.00286836f $X=3.76 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_c_278_n N_Y_c_352_n 0.00710254f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_280_n N_Y_c_354_n 0.0189039f $X=1.56 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_278_n N_Y_c_354_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_c_288_n N_Y_c_358_n 0.0189039f $X=2.4 $Y=2.72 $X2=0 $Y2=0
cc_231 N_VPWR_c_278_n N_Y_c_358_n 0.0122217f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_289_n N_Y_c_379_n 0.0151499f $X=3.76 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_c_278_n N_Y_c_379_n 0.00934584f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_234 N_VPWR_M1012_d Y 0.00468912f $X=3.71 $Y=1.485 $X2=0 $Y2=0
cc_235 N_Y_M1006_s N_VGND_c_419_n 0.00216833f $X=3.29 $Y=0.235 $X2=0 $Y2=0
cc_236 N_Y_c_349_n N_A_408_47#_M1009_d 0.00324009f $X=3.85 $Y=0.77 $X2=0 $Y2=0
cc_237 N_Y_c_349_n N_A_408_47#_c_503_n 0.0119693f $X=3.85 $Y=0.77 $X2=0 $Y2=0
cc_238 N_Y_M1006_s N_A_408_47#_c_504_n 0.00305599f $X=3.29 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_c_349_n N_A_408_47#_c_504_n 0.045199f $X=3.85 $Y=0.77 $X2=0 $Y2=0
cc_240 N_VGND_c_419_n N_A_218_47#_M1005_s 0.00215201f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_241 N_VGND_c_419_n N_A_218_47#_M1000_d 0.00216833f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_242 N_VGND_c_415_n N_A_218_47#_c_472_n 0.0188551f $X=1.56 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_419_n N_A_218_47#_c_472_n 0.0122069f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_c_414_n N_A_218_47#_c_468_n 0.00878993f $X=0.745 $Y=0.38 $X2=0
+ $Y2=0
cc_245 N_VGND_M1008_d N_A_218_47#_c_471_n 0.00285834f $X=1.51 $Y=0.235 $X2=0
+ $Y2=0
cc_246 N_VGND_c_415_n N_A_218_47#_c_471_n 0.00203746f $X=1.56 $Y=0 $X2=0 $Y2=0
cc_247 N_VGND_c_416_n N_A_218_47#_c_471_n 0.0191473f $X=1.645 $Y=0.38 $X2=0
+ $Y2=0
cc_248 N_VGND_c_418_n N_A_218_47#_c_471_n 0.00296114f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_419_n N_A_218_47#_c_471_n 0.00998562f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_c_419_n N_A_408_47#_M1000_s 0.00209344f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_251 N_VGND_c_419_n N_A_408_47#_M1002_s 0.0021521f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_419_n N_A_408_47#_M1009_d 0.00209344f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_416_n N_A_408_47#_c_502_n 0.0166761f $X=1.645 $Y=0.38 $X2=0
+ $Y2=0
cc_254 N_VGND_c_418_n N_A_408_47#_c_502_n 0.0521531f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_419_n N_A_408_47#_c_502_n 0.0329109f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_418_n N_A_408_47#_c_504_n 0.0547682f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_419_n N_A_408_47#_c_504_n 0.0344075f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_418_n N_A_408_47#_c_523_n 0.0114305f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_c_419_n N_A_408_47#_c_523_n 0.00653933f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_260 N_A_218_47#_c_469_n N_A_408_47#_M1000_s 0.00209037f $X=2.135 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_261 N_A_218_47#_c_470_n N_A_408_47#_M1000_s 0.00111257f $X=2.585 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_262 N_A_218_47#_M1000_d N_A_408_47#_c_502_n 0.00305599f $X=2.45 $Y=0.235
+ $X2=0 $Y2=0
cc_263 N_A_218_47#_c_469_n N_A_408_47#_c_502_n 0.0410587f $X=2.135 $Y=0.77 $X2=0
+ $Y2=0
cc_264 N_A_218_47#_c_470_n N_A_408_47#_c_503_n 0.0119693f $X=2.585 $Y=0.72 $X2=0
+ $Y2=0

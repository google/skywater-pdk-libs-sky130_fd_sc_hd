* File: sky130_fd_sc_hd__nor2_2.pex.spice
* Created: Thu Aug 27 14:31:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR2_2%A 1 3 6 8 10 13 15 16 24
c38 16 0 1.24925e-19 $X=0.61 $Y=1.105
c39 13 0 1.19433e-19 $X=0.91 $Y=1.985
r40 22 24 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=0.645 $Y=1.16
+ $X2=0.91 $Y2=1.16
r41 19 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.645 $Y2=1.16
r42 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r43 15 16 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.645 $Y2=1.175
r44 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r45 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r46 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r47 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r48 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r49 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r50 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_2%B 1 3 6 8 10 13 15 16 24
c47 24 0 1.24925e-19 $X=1.75 $Y=1.16
r48 22 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.54 $Y=1.16
+ $X2=1.75 $Y2=1.16
r49 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.54 $Y2=1.16
r50 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.16 $X2=1.54 $Y2=1.16
r51 15 16 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.54 $Y2=1.175
r52 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r54 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r56 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325 $X2=1.33
+ $Y2=1.985
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995 $X2=1.33
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_2%A_27_297# 1 2 3 10 12 14 16 17 18 22
r35 20 22 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.025 $Y=2.295
+ $X2=2.025 $Y2=2
r36 19 29 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=2.38
+ $X2=1.12 $Y2=2.38
r37 18 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.875 $Y=2.38
+ $X2=2.025 $Y2=2.295
r38 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.875 $Y=2.38
+ $X2=1.205 $Y2=2.38
r39 17 29 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.295
+ $X2=1.12 $Y2=2.38
r40 16 27 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.56
r41 16 17 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=2.295
r42 15 25 3.96222 $w=2.1e-07 $l=1.38e-07 $layer=LI1_cond $X=0.365 $Y=1.56
+ $X2=0.227 $Y2=1.56
r43 14 27 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=1.56
+ $X2=1.12 $Y2=1.56
r44 14 15 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.035 $Y=1.56
+ $X2=0.365 $Y2=1.56
r45 10 25 3.01473 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=1.56
r46 10 12 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=2.3
r47 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2
r48 2 29 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r49 2 27 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r50 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r51 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_2%VPWR 1 6 8 10 20 21 24
r29 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r30 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r31 18 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 17 20 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.7 $Y2=2.72
r36 15 17 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.7 $Y2=2.72
r38 10 12 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r39 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r41 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2.72
r42 4 6 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2
r43 1 6 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_2%Y 1 2 3 12 14 15 18 20 23 24 29 31
c59 29 0 1.19433e-19 $X=2.027 $Y=1.555
r60 26 31 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.54 $Y=1.665
+ $X2=1.54 $Y2=1.87
r61 26 29 25.5109 $w=2.18e-07 $l=4.87e-07 $layer=LI1_cond $X=1.54 $Y=1.555
+ $X2=2.027 $Y2=1.555
r62 23 29 0.884026 $w=2.15e-07 $l=1.1e-07 $layer=LI1_cond $X=2.027 $Y=1.445
+ $X2=2.027 $Y2=1.555
r63 22 23 28.9451 $w=2.13e-07 $l=5.4e-07 $layer=LI1_cond $X=2.027 $Y=0.905
+ $X2=2.027 $Y2=1.445
r64 21 24 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.705 $Y=0.82
+ $X2=1.54 $Y2=0.815
r65 20 22 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.92 $Y=0.82
+ $X2=2.027 $Y2=0.905
r66 20 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.92 $Y=0.82
+ $X2=1.705 $Y2=0.82
r67 16 24 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725 $X2=1.54
+ $Y2=0.815
r68 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r69 14 24 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r70 14 15 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r71 10 15 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r72 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725 $X2=0.7
+ $Y2=0.39
r73 3 26 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.62
r74 2 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r75 1 12 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_2%VGND 1 2 3 10 12 16 18 20 23 24 25 31 40
r38 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r39 34 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r40 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r41 31 39 4.33193 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.087
+ $Y2=0
r42 31 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.61
+ $Y2=0
r43 30 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r44 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 27 36 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r46 27 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r47 25 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r48 25 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r49 23 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r50 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r51 22 33 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.61
+ $Y2=0
r52 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r53 18 39 3.10591 $w=2.9e-07 $l=1.13666e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.087 $Y2=0
r54 18 20 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.39
r55 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r56 14 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r57 10 36 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r58 10 12 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r59 3 20 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r60 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r61 1 12 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


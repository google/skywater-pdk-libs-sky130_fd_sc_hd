* File: sky130_fd_sc_hd__nand4bb_4.pex.spice
* Created: Tue Sep  1 19:17:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%A_N 1 3 6 8 9 16
c25 6 0 6.72171e-20 $X=0.47 $Y=1.985
r26 13 16 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r27 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.16
+ $X2=0.215 $Y2=1.53
r28 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r29 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r31 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%B_N 1 3 6 8 9 13 14
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r35 8 9 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.782 $Y=1.19
+ $X2=0.782 $Y2=1.53
r36 8 14 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=0.782 $Y=1.19
+ $X2=0.782 $Y2=1.16
r37 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r38 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r39 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%A_27_47# 1 2 7 9 12 16 20 24 28 30 32 36
+ 40 44 46 47 48 49 53 57 60
c143 20 0 5.15114e-20 $X=2.915 $Y=1.985
r144 60 63 12.3868 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.42 $Y=1.16
+ $X2=2.495 $Y2=1.16
r145 54 60 183.604 $w=3.3e-07 $l=1.05e-06 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=2.42 $Y2=1.16
r146 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r147 51 53 23.2347 $w=3.08e-07 $l=6.25e-07 $layer=LI1_cond $X=1.3 $Y=1.785
+ $X2=1.3 $Y2=1.16
r148 50 53 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=1.3 $Y=0.805
+ $X2=1.3 $Y2=1.16
r149 48 51 7.28659 $w=1.95e-07 $l=1.97636e-07 $layer=LI1_cond $X=1.145 $Y=1.882
+ $X2=1.3 $Y2=1.785
r150 48 49 44.0793 $w=1.93e-07 $l=7.75e-07 $layer=LI1_cond $X=1.145 $Y=1.882
+ $X2=0.37 $Y2=1.882
r151 46 50 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=1.145 $Y=0.72
+ $X2=1.3 $Y2=0.805
r152 46 47 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.145 $Y=0.72
+ $X2=0.345 $Y2=0.72
r153 42 49 7.13288 $w=1.95e-07 $l=1.85642e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.37 $Y2=1.882
r154 42 44 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.227 $Y=1.98
+ $X2=0.227 $Y2=2.275
r155 38 47 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r156 38 40 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.46
r157 30 36 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.755 $Y=1.295
+ $X2=3.755 $Y2=1.985
r158 30 32 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.755 $Y=1.025
+ $X2=3.755 $Y2=0.56
r159 22 30 73.3478 $w=2.76e-07 $l=4.2e-07 $layer=POLY_cond $X=3.335 $Y=1.16
+ $X2=3.755 $Y2=1.16
r160 22 57 37.5471 $w=2.76e-07 $l=2.15e-07 $layer=POLY_cond $X=3.335 $Y=1.16
+ $X2=3.12 $Y2=1.16
r161 22 28 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.335 $Y=1.295
+ $X2=3.335 $Y2=1.985
r162 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.335 $Y=1.025
+ $X2=3.335 $Y2=0.56
r163 14 57 35.8007 $w=2.76e-07 $l=2.05e-07 $layer=POLY_cond $X=2.915 $Y=1.16
+ $X2=3.12 $Y2=1.16
r164 14 63 73.3478 $w=2.76e-07 $l=4.2e-07 $layer=POLY_cond $X=2.915 $Y=1.16
+ $X2=2.495 $Y2=1.16
r165 14 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.915 $Y=1.295
+ $X2=2.915 $Y2=1.985
r166 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.915 $Y=1.025
+ $X2=2.915 $Y2=0.56
r167 10 63 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.325
+ $X2=2.495 $Y2=1.16
r168 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.495 $Y=1.325
+ $X2=2.495 $Y2=1.985
r169 7 63 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=0.995
+ $X2=2.495 $Y2=1.16
r170 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.495 $Y=0.995
+ $X2=2.495 $Y2=0.56
r171 2 44 600 $w=1.7e-07 $l=8.50206e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.275
r172 1 40 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%A_193_47# 1 2 9 13 17 21 25 29 33 37 39 43
+ 48 50 52 53 54 57 60 72 73
c137 60 0 1.47729e-19 $X=4.365 $Y=1.19
c138 57 0 5.15114e-20 $X=2.065 $Y=1.19
c139 39 0 6.72171e-20 $X=1.625 $Y=2.307
r140 71 73 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=5.225 $Y=1.16
+ $X2=5.435 $Y2=1.16
r141 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.225
+ $Y=1.16 $X2=5.225 $Y2=1.16
r142 69 71 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=5.015 $Y=1.16
+ $X2=5.225 $Y2=1.16
r143 68 69 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.595 $Y=1.16
+ $X2=5.015 $Y2=1.16
r144 66 68 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=4.39 $Y=1.16
+ $X2=4.595 $Y2=1.16
r145 63 66 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=4.175 $Y=1.16
+ $X2=4.39 $Y2=1.16
r146 61 72 47.6909 $w=1.98e-07 $l=8.6e-07 $layer=LI1_cond $X=4.365 $Y=1.175
+ $X2=5.225 $Y2=1.175
r147 61 66 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.39
+ $Y=1.16 $X2=4.39 $Y2=1.16
r148 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.365 $Y=1.19
+ $X2=4.365 $Y2=1.19
r149 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.065 $Y=1.19
+ $X2=2.065 $Y2=1.19
r150 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.21 $Y=1.19
+ $X2=2.065 $Y2=1.19
r151 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.22 $Y=1.19
+ $X2=4.365 $Y2=1.19
r152 53 54 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=4.22 $Y=1.19
+ $X2=2.21 $Y2=1.19
r153 51 57 13.5287 $w=2.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.795 $Y=1.19
+ $X2=2.065 $Y2=1.19
r154 51 52 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=1.19
+ $X2=1.71 $Y2=1.19
r155 49 52 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.71 $Y=1.305
+ $X2=1.71 $Y2=1.19
r156 49 50 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.71 $Y=1.305
+ $X2=1.71 $Y2=2.15
r157 48 52 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.71 $Y=1.075
+ $X2=1.71 $Y2=1.19
r158 47 48 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.71 $Y=0.465
+ $X2=1.71 $Y2=1.075
r159 43 47 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.625 $Y=0.36
+ $X2=1.71 $Y2=0.465
r160 43 45 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=1.625 $Y=0.36
+ $X2=1.18 $Y2=0.36
r161 39 50 7.64049 $w=3.15e-07 $l=1.94921e-07 $layer=LI1_cond $X=1.625 $Y=2.307
+ $X2=1.71 $Y2=2.15
r162 39 41 19.2074 $w=3.13e-07 $l=5.25e-07 $layer=LI1_cond $X=1.625 $Y=2.307
+ $X2=1.1 $Y2=2.307
r163 35 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.435 $Y=1.295
+ $X2=5.435 $Y2=1.16
r164 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.435 $Y=1.295
+ $X2=5.435 $Y2=1.985
r165 31 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.435 $Y=1.025
+ $X2=5.435 $Y2=1.16
r166 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.435 $Y=1.025
+ $X2=5.435 $Y2=0.56
r167 27 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.015 $Y=1.295
+ $X2=5.015 $Y2=1.16
r168 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.015 $Y=1.295
+ $X2=5.015 $Y2=1.985
r169 23 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.015 $Y=1.025
+ $X2=5.015 $Y2=1.16
r170 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.015 $Y=1.025
+ $X2=5.015 $Y2=0.56
r171 19 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.595 $Y=1.295
+ $X2=4.595 $Y2=1.16
r172 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.595 $Y=1.295
+ $X2=4.595 $Y2=1.985
r173 15 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.595 $Y=1.025
+ $X2=4.595 $Y2=1.16
r174 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.595 $Y=1.025
+ $X2=4.595 $Y2=0.56
r175 11 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.175 $Y=1.295
+ $X2=4.175 $Y2=1.16
r176 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.175 $Y=1.295
+ $X2=4.175 $Y2=1.985
r177 7 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.175 $Y=1.025
+ $X2=4.175 $Y2=1.16
r178 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.175 $Y=1.025
+ $X2=4.175 $Y2=0.56
r179 2 41 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.33
r180 1 45 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.18 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%C 3 7 11 15 19 23 27 31 33 34 35 36 41 51
+ 52
r82 50 52 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=7.745 $Y=1.16
+ $X2=7.955 $Y2=1.16
r83 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.745
+ $Y=1.16 $X2=7.745 $Y2=1.16
r84 48 50 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=7.535 $Y=1.16
+ $X2=7.745 $Y2=1.16
r85 47 48 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.115 $Y=1.16
+ $X2=7.535 $Y2=1.16
r86 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.695 $Y=1.16
+ $X2=7.115 $Y2=1.16
r87 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.455
+ $Y=1.16 $X2=6.455 $Y2=1.16
r88 41 46 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.62 $Y=1.16
+ $X2=6.695 $Y2=1.16
r89 41 43 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.62 $Y=1.16
+ $X2=6.455 $Y2=1.16
r90 36 51 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=7.585 $Y=1.175
+ $X2=7.745 $Y2=1.175
r91 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=7.125 $Y=1.175
+ $X2=7.585 $Y2=1.175
r92 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.665 $Y=1.175
+ $X2=7.125 $Y2=1.175
r93 34 44 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=6.665 $Y=1.175
+ $X2=6.455 $Y2=1.175
r94 33 44 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=6.205 $Y=1.175
+ $X2=6.455 $Y2=1.175
r95 29 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.955 $Y=1.295
+ $X2=7.955 $Y2=1.16
r96 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.955 $Y=1.295
+ $X2=7.955 $Y2=1.985
r97 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.955 $Y=1.025
+ $X2=7.955 $Y2=1.16
r98 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.955 $Y=1.025
+ $X2=7.955 $Y2=0.56
r99 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.535 $Y=1.295
+ $X2=7.535 $Y2=1.16
r100 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.535 $Y=1.295
+ $X2=7.535 $Y2=1.985
r101 17 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.535 $Y=1.025
+ $X2=7.535 $Y2=1.16
r102 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.535 $Y=1.025
+ $X2=7.535 $Y2=0.56
r103 13 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.115 $Y=1.295
+ $X2=7.115 $Y2=1.16
r104 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.115 $Y=1.295
+ $X2=7.115 $Y2=1.985
r105 9 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.115 $Y=1.025
+ $X2=7.115 $Y2=1.16
r106 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.115 $Y=1.025
+ $X2=7.115 $Y2=0.56
r107 5 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.695 $Y=1.295
+ $X2=6.695 $Y2=1.16
r108 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.695 $Y=1.295
+ $X2=6.695 $Y2=1.985
r109 1 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.695 $Y=1.025
+ $X2=6.695 $Y2=1.16
r110 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.695 $Y=1.025
+ $X2=6.695 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%D 3 7 11 15 19 23 27 31 33 34 35 36 41 43
r77 41 52 12.7139 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=9.71 $Y=1.16
+ $X2=9.635 $Y2=1.16
r78 41 43 27.9249 $w=2.9e-07 $l=1.35e-07 $layer=POLY_cond $X=9.71 $Y=1.16
+ $X2=9.845 $Y2=1.16
r79 36 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.845
+ $Y=1.16 $X2=9.845 $Y2=1.16
r80 35 36 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=9.425 $Y=1.175
+ $X2=9.845 $Y2=1.175
r81 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=8.965 $Y=1.175
+ $X2=9.425 $Y2=1.175
r82 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=8.505 $Y=1.175
+ $X2=8.965 $Y2=1.175
r83 33 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.585
+ $Y=1.16 $X2=8.585 $Y2=1.16
r84 29 52 16.6763 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=9.635 $Y=1.305
+ $X2=9.635 $Y2=1.16
r85 29 31 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.635 $Y=1.305
+ $X2=9.635 $Y2=1.985
r86 25 52 16.6763 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=9.635 $Y=1.015
+ $X2=9.635 $Y2=1.16
r87 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.635 $Y=1.015
+ $X2=9.635 $Y2=0.56
r88 17 52 74.4265 $w=2.72e-07 $l=4.2e-07 $layer=POLY_cond $X=9.215 $Y=1.16
+ $X2=9.635 $Y2=1.16
r89 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.215 $Y=1.295
+ $X2=9.215 $Y2=1.985
r90 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.215 $Y=1.025
+ $X2=9.215 $Y2=0.56
r91 9 17 74.4265 $w=2.72e-07 $l=4.2e-07 $layer=POLY_cond $X=8.795 $Y=1.16
+ $X2=9.215 $Y2=1.16
r92 9 48 37.2132 $w=2.72e-07 $l=2.1e-07 $layer=POLY_cond $X=8.795 $Y=1.16
+ $X2=8.585 $Y2=1.16
r93 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.795 $Y=1.295
+ $X2=8.795 $Y2=1.985
r94 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.795 $Y=1.025
+ $X2=8.795 $Y2=0.56
r95 1 48 37.2132 $w=2.72e-07 $l=2.1e-07 $layer=POLY_cond $X=8.375 $Y=1.16
+ $X2=8.585 $Y2=1.16
r96 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.375 $Y=1.295
+ $X2=8.375 $Y2=1.985
r97 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.375 $Y=1.025
+ $X2=8.375 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 47
+ 51 55 59 63 65 69 71 73 77 78 80 81 83 84 85 86 87 89 113 119 122 125 129 135
+ 137 141
r150 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r151 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r152 134 135 11.6744 $w=9.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.32
+ $X2=6.54 $Y2=2.32
r153 131 134 3.08144 $w=9.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.21 $Y=2.32
+ $X2=6.455 $Y2=2.32
r154 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r155 128 131 6.47732 $w=9.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.695 $Y=2.32
+ $X2=6.21 $Y2=2.32
r156 128 129 11.6744 $w=9.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=2.32
+ $X2=5.61 $Y2=2.32
r157 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r158 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r159 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r160 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r161 117 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r162 117 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r163 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r164 114 137 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.09 $Y=2.72
+ $X2=9.005 $Y2=2.72
r165 114 116 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.09 $Y=2.72
+ $X2=9.43 $Y2=2.72
r166 113 140 4.27912 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=9.76 $Y=2.72
+ $X2=9.94 $Y2=2.72
r167 113 116 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.76 $Y=2.72
+ $X2=9.43 $Y2=2.72
r168 112 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r169 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r170 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r171 109 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.21 $Y2=2.72
r172 108 135 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.13 $Y=2.72
+ $X2=6.54 $Y2=2.72
r173 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r174 105 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r175 104 129 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=5.61 $Y2=2.72
r176 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r177 101 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r178 101 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r179 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r180 98 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=2.72
+ $X2=3.965 $Y2=2.72
r181 98 100 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.05 $Y=2.72
+ $X2=4.37 $Y2=2.72
r182 97 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r183 97 120 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r185 94 119 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.652 $Y2=2.72
r186 94 96 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=2.07 $Y2=2.72
r187 89 119 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.652 $Y2=2.72
r188 89 91 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r189 87 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r190 87 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r191 85 111 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=8.08 $Y=2.72
+ $X2=8.05 $Y2=2.72
r192 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.08 $Y=2.72
+ $X2=8.165 $Y2=2.72
r193 83 108 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.24 $Y=2.72
+ $X2=7.13 $Y2=2.72
r194 83 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=2.72
+ $X2=7.325 $Y2=2.72
r195 82 111 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=7.41 $Y=2.72
+ $X2=8.05 $Y2=2.72
r196 82 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=2.72
+ $X2=7.325 $Y2=2.72
r197 80 100 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=4.37 $Y2=2.72
r198 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=4.805 $Y2=2.72
r199 79 104 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.89 $Y=2.72
+ $X2=5.29 $Y2=2.72
r200 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.89 $Y=2.72
+ $X2=4.805 $Y2=2.72
r201 77 96 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.07 $Y2=2.72
r202 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.285 $Y2=2.72
r203 73 76 28.4968 $w=2.73e-07 $l=6.8e-07 $layer=LI1_cond $X=9.897 $Y=1.66
+ $X2=9.897 $Y2=2.34
r204 71 140 3.04293 $w=2.75e-07 $l=1.04307e-07 $layer=LI1_cond $X=9.897 $Y=2.635
+ $X2=9.94 $Y2=2.72
r205 71 76 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=9.897 $Y=2.635
+ $X2=9.897 $Y2=2.34
r206 67 137 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=2.635
+ $X2=9.005 $Y2=2.72
r207 67 69 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.005 $Y=2.635
+ $X2=9.005 $Y2=2
r208 66 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.25 $Y=2.72
+ $X2=8.165 $Y2=2.72
r209 65 137 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.92 $Y=2.72
+ $X2=9.005 $Y2=2.72
r210 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.92 $Y=2.72
+ $X2=8.25 $Y2=2.72
r211 61 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.165 $Y=2.635
+ $X2=8.165 $Y2=2.72
r212 61 63 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.165 $Y=2.635
+ $X2=8.165 $Y2=2
r213 57 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=2.635
+ $X2=7.325 $Y2=2.72
r214 57 59 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.325 $Y=2.635
+ $X2=7.325 $Y2=2
r215 53 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.805 $Y=2.635
+ $X2=4.805 $Y2=2.72
r216 53 55 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.805 $Y=2.635
+ $X2=4.805 $Y2=2
r217 49 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=2.635
+ $X2=3.965 $Y2=2.72
r218 49 51 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.965 $Y=2.635
+ $X2=3.965 $Y2=2
r219 48 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.21 $Y=2.72
+ $X2=3.085 $Y2=2.72
r220 47 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=2.72
+ $X2=3.965 $Y2=2.72
r221 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.88 $Y=2.72
+ $X2=3.21 $Y2=2.72
r222 43 122 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=2.635
+ $X2=3.085 $Y2=2.72
r223 43 45 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.085 $Y=2.635
+ $X2=3.085 $Y2=2
r224 42 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=2.72
+ $X2=2.285 $Y2=2.72
r225 41 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.96 $Y=2.72
+ $X2=3.085 $Y2=2.72
r226 41 42 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.96 $Y=2.72
+ $X2=2.37 $Y2=2.72
r227 37 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.285 $Y=1.66
+ $X2=2.285 $Y2=2.34
r228 35 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=2.635
+ $X2=2.285 $Y2=2.72
r229 35 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.285 $Y=2.635
+ $X2=2.285 $Y2=2.34
r230 31 119 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.652 $Y=2.635
+ $X2=0.652 $Y2=2.72
r231 31 33 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=0.652 $Y=2.635
+ $X2=0.652 $Y2=2.36
r232 10 76 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.71
+ $Y=1.485 $X2=9.845 $Y2=2.34
r233 10 73 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.71
+ $Y=1.485 $X2=9.845 $Y2=1.66
r234 9 69 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.87
+ $Y=1.485 $X2=9.005 $Y2=2
r235 8 63 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.03
+ $Y=1.485 $X2=8.165 $Y2=2
r236 7 59 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.19
+ $Y=1.485 $X2=7.325 $Y2=2
r237 6 134 200 $w=1.7e-07 $l=1.17461e-06 $layer=licon1_PDIFF $count=3 $X=5.51
+ $Y=1.485 $X2=6.455 $Y2=2
r238 6 128 200 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=3 $X=5.51
+ $Y=1.485 $X2=5.695 $Y2=2
r239 5 55 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.67
+ $Y=1.485 $X2=4.805 $Y2=2
r240 4 51 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.83
+ $Y=1.485 $X2=3.965 $Y2=2
r241 3 45 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.99
+ $Y=1.485 $X2=3.125 $Y2=2
r242 2 40 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=1.485 $X2=2.285 $Y2=2.34
r243 2 37 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=1.485 $X2=2.285 $Y2=1.66
r244 1 33 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%Y 1 2 3 4 5 6 7 8 9 10 31 39 41 42 45 49
+ 51 55 57 61 63 67 69 73 75 77 79 81 83 85 87 89 91 94 95 101
c176 101 0 1.25381e-19 $X=3.845 $Y=0.905
r177 95 110 15.7151 $w=2.18e-07 $l=3e-07 $layer=LI1_cond $X=3.845 $Y=1.555
+ $X2=3.545 $Y2=1.555
r178 94 101 3.17836 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=0.78
+ $X2=3.845 $Y2=0.905
r179 94 95 15.2768 $w=4.58e-07 $l=5.25e-07 $layer=LI1_cond $X=3.845 $Y=0.92
+ $X2=3.845 $Y2=1.445
r180 94 101 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=3.845 $Y=0.92
+ $X2=3.845 $Y2=0.905
r181 81 95 8.06961 $w=3.88e-07 $l=2.3e-07 $layer=LI1_cond $X=4.22 $Y=1.555
+ $X2=3.99 $Y2=1.555
r182 81 83 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.22 $Y=1.555
+ $X2=4.385 $Y2=1.555
r183 77 93 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=9.425 $Y=1.665
+ $X2=9.425 $Y2=1.555
r184 77 79 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.425 $Y=1.665
+ $X2=9.425 $Y2=2.34
r185 76 91 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=8.75 $Y=1.555
+ $X2=8.585 $Y2=1.555
r186 75 93 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=9.26 $Y=1.555
+ $X2=9.425 $Y2=1.555
r187 75 76 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=9.26 $Y=1.555
+ $X2=8.75 $Y2=1.555
r188 71 91 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=8.585 $Y=1.665
+ $X2=8.585 $Y2=1.555
r189 71 73 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.585 $Y=1.665
+ $X2=8.585 $Y2=2.34
r190 70 89 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.91 $Y=1.555
+ $X2=7.745 $Y2=1.555
r191 69 91 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=8.42 $Y=1.555
+ $X2=8.585 $Y2=1.555
r192 69 70 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=8.42 $Y=1.555
+ $X2=7.91 $Y2=1.555
r193 65 89 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=7.745 $Y=1.665
+ $X2=7.745 $Y2=1.555
r194 65 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.745 $Y=1.665
+ $X2=7.745 $Y2=2.34
r195 64 87 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.07 $Y=1.555
+ $X2=6.905 $Y2=1.555
r196 63 89 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.58 $Y=1.555
+ $X2=7.745 $Y2=1.555
r197 63 64 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=7.58 $Y=1.555
+ $X2=7.07 $Y2=1.555
r198 59 87 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.905 $Y=1.665
+ $X2=6.905 $Y2=1.555
r199 59 61 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.905 $Y=1.665
+ $X2=6.905 $Y2=2.34
r200 58 85 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.39 $Y=1.555
+ $X2=5.225 $Y2=1.555
r201 57 87 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=1.555
+ $X2=6.905 $Y2=1.555
r202 57 58 70.7181 $w=2.18e-07 $l=1.35e-06 $layer=LI1_cond $X=6.74 $Y=1.555
+ $X2=5.39 $Y2=1.555
r203 53 85 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=5.225 $Y=1.665
+ $X2=5.225 $Y2=1.555
r204 53 55 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.225 $Y=1.665
+ $X2=5.225 $Y2=2.34
r205 52 83 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.55 $Y=1.555
+ $X2=4.385 $Y2=1.555
r206 51 85 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.06 $Y=1.555
+ $X2=5.225 $Y2=1.555
r207 51 52 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=5.06 $Y=1.555
+ $X2=4.55 $Y2=1.555
r208 47 83 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.385 $Y=1.665
+ $X2=4.385 $Y2=1.555
r209 47 49 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.385 $Y=1.665
+ $X2=4.385 $Y2=2.34
r210 45 110 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.545 $Y=2.34
+ $X2=3.545 $Y2=1.665
r211 41 110 8.64332 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=1.555
+ $X2=3.545 $Y2=1.555
r212 41 42 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=3.38 $Y=1.555
+ $X2=2.79 $Y2=1.555
r213 37 42 6.85268 $w=2.2e-07 $l=1.71391e-07 $layer=LI1_cond $X=2.665 $Y=1.665
+ $X2=2.79 $Y2=1.555
r214 37 39 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=2.665 $Y=1.665
+ $X2=2.665 $Y2=1.785
r215 33 36 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=2.705 $Y=0.78
+ $X2=3.545 $Y2=0.78
r216 31 94 3.6869 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=3.7 $Y=0.78
+ $X2=3.845 $Y2=0.78
r217 31 36 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.7 $Y=0.78
+ $X2=3.545 $Y2=0.78
r218 10 93 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.29
+ $Y=1.485 $X2=9.425 $Y2=1.66
r219 10 79 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.29
+ $Y=1.485 $X2=9.425 $Y2=2.34
r220 9 91 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.45
+ $Y=1.485 $X2=8.585 $Y2=1.66
r221 9 73 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.45
+ $Y=1.485 $X2=8.585 $Y2=2.34
r222 8 89 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.61
+ $Y=1.485 $X2=7.745 $Y2=1.66
r223 8 67 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.61
+ $Y=1.485 $X2=7.745 $Y2=2.34
r224 7 87 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.485 $X2=6.905 $Y2=1.66
r225 7 61 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.485 $X2=6.905 $Y2=2.34
r226 6 85 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=1.485 $X2=5.225 $Y2=1.66
r227 6 55 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=1.485 $X2=5.225 $Y2=2.34
r228 5 83 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.25
+ $Y=1.485 $X2=4.385 $Y2=1.66
r229 5 49 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.25
+ $Y=1.485 $X2=4.385 $Y2=2.34
r230 4 110 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.485 $X2=3.545 $Y2=1.66
r231 4 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.485 $X2=3.545 $Y2=2.34
r232 3 39 300 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_PDIFF $count=2 $X=2.57
+ $Y=1.485 $X2=2.705 $Y2=1.785
r233 2 36 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.235 $X2=3.545 $Y2=0.74
r234 1 33 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.235 $X2=2.705 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48
+ 51 54
r102 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r103 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r104 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r105 45 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0 $X2=9.43
+ $Y2=0
r106 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r107 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.59 $Y=0 $X2=9.425
+ $Y2=0
r108 42 44 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.59 $Y=0 $X2=9.89
+ $Y2=0
r109 41 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.43
+ $Y2=0
r110 41 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=8.51
+ $Y2=0
r111 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r112 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.75 $Y=0 $X2=8.585
+ $Y2=0
r113 38 40 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.75 $Y=0 $X2=8.97
+ $Y2=0
r114 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.26 $Y=0 $X2=9.425
+ $Y2=0
r115 37 40 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.26 $Y=0 $X2=8.97
+ $Y2=0
r116 36 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.51
+ $Y2=0
r117 35 36 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r118 33 36 1.96334 $w=4.8e-07 $l=6.9e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=8.05
+ $Y2=0
r119 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r120 32 35 450.16 $w=1.68e-07 $l=6.9e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=8.05
+ $Y2=0
r121 32 33 1.1625 $w=1.7e-07 $l=1.36e-06 $layer=mcon $count=8 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r122 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r123 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r124 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.42 $Y=0 $X2=8.585
+ $Y2=0
r125 29 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.42 $Y=0 $X2=8.05
+ $Y2=0
r126 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r127 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r128 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r129 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r130 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.425 $Y=0.085
+ $X2=9.425 $Y2=0
r131 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=9.425 $Y=0.085
+ $X2=9.425 $Y2=0.4
r132 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.585 $Y=0.085
+ $X2=8.585 $Y2=0
r133 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=8.585 $Y=0.085
+ $X2=8.585 $Y2=0.4
r134 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r135 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r136 3 20 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=9.29
+ $Y=0.235 $X2=9.425 $Y2=0.4
r137 2 16 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.45
+ $Y=0.235 $X2=8.585 $Y2=0.4
r138 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%A_432_47# 1 2 3 4 5 18 20 28
r43 26 28 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=4.805 $Y=0.37
+ $X2=5.645 $Y2=0.37
r44 24 26 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=3.965 $Y=0.37
+ $X2=4.805 $Y2=0.37
r45 22 24 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=3.125 $Y=0.37
+ $X2=3.965 $Y2=0.37
r46 20 22 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=2.37 $Y=0.37
+ $X2=3.125 $Y2=0.37
r47 16 20 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.285 $Y=0.485
+ $X2=2.37 $Y2=0.37
r48 16 18 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.285 $Y=0.485
+ $X2=2.285 $Y2=0.74
r49 5 28 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.51
+ $Y=0.235 $X2=5.645 $Y2=0.4
r50 4 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.235 $X2=4.805 $Y2=0.4
r51 3 24 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.83
+ $Y=0.235 $X2=3.965 $Y2=0.4
r52 2 22 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.235 $X2=3.125 $Y2=0.4
r53 1 18 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=2.16
+ $Y=0.235 $X2=2.285 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%A_850_47# 1 2 3 4 13 19 22 23 27 29
r53 25 27 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=6.905 $Y=0.37
+ $X2=7.745 $Y2=0.37
r54 23 25 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=6.15 $Y=0.37
+ $X2=6.905 $Y2=0.37
r55 21 23 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.065 $Y=0.485
+ $X2=6.15 $Y2=0.37
r56 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.065 $Y=0.485
+ $X2=6.065 $Y2=0.735
r57 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.98 $Y=0.82
+ $X2=6.065 $Y2=0.735
r58 19 29 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.98 $Y=0.82 $X2=5.39
+ $Y2=0.82
r59 15 18 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=4.385 $Y=0.78
+ $X2=5.225 $Y2=0.78
r60 13 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.265 $Y=0.78
+ $X2=5.39 $Y2=0.78
r61 13 18 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=5.265 $Y=0.78
+ $X2=5.225 $Y2=0.78
r62 4 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.61
+ $Y=0.235 $X2=7.745 $Y2=0.4
r63 3 25 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.235 $X2=6.905 $Y2=0.4
r64 2 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.235 $X2=5.225 $Y2=0.74
r65 1 15 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.25
+ $Y=0.235 $X2=4.385 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_4%A_1266_47# 1 2 3 4 5 26
r37 24 26 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=9.005 $Y=0.78
+ $X2=9.845 $Y2=0.78
r38 22 24 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=8.165 $Y=0.78
+ $X2=9.005 $Y2=0.78
r39 20 22 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=7.325 $Y=0.78
+ $X2=8.165 $Y2=0.78
r40 17 20 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=6.485 $Y=0.78
+ $X2=7.325 $Y2=0.78
r41 5 26 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=9.71
+ $Y=0.235 $X2=9.845 $Y2=0.74
r42 4 24 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=8.87
+ $Y=0.235 $X2=9.005 $Y2=0.74
r43 3 22 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=8.03
+ $Y=0.235 $X2=8.165 $Y2=0.74
r44 2 20 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=7.19
+ $Y=0.235 $X2=7.325 $Y2=0.74
r45 1 17 182 $w=1.7e-07 $l=5.77321e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.235 $X2=6.485 $Y2=0.74
.ends


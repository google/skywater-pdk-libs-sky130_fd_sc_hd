* File: sky130_fd_sc_hd__xor3_4.pxi.spice
* Created: Thu Aug 27 14:50:21 2020
* 
x_PM_SKY130_FD_SC_HD__XOR3_4%A_79_21# N_A_79_21#_M1007_d N_A_79_21#_M1010_d
+ N_A_79_21#_c_178_n N_A_79_21#_M1012_g N_A_79_21#_M1000_g N_A_79_21#_c_179_n
+ N_A_79_21#_M1017_g N_A_79_21#_M1003_g N_A_79_21#_c_180_n N_A_79_21#_M1018_g
+ N_A_79_21#_M1016_g N_A_79_21#_c_181_n N_A_79_21#_M1025_g N_A_79_21#_M1023_g
+ N_A_79_21#_c_182_n N_A_79_21#_c_192_n N_A_79_21#_c_198_p N_A_79_21#_c_230_p
+ N_A_79_21#_c_203_p N_A_79_21#_c_183_n N_A_79_21#_c_193_n N_A_79_21#_c_194_n
+ N_A_79_21#_c_195_n N_A_79_21#_c_184_n N_A_79_21#_c_185_n N_A_79_21#_c_209_p
+ N_A_79_21#_c_186_n N_A_79_21#_c_187_n PM_SKY130_FD_SC_HD__XOR3_4%A_79_21#
x_PM_SKY130_FD_SC_HD__XOR3_4%C N_C_c_327_n N_C_M1002_g N_C_c_321_n N_C_M1021_g
+ N_C_c_322_n N_C_M1010_g N_C_c_323_n N_C_M1007_g N_C_c_324_n C N_C_c_325_n
+ N_C_c_326_n PM_SKY130_FD_SC_HD__XOR3_4%C
x_PM_SKY130_FD_SC_HD__XOR3_4%A_480_297# N_A_480_297#_M1021_d
+ N_A_480_297#_M1002_d N_A_480_297#_M1024_g N_A_480_297#_M1026_g
+ N_A_480_297#_c_401_n N_A_480_297#_c_388_n N_A_480_297#_c_394_n
+ N_A_480_297#_c_395_n N_A_480_297#_c_389_n N_A_480_297#_c_390_n
+ N_A_480_297#_c_391_n PM_SKY130_FD_SC_HD__XOR3_4%A_480_297#
x_PM_SKY130_FD_SC_HD__XOR3_4%A_1031_297# N_A_1031_297#_M1027_d
+ N_A_1031_297#_M1005_d N_A_1031_297#_M1004_g N_A_1031_297#_M1014_g
+ N_A_1031_297#_c_466_n N_A_1031_297#_M1009_g N_A_1031_297#_c_468_n
+ N_A_1031_297#_M1022_g N_A_1031_297#_c_469_n N_A_1031_297#_c_470_n
+ N_A_1031_297#_c_483_n N_A_1031_297#_c_471_n N_A_1031_297#_c_472_n
+ N_A_1031_297#_c_487_p N_A_1031_297#_c_473_n N_A_1031_297#_c_474_n
+ N_A_1031_297#_c_475_n N_A_1031_297#_c_476_n N_A_1031_297#_c_477_n
+ N_A_1031_297#_c_478_n PM_SKY130_FD_SC_HD__XOR3_4%A_1031_297#
x_PM_SKY130_FD_SC_HD__XOR3_4%B N_B_M1005_g N_B_M1027_g N_B_c_635_n N_B_c_636_n
+ N_B_M1001_g N_B_M1020_g N_B_c_645_n N_B_c_646_n N_B_M1008_g N_B_M1011_g
+ N_B_c_639_n N_B_c_640_n N_B_c_641_n N_B_c_650_n B N_B_c_642_n
+ PM_SKY130_FD_SC_HD__XOR3_4%B
x_PM_SKY130_FD_SC_HD__XOR3_4%A N_A_M1019_g N_A_M1013_g A N_A_c_754_n N_A_c_755_n
+ N_A_c_756_n PM_SKY130_FD_SC_HD__XOR3_4%A
x_PM_SKY130_FD_SC_HD__XOR3_4%A_1135_365# N_A_1135_365#_M1001_s
+ N_A_1135_365#_M1022_d N_A_1135_365#_M1020_s N_A_1135_365#_M1009_d
+ N_A_1135_365#_M1006_g N_A_1135_365#_M1015_g N_A_1135_365#_c_797_n
+ N_A_1135_365#_c_807_n N_A_1135_365#_c_798_n N_A_1135_365#_c_799_n
+ N_A_1135_365#_c_800_n N_A_1135_365#_c_808_n N_A_1135_365#_c_801_n
+ N_A_1135_365#_c_819_n N_A_1135_365#_c_802_n N_A_1135_365#_c_803_n
+ N_A_1135_365#_c_832_n N_A_1135_365#_c_833_n N_A_1135_365#_c_804_n
+ PM_SKY130_FD_SC_HD__XOR3_4%A_1135_365#
x_PM_SKY130_FD_SC_HD__XOR3_4%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1023_s
+ N_VPWR_M1005_s N_VPWR_M1013_d N_VPWR_c_931_n N_VPWR_c_932_n N_VPWR_c_933_n
+ N_VPWR_c_934_n N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n VPWR
+ N_VPWR_c_938_n N_VPWR_c_939_n N_VPWR_c_940_n N_VPWR_c_941_n N_VPWR_c_942_n
+ N_VPWR_c_930_n N_VPWR_c_944_n N_VPWR_c_945_n N_VPWR_c_946_n N_VPWR_c_947_n
+ N_VPWR_X30_noxref_CONDUCTOR VPWR PM_SKY130_FD_SC_HD__XOR3_4%VPWR
x_PM_SKY130_FD_SC_HD__XOR3_4%X N_X_M1012_s N_X_M1018_s N_X_M1000_d N_X_M1016_d
+ N_X_c_1096_p N_X_c_1081_n N_X_c_1049_n N_X_c_1050_n N_X_c_1051_n N_X_c_1094_p
+ N_X_c_1083_n N_X_c_1052_n X N_X_c_1054_n PM_SKY130_FD_SC_HD__XOR3_4%X
x_PM_SKY130_FD_SC_HD__XOR3_4%A_602_325# N_A_602_325#_M1026_d
+ N_A_602_325#_M1008_d N_A_602_325#_M1010_s N_A_602_325#_M1020_d
+ N_A_602_325#_c_1106_n N_A_602_325#_c_1127_n N_A_602_325#_c_1104_n
+ N_A_602_325#_c_1108_n N_A_602_325#_c_1146_n N_A_602_325#_c_1109_n
+ N_A_602_325#_c_1105_n N_A_602_325#_c_1232_p N_A_602_325#_c_1157_n
+ N_A_602_325#_c_1176_n N_A_602_325#_c_1111_n N_A_602_325#_c_1112_n
+ N_A_602_325#_c_1113_n N_A_602_325#_c_1114_n
+ PM_SKY130_FD_SC_HD__XOR3_4%A_602_325#
x_PM_SKY130_FD_SC_HD__XOR3_4%A_608_49# N_A_608_49#_M1007_s N_A_608_49#_M1001_d
+ N_A_608_49#_M1024_d N_A_608_49#_M1011_d N_A_608_49#_c_1246_n
+ N_A_608_49#_c_1269_n N_A_608_49#_c_1247_n N_A_608_49#_c_1270_n
+ N_A_608_49#_c_1253_n N_A_608_49#_c_1254_n N_A_608_49#_c_1255_n
+ N_A_608_49#_c_1248_n N_A_608_49#_c_1249_n N_A_608_49#_c_1257_n
+ N_A_608_49#_c_1258_n N_A_608_49#_c_1259_n N_A_608_49#_c_1260_n
+ N_A_608_49#_c_1250_n N_A_608_49#_c_1262_n N_A_608_49#_c_1305_n
+ N_A_608_49#_c_1263_n N_A_608_49#_c_1251_n N_A_608_49#_c_1264_n
+ N_A_608_49#_c_1252_n N_A_608_49#_c_1331_n PM_SKY130_FD_SC_HD__XOR3_4%A_608_49#
x_PM_SKY130_FD_SC_HD__XOR3_4%A_1402_49# N_A_1402_49#_M1004_d
+ N_A_1402_49#_M1006_d N_A_1402_49#_M1014_d N_A_1402_49#_M1015_d
+ N_A_1402_49#_c_1425_n N_A_1402_49#_c_1437_n N_A_1402_49#_c_1429_n
+ N_A_1402_49#_c_1426_n N_A_1402_49#_c_1438_n N_A_1402_49#_c_1431_n
+ N_A_1402_49#_c_1427_n PM_SKY130_FD_SC_HD__XOR3_4%A_1402_49#
x_PM_SKY130_FD_SC_HD__XOR3_4%VGND N_VGND_M1012_d N_VGND_M1017_d N_VGND_M1025_d
+ N_VGND_M1027_s N_VGND_M1019_d N_VGND_c_1487_n N_VGND_c_1488_n N_VGND_c_1489_n
+ N_VGND_c_1490_n N_VGND_c_1491_n N_VGND_c_1492_n N_VGND_c_1493_n
+ N_VGND_c_1494_n N_VGND_c_1495_n N_VGND_c_1496_n N_VGND_c_1497_n
+ N_VGND_c_1498_n VGND N_VGND_c_1499_n N_VGND_c_1500_n N_VGND_c_1501_n
+ N_VGND_c_1502_n VGND PM_SKY130_FD_SC_HD__XOR3_4%VGND
cc_1 VNB N_A_79_21#_c_178_n 0.0219679f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_179_n 0.0153756f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_180_n 0.0147974f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_181_n 0.0196823f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_182_n 0.00120878f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_6 VNB N_A_79_21#_c_183_n 7.26786e-19 $X=-0.19 $Y=-0.24 $X2=2.365 $Y2=0.34
cc_7 VNB N_A_79_21#_c_184_n 0.00421536f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=0.865
cc_8 VNB N_A_79_21#_c_185_n 8.29908e-19 $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.325
cc_9 VNB N_A_79_21#_c_186_n 0.0141957f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.355
cc_10 VNB N_A_79_21#_c_187_n 0.0885362f $X=-0.19 $Y=-0.24 $X2=1.83 $Y2=1.16
cc_11 VNB N_C_c_321_n 0.0204568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_C_c_322_n 0.0439409f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_C_c_323_n 0.0215718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_C_c_324_n 0.0154613f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_15 VNB N_C_c_325_n 0.0112837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_C_c_326_n 0.00240757f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_17 VNB N_A_480_297#_c_388_n 0.0024607f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_18 VNB N_A_480_297#_c_389_n 0.00597091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_480_297#_c_390_n 0.0247988f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_20 VNB N_A_480_297#_c_391_n 0.0215524f $X=-0.19 $Y=-0.24 $X2=1.83 $Y2=1.325
cc_21 VNB N_A_1031_297#_M1004_g 0.0355962f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_22 VNB N_A_1031_297#_c_466_n 0.0259644f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_23 VNB N_A_1031_297#_M1009_g 0.00127227f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.325
cc_24 VNB N_A_1031_297#_c_468_n 0.018065f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_25 VNB N_A_1031_297#_c_469_n 0.0291425f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_26 VNB N_A_1031_297#_c_470_n 0.0141001f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_27 VNB N_A_1031_297#_c_471_n 0.0021604f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.077
cc_28 VNB N_A_1031_297#_c_472_n 0.00834501f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.16
cc_29 VNB N_A_1031_297#_c_473_n 0.0124845f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_30 VNB N_A_1031_297#_c_474_n 5.88857e-19 $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.325
cc_31 VNB N_A_1031_297#_c_475_n 0.0027253f $X=-0.19 $Y=-0.24 $X2=2.365 $Y2=0.34
cc_32 VNB N_A_1031_297#_c_476_n 9.00189e-19 $X=-0.19 $Y=-0.24 $X2=2.46 $Y2=2.235
cc_33 VNB N_A_1031_297#_c_477_n 0.00544296f $X=-0.19 $Y=-0.24 $X2=2.545 $Y2=2.32
cc_34 VNB N_A_1031_297#_c_478_n 0.00247748f $X=-0.19 $Y=-0.24 $X2=3.595 $Y2=0.37
cc_35 VNB N_B_M1005_g 0.00410984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_B_M1027_g 0.029876f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_37 VNB N_B_c_635_n 0.0515413f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_38 VNB N_B_c_636_n 0.0167238f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.325
cc_39 VNB N_B_M1001_g 0.0285283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_B_M1020_g 0.00419891f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_41 VNB N_B_c_639_n 0.00493047f $X=-0.19 $Y=-0.24 $X2=1.83 $Y2=1.325
cc_42 VNB N_B_c_640_n 7.60368e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_B_c_641_n 0.0267383f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.077
cc_44 VNB N_B_c_642_n 0.0206335f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.875
cc_45 VNB N_A_c_754_n 0.0201493f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.985
cc_46 VNB N_A_c_755_n 0.00393727f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.985
cc_47 VNB N_A_c_756_n 0.0177121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1135_365#_c_797_n 0.00636967f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_49 VNB N_A_1135_365#_c_798_n 0.00264442f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_50 VNB N_A_1135_365#_c_799_n 0.00179065f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_51 VNB N_A_1135_365#_c_800_n 0.00310506f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_52 VNB N_A_1135_365#_c_801_n 0.0230746f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.213
cc_53 VNB N_A_1135_365#_c_802_n 0.00195542f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_54 VNB N_A_1135_365#_c_803_n 0.00471664f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.875
cc_55 VNB N_A_1135_365#_c_804_n 0.0197295f $X=-0.19 $Y=-0.24 $X2=2.46 $Y2=2.045
cc_56 VNB N_VPWR_c_930_n 0.421552f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_57 VNB N_X_c_1049_n 0.00215131f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_58 VNB N_X_c_1050_n 0.00339489f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_59 VNB N_X_c_1051_n 0.0013034f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.325
cc_60 VNB N_X_c_1052_n 0.00146796f $X=-0.19 $Y=-0.24 $X2=1.83 $Y2=1.985
cc_61 VNB N_A_602_325#_c_1104_n 0.00944527f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_62 VNB N_A_602_325#_c_1105_n 0.00928634f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_63 VNB N_A_608_49#_c_1246_n 0.00251794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_608_49#_c_1247_n 0.00844142f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_65 VNB N_A_608_49#_c_1248_n 0.0131922f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.985
cc_66 VNB N_A_608_49#_c_1249_n 0.00250766f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_67 VNB N_A_608_49#_c_1250_n 0.0023252f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.213
cc_68 VNB N_A_608_49#_c_1251_n 0.0107882f $X=-0.19 $Y=-0.24 $X2=2.545 $Y2=2.32
cc_69 VNB N_A_608_49#_c_1252_n 3.20957e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1402_49#_c_1425_n 0.00783929f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_71 VNB N_A_1402_49#_c_1426_n 0.03052f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.985
cc_72 VNB N_A_1402_49#_c_1427_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.213
cc_73 VNB N_VGND_c_1487_n 0.0110259f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_74 VNB N_VGND_c_1488_n 0.00411685f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.985
cc_75 VNB N_VGND_c_1489_n 3.29525e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_76 VNB N_VGND_c_1490_n 0.00411685f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=1.985
cc_77 VNB N_VGND_c_1491_n 0.00642922f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_78 VNB N_VGND_c_1492_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1493_n 0.0156235f $X=-0.19 $Y=-0.24 $X2=1.932 $Y2=1.16
cc_80 VNB N_VGND_c_1494_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_81 VNB N_VGND_c_1495_n 0.0686407f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.325
cc_82 VNB N_VGND_c_1496_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.875
cc_83 VNB N_VGND_c_1497_n 0.100207f $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=1.96
cc_84 VNB N_VGND_c_1498_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=2.28 $Y2=0.425
cc_85 VNB N_VGND_c_1499_n 0.0156249f $X=-0.19 $Y=-0.24 $X2=2.365 $Y2=0.34
cc_86 VNB N_VGND_c_1500_n 0.0296912f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.16
cc_87 VNB N_VGND_c_1501_n 0.516355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1502_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VPB N_A_79_21#_M1000_g 0.0259656f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.985
cc_90 VPB N_A_79_21#_M1003_g 0.0178265f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_91 VPB N_A_79_21#_M1016_g 0.0174234f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.985
cc_92 VPB N_A_79_21#_M1023_g 0.0200768f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.985
cc_93 VPB N_A_79_21#_c_192_n 0.00142563f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.875
cc_94 VPB N_A_79_21#_c_193_n 0.00374454f $X=-0.19 $Y=1.305 $X2=2.46 $Y2=2.235
cc_95 VPB N_A_79_21#_c_194_n 0.00116793f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=2.32
cc_96 VPB N_A_79_21#_c_195_n 0.012572f $X=-0.19 $Y=1.305 $X2=3.6 $Y2=2.32
cc_97 VPB N_A_79_21#_c_187_n 0.0210648f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.16
cc_98 VPB N_C_c_327_n 0.0326256f $X=-0.19 $Y=1.305 $X2=3.46 $Y2=0.245
cc_99 VPB N_C_c_322_n 0.0194051f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_100 VPB N_C_M1010_g 0.0316695f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.985
cc_101 VPB N_C_c_324_n 8.48743e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_102 VPB N_C_c_325_n 0.00399716f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_C_c_326_n 6.20084e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_104 VPB N_A_480_297#_M1024_g 0.0309169f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_105 VPB N_A_480_297#_c_388_n 0.00355478f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_106 VPB N_A_480_297#_c_394_n 0.0168369f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_107 VPB N_A_480_297#_c_395_n 0.00230347f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_108 VPB N_A_480_297#_c_389_n 9.94335e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_480_297#_c_390_n 0.00516672f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_110 VPB N_A_1031_297#_M1014_g 0.024826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_1031_297#_M1009_g 0.0307087f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.325
cc_112 VPB N_A_1031_297#_c_469_n 0.0105812f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_113 VPB N_A_1031_297#_c_470_n 9.09687e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_114 VPB N_A_1031_297#_c_483_n 0.0079496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_1031_297#_c_478_n 0.00295841f $X=-0.19 $Y=1.305 $X2=3.595
+ $Y2=0.37
cc_116 VPB N_B_M1005_g 0.0262931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_B_M1020_g 0.0236344f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_118 VPB N_B_c_645_n 0.110749f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_119 VPB N_B_c_646_n 0.0129123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_B_M1011_g 0.0314866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_B_c_640_n 9.25804e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_B_c_641_n 0.00514585f $X=-0.19 $Y=1.305 $X2=1.932 $Y2=1.077
cc_123 VPB N_B_c_650_n 0.00168086f $X=-0.19 $Y=1.305 $X2=1.932 $Y2=1.16
cc_124 VPB B 0.00780431f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.16
cc_125 VPB N_A_M1013_g 0.0204714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_c_754_n 0.00439035f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.985
cc_127 VPB N_A_c_755_n 0.00141167f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.985
cc_128 VPB N_A_1135_365#_M1015_g 0.0215569f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_129 VPB N_A_1135_365#_c_797_n 0.00274605f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_130 VPB N_A_1135_365#_c_807_n 0.00177722f $X=-0.19 $Y=1.305 $X2=1.41
+ $Y2=1.325
cc_131 VPB N_A_1135_365#_c_808_n 0.0015591f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.325
cc_132 VPB N_A_1135_365#_c_801_n 0.00472052f $X=-0.19 $Y=1.305 $X2=1.932
+ $Y2=1.213
cc_133 VPB N_VPWR_c_931_n 0.00411685f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.985
cc_134 VPB N_VPWR_c_932_n 3.15634e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_135 VPB N_VPWR_c_933_n 0.00704036f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.985
cc_136 VPB N_VPWR_c_934_n 0.00798922f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_137 VPB N_VPWR_c_935_n 0.00280379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_936_n 0.0108943f $X=-0.19 $Y=1.305 $X2=1.932 $Y2=1.16
cc_139 VPB N_VPWR_c_937_n 0.00324376f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.16
cc_140 VPB N_VPWR_c_938_n 0.015582f $X=-0.19 $Y=1.305 $X2=2.28 $Y2=0.425
cc_141 VPB N_VPWR_c_939_n 0.0119895f $X=-0.19 $Y=1.305 $X2=2.46 $Y2=2.045
cc_142 VPB N_VPWR_c_940_n 0.0609097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_941_n 0.0908898f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_144 VPB N_VPWR_c_942_n 0.0257148f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.16
cc_145 VPB N_VPWR_c_930_n 0.0905617f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.16
cc_146 VPB N_VPWR_c_944_n 0.0043639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_945_n 0.00507404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_946_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_947_n 0.00507043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_X_c_1051_n 0.00111309f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.325
cc_151 VPB N_X_c_1054_n 0.00733254f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.96
cc_152 VPB N_A_602_325#_c_1106_n 0.00424071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_602_325#_c_1104_n 0.00160434f $X=-0.19 $Y=1.305 $X2=1.31
+ $Y2=0.995
cc_154 VPB N_A_602_325#_c_1108_n 0.00264019f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_155 VPB N_A_602_325#_c_1109_n 6.69494e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_602_325#_c_1105_n 0.00210227f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_157 VPB N_A_602_325#_c_1111_n 0.0149758f $X=-0.19 $Y=1.305 $X2=1.932 $Y2=1.16
cc_158 VPB N_A_602_325#_c_1112_n 0.00318498f $X=-0.19 $Y=1.305 $X2=1.905
+ $Y2=1.16
cc_159 VPB N_A_602_325#_c_1113_n 0.00143878f $X=-0.19 $Y=1.305 $X2=2.28
+ $Y2=0.425
cc_160 VPB N_A_602_325#_c_1114_n 0.0205487f $X=-0.19 $Y=1.305 $X2=2.46 $Y2=2.045
cc_161 VPB N_A_608_49#_c_1253_n 0.00262503f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_162 VPB N_A_608_49#_c_1254_n 0.00579762f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_163 VPB N_A_608_49#_c_1255_n 8.62166e-19 $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.325
cc_164 VPB N_A_608_49#_c_1249_n 0.00842441f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_165 VPB N_A_608_49#_c_1257_n 0.00305847f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_166 VPB N_A_608_49#_c_1258_n 0.00300854f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.985
cc_167 VPB N_A_608_49#_c_1259_n 0.0104459f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.985
cc_168 VPB N_A_608_49#_c_1260_n 0.00185607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_608_49#_c_1250_n 0.00156022f $X=-0.19 $Y=1.305 $X2=1.932
+ $Y2=1.213
cc_170 VPB N_A_608_49#_c_1262_n 0.0239398f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.16
cc_171 VPB N_A_608_49#_c_1263_n 0.00221054f $X=-0.19 $Y=1.305 $X2=2.46 $Y2=2.045
cc_172 VPB N_A_608_49#_c_1264_n 2.86933e-19 $X=-0.19 $Y=1.305 $X2=3.6 $Y2=2.32
cc_173 VPB N_A_1402_49#_c_1425_n 0.00467504f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_174 VPB N_A_1402_49#_c_1429_n 0.0141756f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_175 VPB N_A_1402_49#_c_1426_n 0.0226382f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.985
cc_176 VPB N_A_1402_49#_c_1431_n 0.00987855f $X=-0.19 $Y=1.305 $X2=1.83
+ $Y2=1.325
cc_177 N_A_79_21#_M1023_g N_C_c_327_n 0.0289838f $X=1.83 $Y=1.985 $X2=-0.19
+ $Y2=-0.24
cc_178 N_A_79_21#_c_198_p N_C_c_327_n 0.0160133f $X=2.375 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A_79_21#_c_193_n N_C_c_327_n 0.00682238f $X=2.46 $Y=2.235 $X2=-0.19
+ $Y2=-0.24
cc_180 N_A_79_21#_c_194_n N_C_c_327_n 0.00601016f $X=2.545 $Y=2.32 $X2=-0.19
+ $Y2=-0.24
cc_181 N_A_79_21#_c_185_n N_C_c_327_n 0.00441806f $X=1.932 $Y=1.325 $X2=-0.19
+ $Y2=-0.24
cc_182 N_A_79_21#_c_181_n N_C_c_321_n 0.00846978f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_79_21#_c_203_p N_C_c_321_n 0.0110915f $X=2.28 $Y=0.695 $X2=0 $Y2=0
cc_184 N_A_79_21#_c_183_n N_C_c_321_n 0.00168073f $X=2.365 $Y=0.34 $X2=0 $Y2=0
cc_185 N_A_79_21#_c_184_n N_C_c_321_n 0.00723761f $X=1.932 $Y=0.865 $X2=0 $Y2=0
cc_186 N_A_79_21#_c_186_n N_C_c_321_n 0.0106199f $X=3.41 $Y=0.355 $X2=0 $Y2=0
cc_187 N_A_79_21#_c_186_n N_C_c_322_n 0.00677049f $X=3.41 $Y=0.355 $X2=0 $Y2=0
cc_188 N_A_79_21#_c_195_n N_C_M1010_g 0.0100647f $X=3.6 $Y=2.32 $X2=0 $Y2=0
cc_189 N_A_79_21#_c_209_p N_C_c_323_n 0.00326397f $X=3.595 $Y=0.37 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_186_n N_C_c_323_n 0.00805634f $X=3.41 $Y=0.355 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_182_n N_C_c_324_n 0.00441806f $X=1.905 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_184_n N_C_c_324_n 0.00381961f $X=1.932 $Y=0.865 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_187_n N_C_c_324_n 0.0220966f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_79_21#_c_186_n N_C_c_326_n 0.00331115f $X=3.41 $Y=0.355 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_198_p N_A_480_297#_M1002_d 0.00412091f $X=2.375 $Y=1.96
+ $X2=0 $Y2=0
cc_196 N_A_79_21#_c_193_n N_A_480_297#_M1002_d 0.00259446f $X=2.46 $Y=2.235
+ $X2=0 $Y2=0
cc_197 N_A_79_21#_c_195_n N_A_480_297#_M1024_g 0.00829016f $X=3.6 $Y=2.32 $X2=0
+ $Y2=0
cc_198 N_A_79_21#_c_192_n N_A_480_297#_c_401_n 0.00809404f $X=1.96 $Y=1.875
+ $X2=0 $Y2=0
cc_199 N_A_79_21#_c_198_p N_A_480_297#_c_401_n 0.00924302f $X=2.375 $Y=1.96
+ $X2=0 $Y2=0
cc_200 N_A_79_21#_c_195_n N_A_480_297#_c_401_n 0.00596778f $X=3.6 $Y=2.32 $X2=0
+ $Y2=0
cc_201 N_A_79_21#_c_182_n N_A_480_297#_c_388_n 0.01542f $X=1.905 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_79_21#_c_184_n N_A_480_297#_c_388_n 0.00696916f $X=1.932 $Y=0.865
+ $X2=0 $Y2=0
cc_203 N_A_79_21#_c_186_n N_A_480_297#_c_388_n 0.0127861f $X=3.41 $Y=0.355 $X2=0
+ $Y2=0
cc_204 N_A_79_21#_c_187_n N_A_480_297#_c_388_n 2.85707e-19 $X=1.83 $Y=1.16 $X2=0
+ $Y2=0
cc_205 N_A_79_21#_M1010_d N_A_480_297#_c_394_n 0.0030509f $X=3.42 $Y=1.625 $X2=0
+ $Y2=0
cc_206 N_A_79_21#_c_195_n N_A_480_297#_c_394_n 0.00613544f $X=3.6 $Y=2.32 $X2=0
+ $Y2=0
cc_207 N_A_79_21#_c_209_p N_A_480_297#_c_391_n 0.00171346f $X=3.595 $Y=0.37
+ $X2=0 $Y2=0
cc_208 N_A_79_21#_c_192_n N_VPWR_M1023_s 0.00455049f $X=1.96 $Y=1.875 $X2=0
+ $Y2=0
cc_209 N_A_79_21#_c_198_p N_VPWR_M1023_s 0.00712267f $X=2.375 $Y=1.96 $X2=0
+ $Y2=0
cc_210 N_A_79_21#_c_230_p N_VPWR_M1023_s 8.79014e-19 $X=2.045 $Y=1.96 $X2=0
+ $Y2=0
cc_211 N_A_79_21#_M1000_g N_VPWR_c_931_n 0.0030732f $X=0.57 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_79_21#_M1000_g N_VPWR_c_932_n 5.53539e-19 $X=0.57 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A_79_21#_M1003_g N_VPWR_c_932_n 0.00724679f $X=0.99 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_79_21#_M1016_g N_VPWR_c_932_n 0.00706138f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_79_21#_M1023_g N_VPWR_c_932_n 5.20591e-19 $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_79_21#_M1016_g N_VPWR_c_933_n 5.20591e-19 $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_79_21#_M1023_g N_VPWR_c_933_n 0.00816288f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_79_21#_c_198_p N_VPWR_c_933_n 0.0119458f $X=2.375 $Y=1.96 $X2=0 $Y2=0
cc_219 N_A_79_21#_c_230_p N_VPWR_c_933_n 0.00931978f $X=2.045 $Y=1.96 $X2=0
+ $Y2=0
cc_220 N_A_79_21#_c_193_n N_VPWR_c_933_n 0.00147602f $X=2.46 $Y=2.235 $X2=0
+ $Y2=0
cc_221 N_A_79_21#_c_194_n N_VPWR_c_933_n 0.0142636f $X=2.545 $Y=2.32 $X2=0 $Y2=0
cc_222 N_A_79_21#_M1000_g N_VPWR_c_938_n 0.00585385f $X=0.57 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_79_21#_M1003_g N_VPWR_c_938_n 0.00343856f $X=0.99 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_79_21#_M1016_g N_VPWR_c_939_n 0.00343856f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_M1023_g N_VPWR_c_939_n 0.0046653f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A_79_21#_c_198_p N_VPWR_c_940_n 0.00224897f $X=2.375 $Y=1.96 $X2=0
+ $Y2=0
cc_227 N_A_79_21#_c_194_n N_VPWR_c_940_n 0.00859029f $X=2.545 $Y=2.32 $X2=0
+ $Y2=0
cc_228 N_A_79_21#_c_195_n N_VPWR_c_940_n 0.05948f $X=3.6 $Y=2.32 $X2=0 $Y2=0
cc_229 N_A_79_21#_M1000_g N_VPWR_c_930_n 0.0115744f $X=0.57 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_79_21#_M1003_g N_VPWR_c_930_n 0.00402014f $X=0.99 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_79_21#_M1016_g N_VPWR_c_930_n 0.00402014f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_79_21#_M1023_g N_VPWR_c_930_n 0.00789179f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_79_21#_c_198_p N_VPWR_c_930_n 0.00522413f $X=2.375 $Y=1.96 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_c_230_p N_VPWR_c_930_n 7.79838e-19 $X=2.045 $Y=1.96 $X2=0
+ $Y2=0
cc_235 N_A_79_21#_c_194_n N_VPWR_c_930_n 0.00628099f $X=2.545 $Y=2.32 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_c_195_n N_VPWR_c_930_n 0.0478867f $X=3.6 $Y=2.32 $X2=0 $Y2=0
cc_237 N_A_79_21#_c_179_n N_X_c_1049_n 0.015023f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_79_21#_c_187_n N_X_c_1049_n 0.00172753f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_79_21#_c_178_n N_X_c_1050_n 0.00177707f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_79_21#_c_187_n N_X_c_1050_n 0.00424401f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_79_21#_c_179_n N_X_c_1051_n 0.0016611f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_79_21#_M1003_g N_X_c_1051_n 0.00310503f $X=0.99 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_79_21#_c_180_n N_X_c_1051_n 0.00167131f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_79_21#_M1016_g N_X_c_1051_n 0.00328854f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_79_21#_c_181_n N_X_c_1051_n 5.48297e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_79_21#_M1023_g N_X_c_1051_n 3.64492e-19 $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_79_21#_c_182_n N_X_c_1051_n 0.00900539f $X=1.905 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_79_21#_c_192_n N_X_c_1051_n 0.00363351f $X=1.96 $Y=1.875 $X2=0 $Y2=0
cc_249 N_A_79_21#_c_184_n N_X_c_1051_n 0.00590785f $X=1.932 $Y=0.865 $X2=0 $Y2=0
cc_250 N_A_79_21#_c_187_n N_X_c_1051_n 0.0358922f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_79_21#_c_180_n N_X_c_1052_n 0.0113198f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_79_21#_c_181_n N_X_c_1052_n 9.34976e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_79_21#_c_184_n N_X_c_1052_n 0.00490428f $X=1.932 $Y=0.865 $X2=0 $Y2=0
cc_254 N_A_79_21#_c_187_n N_X_c_1052_n 0.00317726f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_79_21#_M1000_g N_X_c_1054_n 0.00139912f $X=0.57 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A_79_21#_M1003_g N_X_c_1054_n 0.0226257f $X=0.99 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A_79_21#_M1016_g N_X_c_1054_n 0.0205164f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_79_21#_M1023_g N_X_c_1054_n 2.84824e-19 $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A_79_21#_c_192_n N_X_c_1054_n 0.0161322f $X=1.96 $Y=1.875 $X2=0 $Y2=0
cc_260 N_A_79_21#_c_187_n N_X_c_1054_n 0.00721115f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_79_21#_c_195_n N_A_602_325#_M1010_s 0.00506904f $X=3.6 $Y=2.32 $X2=0
+ $Y2=0
cc_262 N_A_79_21#_M1010_d N_A_602_325#_c_1106_n 0.00585874f $X=3.42 $Y=1.625
+ $X2=0 $Y2=0
cc_263 N_A_79_21#_c_198_p N_A_602_325#_c_1106_n 0.00822485f $X=2.375 $Y=1.96
+ $X2=0 $Y2=0
cc_264 N_A_79_21#_c_193_n N_A_602_325#_c_1106_n 9.31402e-19 $X=2.46 $Y=2.235
+ $X2=0 $Y2=0
cc_265 N_A_79_21#_c_195_n N_A_602_325#_c_1106_n 0.0580862f $X=3.6 $Y=2.32 $X2=0
+ $Y2=0
cc_266 N_A_79_21#_c_186_n N_A_608_49#_M1007_s 0.00521002f $X=3.41 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_267 N_A_79_21#_M1007_d N_A_608_49#_c_1246_n 0.0113061f $X=3.46 $Y=0.245 $X2=0
+ $Y2=0
cc_268 N_A_79_21#_c_209_p N_A_608_49#_c_1246_n 0.017564f $X=3.595 $Y=0.37 $X2=0
+ $Y2=0
cc_269 N_A_79_21#_c_186_n N_A_608_49#_c_1246_n 0.0188825f $X=3.41 $Y=0.355 $X2=0
+ $Y2=0
cc_270 N_A_79_21#_c_209_p N_A_608_49#_c_1269_n 0.00213283f $X=3.595 $Y=0.37
+ $X2=0 $Y2=0
cc_271 N_A_79_21#_c_209_p N_A_608_49#_c_1270_n 0.0147712f $X=3.595 $Y=0.37 $X2=0
+ $Y2=0
cc_272 N_A_79_21#_c_195_n N_A_608_49#_c_1263_n 0.0117643f $X=3.6 $Y=2.32 $X2=0
+ $Y2=0
cc_273 N_A_79_21#_c_203_p N_VGND_M1025_d 0.00354015f $X=2.28 $Y=0.695 $X2=0
+ $Y2=0
cc_274 N_A_79_21#_c_183_n N_VGND_M1025_d 0.00229493f $X=2.365 $Y=0.34 $X2=0
+ $Y2=0
cc_275 N_A_79_21#_c_184_n N_VGND_M1025_d 0.0175425f $X=1.932 $Y=0.865 $X2=0
+ $Y2=0
cc_276 N_A_79_21#_c_178_n N_VGND_c_1488_n 0.0030732f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_A_79_21#_c_178_n N_VGND_c_1489_n 8.41733e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_A_79_21#_c_179_n N_VGND_c_1489_n 0.00764331f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A_79_21#_c_180_n N_VGND_c_1489_n 0.00764213f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_79_21#_c_181_n N_VGND_c_1489_n 8.41733e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_79_21#_c_187_n N_VGND_c_1489_n 2.50736e-19 $X=1.83 $Y=1.16 $X2=0
+ $Y2=0
cc_282 N_A_79_21#_c_181_n N_VGND_c_1490_n 0.0030732f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_79_21#_c_203_p N_VGND_c_1490_n 0.00722697f $X=2.28 $Y=0.695 $X2=0
+ $Y2=0
cc_284 N_A_79_21#_c_183_n N_VGND_c_1490_n 0.0138309f $X=2.365 $Y=0.34 $X2=0
+ $Y2=0
cc_285 N_A_79_21#_c_184_n N_VGND_c_1490_n 0.0134844f $X=1.932 $Y=0.865 $X2=0
+ $Y2=0
cc_286 N_A_79_21#_c_187_n N_VGND_c_1490_n 7.03008e-19 $X=1.83 $Y=1.16 $X2=0
+ $Y2=0
cc_287 N_A_79_21#_c_180_n N_VGND_c_1493_n 0.00342148f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_79_21#_c_181_n N_VGND_c_1493_n 0.00585385f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_A_79_21#_c_183_n N_VGND_c_1495_n 0.0119943f $X=2.365 $Y=0.34 $X2=0
+ $Y2=0
cc_290 N_A_79_21#_c_184_n N_VGND_c_1495_n 0.00264854f $X=1.932 $Y=0.865 $X2=0
+ $Y2=0
cc_291 N_A_79_21#_c_186_n N_VGND_c_1495_n 0.085762f $X=3.41 $Y=0.355 $X2=0 $Y2=0
cc_292 N_A_79_21#_c_178_n N_VGND_c_1499_n 0.00585385f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_79_21#_c_179_n N_VGND_c_1499_n 0.00342263f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_79_21#_c_178_n N_VGND_c_1501_n 0.0115672f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A_79_21#_c_179_n N_VGND_c_1501_n 0.00403605f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_79_21#_c_180_n N_VGND_c_1501_n 0.00403408f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_79_21#_c_181_n N_VGND_c_1501_n 0.0119391f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_79_21#_c_183_n N_VGND_c_1501_n 0.00652842f $X=2.365 $Y=0.34 $X2=0
+ $Y2=0
cc_299 N_A_79_21#_c_184_n N_VGND_c_1501_n 0.00535855f $X=1.932 $Y=0.865 $X2=0
+ $Y2=0
cc_300 N_A_79_21#_c_186_n N_VGND_c_1501_n 0.0513053f $X=3.41 $Y=0.355 $X2=0
+ $Y2=0
cc_301 N_C_M1010_g N_A_480_297#_M1024_g 0.0343211f $X=3.345 $Y=2.045 $X2=0 $Y2=0
cc_302 N_C_c_325_n N_A_480_297#_M1024_g 9.62949e-19 $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_303 N_C_c_327_n N_A_480_297#_c_401_n 0.00408567f $X=2.325 $Y=1.325 $X2=0
+ $Y2=0
cc_304 N_C_c_322_n N_A_480_297#_c_401_n 0.00196902f $X=3.27 $Y=1.16 $X2=0 $Y2=0
cc_305 N_C_c_327_n N_A_480_297#_c_388_n 0.00401632f $X=2.325 $Y=1.325 $X2=0
+ $Y2=0
cc_306 N_C_c_321_n N_A_480_297#_c_388_n 0.00286897f $X=2.415 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_C_c_322_n N_A_480_297#_c_388_n 0.0220261f $X=3.27 $Y=1.16 $X2=0 $Y2=0
cc_308 N_C_c_323_n N_A_480_297#_c_388_n 0.00307699f $X=3.385 $Y=0.985 $X2=0
+ $Y2=0
cc_309 N_C_c_325_n N_A_480_297#_c_388_n 0.00478624f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_310 N_C_c_326_n N_A_480_297#_c_388_n 0.0248423f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_311 N_C_c_322_n N_A_480_297#_c_394_n 0.0126513f $X=3.27 $Y=1.16 $X2=0 $Y2=0
cc_312 N_C_M1010_g N_A_480_297#_c_394_n 0.0133707f $X=3.345 $Y=2.045 $X2=0 $Y2=0
cc_313 N_C_c_325_n N_A_480_297#_c_394_n 0.00117647f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_314 N_C_c_326_n N_A_480_297#_c_394_n 0.0403344f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_315 N_C_M1010_g N_A_480_297#_c_395_n 0.00345696f $X=3.345 $Y=2.045 $X2=0
+ $Y2=0
cc_316 N_C_c_325_n N_A_480_297#_c_395_n 6.06227e-19 $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_317 N_C_c_325_n N_A_480_297#_c_389_n 0.0010244f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_318 N_C_c_326_n N_A_480_297#_c_389_n 0.0292232f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_319 N_C_c_325_n N_A_480_297#_c_390_n 0.0153962f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_320 N_C_c_326_n N_A_480_297#_c_390_n 0.00111895f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_321 N_C_c_323_n N_A_480_297#_c_391_n 0.0223998f $X=3.385 $Y=0.985 $X2=0 $Y2=0
cc_322 N_C_c_325_n N_A_480_297#_c_391_n 3.54366e-19 $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_323 N_C_c_327_n N_VPWR_c_933_n 0.00188658f $X=2.325 $Y=1.325 $X2=0 $Y2=0
cc_324 N_C_c_327_n N_VPWR_c_940_n 0.00404465f $X=2.325 $Y=1.325 $X2=0 $Y2=0
cc_325 N_C_M1010_g N_VPWR_c_940_n 0.00356303f $X=3.345 $Y=2.045 $X2=0 $Y2=0
cc_326 N_C_c_327_n N_VPWR_c_930_n 0.00522107f $X=2.325 $Y=1.325 $X2=0 $Y2=0
cc_327 N_C_M1010_g N_VPWR_c_930_n 0.00649631f $X=3.345 $Y=2.045 $X2=0 $Y2=0
cc_328 N_C_c_327_n N_A_602_325#_c_1106_n 9.5077e-19 $X=2.325 $Y=1.325 $X2=0
+ $Y2=0
cc_329 N_C_M1010_g N_A_602_325#_c_1106_n 0.00901837f $X=3.345 $Y=2.045 $X2=0
+ $Y2=0
cc_330 N_C_c_322_n N_A_608_49#_c_1246_n 0.00531432f $X=3.27 $Y=1.16 $X2=0 $Y2=0
cc_331 N_C_c_323_n N_A_608_49#_c_1246_n 0.00927259f $X=3.385 $Y=0.985 $X2=0
+ $Y2=0
cc_332 N_C_c_326_n N_A_608_49#_c_1246_n 0.0345339f $X=3.33 $Y=1.16 $X2=0 $Y2=0
cc_333 N_C_c_323_n N_A_608_49#_c_1269_n 7.28465e-19 $X=3.385 $Y=0.985 $X2=0
+ $Y2=0
cc_334 N_C_c_321_n N_VGND_c_1490_n 5.13792e-19 $X=2.415 $Y=0.995 $X2=0 $Y2=0
cc_335 N_C_c_321_n N_VGND_c_1495_n 7.9235e-19 $X=2.415 $Y=0.995 $X2=0 $Y2=0
cc_336 N_C_c_323_n N_VGND_c_1495_n 0.00357877f $X=3.385 $Y=0.985 $X2=0 $Y2=0
cc_337 N_C_c_323_n N_VGND_c_1501_n 0.00696677f $X=3.385 $Y=0.985 $X2=0 $Y2=0
cc_338 N_A_480_297#_M1024_g N_VPWR_c_940_n 0.00369158f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_339 N_A_480_297#_M1024_g N_VPWR_c_930_n 0.00664398f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_340 N_A_480_297#_c_394_n N_A_602_325#_M1010_s 0.00261724f $X=3.685 $Y=1.62
+ $X2=0 $Y2=0
cc_341 N_A_480_297#_M1024_g N_A_602_325#_c_1106_n 0.0137617f $X=3.875 $Y=2.045
+ $X2=0 $Y2=0
cc_342 N_A_480_297#_c_394_n N_A_602_325#_c_1106_n 0.0528429f $X=3.685 $Y=1.62
+ $X2=0 $Y2=0
cc_343 N_A_480_297#_c_389_n N_A_602_325#_c_1106_n 0.00388885f $X=3.875 $Y=1.16
+ $X2=0 $Y2=0
cc_344 N_A_480_297#_c_390_n N_A_602_325#_c_1106_n 0.0010905f $X=3.875 $Y=1.16
+ $X2=0 $Y2=0
cc_345 N_A_480_297#_M1024_g N_A_602_325#_c_1127_n 0.00740594f $X=3.875 $Y=2.045
+ $X2=0 $Y2=0
cc_346 N_A_480_297#_c_394_n N_A_602_325#_c_1127_n 7.49507e-19 $X=3.685 $Y=1.62
+ $X2=0 $Y2=0
cc_347 N_A_480_297#_M1024_g N_A_602_325#_c_1104_n 8.85667e-19 $X=3.875 $Y=2.045
+ $X2=0 $Y2=0
cc_348 N_A_480_297#_c_395_n N_A_602_325#_c_1104_n 0.00180217f $X=3.77 $Y=1.535
+ $X2=0 $Y2=0
cc_349 N_A_480_297#_c_389_n N_A_602_325#_c_1104_n 0.0223427f $X=3.875 $Y=1.16
+ $X2=0 $Y2=0
cc_350 N_A_480_297#_c_390_n N_A_602_325#_c_1104_n 0.00197942f $X=3.875 $Y=1.16
+ $X2=0 $Y2=0
cc_351 N_A_480_297#_c_391_n N_A_602_325#_c_1104_n 0.00661331f $X=3.875 $Y=0.995
+ $X2=0 $Y2=0
cc_352 N_A_480_297#_c_394_n N_A_602_325#_c_1112_n 4.43984e-19 $X=3.685 $Y=1.62
+ $X2=0 $Y2=0
cc_353 N_A_480_297#_c_395_n N_A_602_325#_c_1112_n 6.14306e-19 $X=3.77 $Y=1.535
+ $X2=0 $Y2=0
cc_354 N_A_480_297#_M1024_g N_A_602_325#_c_1114_n 0.00655666f $X=3.875 $Y=2.045
+ $X2=0 $Y2=0
cc_355 N_A_480_297#_c_394_n N_A_602_325#_c_1114_n 0.0135143f $X=3.685 $Y=1.62
+ $X2=0 $Y2=0
cc_356 N_A_480_297#_c_395_n N_A_602_325#_c_1114_n 0.00587493f $X=3.77 $Y=1.535
+ $X2=0 $Y2=0
cc_357 N_A_480_297#_c_389_n N_A_602_325#_c_1114_n 0.00232363f $X=3.875 $Y=1.16
+ $X2=0 $Y2=0
cc_358 N_A_480_297#_c_388_n N_A_608_49#_c_1246_n 0.00976986f $X=2.625 $Y=0.76
+ $X2=0 $Y2=0
cc_359 N_A_480_297#_c_389_n N_A_608_49#_c_1246_n 0.024221f $X=3.875 $Y=1.16
+ $X2=0 $Y2=0
cc_360 N_A_480_297#_c_390_n N_A_608_49#_c_1246_n 0.00280181f $X=3.875 $Y=1.16
+ $X2=0 $Y2=0
cc_361 N_A_480_297#_c_391_n N_A_608_49#_c_1246_n 0.0113781f $X=3.875 $Y=0.995
+ $X2=0 $Y2=0
cc_362 N_A_480_297#_c_391_n N_A_608_49#_c_1269_n 0.00862425f $X=3.875 $Y=0.995
+ $X2=0 $Y2=0
cc_363 N_A_480_297#_c_391_n N_A_608_49#_c_1270_n 0.00716742f $X=3.875 $Y=0.995
+ $X2=0 $Y2=0
cc_364 N_A_480_297#_M1024_g N_A_608_49#_c_1253_n 0.00447876f $X=3.875 $Y=2.045
+ $X2=0 $Y2=0
cc_365 N_A_480_297#_M1024_g N_A_608_49#_c_1255_n 7.78208e-19 $X=3.875 $Y=2.045
+ $X2=0 $Y2=0
cc_366 N_A_480_297#_c_391_n N_A_608_49#_c_1248_n 0.00103799f $X=3.875 $Y=0.995
+ $X2=0 $Y2=0
cc_367 N_A_480_297#_M1024_g N_A_608_49#_c_1263_n 0.00335543f $X=3.875 $Y=2.045
+ $X2=0 $Y2=0
cc_368 N_A_480_297#_c_391_n N_VGND_c_1495_n 0.00390499f $X=3.875 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A_480_297#_c_391_n N_VGND_c_1501_n 0.00727536f $X=3.875 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_1031_297#_c_483_n N_B_M1005_g 0.00527417f $X=5.42 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A_1031_297#_c_478_n N_B_M1005_g 0.00476142f $X=5.455 $Y=0.72 $X2=0
+ $Y2=0
cc_372 N_A_1031_297#_c_487_p N_B_M1027_g 0.00352253f $X=5.535 $Y=0.85 $X2=0
+ $Y2=0
cc_373 N_A_1031_297#_c_478_n N_B_M1027_g 0.01361f $X=5.455 $Y=0.72 $X2=0 $Y2=0
cc_374 N_A_1031_297#_c_472_n N_B_c_635_n 0.00436054f $X=6.625 $Y=0.85 $X2=0
+ $Y2=0
cc_375 N_A_1031_297#_c_478_n N_B_c_635_n 0.0122014f $X=5.455 $Y=0.72 $X2=0 $Y2=0
cc_376 N_A_1031_297#_c_483_n N_B_c_636_n 0.00335249f $X=5.42 $Y=1.58 $X2=0 $Y2=0
cc_377 N_A_1031_297#_c_478_n N_B_c_636_n 0.00330956f $X=5.455 $Y=0.72 $X2=0
+ $Y2=0
cc_378 N_A_1031_297#_M1004_g N_B_M1001_g 0.0114571f $X=6.935 $Y=0.455 $X2=0
+ $Y2=0
cc_379 N_A_1031_297#_c_469_n N_B_M1001_g 0.0209986f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_380 N_A_1031_297#_c_471_n N_B_M1001_g 0.00162996f $X=6.747 $Y=0.995 $X2=0
+ $Y2=0
cc_381 N_A_1031_297#_c_472_n N_B_M1001_g 4.27585e-19 $X=6.625 $Y=0.85 $X2=0
+ $Y2=0
cc_382 N_A_1031_297#_c_474_n N_B_M1001_g 6.64234e-19 $X=6.915 $Y=0.85 $X2=0
+ $Y2=0
cc_383 N_A_1031_297#_c_475_n N_B_M1001_g 0.00115919f $X=6.77 $Y=0.85 $X2=0 $Y2=0
cc_384 N_A_1031_297#_M1014_g N_B_M1020_g 0.0137344f $X=6.935 $Y=1.805 $X2=0
+ $Y2=0
cc_385 N_A_1031_297#_M1014_g N_B_c_645_n 0.00881703f $X=6.935 $Y=1.805 $X2=0
+ $Y2=0
cc_386 N_A_1031_297#_M1009_g N_B_M1011_g 0.0403239f $X=8.325 $Y=2.065 $X2=0
+ $Y2=0
cc_387 N_A_1031_297#_c_466_n N_B_c_640_n 0.00114568f $X=8.325 $Y=1.28 $X2=0
+ $Y2=0
cc_388 N_A_1031_297#_c_473_n N_B_c_640_n 0.00555012f $X=8.005 $Y=0.85 $X2=0
+ $Y2=0
cc_389 N_A_1031_297#_c_477_n N_B_c_640_n 0.0211354f $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_390 N_A_1031_297#_c_466_n N_B_c_641_n 0.0189136f $X=8.325 $Y=1.28 $X2=0 $Y2=0
cc_391 N_A_1031_297#_c_470_n N_B_c_641_n 0.00771356f $X=6.935 $Y=1.16 $X2=0
+ $Y2=0
cc_392 N_A_1031_297#_c_473_n N_B_c_641_n 0.00134545f $X=8.005 $Y=0.85 $X2=0
+ $Y2=0
cc_393 N_A_1031_297#_c_477_n N_B_c_641_n 0.00169113f $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_394 N_A_1031_297#_c_466_n B 8.1069e-19 $X=8.325 $Y=1.28 $X2=0 $Y2=0
cc_395 N_A_1031_297#_M1009_g B 0.00593518f $X=8.325 $Y=2.065 $X2=0 $Y2=0
cc_396 N_A_1031_297#_c_473_n B 0.00414594f $X=8.005 $Y=0.85 $X2=0 $Y2=0
cc_397 N_A_1031_297#_c_476_n B 0.00235209f $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_398 N_A_1031_297#_c_477_n B 0.0183366f $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_399 N_A_1031_297#_M1004_g N_B_c_642_n 0.00771356f $X=6.935 $Y=0.455 $X2=0
+ $Y2=0
cc_400 N_A_1031_297#_c_466_n N_B_c_642_n 0.00163786f $X=8.325 $Y=1.28 $X2=0
+ $Y2=0
cc_401 N_A_1031_297#_c_468_n N_B_c_642_n 0.0180222f $X=8.33 $Y=0.945 $X2=0 $Y2=0
cc_402 N_A_1031_297#_c_473_n N_B_c_642_n 0.00749482f $X=8.005 $Y=0.85 $X2=0
+ $Y2=0
cc_403 N_A_1031_297#_c_476_n N_B_c_642_n 0.00142159f $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_404 N_A_1031_297#_c_477_n N_B_c_642_n 0.00206701f $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_405 N_A_1031_297#_M1009_g N_A_M1013_g 0.0404894f $X=8.325 $Y=2.065 $X2=0
+ $Y2=0
cc_406 N_A_1031_297#_c_466_n N_A_c_754_n 0.0176934f $X=8.325 $Y=1.28 $X2=0 $Y2=0
cc_407 N_A_1031_297#_M1009_g N_A_c_754_n 0.00255062f $X=8.325 $Y=2.065 $X2=0
+ $Y2=0
cc_408 N_A_1031_297#_c_477_n N_A_c_754_n 7.00021e-19 $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_409 N_A_1031_297#_c_466_n N_A_c_755_n 0.00129629f $X=8.325 $Y=1.28 $X2=0
+ $Y2=0
cc_410 N_A_1031_297#_M1009_g N_A_c_755_n 5.31842e-19 $X=8.325 $Y=2.065 $X2=0
+ $Y2=0
cc_411 N_A_1031_297#_c_477_n N_A_c_755_n 0.016109f $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_412 N_A_1031_297#_c_468_n N_A_c_756_n 0.0225611f $X=8.33 $Y=0.945 $X2=0 $Y2=0
cc_413 N_A_1031_297#_c_477_n N_A_c_756_n 2.68453e-19 $X=8.15 $Y=0.85 $X2=0 $Y2=0
cc_414 N_A_1031_297#_c_472_n N_A_1135_365#_M1001_s 9.5256e-19 $X=6.625 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_415 N_A_1031_297#_c_483_n N_A_1135_365#_c_797_n 0.019709f $X=5.42 $Y=1.58
+ $X2=0 $Y2=0
cc_416 N_A_1031_297#_c_472_n N_A_1135_365#_c_797_n 0.0125056f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_417 N_A_1031_297#_c_487_p N_A_1135_365#_c_797_n 6.70277e-19 $X=5.535 $Y=0.85
+ $X2=0 $Y2=0
cc_418 N_A_1031_297#_c_478_n N_A_1135_365#_c_797_n 0.0609172f $X=5.455 $Y=0.72
+ $X2=0 $Y2=0
cc_419 N_A_1031_297#_M1009_g N_A_1135_365#_c_807_n 0.00235326f $X=8.325 $Y=2.065
+ $X2=0 $Y2=0
cc_420 N_A_1031_297#_c_468_n N_A_1135_365#_c_799_n 0.00164439f $X=8.33 $Y=0.945
+ $X2=0 $Y2=0
cc_421 N_A_1031_297#_c_476_n N_A_1135_365#_c_799_n 0.00485657f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_422 N_A_1031_297#_c_477_n N_A_1135_365#_c_799_n 0.00616889f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_423 N_A_1031_297#_M1004_g N_A_1135_365#_c_819_n 0.00602851f $X=6.935 $Y=0.455
+ $X2=0 $Y2=0
cc_424 N_A_1031_297#_c_468_n N_A_1135_365#_c_819_n 0.00716191f $X=8.33 $Y=0.945
+ $X2=0 $Y2=0
cc_425 N_A_1031_297#_c_471_n N_A_1135_365#_c_819_n 3.7129e-19 $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_426 N_A_1031_297#_c_472_n N_A_1135_365#_c_819_n 0.049102f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_427 N_A_1031_297#_c_473_n N_A_1135_365#_c_819_n 0.0873524f $X=8.005 $Y=0.85
+ $X2=0 $Y2=0
cc_428 N_A_1031_297#_c_474_n N_A_1135_365#_c_819_n 0.0265257f $X=6.915 $Y=0.85
+ $X2=0 $Y2=0
cc_429 N_A_1031_297#_c_475_n N_A_1135_365#_c_819_n 0.00319269f $X=6.77 $Y=0.85
+ $X2=0 $Y2=0
cc_430 N_A_1031_297#_c_476_n N_A_1135_365#_c_819_n 0.0265508f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_431 N_A_1031_297#_c_477_n N_A_1135_365#_c_819_n 0.00472786f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_432 N_A_1031_297#_c_472_n N_A_1135_365#_c_802_n 0.0261136f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_433 N_A_1031_297#_c_478_n N_A_1135_365#_c_802_n 0.00675389f $X=5.455 $Y=0.72
+ $X2=0 $Y2=0
cc_434 N_A_1031_297#_c_472_n N_A_1135_365#_c_803_n 0.00122177f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_435 N_A_1031_297#_c_478_n N_A_1135_365#_c_803_n 0.0117267f $X=5.455 $Y=0.72
+ $X2=0 $Y2=0
cc_436 N_A_1031_297#_c_468_n N_A_1135_365#_c_832_n 0.00153367f $X=8.33 $Y=0.945
+ $X2=0 $Y2=0
cc_437 N_A_1031_297#_c_468_n N_A_1135_365#_c_833_n 0.0077529f $X=8.33 $Y=0.945
+ $X2=0 $Y2=0
cc_438 N_A_1031_297#_M1009_g N_VPWR_c_941_n 0.00362032f $X=8.325 $Y=2.065 $X2=0
+ $Y2=0
cc_439 N_A_1031_297#_M1005_d N_VPWR_c_930_n 0.00286702f $X=5.155 $Y=1.485 $X2=0
+ $Y2=0
cc_440 N_A_1031_297#_M1009_g N_VPWR_c_930_n 0.00570414f $X=8.325 $Y=2.065 $X2=0
+ $Y2=0
cc_441 N_A_1031_297#_c_473_n N_A_602_325#_M1008_d 0.00109392f $X=8.005 $Y=0.85
+ $X2=0 $Y2=0
cc_442 N_A_1031_297#_c_476_n N_A_602_325#_M1008_d 7.4435e-19 $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_443 N_A_1031_297#_c_477_n N_A_602_325#_M1008_d 0.00406077f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_444 N_A_1031_297#_c_469_n N_A_602_325#_c_1108_n 0.00894291f $X=6.86 $Y=1.16
+ $X2=0 $Y2=0
cc_445 N_A_1031_297#_c_471_n N_A_602_325#_c_1108_n 0.0270839f $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_446 N_A_1031_297#_c_472_n N_A_602_325#_c_1108_n 5.63647e-19 $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_447 N_A_1031_297#_M1014_g N_A_602_325#_c_1146_n 0.00368795f $X=6.935 $Y=1.805
+ $X2=0 $Y2=0
cc_448 N_A_1031_297#_M1014_g N_A_602_325#_c_1109_n 0.01555f $X=6.935 $Y=1.805
+ $X2=0 $Y2=0
cc_449 N_A_1031_297#_c_469_n N_A_602_325#_c_1109_n 7.42472e-19 $X=6.86 $Y=1.16
+ $X2=0 $Y2=0
cc_450 N_A_1031_297#_c_471_n N_A_602_325#_c_1109_n 0.00152864f $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_451 N_A_1031_297#_c_473_n N_A_602_325#_c_1109_n 0.00288457f $X=8.005 $Y=0.85
+ $X2=0 $Y2=0
cc_452 N_A_1031_297#_c_474_n N_A_602_325#_c_1109_n 6.69145e-19 $X=6.915 $Y=0.85
+ $X2=0 $Y2=0
cc_453 N_A_1031_297#_M1004_g N_A_602_325#_c_1105_n 0.0170984f $X=6.935 $Y=0.455
+ $X2=0 $Y2=0
cc_454 N_A_1031_297#_c_471_n N_A_602_325#_c_1105_n 0.0210201f $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_455 N_A_1031_297#_c_473_n N_A_602_325#_c_1105_n 0.0170211f $X=8.005 $Y=0.85
+ $X2=0 $Y2=0
cc_456 N_A_1031_297#_c_474_n N_A_602_325#_c_1105_n 0.00240264f $X=6.915 $Y=0.85
+ $X2=0 $Y2=0
cc_457 N_A_1031_297#_c_475_n N_A_602_325#_c_1105_n 0.0233729f $X=6.77 $Y=0.85
+ $X2=0 $Y2=0
cc_458 N_A_1031_297#_c_468_n N_A_602_325#_c_1157_n 0.00328526f $X=8.33 $Y=0.945
+ $X2=0 $Y2=0
cc_459 N_A_1031_297#_c_473_n N_A_602_325#_c_1157_n 0.00149151f $X=8.005 $Y=0.85
+ $X2=0 $Y2=0
cc_460 N_A_1031_297#_c_476_n N_A_602_325#_c_1157_n 3.55136e-19 $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_461 N_A_1031_297#_c_477_n N_A_602_325#_c_1157_n 0.00528249f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_462 N_A_1031_297#_c_483_n N_A_602_325#_c_1111_n 0.0236641f $X=5.42 $Y=1.58
+ $X2=0 $Y2=0
cc_463 N_A_1031_297#_c_471_n N_A_602_325#_c_1111_n 8.37577e-19 $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_464 N_A_1031_297#_c_472_n N_A_602_325#_c_1111_n 0.0484178f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_465 N_A_1031_297#_c_487_p N_A_602_325#_c_1111_n 0.0124517f $X=5.535 $Y=0.85
+ $X2=0 $Y2=0
cc_466 N_A_1031_297#_c_478_n N_A_602_325#_c_1111_n 0.00191432f $X=5.455 $Y=0.72
+ $X2=0 $Y2=0
cc_467 N_A_1031_297#_M1014_g N_A_602_325#_c_1113_n 0.00414596f $X=6.935 $Y=1.805
+ $X2=0 $Y2=0
cc_468 N_A_1031_297#_c_469_n N_A_602_325#_c_1113_n 0.00431105f $X=6.86 $Y=1.16
+ $X2=0 $Y2=0
cc_469 N_A_1031_297#_c_471_n N_A_602_325#_c_1113_n 0.00243787f $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_470 N_A_1031_297#_c_474_n N_A_602_325#_c_1113_n 0.0153495f $X=6.915 $Y=0.85
+ $X2=0 $Y2=0
cc_471 N_A_1031_297#_c_472_n N_A_608_49#_M1001_d 0.00139415f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_472 N_A_1031_297#_c_474_n N_A_608_49#_M1001_d 5.07779e-19 $X=6.915 $Y=0.85
+ $X2=0 $Y2=0
cc_473 N_A_1031_297#_c_475_n N_A_608_49#_M1001_d 0.00574398f $X=6.77 $Y=0.85
+ $X2=0 $Y2=0
cc_474 N_A_1031_297#_c_487_p N_A_608_49#_c_1248_n 0.00200331f $X=5.535 $Y=0.85
+ $X2=0 $Y2=0
cc_475 N_A_1031_297#_c_478_n N_A_608_49#_c_1248_n 0.00355568f $X=5.455 $Y=0.72
+ $X2=0 $Y2=0
cc_476 N_A_1031_297#_c_483_n N_A_608_49#_c_1249_n 0.0142825f $X=5.42 $Y=1.58
+ $X2=0 $Y2=0
cc_477 N_A_1031_297#_c_478_n N_A_608_49#_c_1249_n 0.00999923f $X=5.455 $Y=0.72
+ $X2=0 $Y2=0
cc_478 N_A_1031_297#_M1005_d N_A_608_49#_c_1257_n 0.00530614f $X=5.155 $Y=1.485
+ $X2=0 $Y2=0
cc_479 N_A_1031_297#_c_483_n N_A_608_49#_c_1257_n 0.0250069f $X=5.42 $Y=1.58
+ $X2=0 $Y2=0
cc_480 N_A_1031_297#_M1005_d N_A_608_49#_c_1258_n 0.00285479f $X=5.155 $Y=1.485
+ $X2=0 $Y2=0
cc_481 N_A_1031_297#_M1005_d N_A_608_49#_c_1260_n 0.00268234f $X=5.155 $Y=1.485
+ $X2=0 $Y2=0
cc_482 N_A_1031_297#_M1014_g N_A_608_49#_c_1250_n 0.0018148f $X=6.935 $Y=1.805
+ $X2=0 $Y2=0
cc_483 N_A_1031_297#_c_469_n N_A_608_49#_c_1250_n 7.37003e-19 $X=6.86 $Y=1.16
+ $X2=0 $Y2=0
cc_484 N_A_1031_297#_c_471_n N_A_608_49#_c_1250_n 0.0197915f $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_485 N_A_1031_297#_c_472_n N_A_608_49#_c_1250_n 0.00614388f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_486 N_A_1031_297#_c_474_n N_A_608_49#_c_1250_n 0.00109882f $X=6.915 $Y=0.85
+ $X2=0 $Y2=0
cc_487 N_A_1031_297#_c_475_n N_A_608_49#_c_1250_n 0.00311414f $X=6.77 $Y=0.85
+ $X2=0 $Y2=0
cc_488 N_A_1031_297#_M1014_g N_A_608_49#_c_1262_n 0.00215111f $X=6.935 $Y=1.805
+ $X2=0 $Y2=0
cc_489 N_A_1031_297#_M1009_g N_A_608_49#_c_1262_n 0.00693683f $X=8.325 $Y=2.065
+ $X2=0 $Y2=0
cc_490 N_A_1031_297#_M1004_g N_A_608_49#_c_1305_n 0.00229256f $X=6.935 $Y=0.455
+ $X2=0 $Y2=0
cc_491 N_A_1031_297#_c_475_n N_A_608_49#_c_1305_n 0.00181204f $X=6.77 $Y=0.85
+ $X2=0 $Y2=0
cc_492 N_A_1031_297#_c_478_n N_A_608_49#_c_1251_n 0.0067792f $X=5.455 $Y=0.72
+ $X2=0 $Y2=0
cc_493 N_A_1031_297#_c_469_n N_A_608_49#_c_1252_n 2.22283e-19 $X=6.86 $Y=1.16
+ $X2=0 $Y2=0
cc_494 N_A_1031_297#_c_471_n N_A_608_49#_c_1252_n 0.00265833f $X=6.747 $Y=0.995
+ $X2=0 $Y2=0
cc_495 N_A_1031_297#_c_472_n N_A_608_49#_c_1252_n 0.0150436f $X=6.625 $Y=0.85
+ $X2=0 $Y2=0
cc_496 N_A_1031_297#_c_474_n N_A_608_49#_c_1252_n 0.0013346f $X=6.915 $Y=0.85
+ $X2=0 $Y2=0
cc_497 N_A_1031_297#_c_475_n N_A_608_49#_c_1252_n 0.014091f $X=6.77 $Y=0.85
+ $X2=0 $Y2=0
cc_498 N_A_1031_297#_c_473_n N_A_1402_49#_M1004_d 0.00166227f $X=8.005 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_499 N_A_1031_297#_M1014_g N_A_1402_49#_c_1425_n 0.00785518f $X=6.935 $Y=1.805
+ $X2=0 $Y2=0
cc_500 N_A_1031_297#_c_473_n N_A_1402_49#_c_1425_n 0.0179438f $X=8.005 $Y=0.85
+ $X2=0 $Y2=0
cc_501 N_A_1031_297#_c_476_n N_A_1402_49#_c_1425_n 0.00214961f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_502 N_A_1031_297#_c_477_n N_A_1402_49#_c_1425_n 0.00583126f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_503 N_A_1031_297#_M1014_g N_A_1402_49#_c_1437_n 0.00421122f $X=6.935 $Y=1.805
+ $X2=0 $Y2=0
cc_504 N_A_1031_297#_M1009_g N_A_1402_49#_c_1438_n 0.0138456f $X=8.325 $Y=2.065
+ $X2=0 $Y2=0
cc_505 N_A_1031_297#_c_477_n N_A_1402_49#_c_1438_n 0.00161448f $X=8.15 $Y=0.85
+ $X2=0 $Y2=0
cc_506 N_A_1031_297#_c_487_p N_VGND_c_1491_n 0.00444564f $X=5.535 $Y=0.85 $X2=0
+ $Y2=0
cc_507 N_A_1031_297#_M1004_g N_VGND_c_1497_n 0.00575161f $X=6.935 $Y=0.455 $X2=0
+ $Y2=0
cc_508 N_A_1031_297#_c_468_n N_VGND_c_1497_n 0.00585385f $X=8.33 $Y=0.945 $X2=0
+ $Y2=0
cc_509 N_A_1031_297#_c_475_n N_VGND_c_1497_n 0.00316593f $X=6.77 $Y=0.85 $X2=0
+ $Y2=0
cc_510 N_A_1031_297#_c_477_n N_VGND_c_1497_n 7.70543e-19 $X=8.15 $Y=0.85 $X2=0
+ $Y2=0
cc_511 N_A_1031_297#_c_478_n N_VGND_c_1497_n 0.0072215f $X=5.455 $Y=0.72 $X2=0
+ $Y2=0
cc_512 N_A_1031_297#_M1027_d N_VGND_c_1501_n 0.00194539f $X=5.32 $Y=0.235 $X2=0
+ $Y2=0
cc_513 N_A_1031_297#_M1004_g N_VGND_c_1501_n 0.00663327f $X=6.935 $Y=0.455 $X2=0
+ $Y2=0
cc_514 N_A_1031_297#_c_468_n N_VGND_c_1501_n 0.00607914f $X=8.33 $Y=0.945 $X2=0
+ $Y2=0
cc_515 N_A_1031_297#_c_472_n N_VGND_c_1501_n 0.00899211f $X=6.625 $Y=0.85 $X2=0
+ $Y2=0
cc_516 N_A_1031_297#_c_487_p N_VGND_c_1501_n 0.0148507f $X=5.535 $Y=0.85 $X2=0
+ $Y2=0
cc_517 N_A_1031_297#_c_478_n N_VGND_c_1501_n 0.00376241f $X=5.455 $Y=0.72 $X2=0
+ $Y2=0
cc_518 B N_A_M1013_g 2.12214e-19 $X=8.065 $Y=1.445 $X2=0 $Y2=0
cc_519 N_B_c_640_n N_A_c_755_n 0.00135728f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_520 N_B_M1005_g N_A_1135_365#_c_797_n 0.00405425f $X=5.08 $Y=1.985 $X2=0
+ $Y2=0
cc_521 N_B_M1027_g N_A_1135_365#_c_797_n 0.00120086f $X=5.245 $Y=0.56 $X2=0
+ $Y2=0
cc_522 N_B_c_635_n N_A_1135_365#_c_797_n 0.0146445f $X=6.1 $Y=1.16 $X2=0 $Y2=0
cc_523 N_B_M1001_g N_A_1135_365#_c_797_n 0.00472628f $X=6.175 $Y=0.565 $X2=0
+ $Y2=0
cc_524 N_B_M1020_g N_A_1135_365#_c_797_n 0.00560683f $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_525 B N_A_1135_365#_c_807_n 0.0103993f $X=8.065 $Y=1.445 $X2=0 $Y2=0
cc_526 N_B_M1001_g N_A_1135_365#_c_819_n 0.00165623f $X=6.175 $Y=0.565 $X2=0
+ $Y2=0
cc_527 N_B_c_642_n N_A_1135_365#_c_819_n 0.00325031f $X=7.79 $Y=0.995 $X2=0
+ $Y2=0
cc_528 N_B_M1027_g N_A_1135_365#_c_802_n 4.1997e-19 $X=5.245 $Y=0.56 $X2=0 $Y2=0
cc_529 N_B_M1001_g N_A_1135_365#_c_802_n 9.47409e-19 $X=6.175 $Y=0.565 $X2=0
+ $Y2=0
cc_530 N_B_M1027_g N_A_1135_365#_c_803_n 0.00326325f $X=5.245 $Y=0.56 $X2=0
+ $Y2=0
cc_531 N_B_c_635_n N_A_1135_365#_c_803_n 0.00234074f $X=6.1 $Y=1.16 $X2=0 $Y2=0
cc_532 N_B_M1001_g N_A_1135_365#_c_803_n 0.00457137f $X=6.175 $Y=0.565 $X2=0
+ $Y2=0
cc_533 N_B_M1005_g N_VPWR_c_934_n 0.0112156f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_534 N_B_M1005_g N_VPWR_c_941_n 0.00341689f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_535 N_B_c_646_n N_VPWR_c_941_n 0.0381737f $X=6.25 $Y=2.54 $X2=0 $Y2=0
cc_536 N_B_M1005_g N_VPWR_c_930_n 0.00540327f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_537 N_B_c_645_n N_VPWR_c_930_n 0.0391964f $X=7.735 $Y=2.54 $X2=0 $Y2=0
cc_538 N_B_c_646_n N_VPWR_c_930_n 0.0059249f $X=6.25 $Y=2.54 $X2=0 $Y2=0
cc_539 N_B_M1020_g N_A_602_325#_c_1108_n 0.00130858f $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_540 N_B_M1020_g N_A_602_325#_c_1146_n 0.00396146f $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_541 N_B_c_642_n N_A_602_325#_c_1105_n 0.0026019f $X=7.79 $Y=0.995 $X2=0 $Y2=0
cc_542 N_B_c_640_n N_A_602_325#_c_1157_n 0.00216976f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_543 N_B_c_641_n N_A_602_325#_c_1157_n 0.00134398f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_544 N_B_c_642_n N_A_602_325#_c_1157_n 0.00498906f $X=7.79 $Y=0.995 $X2=0
+ $Y2=0
cc_545 N_B_c_642_n N_A_602_325#_c_1176_n 0.00521263f $X=7.79 $Y=0.995 $X2=0
+ $Y2=0
cc_546 N_B_M1005_g N_A_602_325#_c_1111_n 0.00511313f $X=5.08 $Y=1.985 $X2=0
+ $Y2=0
cc_547 N_B_c_635_n N_A_602_325#_c_1111_n 0.0041572f $X=6.1 $Y=1.16 $X2=0 $Y2=0
cc_548 N_B_M1020_g N_A_602_325#_c_1111_n 0.00184208f $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_549 N_B_M1020_g N_A_602_325#_c_1113_n 4.42823e-19 $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_550 N_B_M1005_g N_A_608_49#_c_1253_n 0.00287704f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_551 N_B_M1027_g N_A_608_49#_c_1248_n 0.00325845f $X=5.245 $Y=0.56 $X2=0 $Y2=0
cc_552 N_B_c_636_n N_A_608_49#_c_1249_n 0.0176408f $X=5.32 $Y=1.16 $X2=0 $Y2=0
cc_553 N_B_M1005_g N_A_608_49#_c_1257_n 0.0156612f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_554 N_B_M1005_g N_A_608_49#_c_1258_n 0.00631689f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_555 N_B_M1020_g N_A_608_49#_c_1258_n 9.23301e-19 $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_556 N_B_M1005_g N_A_608_49#_c_1260_n 0.00361658f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_557 N_B_c_635_n N_A_608_49#_c_1250_n 0.00249998f $X=6.1 $Y=1.16 $X2=0 $Y2=0
cc_558 N_B_M1001_g N_A_608_49#_c_1250_n 0.00670076f $X=6.175 $Y=0.565 $X2=0
+ $Y2=0
cc_559 N_B_M1020_g N_A_608_49#_c_1250_n 0.0381078f $X=6.175 $Y=1.905 $X2=0 $Y2=0
cc_560 N_B_c_639_n N_A_608_49#_c_1250_n 0.0027414f $X=6.175 $Y=1.16 $X2=0 $Y2=0
cc_561 N_B_M1020_g N_A_608_49#_c_1262_n 0.00411041f $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_562 N_B_c_645_n N_A_608_49#_c_1262_n 0.0278445f $X=7.735 $Y=2.54 $X2=0 $Y2=0
cc_563 N_B_M1011_g N_A_608_49#_c_1262_n 0.0122992f $X=7.81 $Y=1.965 $X2=0 $Y2=0
cc_564 N_B_M1001_g N_A_608_49#_c_1305_n 5.18677e-19 $X=6.175 $Y=0.565 $X2=0
+ $Y2=0
cc_565 N_B_M1027_g N_A_608_49#_c_1251_n 9.56267e-19 $X=5.245 $Y=0.56 $X2=0 $Y2=0
cc_566 N_B_c_636_n N_A_608_49#_c_1251_n 0.00382072f $X=5.32 $Y=1.16 $X2=0 $Y2=0
cc_567 N_B_M1001_g N_A_608_49#_c_1252_n 0.0108816f $X=6.175 $Y=0.565 $X2=0 $Y2=0
cc_568 N_B_M1020_g N_A_608_49#_c_1331_n 0.00778069f $X=6.175 $Y=1.905 $X2=0
+ $Y2=0
cc_569 N_B_M1011_g N_A_1402_49#_c_1425_n 0.0107026f $X=7.81 $Y=1.965 $X2=0 $Y2=0
cc_570 N_B_c_640_n N_A_1402_49#_c_1425_n 0.0325983f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_571 N_B_c_650_n N_A_1402_49#_c_1425_n 0.0141708f $X=7.875 $Y=1.53 $X2=0 $Y2=0
cc_572 N_B_c_642_n N_A_1402_49#_c_1425_n 0.0103225f $X=7.79 $Y=0.995 $X2=0 $Y2=0
cc_573 N_B_M1011_g N_A_1402_49#_c_1438_n 0.0096343f $X=7.81 $Y=1.965 $X2=0 $Y2=0
cc_574 N_B_c_641_n N_A_1402_49#_c_1438_n 0.00103367f $X=7.79 $Y=1.16 $X2=0 $Y2=0
cc_575 N_B_c_650_n N_A_1402_49#_c_1438_n 0.00720786f $X=7.875 $Y=1.53 $X2=0
+ $Y2=0
cc_576 B N_A_1402_49#_c_1438_n 0.0164129f $X=8.065 $Y=1.445 $X2=0 $Y2=0
cc_577 N_B_M1027_g N_VGND_c_1491_n 0.00438629f $X=5.245 $Y=0.56 $X2=0 $Y2=0
cc_578 N_B_c_636_n N_VGND_c_1491_n 0.00519988f $X=5.32 $Y=1.16 $X2=0 $Y2=0
cc_579 N_B_M1027_g N_VGND_c_1497_n 0.00560495f $X=5.245 $Y=0.56 $X2=0 $Y2=0
cc_580 N_B_M1001_g N_VGND_c_1497_n 0.00414252f $X=6.175 $Y=0.565 $X2=0 $Y2=0
cc_581 N_B_c_642_n N_VGND_c_1497_n 0.00357877f $X=7.79 $Y=0.995 $X2=0 $Y2=0
cc_582 N_B_M1027_g N_VGND_c_1501_n 0.0109355f $X=5.245 $Y=0.56 $X2=0 $Y2=0
cc_583 N_B_M1001_g N_VGND_c_1501_n 0.00707752f $X=6.175 $Y=0.565 $X2=0 $Y2=0
cc_584 N_B_c_642_n N_VGND_c_1501_n 0.00596272f $X=7.79 $Y=0.995 $X2=0 $Y2=0
cc_585 N_A_M1013_g N_A_1135_365#_M1015_g 0.0384393f $X=8.83 $Y=1.985 $X2=0 $Y2=0
cc_586 N_A_M1013_g N_A_1135_365#_c_807_n 0.0100313f $X=8.83 $Y=1.985 $X2=0 $Y2=0
cc_587 N_A_c_754_n N_A_1135_365#_c_807_n 0.00302292f $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_588 N_A_c_755_n N_A_1135_365#_c_807_n 0.0269201f $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_589 N_A_c_755_n N_A_1135_365#_c_798_n 0.0106752f $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_590 N_A_c_756_n N_A_1135_365#_c_798_n 0.00868878f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_591 N_A_c_754_n N_A_1135_365#_c_799_n 0.00357599f $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_592 N_A_c_755_n N_A_1135_365#_c_799_n 0.0204454f $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_593 N_A_c_756_n N_A_1135_365#_c_799_n 0.00178341f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_594 N_A_c_754_n N_A_1135_365#_c_800_n 7.09491e-19 $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_595 N_A_c_755_n N_A_1135_365#_c_800_n 0.0206309f $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_596 N_A_c_756_n N_A_1135_365#_c_800_n 0.00351546f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_597 N_A_M1013_g N_A_1135_365#_c_808_n 0.00340346f $X=8.83 $Y=1.985 $X2=0
+ $Y2=0
cc_598 N_A_c_754_n N_A_1135_365#_c_801_n 0.0211645f $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_599 N_A_c_755_n N_A_1135_365#_c_801_n 8.25692e-19 $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_600 N_A_c_755_n N_A_1135_365#_c_832_n 9.51454e-19 $X=8.75 $Y=1.16 $X2=0 $Y2=0
cc_601 N_A_c_756_n N_A_1135_365#_c_833_n 0.00811137f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_602 N_A_c_756_n N_A_1135_365#_c_804_n 0.0209318f $X=8.76 $Y=0.995 $X2=0 $Y2=0
cc_603 N_A_M1013_g N_VPWR_c_935_n 0.00317431f $X=8.83 $Y=1.985 $X2=0 $Y2=0
cc_604 N_A_M1013_g N_VPWR_c_941_n 0.00422112f $X=8.83 $Y=1.985 $X2=0 $Y2=0
cc_605 N_A_M1013_g N_VPWR_c_930_n 0.00591637f $X=8.83 $Y=1.985 $X2=0 $Y2=0
cc_606 N_A_M1013_g N_A_608_49#_c_1262_n 0.00152622f $X=8.83 $Y=1.985 $X2=0 $Y2=0
cc_607 N_A_M1013_g N_A_1402_49#_c_1438_n 0.0126206f $X=8.83 $Y=1.985 $X2=0 $Y2=0
cc_608 N_A_c_756_n N_VGND_c_1492_n 0.00447435f $X=8.76 $Y=0.995 $X2=0 $Y2=0
cc_609 N_A_c_756_n N_VGND_c_1497_n 0.0042601f $X=8.76 $Y=0.995 $X2=0 $Y2=0
cc_610 N_A_c_756_n N_VGND_c_1501_n 0.00622026f $X=8.76 $Y=0.995 $X2=0 $Y2=0
cc_611 N_A_1135_365#_c_807_n N_VPWR_M1013_d 0.00502786f $X=9.105 $Y=1.6 $X2=0
+ $Y2=0
cc_612 N_A_1135_365#_M1015_g N_VPWR_c_935_n 0.0080626f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_613 N_A_1135_365#_M1015_g N_VPWR_c_942_n 0.00337001f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_614 N_A_1135_365#_M1009_d N_VPWR_c_930_n 0.00382772f $X=8.4 $Y=1.645 $X2=0
+ $Y2=0
cc_615 N_A_1135_365#_M1015_g N_VPWR_c_930_n 0.00523175f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_616 N_A_1135_365#_c_819_n N_A_602_325#_M1008_d 0.00332817f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_617 N_A_1135_365#_c_819_n N_A_602_325#_c_1105_n 0.0145847f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_618 N_A_1135_365#_c_819_n N_A_602_325#_c_1157_n 0.0145995f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_619 N_A_1135_365#_c_832_n N_A_602_325#_c_1157_n 0.00126391f $X=8.61 $Y=0.51
+ $X2=0 $Y2=0
cc_620 N_A_1135_365#_c_833_n N_A_602_325#_c_1157_n 0.00765914f $X=8.61 $Y=0.51
+ $X2=0 $Y2=0
cc_621 N_A_1135_365#_c_819_n N_A_602_325#_c_1176_n 0.0119237f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_622 N_A_1135_365#_M1020_s N_A_602_325#_c_1111_n 0.00840572f $X=5.675 $Y=1.825
+ $X2=0 $Y2=0
cc_623 N_A_1135_365#_c_797_n N_A_602_325#_c_1111_n 0.0184168f $X=5.8 $Y=1.94
+ $X2=0 $Y2=0
cc_624 N_A_1135_365#_c_819_n N_A_608_49#_M1001_d 0.00519015f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_625 N_A_1135_365#_c_797_n N_A_608_49#_c_1257_n 0.0138372f $X=5.8 $Y=1.94
+ $X2=0 $Y2=0
cc_626 N_A_1135_365#_c_797_n N_A_608_49#_c_1258_n 0.0028603f $X=5.8 $Y=1.94
+ $X2=0 $Y2=0
cc_627 N_A_1135_365#_M1020_s N_A_608_49#_c_1259_n 0.0100815f $X=5.675 $Y=1.825
+ $X2=0 $Y2=0
cc_628 N_A_1135_365#_c_797_n N_A_608_49#_c_1259_n 0.0128549f $X=5.8 $Y=1.94
+ $X2=0 $Y2=0
cc_629 N_A_1135_365#_c_797_n N_A_608_49#_c_1250_n 0.0619827f $X=5.8 $Y=1.94
+ $X2=0 $Y2=0
cc_630 N_A_1135_365#_M1009_d N_A_608_49#_c_1262_n 0.0024914f $X=8.4 $Y=1.645
+ $X2=0 $Y2=0
cc_631 N_A_1135_365#_c_819_n N_A_608_49#_c_1305_n 0.0121773f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_632 N_A_1135_365#_c_802_n N_A_608_49#_c_1305_n 0.001476f $X=5.995 $Y=0.51
+ $X2=0 $Y2=0
cc_633 N_A_1135_365#_c_803_n N_A_608_49#_c_1305_n 0.00942559f $X=5.85 $Y=0.51
+ $X2=0 $Y2=0
cc_634 N_A_1135_365#_c_797_n N_A_608_49#_c_1252_n 0.0112297f $X=5.8 $Y=1.94
+ $X2=0 $Y2=0
cc_635 N_A_1135_365#_c_819_n N_A_608_49#_c_1252_n 0.00287405f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_636 N_A_1135_365#_c_803_n N_A_608_49#_c_1252_n 0.0022251f $X=5.85 $Y=0.51
+ $X2=0 $Y2=0
cc_637 N_A_1135_365#_c_819_n N_A_1402_49#_M1004_d 0.00653094f $X=8.465 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_638 N_A_1135_365#_c_819_n N_A_1402_49#_c_1425_n 0.00162336f $X=8.465 $Y=0.51
+ $X2=0 $Y2=0
cc_639 N_A_1135_365#_M1015_g N_A_1402_49#_c_1426_n 0.0118718f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_640 N_A_1135_365#_c_807_n N_A_1402_49#_c_1426_n 0.0130582f $X=9.105 $Y=1.6
+ $X2=0 $Y2=0
cc_641 N_A_1135_365#_c_800_n N_A_1402_49#_c_1426_n 0.0400001f $X=9.19 $Y=1.325
+ $X2=0 $Y2=0
cc_642 N_A_1135_365#_c_808_n N_A_1402_49#_c_1426_n 0.00963437f $X=9.19 $Y=1.495
+ $X2=0 $Y2=0
cc_643 N_A_1135_365#_c_801_n N_A_1402_49#_c_1426_n 0.00752814f $X=9.25 $Y=1.16
+ $X2=0 $Y2=0
cc_644 N_A_1135_365#_c_804_n N_A_1402_49#_c_1426_n 0.0100973f $X=9.25 $Y=0.995
+ $X2=0 $Y2=0
cc_645 N_A_1135_365#_M1009_d N_A_1402_49#_c_1438_n 0.00689243f $X=8.4 $Y=1.645
+ $X2=0 $Y2=0
cc_646 N_A_1135_365#_c_807_n N_A_1402_49#_c_1438_n 0.0341401f $X=9.105 $Y=1.6
+ $X2=0 $Y2=0
cc_647 N_A_1135_365#_M1015_g N_A_1402_49#_c_1431_n 0.0123928f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_648 N_A_1135_365#_c_807_n N_A_1402_49#_c_1431_n 0.0046677f $X=9.105 $Y=1.6
+ $X2=0 $Y2=0
cc_649 N_A_1135_365#_c_800_n N_A_1402_49#_c_1431_n 0.0016745f $X=9.19 $Y=1.325
+ $X2=0 $Y2=0
cc_650 N_A_1135_365#_c_798_n N_VGND_M1019_d 0.00176133f $X=9.105 $Y=0.82 $X2=0
+ $Y2=0
cc_651 N_A_1135_365#_c_800_n N_VGND_M1019_d 5.72954e-19 $X=9.19 $Y=1.325 $X2=0
+ $Y2=0
cc_652 N_A_1135_365#_c_802_n N_VGND_c_1491_n 7.53702e-19 $X=5.995 $Y=0.51 $X2=0
+ $Y2=0
cc_653 N_A_1135_365#_c_798_n N_VGND_c_1492_n 0.00851939f $X=9.105 $Y=0.82 $X2=0
+ $Y2=0
cc_654 N_A_1135_365#_c_800_n N_VGND_c_1492_n 0.00459507f $X=9.19 $Y=1.325 $X2=0
+ $Y2=0
cc_655 N_A_1135_365#_c_801_n N_VGND_c_1492_n 2.05208e-19 $X=9.25 $Y=1.16 $X2=0
+ $Y2=0
cc_656 N_A_1135_365#_c_832_n N_VGND_c_1492_n 0.00113301f $X=8.61 $Y=0.51 $X2=0
+ $Y2=0
cc_657 N_A_1135_365#_c_833_n N_VGND_c_1492_n 0.0155694f $X=8.61 $Y=0.51 $X2=0
+ $Y2=0
cc_658 N_A_1135_365#_c_804_n N_VGND_c_1492_n 0.00274672f $X=9.25 $Y=0.995 $X2=0
+ $Y2=0
cc_659 N_A_1135_365#_c_798_n N_VGND_c_1497_n 0.0024589f $X=9.105 $Y=0.82 $X2=0
+ $Y2=0
cc_660 N_A_1135_365#_c_819_n N_VGND_c_1497_n 0.00505812f $X=8.465 $Y=0.51 $X2=0
+ $Y2=0
cc_661 N_A_1135_365#_c_802_n N_VGND_c_1497_n 2.49898e-19 $X=5.995 $Y=0.51 $X2=0
+ $Y2=0
cc_662 N_A_1135_365#_c_803_n N_VGND_c_1497_n 0.024795f $X=5.85 $Y=0.51 $X2=0
+ $Y2=0
cc_663 N_A_1135_365#_c_832_n N_VGND_c_1497_n 3.63685e-19 $X=8.61 $Y=0.51 $X2=0
+ $Y2=0
cc_664 N_A_1135_365#_c_833_n N_VGND_c_1497_n 0.0143515f $X=8.61 $Y=0.51 $X2=0
+ $Y2=0
cc_665 N_A_1135_365#_c_800_n N_VGND_c_1500_n 0.00123845f $X=9.19 $Y=1.325 $X2=0
+ $Y2=0
cc_666 N_A_1135_365#_c_804_n N_VGND_c_1500_n 0.00526859f $X=9.25 $Y=0.995 $X2=0
+ $Y2=0
cc_667 N_A_1135_365#_M1022_d N_VGND_c_1501_n 0.00190368f $X=8.405 $Y=0.235 $X2=0
+ $Y2=0
cc_668 N_A_1135_365#_c_798_n N_VGND_c_1501_n 0.00531107f $X=9.105 $Y=0.82 $X2=0
+ $Y2=0
cc_669 N_A_1135_365#_c_800_n N_VGND_c_1501_n 0.00298021f $X=9.19 $Y=1.325 $X2=0
+ $Y2=0
cc_670 N_A_1135_365#_c_819_n N_VGND_c_1501_n 0.215427f $X=8.465 $Y=0.51 $X2=0
+ $Y2=0
cc_671 N_A_1135_365#_c_802_n N_VGND_c_1501_n 0.0285546f $X=5.995 $Y=0.51 $X2=0
+ $Y2=0
cc_672 N_A_1135_365#_c_803_n N_VGND_c_1501_n 0.00391709f $X=5.85 $Y=0.51 $X2=0
+ $Y2=0
cc_673 N_A_1135_365#_c_832_n N_VGND_c_1501_n 0.0285254f $X=8.61 $Y=0.51 $X2=0
+ $Y2=0
cc_674 N_A_1135_365#_c_833_n N_VGND_c_1501_n 0.00348354f $X=8.61 $Y=0.51 $X2=0
+ $Y2=0
cc_675 N_A_1135_365#_c_804_n N_VGND_c_1501_n 0.0101408f $X=9.25 $Y=0.995 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_930_n N_X_M1000_d 0.00562358f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_677 N_VPWR_c_930_n N_X_M1016_d 0.00562358f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_678 N_VPWR_c_938_n N_X_c_1081_n 0.0113958f $X=1.035 $Y=2.72 $X2=0 $Y2=0
cc_679 N_VPWR_c_930_n N_X_c_1081_n 0.00646998f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_680 N_VPWR_c_939_n N_X_c_1083_n 0.0113958f $X=1.875 $Y=2.72 $X2=0 $Y2=0
cc_681 N_VPWR_c_930_n N_X_c_1083_n 0.00646998f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_682 N_VPWR_M1003_s N_X_c_1054_n 0.00167227f $X=1.065 $Y=1.485 $X2=0 $Y2=0
cc_683 N_VPWR_c_932_n N_X_c_1054_n 0.0178491f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_684 N_VPWR_c_938_n N_X_c_1054_n 0.00194746f $X=1.035 $Y=2.72 $X2=0 $Y2=0
cc_685 N_VPWR_c_939_n N_X_c_1054_n 0.00195299f $X=1.875 $Y=2.72 $X2=0 $Y2=0
cc_686 N_VPWR_c_930_n N_X_c_1054_n 0.00728868f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_687 N_VPWR_c_940_n N_A_602_325#_c_1106_n 0.00328201f $X=4.705 $Y=2.72 $X2=0
+ $Y2=0
cc_688 N_VPWR_c_930_n N_A_602_325#_c_1106_n 0.00795134f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_689 N_VPWR_M1005_s N_A_602_325#_c_1111_n 0.00100785f $X=4.745 $Y=1.485 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_930_n N_A_608_49#_M1011_d 0.00233026f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_934_n N_A_608_49#_c_1254_n 0.00147971f $X=4.87 $Y=2.32 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_940_n N_A_608_49#_c_1254_n 0.00296166f $X=4.705 $Y=2.72 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_930_n N_A_608_49#_c_1254_n 0.00485654f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_694 N_VPWR_M1005_s N_A_608_49#_c_1249_n 0.00648805f $X=4.745 $Y=1.485 $X2=0
+ $Y2=0
cc_695 N_VPWR_M1005_s N_A_608_49#_c_1257_n 0.00130442f $X=4.745 $Y=1.485 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_934_n N_A_608_49#_c_1257_n 0.00607843f $X=4.87 $Y=2.32 $X2=0
+ $Y2=0
cc_697 N_VPWR_c_941_n N_A_608_49#_c_1257_n 0.00503515f $X=8.915 $Y=2.72 $X2=0
+ $Y2=0
cc_698 N_VPWR_c_930_n N_A_608_49#_c_1257_n 0.00935628f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_934_n N_A_608_49#_c_1258_n 0.00173147f $X=4.87 $Y=2.32 $X2=0
+ $Y2=0
cc_700 N_VPWR_c_941_n N_A_608_49#_c_1259_n 0.0305955f $X=8.915 $Y=2.72 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_930_n N_A_608_49#_c_1259_n 0.0196786f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_934_n N_A_608_49#_c_1260_n 0.00833535f $X=4.87 $Y=2.32 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_941_n N_A_608_49#_c_1260_n 0.0105745f $X=8.915 $Y=2.72 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_930_n N_A_608_49#_c_1260_n 0.00644066f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_705 N_VPWR_c_941_n N_A_608_49#_c_1262_n 0.123059f $X=8.915 $Y=2.72 $X2=0
+ $Y2=0
cc_706 N_VPWR_c_930_n N_A_608_49#_c_1262_n 0.074231f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_707 N_VPWR_c_934_n N_A_608_49#_c_1263_n 0.0142739f $X=4.87 $Y=2.32 $X2=0
+ $Y2=0
cc_708 N_VPWR_c_940_n N_A_608_49#_c_1263_n 0.0186431f $X=4.705 $Y=2.72 $X2=0
+ $Y2=0
cc_709 N_VPWR_c_930_n N_A_608_49#_c_1263_n 0.0145279f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_710 N_VPWR_M1005_s N_A_608_49#_c_1264_n 0.00234468f $X=4.745 $Y=1.485 $X2=0
+ $Y2=0
cc_711 N_VPWR_c_934_n N_A_608_49#_c_1264_n 0.0143988f $X=4.87 $Y=2.32 $X2=0
+ $Y2=0
cc_712 N_VPWR_c_930_n N_A_608_49#_c_1264_n 8.22076e-19 $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_713 N_VPWR_c_941_n N_A_608_49#_c_1331_n 0.010266f $X=8.915 $Y=2.72 $X2=0
+ $Y2=0
cc_714 N_VPWR_c_930_n N_A_608_49#_c_1331_n 0.005802f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_715 N_VPWR_c_930_n N_A_1402_49#_M1015_d 0.00226128f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_716 N_VPWR_c_942_n N_A_1402_49#_c_1429_n 0.0172026f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_717 N_VPWR_c_930_n N_A_1402_49#_c_1429_n 0.00977915f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_718 N_VPWR_M1013_d N_A_1402_49#_c_1438_n 0.00432135f $X=8.905 $Y=1.485 $X2=0
+ $Y2=0
cc_719 N_VPWR_c_935_n N_A_1402_49#_c_1438_n 0.0169172f $X=9.08 $Y=2.36 $X2=0
+ $Y2=0
cc_720 N_VPWR_c_941_n N_A_1402_49#_c_1438_n 0.00751819f $X=8.915 $Y=2.72 $X2=0
+ $Y2=0
cc_721 N_VPWR_c_930_n N_A_1402_49#_c_1438_n 0.0154111f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_722 N_VPWR_c_942_n N_A_1402_49#_c_1431_n 0.00261604f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_723 N_VPWR_c_930_n N_A_1402_49#_c_1431_n 0.00438473f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_724 N_X_c_1049_n N_VGND_M1017_d 9.03344e-19 $X=1.105 $Y=0.792 $X2=0 $Y2=0
cc_725 N_X_c_1052_n N_VGND_M1017_d 8.2611e-19 $X=1.105 $Y=0.66 $X2=0 $Y2=0
cc_726 N_X_c_1049_n N_VGND_c_1489_n 0.00763326f $X=1.105 $Y=0.792 $X2=0 $Y2=0
cc_727 N_X_c_1052_n N_VGND_c_1489_n 0.00746531f $X=1.105 $Y=0.66 $X2=0 $Y2=0
cc_728 N_X_c_1094_p N_VGND_c_1493_n 0.00694438f $X=1.52 $Y=0.56 $X2=0 $Y2=0
cc_729 N_X_c_1052_n N_VGND_c_1493_n 0.00247993f $X=1.105 $Y=0.66 $X2=0 $Y2=0
cc_730 N_X_c_1096_p N_VGND_c_1499_n 0.00697776f $X=0.68 $Y=0.56 $X2=0 $Y2=0
cc_731 N_X_c_1049_n N_VGND_c_1499_n 0.00234972f $X=1.105 $Y=0.792 $X2=0 $Y2=0
cc_732 N_X_M1012_s N_VGND_c_1501_n 0.00419147f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_733 N_X_M1018_s N_VGND_c_1501_n 0.00419074f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_734 N_X_c_1096_p N_VGND_c_1501_n 0.00611294f $X=0.68 $Y=0.56 $X2=0 $Y2=0
cc_735 N_X_c_1049_n N_VGND_c_1501_n 0.00500079f $X=1.105 $Y=0.792 $X2=0 $Y2=0
cc_736 N_X_c_1094_p N_VGND_c_1501_n 0.00609811f $X=1.52 $Y=0.56 $X2=0 $Y2=0
cc_737 N_X_c_1052_n N_VGND_c_1501_n 0.00521842f $X=1.105 $Y=0.66 $X2=0 $Y2=0
cc_738 N_A_602_325#_c_1106_n N_A_608_49#_M1024_d 0.00570726f $X=4.025 $Y=1.98
+ $X2=0 $Y2=0
cc_739 N_A_602_325#_c_1127_n N_A_608_49#_M1024_d 0.00664959f $X=4.11 $Y=1.895
+ $X2=0 $Y2=0
cc_740 N_A_602_325#_c_1114_n N_A_608_49#_M1024_d 0.00687512f $X=4.355 $Y=1.535
+ $X2=0 $Y2=0
cc_741 N_A_602_325#_M1026_d N_A_608_49#_c_1246_n 0.00334341f $X=4.01 $Y=0.245
+ $X2=0 $Y2=0
cc_742 N_A_602_325#_c_1104_n N_A_608_49#_c_1246_n 0.0138308f $X=4.355 $Y=0.76
+ $X2=0 $Y2=0
cc_743 N_A_602_325#_M1026_d N_A_608_49#_c_1269_n 0.00347935f $X=4.01 $Y=0.245
+ $X2=0 $Y2=0
cc_744 N_A_602_325#_c_1104_n N_A_608_49#_c_1269_n 0.00432164f $X=4.355 $Y=0.76
+ $X2=0 $Y2=0
cc_745 N_A_602_325#_M1026_d N_A_608_49#_c_1247_n 0.0175141f $X=4.01 $Y=0.245
+ $X2=0 $Y2=0
cc_746 N_A_602_325#_c_1104_n N_A_608_49#_c_1247_n 0.0128008f $X=4.355 $Y=0.76
+ $X2=0 $Y2=0
cc_747 N_A_602_325#_M1026_d N_A_608_49#_c_1270_n 3.2099e-19 $X=4.01 $Y=0.245
+ $X2=0 $Y2=0
cc_748 N_A_602_325#_c_1111_n N_A_608_49#_c_1254_n 0.00437461f $X=6.625 $Y=1.53
+ $X2=0 $Y2=0
cc_749 N_A_602_325#_c_1112_n N_A_608_49#_c_1254_n 0.00277011f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_750 N_A_602_325#_c_1114_n N_A_608_49#_c_1254_n 0.00125154f $X=4.355 $Y=1.535
+ $X2=0 $Y2=0
cc_751 N_A_602_325#_c_1106_n N_A_608_49#_c_1255_n 0.0153275f $X=4.025 $Y=1.98
+ $X2=0 $Y2=0
cc_752 N_A_602_325#_c_1112_n N_A_608_49#_c_1255_n 0.00119193f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_753 N_A_602_325#_c_1114_n N_A_608_49#_c_1255_n 0.0114314f $X=4.355 $Y=1.535
+ $X2=0 $Y2=0
cc_754 N_A_602_325#_c_1104_n N_A_608_49#_c_1248_n 0.0327079f $X=4.355 $Y=0.76
+ $X2=0 $Y2=0
cc_755 N_A_602_325#_c_1127_n N_A_608_49#_c_1249_n 0.00649967f $X=4.11 $Y=1.895
+ $X2=0 $Y2=0
cc_756 N_A_602_325#_c_1104_n N_A_608_49#_c_1249_n 0.00889026f $X=4.355 $Y=0.76
+ $X2=0 $Y2=0
cc_757 N_A_602_325#_c_1111_n N_A_608_49#_c_1249_n 0.0221806f $X=6.625 $Y=1.53
+ $X2=0 $Y2=0
cc_758 N_A_602_325#_c_1112_n N_A_608_49#_c_1249_n 0.00275249f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_759 N_A_602_325#_c_1114_n N_A_608_49#_c_1249_n 0.0233324f $X=4.355 $Y=1.535
+ $X2=0 $Y2=0
cc_760 N_A_602_325#_c_1111_n N_A_608_49#_c_1257_n 0.0108493f $X=6.625 $Y=1.53
+ $X2=0 $Y2=0
cc_761 N_A_602_325#_c_1108_n N_A_608_49#_c_1250_n 0.0118725f $X=6.622 $Y=1.615
+ $X2=0 $Y2=0
cc_762 N_A_602_325#_c_1146_n N_A_608_49#_c_1250_n 0.0322664f $X=6.59 $Y=1.62
+ $X2=0 $Y2=0
cc_763 N_A_602_325#_c_1111_n N_A_608_49#_c_1250_n 0.0192027f $X=6.625 $Y=1.53
+ $X2=0 $Y2=0
cc_764 N_A_602_325#_c_1113_n N_A_608_49#_c_1250_n 0.00134009f $X=6.77 $Y=1.53
+ $X2=0 $Y2=0
cc_765 N_A_602_325#_M1020_d N_A_608_49#_c_1262_n 0.00904513f $X=6.25 $Y=1.485
+ $X2=0 $Y2=0
cc_766 N_A_602_325#_c_1146_n N_A_608_49#_c_1262_n 0.0235166f $X=6.59 $Y=1.62
+ $X2=0 $Y2=0
cc_767 N_A_602_325#_c_1109_n N_A_608_49#_c_1262_n 0.00873322f $X=7.025 $Y=1.53
+ $X2=0 $Y2=0
cc_768 N_A_602_325#_c_1105_n N_A_608_49#_c_1305_n 0.0028148f $X=7.11 $Y=1.445
+ $X2=0 $Y2=0
cc_769 N_A_602_325#_c_1106_n N_A_608_49#_c_1263_n 0.0049241f $X=4.025 $Y=1.98
+ $X2=0 $Y2=0
cc_770 N_A_602_325#_c_1112_n N_A_608_49#_c_1263_n 2.48159e-19 $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_771 N_A_602_325#_c_1114_n N_A_608_49#_c_1263_n 0.00535873f $X=4.355 $Y=1.535
+ $X2=0 $Y2=0
cc_772 N_A_602_325#_c_1104_n N_A_608_49#_c_1251_n 0.0133806f $X=4.355 $Y=0.76
+ $X2=0 $Y2=0
cc_773 N_A_602_325#_c_1111_n N_A_608_49#_c_1251_n 0.0053051f $X=6.625 $Y=1.53
+ $X2=0 $Y2=0
cc_774 N_A_602_325#_c_1112_n N_A_608_49#_c_1251_n 2.6396e-19 $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_775 N_A_602_325#_c_1108_n N_A_608_49#_c_1252_n 2.53366e-19 $X=6.622 $Y=1.615
+ $X2=0 $Y2=0
cc_776 N_A_602_325#_c_1111_n N_A_608_49#_c_1252_n 2.04046e-19 $X=6.625 $Y=1.53
+ $X2=0 $Y2=0
cc_777 N_A_602_325#_c_1105_n N_A_1402_49#_M1004_d 0.00729398f $X=7.11 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_778 N_A_602_325#_c_1232_p N_A_1402_49#_M1004_d 0.0024562f $X=7.195 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_779 N_A_602_325#_c_1176_n N_A_1402_49#_M1004_d 0.0107136f $X=7.705 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_780 N_A_602_325#_c_1109_n N_A_1402_49#_M1014_d 0.00414782f $X=7.025 $Y=1.53
+ $X2=0 $Y2=0
cc_781 N_A_602_325#_c_1146_n N_A_1402_49#_c_1425_n 0.00487817f $X=6.59 $Y=1.62
+ $X2=0 $Y2=0
cc_782 N_A_602_325#_c_1109_n N_A_1402_49#_c_1425_n 0.0134336f $X=7.025 $Y=1.53
+ $X2=0 $Y2=0
cc_783 N_A_602_325#_c_1105_n N_A_1402_49#_c_1425_n 0.0622566f $X=7.11 $Y=1.445
+ $X2=0 $Y2=0
cc_784 N_A_602_325#_c_1176_n N_A_1402_49#_c_1425_n 0.0106102f $X=7.705 $Y=0.36
+ $X2=0 $Y2=0
cc_785 N_A_602_325#_c_1113_n N_A_1402_49#_c_1425_n 0.0013871f $X=6.77 $Y=1.53
+ $X2=0 $Y2=0
cc_786 N_A_602_325#_c_1111_n N_VGND_c_1491_n 0.00565637f $X=6.625 $Y=1.53 $X2=0
+ $Y2=0
cc_787 N_A_602_325#_c_1232_p N_VGND_c_1497_n 0.0104913f $X=7.195 $Y=0.34 $X2=0
+ $Y2=0
cc_788 N_A_602_325#_c_1176_n N_VGND_c_1497_n 0.0586043f $X=7.705 $Y=0.36 $X2=0
+ $Y2=0
cc_789 N_A_602_325#_M1008_d N_VGND_c_1501_n 0.00184103f $X=7.805 $Y=0.245 $X2=0
+ $Y2=0
cc_790 N_A_602_325#_c_1232_p N_VGND_c_1501_n 0.00184693f $X=7.195 $Y=0.34 $X2=0
+ $Y2=0
cc_791 N_A_602_325#_c_1176_n N_VGND_c_1501_n 0.0092581f $X=7.705 $Y=0.36 $X2=0
+ $Y2=0
cc_792 N_A_608_49#_c_1262_n N_A_1402_49#_M1014_d 0.0055303f $X=8.105 $Y=2.36
+ $X2=0 $Y2=0
cc_793 N_A_608_49#_c_1262_n N_A_1402_49#_c_1437_n 0.0129278f $X=8.105 $Y=2.36
+ $X2=0 $Y2=0
cc_794 N_A_608_49#_M1011_d N_A_1402_49#_c_1438_n 0.00612338f $X=7.885 $Y=1.645
+ $X2=0 $Y2=0
cc_795 N_A_608_49#_c_1262_n N_A_1402_49#_c_1438_n 0.0467387f $X=8.105 $Y=2.36
+ $X2=0 $Y2=0
cc_796 N_A_608_49#_c_1247_n N_VGND_c_1491_n 0.0141315f $X=4.61 $Y=0.34 $X2=0
+ $Y2=0
cc_797 N_A_608_49#_c_1248_n N_VGND_c_1491_n 0.0335332f $X=4.695 $Y=1.035 $X2=0
+ $Y2=0
cc_798 N_A_608_49#_c_1246_n N_VGND_c_1495_n 0.00233735f $X=3.93 $Y=0.74 $X2=0
+ $Y2=0
cc_799 N_A_608_49#_c_1247_n N_VGND_c_1495_n 0.0445697f $X=4.61 $Y=0.34 $X2=0
+ $Y2=0
cc_800 N_A_608_49#_c_1270_n N_VGND_c_1495_n 0.0096984f $X=4.1 $Y=0.34 $X2=0
+ $Y2=0
cc_801 N_A_608_49#_c_1305_n N_VGND_c_1497_n 0.00800682f $X=6.385 $Y=0.545 $X2=0
+ $Y2=0
cc_802 N_A_608_49#_c_1252_n N_VGND_c_1497_n 0.00225825f $X=6.16 $Y=0.772 $X2=0
+ $Y2=0
cc_803 N_A_608_49#_c_1246_n N_VGND_c_1501_n 0.00612861f $X=3.93 $Y=0.74 $X2=0
+ $Y2=0
cc_804 N_A_608_49#_c_1247_n N_VGND_c_1501_n 0.0255342f $X=4.61 $Y=0.34 $X2=0
+ $Y2=0
cc_805 N_A_608_49#_c_1270_n N_VGND_c_1501_n 0.00615131f $X=4.1 $Y=0.34 $X2=0
+ $Y2=0
cc_806 N_A_608_49#_c_1305_n N_VGND_c_1501_n 0.0018012f $X=6.385 $Y=0.545 $X2=0
+ $Y2=0
cc_807 N_A_1402_49#_c_1427_n N_VGND_c_1500_n 0.0170867f $X=9.59 $Y=0.42 $X2=0
+ $Y2=0
cc_808 N_A_1402_49#_M1006_d N_VGND_c_1501_n 0.00379446f $X=9.365 $Y=0.235 $X2=0
+ $Y2=0
cc_809 N_A_1402_49#_c_1427_n N_VGND_c_1501_n 0.00982816f $X=9.59 $Y=0.42 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__nor2_8.pxi.spice
* Created: Tue Sep  1 19:17:53 2020
* 
x_PM_SKY130_FD_SC_HD__NOR2_8%A N_A_c_113_n N_A_M1004_g N_A_M1001_g N_A_c_114_n
+ N_A_M1006_g N_A_M1003_g N_A_c_115_n N_A_M1008_g N_A_M1009_g N_A_c_116_n
+ N_A_M1011_g N_A_M1010_g N_A_c_117_n N_A_M1012_g N_A_M1014_g N_A_c_118_n
+ N_A_M1013_g N_A_M1019_g N_A_c_119_n N_A_M1017_g N_A_M1020_g N_A_c_120_n
+ N_A_M1021_g N_A_M1029_g A N_A_c_121_n N_A_c_122_n PM_SKY130_FD_SC_HD__NOR2_8%A
x_PM_SKY130_FD_SC_HD__NOR2_8%B N_B_c_255_n N_B_M1007_g N_B_M1000_g N_B_c_256_n
+ N_B_M1015_g N_B_M1002_g N_B_c_257_n N_B_M1018_g N_B_M1005_g N_B_c_258_n
+ N_B_M1023_g N_B_M1016_g N_B_c_259_n N_B_M1024_g N_B_M1022_g N_B_c_260_n
+ N_B_M1025_g N_B_M1027_g N_B_c_261_n N_B_M1026_g N_B_M1030_g N_B_c_262_n
+ N_B_M1028_g N_B_M1031_g B N_B_c_275_n N_B_c_263_n PM_SKY130_FD_SC_HD__NOR2_8%B
x_PM_SKY130_FD_SC_HD__NOR2_8%A_27_297# N_A_27_297#_M1001_d N_A_27_297#_M1003_d
+ N_A_27_297#_M1010_d N_A_27_297#_M1019_d N_A_27_297#_M1029_d
+ N_A_27_297#_M1002_s N_A_27_297#_M1016_s N_A_27_297#_M1027_s
+ N_A_27_297#_M1031_s N_A_27_297#_c_398_n N_A_27_297#_c_399_n
+ N_A_27_297#_c_400_n N_A_27_297#_c_449_p N_A_27_297#_c_401_n
+ N_A_27_297#_c_450_p N_A_27_297#_c_402_n N_A_27_297#_c_451_p
+ N_A_27_297#_c_403_n N_A_27_297#_c_404_n N_A_27_297#_c_453_p
+ N_A_27_297#_c_433_n N_A_27_297#_c_489_p N_A_27_297#_c_435_n
+ N_A_27_297#_c_493_p N_A_27_297#_c_437_n N_A_27_297#_c_496_p
+ N_A_27_297#_c_439_n N_A_27_297#_c_499_p N_A_27_297#_c_405_n
+ N_A_27_297#_c_406_n N_A_27_297#_c_407_n N_A_27_297#_c_458_p
+ N_A_27_297#_c_459_p N_A_27_297#_c_460_p PM_SKY130_FD_SC_HD__NOR2_8%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR2_8%VPWR N_VPWR_M1001_s N_VPWR_M1009_s N_VPWR_M1014_s
+ N_VPWR_M1020_s N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n
+ N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_510_n
+ N_VPWR_c_511_n VPWR N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_501_n
+ N_VPWR_c_515_n PM_SKY130_FD_SC_HD__NOR2_8%VPWR
x_PM_SKY130_FD_SC_HD__NOR2_8%Y N_Y_M1004_d N_Y_M1008_d N_Y_M1012_d N_Y_M1017_d
+ N_Y_M1007_d N_Y_M1018_d N_Y_M1024_d N_Y_M1026_d N_Y_M1000_d N_Y_M1005_d
+ N_Y_M1022_d N_Y_M1030_d N_Y_c_624_n N_Y_c_601_n N_Y_c_602_n N_Y_c_635_n
+ N_Y_c_603_n N_Y_c_643_n N_Y_c_604_n N_Y_c_651_n N_Y_c_605_n N_Y_c_656_n
+ N_Y_c_744_n N_Y_c_617_n N_Y_c_618_n N_Y_c_606_n N_Y_c_686_n N_Y_c_748_n
+ N_Y_c_619_n N_Y_c_607_n N_Y_c_698_n N_Y_c_751_n N_Y_c_620_n N_Y_c_608_n
+ N_Y_c_710_n N_Y_c_754_n N_Y_c_609_n N_Y_c_610_n N_Y_c_611_n N_Y_c_612_n
+ N_Y_c_613_n N_Y_c_621_n N_Y_c_614_n N_Y_c_622_n N_Y_c_615_n Y
+ PM_SKY130_FD_SC_HD__NOR2_8%Y
x_PM_SKY130_FD_SC_HD__NOR2_8%VGND N_VGND_M1004_s N_VGND_M1006_s N_VGND_M1011_s
+ N_VGND_M1013_s N_VGND_M1021_s N_VGND_M1015_s N_VGND_M1023_s N_VGND_M1025_s
+ N_VGND_M1028_s N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n
+ N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n
+ N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n
+ N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n
+ N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n
+ VGND N_VGND_c_850_n N_VGND_c_851_n N_VGND_c_852_n
+ PM_SKY130_FD_SC_HD__NOR2_8%VGND
cc_1 VNB N_A_c_113_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_114_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_A_c_115_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_A_c_116_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB N_A_c_117_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.995
cc_6 VNB N_A_c_118_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.995
cc_7 VNB N_A_c_119_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=0.995
cc_8 VNB N_A_c_120_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.995
cc_9 VNB N_A_c_121_n 0.0124434f $X=-0.19 $Y=-0.24 $X2=3.32 $Y2=1.16
cc_10 VNB N_A_c_122_n 0.132922f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=1.16
cc_11 VNB N_B_c_255_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_12 VNB N_B_c_256_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_13 VNB N_B_c_257_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_14 VNB N_B_c_258_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_15 VNB N_B_c_259_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.995
cc_16 VNB N_B_c_260_n 0.0157999f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.995
cc_17 VNB N_B_c_261_n 0.0157944f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=0.995
cc_18 VNB N_B_c_262_n 0.019415f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.995
cc_19 VNB N_B_c_263_n 0.131229f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=1.16
cc_20 VNB N_VPWR_c_501_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_601_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=1.985
cc_22 VNB N_Y_c_602_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_603_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.985
cc_24 VNB N_Y_c_604_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=1.325
cc_25 VNB N_Y_c_605_n 0.00414888f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_26 VNB N_Y_c_606_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=3.32 $Y2=1.16
cc_27 VNB N_Y_c_607_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_608_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_609_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_610_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_611_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_612_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_613_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_614_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_615_n 0.0127619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB Y 0.019785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_826_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_827_n 0.0346469f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.56
cc_39 VNB N_VGND_c_828_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.985
cc_40 VNB N_VGND_c_829_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.56
cc_41 VNB N_VGND_c_830_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_831_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.325
cc_43 VNB N_VGND_c_832_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.995
cc_44 VNB N_VGND_c_833_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.56
cc_45 VNB N_VGND_c_834_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_835_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_836_n 0.0124313f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_48 VNB N_VGND_c_837_n 0.0181289f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_49 VNB N_VGND_c_838_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.16
cc_50 VNB N_VGND_c_839_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=1.16
cc_51 VNB N_VGND_c_840_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=3.32 $Y2=1.16
cc_52 VNB N_VGND_c_841_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=3.32 $Y2=1.16
cc_53 VNB N_VGND_c_842_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=1.16
cc_54 VNB N_VGND_c_843_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_844_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_845_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.175
cc_57 VNB N_VGND_c_846_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_847_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=3.32 $Y2=1.175
cc_59 VNB N_VGND_c_848_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_849_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_850_n 0.0166671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_851_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_852_n 0.351543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VPB N_A_M1001_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_65 VPB N_A_M1003_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_66 VPB N_A_M1009_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_67 VPB N_A_M1010_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_68 VPB N_A_M1014_g 0.0182218f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_69 VPB N_A_M1019_g 0.0182218f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=1.985
cc_70 VPB N_A_M1020_g 0.0182218f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.985
cc_71 VPB N_A_M1029_g 0.0185038f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=1.985
cc_72 VPB N_A_c_122_n 0.0229655f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=1.16
cc_73 VPB N_B_M1000_g 0.018815f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_74 VPB N_B_M1002_g 0.018138f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_75 VPB N_B_M1005_g 0.018138f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_76 VPB N_B_M1016_g 0.018138f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_77 VPB N_B_M1022_g 0.018138f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_78 VPB N_B_M1027_g 0.0181374f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=1.985
cc_79 VPB N_B_M1030_g 0.0181277f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.985
cc_80 VPB N_B_M1031_g 0.022286f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=1.985
cc_81 VPB N_B_c_263_n 0.0223627f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=1.16
cc_82 VPB N_A_27_297#_c_398_n 0.0136149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_297#_c_399_n 0.0312291f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.56
cc_84 VPB N_A_27_297#_c_400_n 0.00240424f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.325
cc_85 VPB N_A_27_297#_c_401_n 0.00240424f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.56
cc_86 VPB N_A_27_297#_c_402_n 0.00240424f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=0.56
cc_87 VPB N_A_27_297#_c_403_n 0.00240424f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=0.995
cc_88 VPB N_A_27_297#_c_404_n 0.00408164f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=0.56
cc_89 VPB N_A_27_297#_c_405_n 0.0020852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_27_297#_c_406_n 0.0020852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_27_297#_c_407_n 0.0020852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_502_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.995
cc_93 VPB N_VPWR_c_503_n 0.00393015f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_94 VPB N_VPWR_c_504_n 0.00393015f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_95 VPB N_VPWR_c_505_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_96 VPB N_VPWR_c_506_n 0.0163782f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.56
cc_97 VPB N_VPWR_c_507_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.56
cc_98 VPB N_VPWR_c_508_n 0.0163782f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_99 VPB N_VPWR_c_509_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.985
cc_100 VPB N_VPWR_c_510_n 0.0163782f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.995
cc_101 VPB N_VPWR_c_511_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.56
cc_102 VPB N_VPWR_c_512_n 0.0174963f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=1.985
cc_103 VPB N_VPWR_c_513_n 0.09497f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_104 VPB N_VPWR_c_501_n 0.0496856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_515_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_106 VPB N_Y_c_617_n 0.00234891f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.16
cc_107 VPB N_Y_c_618_n 0.0023869f $X=-0.19 $Y=1.305 $X2=3.32 $Y2=1.16
cc_108 VPB N_Y_c_619_n 0.00234891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_Y_c_620_n 0.00234891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_Y_c_621_n 0.00202537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_Y_c_622_n 0.00202537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB Y 0.0237382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 N_A_c_120_n N_B_c_255_n 0.0197043f $X=3.43 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_114 N_A_M1029_g N_B_M1000_g 0.0197043f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_c_121_n N_B_c_275_n 0.0124677f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_c_122_n N_B_c_275_n 2.30564e-19 $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_c_121_n N_B_c_263_n 0.00158796f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_c_122_n N_B_c_263_n 0.0197043f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_c_121_n N_A_27_297#_c_398_n 0.0036906f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_M1001_g N_A_27_297#_c_400_n 0.0147898f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_M1003_g N_A_27_297#_c_400_n 0.0145398f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_c_121_n N_A_27_297#_c_400_n 0.0404071f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_c_122_n N_A_27_297#_c_400_n 0.00213789f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_M1009_g N_A_27_297#_c_401_n 0.0145398f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_M1010_g N_A_27_297#_c_401_n 0.0145398f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_c_121_n N_A_27_297#_c_401_n 0.0403683f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_c_122_n N_A_27_297#_c_401_n 0.00213789f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_M1014_g N_A_27_297#_c_402_n 0.0145398f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_M1019_g N_A_27_297#_c_402_n 0.0145398f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_c_121_n N_A_27_297#_c_402_n 0.0403683f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_122_n N_A_27_297#_c_402_n 0.00213789f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_M1020_g N_A_27_297#_c_403_n 0.0144851f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_M1029_g N_A_27_297#_c_403_n 0.0144814f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_c_121_n N_A_27_297#_c_403_n 0.0404071f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_122_n N_A_27_297#_c_403_n 0.00213789f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_121_n N_A_27_297#_c_404_n 0.0012302f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_121_n N_A_27_297#_c_405_n 0.0195324f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_122_n N_A_27_297#_c_405_n 0.00221654f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_c_121_n N_A_27_297#_c_406_n 0.0195324f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_c_122_n N_A_27_297#_c_406_n 0.00221654f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_c_121_n N_A_27_297#_c_407_n 0.0195324f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_c_122_n N_A_27_297#_c_407_n 0.00221654f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_M1001_g N_VPWR_c_502_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1003_g N_VPWR_c_502_n 0.00157837f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1009_g N_VPWR_c_503_n 0.00157837f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1010_g N_VPWR_c_503_n 0.00157837f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1014_g N_VPWR_c_504_n 0.00157837f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1019_g N_VPWR_c_504_n 0.00157837f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1020_g N_VPWR_c_505_n 0.00157837f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1029_g N_VPWR_c_505_n 0.00302074f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_M1003_g N_VPWR_c_506_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1009_g N_VPWR_c_506_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_M1010_g N_VPWR_c_508_n 0.00585385f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_M1014_g N_VPWR_c_508_n 0.00585385f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1019_g N_VPWR_c_510_n 0.00585385f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1020_g N_VPWR_c_510_n 0.00585385f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_M1001_g N_VPWR_c_512_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_M1029_g N_VPWR_c_513_n 0.00585385f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_M1001_g N_VPWR_c_501_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_M1003_g N_VPWR_c_501_n 0.0104367f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_M1009_g N_VPWR_c_501_n 0.0104367f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_M1010_g N_VPWR_c_501_n 0.0104367f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_M1014_g N_VPWR_c_501_n 0.0104367f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_M1019_g N_VPWR_c_501_n 0.0104367f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_M1020_g N_VPWR_c_501_n 0.0104367f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_M1029_g N_VPWR_c_501_n 0.010464f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_c_113_n N_Y_c_624_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_114_n N_Y_c_624_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_115_n N_Y_c_624_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_c_114_n N_Y_c_601_n 0.00870364f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_c_115_n N_Y_c_601_n 0.00870364f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_121_n N_Y_c_601_n 0.036111f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_122_n N_Y_c_601_n 0.00222133f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_c_113_n N_Y_c_602_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_c_114_n N_Y_c_602_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_121_n N_Y_c_602_n 0.0265405f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_c_122_n N_Y_c_602_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_114_n N_Y_c_635_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_115_n N_Y_c_635_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_116_n N_Y_c_635_n 0.00630972f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_117_n N_Y_c_635_n 5.22228e-19 $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_c_116_n N_Y_c_603_n 0.00870364f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_117_n N_Y_c_603_n 0.00870364f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_c_121_n N_Y_c_603_n 0.036111f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_c_122_n N_Y_c_603_n 0.00222133f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_116_n N_Y_c_643_n 5.22228e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_117_n N_Y_c_643_n 0.00630972f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_118_n N_Y_c_643_n 0.00630972f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_119_n N_Y_c_643_n 5.22228e-19 $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_118_n N_Y_c_604_n 0.00870364f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_119_n N_Y_c_604_n 0.00870364f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_121_n N_Y_c_604_n 0.036111f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_c_122_n N_Y_c_604_n 0.00222133f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_c_118_n N_Y_c_651_n 5.22228e-19 $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_119_n N_Y_c_651_n 0.00630972f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_120_n N_Y_c_651_n 0.00630972f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_120_n N_Y_c_605_n 0.00865686f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_c_121_n N_Y_c_605_n 0.0101526f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_c_120_n N_Y_c_656_n 5.22228e-19 $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_115_n N_Y_c_609_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_116_n N_Y_c_609_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_121_n N_Y_c_609_n 0.0265405f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_c_122_n N_Y_c_609_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_c_117_n N_Y_c_610_n 0.00113286f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_c_118_n N_Y_c_610_n 0.00113286f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_c_121_n N_Y_c_610_n 0.0265405f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_c_122_n N_Y_c_610_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_c_119_n N_Y_c_611_n 0.00113286f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_c_120_n N_Y_c_611_n 0.00113286f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_c_121_n N_Y_c_611_n 0.0265405f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_c_122_n N_Y_c_611_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_c_113_n N_VGND_c_827_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_c_114_n N_VGND_c_828_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_115_n N_VGND_c_828_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_c_116_n N_VGND_c_829_n 0.00146448f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_c_117_n N_VGND_c_829_n 0.00146448f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_c_118_n N_VGND_c_830_n 0.00146448f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_c_119_n N_VGND_c_830_n 0.00146448f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_120_n N_VGND_c_831_n 0.00146448f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_113_n N_VGND_c_838_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_c_114_n N_VGND_c_838_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_c_115_n N_VGND_c_840_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_c_116_n N_VGND_c_840_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_c_117_n N_VGND_c_842_n 0.00423334f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_c_118_n N_VGND_c_842_n 0.00423334f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_c_119_n N_VGND_c_844_n 0.00423334f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_c_120_n N_VGND_c_844_n 0.00423334f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_c_113_n N_VGND_c_852_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_c_114_n N_VGND_c_852_n 0.0057163f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_c_115_n N_VGND_c_852_n 0.0057163f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_c_116_n N_VGND_c_852_n 0.0057163f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_c_117_n N_VGND_c_852_n 0.0057163f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_c_118_n N_VGND_c_852_n 0.0057163f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_c_119_n N_VGND_c_852_n 0.0057163f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_c_120_n N_VGND_c_852_n 0.0057435f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B_M1000_g N_A_27_297#_c_404_n 2.57315e-19 $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_237 N_B_M1000_g N_A_27_297#_c_433_n 0.0121747f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_238 N_B_M1002_g N_A_27_297#_c_433_n 0.0121306f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_239 N_B_M1005_g N_A_27_297#_c_435_n 0.0121747f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_240 N_B_M1016_g N_A_27_297#_c_435_n 0.0121747f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_241 N_B_M1022_g N_A_27_297#_c_437_n 0.0121747f $X=5.53 $Y=1.985 $X2=0 $Y2=0
cc_242 N_B_M1027_g N_A_27_297#_c_437_n 0.0121747f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_243 N_B_M1030_g N_A_27_297#_c_439_n 0.0121306f $X=6.37 $Y=1.985 $X2=0 $Y2=0
cc_244 N_B_M1031_g N_A_27_297#_c_439_n 0.0121747f $X=6.79 $Y=1.985 $X2=0 $Y2=0
cc_245 N_B_M1000_g N_VPWR_c_513_n 0.00357877f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_246 N_B_M1002_g N_VPWR_c_513_n 0.00357877f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_247 N_B_M1005_g N_VPWR_c_513_n 0.00357877f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_248 N_B_M1016_g N_VPWR_c_513_n 0.00357877f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B_M1022_g N_VPWR_c_513_n 0.00357877f $X=5.53 $Y=1.985 $X2=0 $Y2=0
cc_250 N_B_M1027_g N_VPWR_c_513_n 0.00357877f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B_M1030_g N_VPWR_c_513_n 0.00357877f $X=6.37 $Y=1.985 $X2=0 $Y2=0
cc_252 N_B_M1031_g N_VPWR_c_513_n 0.00357877f $X=6.79 $Y=1.985 $X2=0 $Y2=0
cc_253 N_B_M1000_g N_VPWR_c_501_n 0.00525237f $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_254 N_B_M1002_g N_VPWR_c_501_n 0.00522516f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B_M1005_g N_VPWR_c_501_n 0.00522516f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_256 N_B_M1016_g N_VPWR_c_501_n 0.00522516f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_257 N_B_M1022_g N_VPWR_c_501_n 0.00522516f $X=5.53 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B_M1027_g N_VPWR_c_501_n 0.00522516f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_259 N_B_M1030_g N_VPWR_c_501_n 0.00522516f $X=6.37 $Y=1.985 $X2=0 $Y2=0
cc_260 N_B_M1031_g N_VPWR_c_501_n 0.00626241f $X=6.79 $Y=1.985 $X2=0 $Y2=0
cc_261 N_B_c_255_n N_Y_c_651_n 5.22228e-19 $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_262 N_B_c_255_n N_Y_c_605_n 0.00942689f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_263 N_B_c_275_n N_Y_c_605_n 0.00651491f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B_c_255_n N_Y_c_656_n 0.00630972f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_265 N_B_c_256_n N_Y_c_656_n 0.00630972f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_266 N_B_c_257_n N_Y_c_656_n 5.22228e-19 $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B_M1002_g N_Y_c_617_n 0.0133089f $X=4.27 $Y=1.985 $X2=0 $Y2=0
cc_268 N_B_M1005_g N_Y_c_617_n 0.0133439f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B_c_275_n N_Y_c_617_n 0.0415099f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B_c_263_n N_Y_c_617_n 0.00214031f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B_M1000_g N_Y_c_618_n 5.90444e-19 $X=3.85 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B_c_275_n N_Y_c_618_n 0.0203891f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B_c_263_n N_Y_c_618_n 0.00222344f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B_c_256_n N_Y_c_606_n 0.00870364f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_275 N_B_c_257_n N_Y_c_606_n 0.00870364f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B_c_275_n N_Y_c_606_n 0.036111f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_277 N_B_c_263_n N_Y_c_606_n 0.00222133f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_278 N_B_c_256_n N_Y_c_686_n 5.22228e-19 $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B_c_257_n N_Y_c_686_n 0.00630972f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B_c_258_n N_Y_c_686_n 0.00630972f $X=5.11 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B_c_259_n N_Y_c_686_n 5.22228e-19 $X=5.53 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B_M1016_g N_Y_c_619_n 0.0133881f $X=5.11 $Y=1.985 $X2=0 $Y2=0
cc_283 N_B_M1022_g N_Y_c_619_n 0.0133881f $X=5.53 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B_c_275_n N_Y_c_619_n 0.0415099f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B_c_263_n N_Y_c_619_n 0.00214031f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B_c_258_n N_Y_c_607_n 0.00870364f $X=5.11 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B_c_259_n N_Y_c_607_n 0.00870364f $X=5.53 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B_c_275_n N_Y_c_607_n 0.036111f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_289 N_B_c_263_n N_Y_c_607_n 0.00222133f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_290 N_B_c_258_n N_Y_c_698_n 5.22228e-19 $X=5.11 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B_c_259_n N_Y_c_698_n 0.00630972f $X=5.53 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B_c_260_n N_Y_c_698_n 0.00630972f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B_c_261_n N_Y_c_698_n 5.22228e-19 $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B_M1027_g N_Y_c_620_n 0.0133881f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_295 N_B_M1030_g N_Y_c_620_n 0.0133881f $X=6.37 $Y=1.985 $X2=0 $Y2=0
cc_296 N_B_c_275_n N_Y_c_620_n 0.0415099f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_297 N_B_c_263_n N_Y_c_620_n 0.00214031f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_298 N_B_c_260_n N_Y_c_608_n 0.00870364f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B_c_261_n N_Y_c_608_n 0.00870364f $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B_c_275_n N_Y_c_608_n 0.036111f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_301 N_B_c_263_n N_Y_c_608_n 0.00222133f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_302 N_B_c_260_n N_Y_c_710_n 5.22228e-19 $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B_c_261_n N_Y_c_710_n 0.00630972f $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B_c_262_n N_Y_c_710_n 0.0109314f $X=6.79 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B_c_255_n N_Y_c_612_n 0.00113286f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B_c_256_n N_Y_c_612_n 0.00113286f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B_c_275_n N_Y_c_612_n 0.0265405f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_308 N_B_c_263_n N_Y_c_612_n 0.00230339f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_309 N_B_c_257_n N_Y_c_613_n 0.00113286f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B_c_258_n N_Y_c_613_n 0.00113286f $X=5.11 $Y=0.995 $X2=0 $Y2=0
cc_311 N_B_c_275_n N_Y_c_613_n 0.0265405f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_312 N_B_c_263_n N_Y_c_613_n 0.00230339f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_313 N_B_c_275_n N_Y_c_621_n 0.0203891f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_314 N_B_c_263_n N_Y_c_621_n 0.00222344f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_315 N_B_c_259_n N_Y_c_614_n 0.00113286f $X=5.53 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B_c_260_n N_Y_c_614_n 0.00113286f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B_c_275_n N_Y_c_614_n 0.0265405f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_318 N_B_c_263_n N_Y_c_614_n 0.00230339f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_319 N_B_c_275_n N_Y_c_622_n 0.0203891f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_320 N_B_c_263_n N_Y_c_622_n 0.00222344f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_321 N_B_c_261_n N_Y_c_615_n 0.00113286f $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B_c_262_n N_Y_c_615_n 0.00967536f $X=6.79 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B_c_275_n N_Y_c_615_n 0.0100214f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_324 N_B_c_263_n N_Y_c_615_n 0.00281533f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_325 N_B_c_261_n Y 9.30556e-19 $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B_M1030_g Y 0.00163049f $X=6.37 $Y=1.985 $X2=0 $Y2=0
cc_327 N_B_c_262_n Y 0.0038166f $X=6.79 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B_M1031_g Y 0.019219f $X=6.79 $Y=1.985 $X2=0 $Y2=0
cc_329 N_B_c_275_n Y 0.0233779f $X=6.355 $Y=1.16 $X2=0 $Y2=0
cc_330 N_B_c_263_n Y 0.0241786f $X=6.79 $Y=1.16 $X2=0 $Y2=0
cc_331 N_B_c_255_n N_VGND_c_831_n 0.00146448f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B_c_256_n N_VGND_c_832_n 0.00146448f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_333 N_B_c_257_n N_VGND_c_832_n 0.00146448f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_334 N_B_c_257_n N_VGND_c_833_n 0.00423334f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B_c_258_n N_VGND_c_833_n 0.00423334f $X=5.11 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B_c_258_n N_VGND_c_834_n 0.00146448f $X=5.11 $Y=0.995 $X2=0 $Y2=0
cc_337 N_B_c_259_n N_VGND_c_834_n 0.00146448f $X=5.53 $Y=0.995 $X2=0 $Y2=0
cc_338 N_B_c_260_n N_VGND_c_835_n 0.00146448f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_339 N_B_c_261_n N_VGND_c_835_n 0.00146448f $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_340 N_B_c_262_n N_VGND_c_837_n 0.0032322f $X=6.79 $Y=0.995 $X2=0 $Y2=0
cc_341 N_B_c_255_n N_VGND_c_846_n 0.00423334f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_342 N_B_c_256_n N_VGND_c_846_n 0.00423334f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_343 N_B_c_259_n N_VGND_c_848_n 0.00423334f $X=5.53 $Y=0.995 $X2=0 $Y2=0
cc_344 N_B_c_260_n N_VGND_c_848_n 0.00423334f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_345 N_B_c_261_n N_VGND_c_850_n 0.00423334f $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_346 N_B_c_262_n N_VGND_c_850_n 0.00423225f $X=6.79 $Y=0.995 $X2=0 $Y2=0
cc_347 N_B_c_255_n N_VGND_c_852_n 0.0057435f $X=3.85 $Y=0.995 $X2=0 $Y2=0
cc_348 N_B_c_256_n N_VGND_c_852_n 0.0057163f $X=4.27 $Y=0.995 $X2=0 $Y2=0
cc_349 N_B_c_257_n N_VGND_c_852_n 0.0057163f $X=4.69 $Y=0.995 $X2=0 $Y2=0
cc_350 N_B_c_258_n N_VGND_c_852_n 0.0057163f $X=5.11 $Y=0.995 $X2=0 $Y2=0
cc_351 N_B_c_259_n N_VGND_c_852_n 0.0057163f $X=5.53 $Y=0.995 $X2=0 $Y2=0
cc_352 N_B_c_260_n N_VGND_c_852_n 0.0057163f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_353 N_B_c_261_n N_VGND_c_852_n 0.0057163f $X=6.37 $Y=0.995 $X2=0 $Y2=0
cc_354 N_B_c_262_n N_VGND_c_852_n 0.00675157f $X=6.79 $Y=0.995 $X2=0 $Y2=0
cc_355 N_A_27_297#_c_400_n N_VPWR_M1001_s 0.00166915f $X=0.995 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_356 N_A_27_297#_c_401_n N_VPWR_M1009_s 0.00166915f $X=1.835 $Y=1.56 $X2=0
+ $Y2=0
cc_357 N_A_27_297#_c_402_n N_VPWR_M1014_s 0.00166915f $X=2.675 $Y=1.56 $X2=0
+ $Y2=0
cc_358 N_A_27_297#_c_403_n N_VPWR_M1020_s 0.00166915f $X=3.515 $Y=1.56 $X2=0
+ $Y2=0
cc_359 N_A_27_297#_c_400_n N_VPWR_c_502_n 0.0128751f $X=0.995 $Y=1.56 $X2=0
+ $Y2=0
cc_360 N_A_27_297#_c_401_n N_VPWR_c_503_n 0.0128751f $X=1.835 $Y=1.56 $X2=0
+ $Y2=0
cc_361 N_A_27_297#_c_402_n N_VPWR_c_504_n 0.0128751f $X=2.675 $Y=1.56 $X2=0
+ $Y2=0
cc_362 N_A_27_297#_c_403_n N_VPWR_c_505_n 0.0128751f $X=3.515 $Y=1.56 $X2=0
+ $Y2=0
cc_363 N_A_27_297#_c_449_p N_VPWR_c_506_n 0.0142343f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_364 N_A_27_297#_c_450_p N_VPWR_c_508_n 0.0142343f $X=1.96 $Y=2.3 $X2=0 $Y2=0
cc_365 N_A_27_297#_c_451_p N_VPWR_c_510_n 0.0142343f $X=2.8 $Y=2.3 $X2=0 $Y2=0
cc_366 N_A_27_297#_c_399_n N_VPWR_c_512_n 0.0204682f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_367 N_A_27_297#_c_453_p N_VPWR_c_513_n 0.0143053f $X=3.64 $Y=2.295 $X2=0
+ $Y2=0
cc_368 N_A_27_297#_c_433_n N_VPWR_c_513_n 0.0330174f $X=4.355 $Y=2.38 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_435_n N_VPWR_c_513_n 0.0330174f $X=5.195 $Y=2.38 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_437_n N_VPWR_c_513_n 0.0330174f $X=6.035 $Y=2.38 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_439_n N_VPWR_c_513_n 0.0489601f $X=6.875 $Y=2.38 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_458_p N_VPWR_c_513_n 0.0143053f $X=4.48 $Y=2.38 $X2=0 $Y2=0
cc_373 N_A_27_297#_c_459_p N_VPWR_c_513_n 0.0143053f $X=5.32 $Y=2.38 $X2=0 $Y2=0
cc_374 N_A_27_297#_c_460_p N_VPWR_c_513_n 0.0143053f $X=6.16 $Y=2.38 $X2=0 $Y2=0
cc_375 N_A_27_297#_M1001_d N_VPWR_c_501_n 0.00260431f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_M1003_d N_VPWR_c_501_n 0.00284632f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_M1010_d N_VPWR_c_501_n 0.00284632f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_M1019_d N_VPWR_c_501_n 0.00284632f $X=2.665 $Y=1.485 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_M1029_d N_VPWR_c_501_n 0.00246446f $X=3.505 $Y=1.485 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_M1002_s N_VPWR_c_501_n 0.00215203f $X=4.345 $Y=1.485 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_M1016_s N_VPWR_c_501_n 0.00215203f $X=5.185 $Y=1.485 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_M1027_s N_VPWR_c_501_n 0.00215203f $X=6.025 $Y=1.485 $X2=0
+ $Y2=0
cc_383 N_A_27_297#_M1031_s N_VPWR_c_501_n 0.00252233f $X=6.865 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_c_399_n N_VPWR_c_501_n 0.0120542f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_385 N_A_27_297#_c_449_p N_VPWR_c_501_n 0.00955092f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_386 N_A_27_297#_c_450_p N_VPWR_c_501_n 0.00955092f $X=1.96 $Y=2.3 $X2=0 $Y2=0
cc_387 N_A_27_297#_c_451_p N_VPWR_c_501_n 0.00955092f $X=2.8 $Y=2.3 $X2=0 $Y2=0
cc_388 N_A_27_297#_c_453_p N_VPWR_c_501_n 0.00962794f $X=3.64 $Y=2.295 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_c_433_n N_VPWR_c_501_n 0.0204627f $X=4.355 $Y=2.38 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_c_435_n N_VPWR_c_501_n 0.0204627f $X=5.195 $Y=2.38 $X2=0
+ $Y2=0
cc_391 N_A_27_297#_c_437_n N_VPWR_c_501_n 0.0204627f $X=6.035 $Y=2.38 $X2=0
+ $Y2=0
cc_392 N_A_27_297#_c_439_n N_VPWR_c_501_n 0.0300907f $X=6.875 $Y=2.38 $X2=0
+ $Y2=0
cc_393 N_A_27_297#_c_458_p N_VPWR_c_501_n 0.00962794f $X=4.48 $Y=2.38 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_459_p N_VPWR_c_501_n 0.00962794f $X=5.32 $Y=2.38 $X2=0
+ $Y2=0
cc_395 N_A_27_297#_c_460_p N_VPWR_c_501_n 0.00962794f $X=6.16 $Y=2.38 $X2=0
+ $Y2=0
cc_396 N_A_27_297#_c_433_n N_Y_M1000_d 0.00312348f $X=4.355 $Y=2.38 $X2=0 $Y2=0
cc_397 N_A_27_297#_c_435_n N_Y_M1005_d 0.00312348f $X=5.195 $Y=2.38 $X2=0 $Y2=0
cc_398 N_A_27_297#_c_437_n N_Y_M1022_d 0.00312348f $X=6.035 $Y=2.38 $X2=0 $Y2=0
cc_399 N_A_27_297#_c_439_n N_Y_M1030_d 0.00312348f $X=6.875 $Y=2.38 $X2=0 $Y2=0
cc_400 N_A_27_297#_c_404_n N_Y_c_605_n 0.0088033f $X=3.64 $Y=1.665 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_433_n N_Y_c_744_n 0.0118865f $X=4.355 $Y=2.38 $X2=0 $Y2=0
cc_402 N_A_27_297#_M1002_s N_Y_c_617_n 0.00165831f $X=4.345 $Y=1.485 $X2=0 $Y2=0
cc_403 N_A_27_297#_c_489_p N_Y_c_617_n 0.0126919f $X=4.48 $Y=1.96 $X2=0 $Y2=0
cc_404 N_A_27_297#_c_404_n N_Y_c_618_n 0.00271526f $X=3.64 $Y=1.665 $X2=0 $Y2=0
cc_405 N_A_27_297#_c_435_n N_Y_c_748_n 0.0118865f $X=5.195 $Y=2.38 $X2=0 $Y2=0
cc_406 N_A_27_297#_M1016_s N_Y_c_619_n 0.00165831f $X=5.185 $Y=1.485 $X2=0 $Y2=0
cc_407 N_A_27_297#_c_493_p N_Y_c_619_n 0.0126919f $X=5.32 $Y=1.96 $X2=0 $Y2=0
cc_408 N_A_27_297#_c_437_n N_Y_c_751_n 0.0118865f $X=6.035 $Y=2.38 $X2=0 $Y2=0
cc_409 N_A_27_297#_M1027_s N_Y_c_620_n 0.00165831f $X=6.025 $Y=1.485 $X2=0 $Y2=0
cc_410 N_A_27_297#_c_496_p N_Y_c_620_n 0.0126919f $X=6.16 $Y=1.96 $X2=0 $Y2=0
cc_411 N_A_27_297#_c_439_n N_Y_c_754_n 0.0118865f $X=6.875 $Y=2.38 $X2=0 $Y2=0
cc_412 N_A_27_297#_M1031_s Y 0.0033792f $X=6.865 $Y=1.485 $X2=0 $Y2=0
cc_413 N_A_27_297#_c_499_p Y 0.0182127f $X=7 $Y=1.96 $X2=0 $Y2=0
cc_414 N_A_27_297#_c_398_n N_VGND_c_827_n 0.0111859f $X=0.247 $Y=1.665 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_501_n N_Y_M1000_d 0.00216833f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_501_n N_Y_M1005_d 0.00216833f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_501_n N_Y_M1022_d 0.00216833f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_c_501_n N_Y_M1030_d 0.00216833f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_419 N_Y_c_601_n N_VGND_M1006_s 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_420 N_Y_c_603_n N_VGND_M1011_s 0.00162089f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_421 N_Y_c_604_n N_VGND_M1013_s 0.00162089f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_422 N_Y_c_605_n N_VGND_M1021_s 0.00162089f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_423 N_Y_c_606_n N_VGND_M1015_s 0.00162089f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_424 N_Y_c_607_n N_VGND_M1023_s 0.00162089f $X=5.575 $Y=0.815 $X2=0 $Y2=0
cc_425 N_Y_c_608_n N_VGND_M1025_s 0.00162089f $X=6.415 $Y=0.815 $X2=0 $Y2=0
cc_426 N_Y_c_615_n N_VGND_M1028_s 0.00290026f $X=6.845 $Y=0.815 $X2=0 $Y2=0
cc_427 N_Y_c_602_n N_VGND_c_827_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_428 N_Y_c_601_n N_VGND_c_828_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_429 N_Y_c_603_n N_VGND_c_829_n 0.0122559f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_430 N_Y_c_604_n N_VGND_c_830_n 0.0122559f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_431 N_Y_c_605_n N_VGND_c_831_n 0.0122559f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_432 N_Y_c_606_n N_VGND_c_832_n 0.0122559f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_433 N_Y_c_606_n N_VGND_c_833_n 0.00198695f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_434 N_Y_c_686_n N_VGND_c_833_n 0.0188551f $X=4.9 $Y=0.39 $X2=0 $Y2=0
cc_435 N_Y_c_607_n N_VGND_c_833_n 0.00198695f $X=5.575 $Y=0.815 $X2=0 $Y2=0
cc_436 N_Y_c_607_n N_VGND_c_834_n 0.0122559f $X=5.575 $Y=0.815 $X2=0 $Y2=0
cc_437 N_Y_c_608_n N_VGND_c_835_n 0.0122559f $X=6.415 $Y=0.815 $X2=0 $Y2=0
cc_438 N_Y_c_615_n N_VGND_c_836_n 0.0011947f $X=6.845 $Y=0.815 $X2=0 $Y2=0
cc_439 N_Y_c_615_n N_VGND_c_837_n 0.0246547f $X=6.845 $Y=0.815 $X2=0 $Y2=0
cc_440 N_Y_c_624_n N_VGND_c_838_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_441 N_Y_c_601_n N_VGND_c_838_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_442 N_Y_c_601_n N_VGND_c_840_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_443 N_Y_c_635_n N_VGND_c_840_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_444 N_Y_c_603_n N_VGND_c_840_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_445 N_Y_c_603_n N_VGND_c_842_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_446 N_Y_c_643_n N_VGND_c_842_n 0.0188551f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_447 N_Y_c_604_n N_VGND_c_842_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_448 N_Y_c_604_n N_VGND_c_844_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_449 N_Y_c_651_n N_VGND_c_844_n 0.0188551f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_450 N_Y_c_605_n N_VGND_c_844_n 0.00198695f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_451 N_Y_c_605_n N_VGND_c_846_n 0.00198695f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_452 N_Y_c_656_n N_VGND_c_846_n 0.0188551f $X=4.06 $Y=0.39 $X2=0 $Y2=0
cc_453 N_Y_c_606_n N_VGND_c_846_n 0.00198695f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_454 N_Y_c_607_n N_VGND_c_848_n 0.00198695f $X=5.575 $Y=0.815 $X2=0 $Y2=0
cc_455 N_Y_c_698_n N_VGND_c_848_n 0.0188551f $X=5.74 $Y=0.39 $X2=0 $Y2=0
cc_456 N_Y_c_608_n N_VGND_c_848_n 0.00198695f $X=6.415 $Y=0.815 $X2=0 $Y2=0
cc_457 N_Y_c_608_n N_VGND_c_850_n 0.00198695f $X=6.415 $Y=0.815 $X2=0 $Y2=0
cc_458 N_Y_c_710_n N_VGND_c_850_n 0.0188614f $X=6.58 $Y=0.39 $X2=0 $Y2=0
cc_459 N_Y_c_615_n N_VGND_c_850_n 0.00215161f $X=6.845 $Y=0.815 $X2=0 $Y2=0
cc_460 N_Y_M1004_d N_VGND_c_852_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_461 N_Y_M1008_d N_VGND_c_852_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_462 N_Y_M1012_d N_VGND_c_852_n 0.00215201f $X=2.245 $Y=0.235 $X2=0 $Y2=0
cc_463 N_Y_M1017_d N_VGND_c_852_n 0.00215201f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_464 N_Y_M1007_d N_VGND_c_852_n 0.00215201f $X=3.925 $Y=0.235 $X2=0 $Y2=0
cc_465 N_Y_M1018_d N_VGND_c_852_n 0.00215201f $X=4.765 $Y=0.235 $X2=0 $Y2=0
cc_466 N_Y_M1024_d N_VGND_c_852_n 0.00215201f $X=5.605 $Y=0.235 $X2=0 $Y2=0
cc_467 N_Y_M1026_d N_VGND_c_852_n 0.00215201f $X=6.445 $Y=0.235 $X2=0 $Y2=0
cc_468 N_Y_c_624_n N_VGND_c_852_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_469 N_Y_c_601_n N_VGND_c_852_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_470 N_Y_c_635_n N_VGND_c_852_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_471 N_Y_c_603_n N_VGND_c_852_n 0.00835832f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_472 N_Y_c_643_n N_VGND_c_852_n 0.0122069f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_473 N_Y_c_604_n N_VGND_c_852_n 0.00835832f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_474 N_Y_c_651_n N_VGND_c_852_n 0.0122069f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_475 N_Y_c_605_n N_VGND_c_852_n 0.00835832f $X=3.895 $Y=0.815 $X2=0 $Y2=0
cc_476 N_Y_c_656_n N_VGND_c_852_n 0.0122069f $X=4.06 $Y=0.39 $X2=0 $Y2=0
cc_477 N_Y_c_606_n N_VGND_c_852_n 0.00835832f $X=4.735 $Y=0.815 $X2=0 $Y2=0
cc_478 N_Y_c_686_n N_VGND_c_852_n 0.0122069f $X=4.9 $Y=0.39 $X2=0 $Y2=0
cc_479 N_Y_c_607_n N_VGND_c_852_n 0.00835832f $X=5.575 $Y=0.815 $X2=0 $Y2=0
cc_480 N_Y_c_698_n N_VGND_c_852_n 0.0122069f $X=5.74 $Y=0.39 $X2=0 $Y2=0
cc_481 N_Y_c_608_n N_VGND_c_852_n 0.00835832f $X=6.415 $Y=0.815 $X2=0 $Y2=0
cc_482 N_Y_c_710_n N_VGND_c_852_n 0.0122084f $X=6.58 $Y=0.39 $X2=0 $Y2=0
cc_483 N_Y_c_615_n N_VGND_c_852_n 0.00739045f $X=6.845 $Y=0.815 $X2=0 $Y2=0

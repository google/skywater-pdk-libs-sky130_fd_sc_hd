# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nand4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 0.995000 2.215000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.300000 1.350000 0.825000 ;
        RECT 1.145000 0.825000 1.350000 0.995000 ;
        RECT 1.145000 0.995000 1.455000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.300000 0.810000 0.995000 ;
        RECT 0.595000 0.995000 0.975000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.995000 0.395000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.795000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 1.795000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.385000 1.665000 1.715000 2.465000 ;
        RECT 1.520000 0.255000 2.215000 0.825000 ;
        RECT 1.625000 0.825000 1.795000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.300000 0.085000 ;
        RECT 0.090000  0.085000 0.425000 0.825000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.300000 2.805000 ;
        RECT 0.085000 1.495000 0.345000 2.635000 ;
        RECT 1.015000 1.835000 1.185000 2.635000 ;
        RECT 1.915000 1.835000 2.195000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__nand4_1
END LIBRARY

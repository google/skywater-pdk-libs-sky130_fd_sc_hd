* File: sky130_fd_sc_hd__sdfstp_4.pxi.spice
* Created: Tue Sep  1 19:30:56 2020
* 
x_PM_SKY130_FD_SC_HD__SDFSTP_4%SCD N_SCD_c_283_n N_SCD_c_287_n N_SCD_c_284_n
+ N_SCD_M1041_g N_SCD_c_288_n N_SCD_M1018_g N_SCD_c_289_n SCD SCD
+ PM_SKY130_FD_SC_HD__SDFSTP_4%SCD
x_PM_SKY130_FD_SC_HD__SDFSTP_4%SCE N_SCE_M1012_g N_SCE_c_317_n N_SCE_M1002_g
+ N_SCE_M1026_g N_SCE_M1013_g SCE N_SCE_c_320_n N_SCE_c_340_n N_SCE_c_356_p
+ N_SCE_c_321_n N_SCE_c_322_n PM_SKY130_FD_SC_HD__SDFSTP_4%SCE
x_PM_SKY130_FD_SC_HD__SDFSTP_4%D N_D_c_424_n N_D_M1019_g N_D_M1004_g D D
+ N_D_c_427_n PM_SKY130_FD_SC_HD__SDFSTP_4%D
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_319_21# N_A_319_21#_M1013_s N_A_319_21#_M1026_s
+ N_A_319_21#_M1031_g N_A_319_21#_M1001_g N_A_319_21#_c_466_n
+ N_A_319_21#_c_467_n N_A_319_21#_c_468_n N_A_319_21#_c_469_n
+ N_A_319_21#_c_470_n N_A_319_21#_c_475_n N_A_319_21#_c_476_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_319_21#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%CLK N_CLK_M1036_g N_CLK_c_541_n N_CLK_M1000_g
+ N_CLK_c_542_n N_CLK_c_547_n N_CLK_c_548_n CLK CLK CLK CLK N_CLK_c_545_n
+ N_CLK_c_546_n PM_SKY130_FD_SC_HD__SDFSTP_4%CLK
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_643_369# N_A_643_369#_M1000_s
+ N_A_643_369#_M1036_s N_A_643_369#_M1029_g N_A_643_369#_c_614_n
+ N_A_643_369#_M1039_g N_A_643_369#_c_615_n N_A_643_369#_c_616_n
+ N_A_643_369#_M1020_g N_A_643_369#_M1038_g N_A_643_369#_M1017_g
+ N_A_643_369#_M1033_g N_A_643_369#_c_618_n N_A_643_369#_c_646_n
+ N_A_643_369#_c_619_n N_A_643_369#_c_634_n N_A_643_369#_c_635_n
+ N_A_643_369#_c_620_n N_A_643_369#_c_621_n N_A_643_369#_c_706_p
+ N_A_643_369#_c_622_n N_A_643_369#_c_623_n N_A_643_369#_c_624_n
+ N_A_643_369#_c_625_n N_A_643_369#_c_626_n N_A_643_369#_c_627_n
+ N_A_643_369#_c_628_n N_A_643_369#_c_629_n N_A_643_369#_c_696_p
+ N_A_643_369#_c_640_n N_A_643_369#_c_641_n N_A_643_369#_c_642_n
+ N_A_643_369#_c_643_n N_A_643_369#_c_752_p N_A_643_369#_c_630_n
+ N_A_643_369#_c_644_n N_A_643_369#_c_645_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_643_369#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_809_369# N_A_809_369#_M1039_d
+ N_A_809_369#_M1029_d N_A_809_369#_c_909_n N_A_809_369#_c_899_n
+ N_A_809_369#_c_910_n N_A_809_369#_M1007_g N_A_809_369#_M1021_g
+ N_A_809_369#_M1044_g N_A_809_369#_c_912_n N_A_809_369#_M1034_g
+ N_A_809_369#_c_914_n N_A_809_369#_c_915_n N_A_809_369#_c_916_n
+ N_A_809_369#_c_1036_p N_A_809_369#_c_902_n N_A_809_369#_c_903_n
+ N_A_809_369#_c_904_n N_A_809_369#_c_905_n N_A_809_369#_c_906_n
+ N_A_809_369#_c_907_n N_A_809_369#_c_908_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_809_369#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_1129_21# N_A_1129_21#_M1008_s
+ N_A_1129_21#_M1005_d N_A_1129_21#_M1023_g N_A_1129_21#_M1040_g
+ N_A_1129_21#_c_1085_n N_A_1129_21#_c_1086_n N_A_1129_21#_c_1079_n
+ N_A_1129_21#_c_1087_n N_A_1129_21#_c_1088_n N_A_1129_21#_c_1080_n
+ N_A_1129_21#_c_1154_p N_A_1129_21#_c_1081_n N_A_1129_21#_c_1082_n
+ N_A_1129_21#_c_1083_n PM_SKY130_FD_SC_HD__SDFSTP_4%A_1129_21#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_997_413# N_A_997_413#_M1020_d
+ N_A_997_413#_M1007_d N_A_997_413#_M1005_g N_A_997_413#_c_1174_n
+ N_A_997_413#_M1008_g N_A_997_413#_M1014_g N_A_997_413#_M1011_g
+ N_A_997_413#_c_1175_n N_A_997_413#_c_1176_n N_A_997_413#_c_1201_n
+ N_A_997_413#_c_1187_n N_A_997_413#_c_1177_n N_A_997_413#_c_1178_n
+ N_A_997_413#_c_1179_n N_A_997_413#_c_1180_n N_A_997_413#_c_1181_n
+ N_A_997_413#_c_1182_n N_A_997_413#_c_1183_n N_A_997_413#_c_1184_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_997_413#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%SET_B N_SET_B_M1030_g N_SET_B_M1043_g
+ N_SET_B_M1025_g N_SET_B_M1042_g N_SET_B_c_1321_n N_SET_B_c_1325_n
+ N_SET_B_c_1326_n N_SET_B_c_1327_n N_SET_B_c_1328_n SET_B N_SET_B_c_1329_n
+ N_SET_B_c_1330_n N_SET_B_c_1331_n N_SET_B_c_1332_n N_SET_B_c_1333_n
+ N_SET_B_c_1334_n N_SET_B_c_1335_n PM_SKY130_FD_SC_HD__SDFSTP_4%SET_B
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_1781_295# N_A_1781_295#_M1010_d
+ N_A_1781_295#_M1015_d N_A_1781_295#_M1006_g N_A_1781_295#_c_1464_n
+ N_A_1781_295#_c_1465_n N_A_1781_295#_M1035_g N_A_1781_295#_c_1456_n
+ N_A_1781_295#_c_1457_n N_A_1781_295#_c_1458_n N_A_1781_295#_c_1459_n
+ N_A_1781_295#_c_1468_n N_A_1781_295#_c_1469_n N_A_1781_295#_c_1460_n
+ N_A_1781_295#_c_1461_n N_A_1781_295#_c_1462_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_1781_295#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_1597_329# N_A_1597_329#_M1044_d
+ N_A_1597_329#_M1017_d N_A_1597_329#_M1025_d N_A_1597_329#_M1010_g
+ N_A_1597_329#_M1015_g N_A_1597_329#_c_1562_n N_A_1597_329#_M1009_g
+ N_A_1597_329#_M1016_g N_A_1597_329#_c_1564_n N_A_1597_329#_c_1565_n
+ N_A_1597_329#_c_1566_n N_A_1597_329#_c_1567_n N_A_1597_329#_c_1588_n
+ N_A_1597_329#_c_1589_n N_A_1597_329#_c_1577_n N_A_1597_329#_c_1578_n
+ N_A_1597_329#_c_1568_n N_A_1597_329#_c_1569_n N_A_1597_329#_c_1570_n
+ N_A_1597_329#_c_1571_n N_A_1597_329#_c_1579_n N_A_1597_329#_c_1580_n
+ N_A_1597_329#_c_1581_n N_A_1597_329#_c_1582_n N_A_1597_329#_c_1583_n
+ N_A_1597_329#_c_1584_n PM_SKY130_FD_SC_HD__SDFSTP_4%A_1597_329#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_2227_47# N_A_2227_47#_M1009_s
+ N_A_2227_47#_M1016_s N_A_2227_47#_c_1717_n N_A_2227_47#_M1022_g
+ N_A_2227_47#_M1003_g N_A_2227_47#_c_1718_n N_A_2227_47#_M1027_g
+ N_A_2227_47#_M1024_g N_A_2227_47#_c_1719_n N_A_2227_47#_M1032_g
+ N_A_2227_47#_M1028_g N_A_2227_47#_c_1720_n N_A_2227_47#_M1037_g
+ N_A_2227_47#_M1045_g N_A_2227_47#_c_1721_n N_A_2227_47#_c_1729_n
+ N_A_2227_47#_c_1722_n N_A_2227_47#_c_1723_n N_A_2227_47#_c_1724_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_2227_47#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_27_369# N_A_27_369#_M1018_s N_A_27_369#_M1001_d
+ N_A_27_369#_c_1810_n N_A_27_369#_c_1811_n N_A_27_369#_c_1812_n
+ N_A_27_369#_c_1818_n N_A_27_369#_c_1825_n N_A_27_369#_c_1813_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_27_369#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%VPWR N_VPWR_M1018_d N_VPWR_M1026_d N_VPWR_M1036_d
+ N_VPWR_M1040_d N_VPWR_M1030_d N_VPWR_M1006_d N_VPWR_M1015_s N_VPWR_M1016_d
+ N_VPWR_M1024_s N_VPWR_M1045_s N_VPWR_c_1852_n N_VPWR_c_1853_n N_VPWR_c_1854_n
+ N_VPWR_c_1855_n N_VPWR_c_1856_n N_VPWR_c_1857_n N_VPWR_c_1858_n
+ N_VPWR_c_1859_n N_VPWR_c_1860_n N_VPWR_c_1861_n N_VPWR_c_1862_n
+ N_VPWR_c_1863_n N_VPWR_c_1864_n N_VPWR_c_1865_n N_VPWR_c_1866_n VPWR
+ N_VPWR_c_1867_n N_VPWR_c_1868_n N_VPWR_c_1869_n N_VPWR_c_1870_n
+ N_VPWR_c_1871_n N_VPWR_c_1872_n N_VPWR_c_1873_n N_VPWR_c_1874_n
+ N_VPWR_c_1875_n N_VPWR_c_1876_n N_VPWR_c_1877_n N_VPWR_c_1878_n
+ N_VPWR_c_1879_n N_VPWR_c_1851_n PM_SKY130_FD_SC_HD__SDFSTP_4%VPWR
x_PM_SKY130_FD_SC_HD__SDFSTP_4%A_181_47# N_A_181_47#_M1012_d N_A_181_47#_M1020_s
+ N_A_181_47#_M1004_d N_A_181_47#_M1007_s N_A_181_47#_c_2073_n
+ N_A_181_47#_c_2061_n N_A_181_47#_c_2066_n N_A_181_47#_c_2067_n
+ N_A_181_47#_c_2062_n N_A_181_47#_c_2077_n N_A_181_47#_c_2063_n
+ N_A_181_47#_c_2064_n N_A_181_47#_c_2069_n N_A_181_47#_c_2070_n
+ N_A_181_47#_c_2065_n N_A_181_47#_c_2072_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%A_181_47#
x_PM_SKY130_FD_SC_HD__SDFSTP_4%Q N_Q_M1022_d N_Q_M1032_d N_Q_M1003_d N_Q_M1028_d
+ N_Q_c_2209_n N_Q_c_2213_n N_Q_c_2216_n N_Q_c_2217_n Q Q Q Q Q Q Q N_Q_c_2226_n
+ Q Q PM_SKY130_FD_SC_HD__SDFSTP_4%Q
x_PM_SKY130_FD_SC_HD__SDFSTP_4%VGND N_VGND_M1041_s N_VGND_M1031_d N_VGND_M1013_d
+ N_VGND_M1000_d N_VGND_M1023_d N_VGND_M1043_d N_VGND_M1042_d N_VGND_M1009_d
+ N_VGND_M1027_s N_VGND_M1037_s N_VGND_c_2250_n N_VGND_c_2251_n N_VGND_c_2252_n
+ N_VGND_c_2253_n N_VGND_c_2254_n N_VGND_c_2255_n N_VGND_c_2256_n
+ N_VGND_c_2257_n N_VGND_c_2258_n N_VGND_c_2259_n N_VGND_c_2260_n
+ N_VGND_c_2261_n VGND N_VGND_c_2262_n N_VGND_c_2263_n N_VGND_c_2264_n
+ N_VGND_c_2265_n N_VGND_c_2266_n N_VGND_c_2267_n N_VGND_c_2268_n
+ N_VGND_c_2269_n N_VGND_c_2270_n N_VGND_c_2271_n N_VGND_c_2272_n
+ N_VGND_c_2273_n N_VGND_c_2274_n N_VGND_c_2275_n
+ PM_SKY130_FD_SC_HD__SDFSTP_4%VGND
cc_1 VNB N_SCD_c_283_n 0.0592907f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.325
cc_2 VNB N_SCD_c_284_n 0.017218f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB SCD 0.0208496f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_SCE_M1012_g 0.030725f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_5 VNB N_SCE_c_317_n 0.0195372f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_6 VNB N_SCE_M1013_g 0.0380569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB SCE 0.00509679f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_8 VNB N_SCE_c_320_n 0.0088747f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_9 VNB N_SCE_c_321_n 0.0281415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_322_n 0.00121095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_D_c_424_n 0.0164669f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.325
cc_12 VNB N_D_M1004_g 0.00862768f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.77
cc_13 VNB D 0.00524595f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_14 VNB N_D_c_427_n 0.0252314f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_15 VNB N_A_319_21#_M1031_g 0.0301667f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_16 VNB N_A_319_21#_c_466_n 0.00865826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_319_21#_c_467_n 0.00437998f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_18 VNB N_A_319_21#_c_468_n 0.0322821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_319_21#_c_469_n 0.0137961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_319_21#_c_470_n 0.00677902f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.53
cc_21 VNB N_CLK_c_541_n 0.0170611f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_22 VNB N_CLK_c_542_n 0.0143095f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_23 VNB CLK 0.0102993f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_24 VNB CLK 0.0136786f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_25 VNB N_CLK_c_545_n 0.0164797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_CLK_c_546_n 0.0133943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_643_369#_c_614_n 0.0171116f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_28 VNB N_A_643_369#_c_615_n 0.051233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_643_369#_c_616_n 0.0170002f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_30 VNB N_A_643_369#_M1033_g 0.0241357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_643_369#_c_618_n 0.00552567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_643_369#_c_619_n 0.00133463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_643_369#_c_620_n 0.00586703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_643_369#_c_621_n 0.00228328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_643_369#_c_622_n 0.00316033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_643_369#_c_623_n 0.0160923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_643_369#_c_624_n 0.00392757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_643_369#_c_625_n 0.025427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_643_369#_c_626_n 0.00902583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_643_369#_c_627_n 3.84112e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_643_369#_c_628_n 0.00443092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_643_369#_c_629_n 0.0279818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_643_369#_c_630_n 0.0110155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_809_369#_c_899_n 0.0426125f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_45 VNB N_A_809_369#_M1021_g 0.0306428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_809_369#_M1044_g 0.0365403f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_47 VNB N_A_809_369#_c_902_n 0.0191288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_809_369#_c_903_n 0.00270322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_809_369#_c_904_n 0.00326418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_809_369#_c_905_n 0.00370222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_809_369#_c_906_n 0.00170987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_809_369#_c_907_n 0.0170178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_809_369#_c_908_n 0.00465628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1129_21#_M1023_g 0.0193358f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_55 VNB N_A_1129_21#_c_1079_n 0.00781478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1129_21#_c_1080_n 0.00452229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1129_21#_c_1081_n 3.23878e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1129_21#_c_1082_n 0.0303054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1129_21#_c_1083_n 0.0126343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_997_413#_c_1174_n 0.0162044f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_61 VNB N_A_997_413#_c_1175_n 0.0205315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_997_413#_c_1176_n 0.00688319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_997_413#_c_1177_n 0.00521515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_997_413#_c_1178_n 0.0147428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_997_413#_c_1179_n 0.01919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_997_413#_c_1180_n 0.00204312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_997_413#_c_1181_n 0.00232092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_997_413#_c_1182_n 0.0218686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_997_413#_c_1183_n 0.0121429f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_997_413#_c_1184_n 0.0192482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_SET_B_M1043_g 0.0359063f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_72 VNB N_SET_B_M1042_g 0.0427416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_SET_B_c_1321_n 0.00599564f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_74 VNB N_A_1781_295#_M1035_g 0.0211658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1781_295#_c_1456_n 0.0063596f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_76 VNB N_A_1781_295#_c_1457_n 0.0011397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1781_295#_c_1458_n 0.0270798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1781_295#_c_1459_n 0.0096039f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.53
cc_79 VNB N_A_1781_295#_c_1460_n 0.0121311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1781_295#_c_1461_n 0.00332436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1781_295#_c_1462_n 5.01057e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1597_329#_c_1562_n 0.0314804f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_83 VNB N_A_1597_329#_M1009_g 0.0311005f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_84 VNB N_A_1597_329#_c_1564_n 0.0128863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1597_329#_c_1565_n 0.0205241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1597_329#_c_1566_n 0.00637671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1597_329#_c_1567_n 0.00260706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1597_329#_c_1568_n 0.00132961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1597_329#_c_1569_n 0.0021216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1597_329#_c_1570_n 0.0100396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1597_329#_c_1571_n 0.0218829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2227_47#_c_1717_n 0.0167001f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_93 VNB N_A_2227_47#_c_1718_n 0.0160018f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_94 VNB N_A_2227_47#_c_1719_n 0.0160039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2227_47#_c_1720_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_2227_47#_c_1721_n 0.00863404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_2227_47#_c_1722_n 0.00377373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_2227_47#_c_1723_n 0.00174595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_2227_47#_c_1724_n 0.0833909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VPWR_c_1851_n 0.573369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_181_47#_c_2061_n 0.00555327f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_102 VNB N_A_181_47#_c_2062_n 0.00327209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_A_181_47#_c_2063_n 0.00180479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_A_181_47#_c_2064_n 0.0012695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_A_181_47#_c_2065_n 0.00260667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB Q 0.00106334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_2250_n 0.00791647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_2251_n 0.00737776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2252_n 3.98222e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2253_n 0.00237268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2254_n 0.0024119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2255_n 0.00468466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2256_n 0.0113527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2257_n 0.0376107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2258_n 0.0278483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2259_n 0.00506925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2260_n 0.0182896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2261_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2262_n 0.0148988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2263_n 0.0132215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2264_n 0.054764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2265_n 0.060881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2266_n 0.0288311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2267_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2268_n 0.0338415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2269_n 0.00664466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2270_n 0.00436611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2271_n 0.0151241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2272_n 0.0177582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2273_n 0.0035381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2274_n 0.00558559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2275_n 0.641238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VPB N_SCD_c_283_n 0.00536633f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.325
cc_134 VPB N_SCD_c_287_n 0.019303f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.62
cc_135 VPB N_SCD_c_288_n 0.0190089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.77
cc_136 VPB N_SCD_c_289_n 0.0259455f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_137 VPB SCD 0.0148037f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_138 VPB N_SCE_c_317_n 0.0133475f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_139 VPB N_SCE_M1002_g 0.0317142f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_140 VPB N_SCE_M1026_g 0.0507543f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_141 VPB SCE 0.00452509f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_142 VPB N_SCE_c_321_n 0.00631733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_SCE_c_322_n 0.00418661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_D_M1004_g 0.0333803f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.77
cc_145 VPB D 0.00602885f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_146 VPB N_A_319_21#_M1001_g 0.0422977f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_147 VPB N_A_319_21#_c_466_n 5.76251e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_319_21#_c_467_n 0.00985028f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_149 VPB N_A_319_21#_c_468_n 0.0147247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_319_21#_c_475_n 0.0040706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_319_21#_c_476_n 0.0119754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_CLK_c_547_n 0.011733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_CLK_c_548_n 0.0312275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB CLK 0.00973579f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_155 VPB CLK 0.0147114f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_156 VPB N_CLK_c_545_n 0.0104614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_643_369#_M1029_g 0.0354172f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.695
cc_158 VPB N_A_643_369#_M1038_g 0.019201f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_159 VPB N_A_643_369#_M1017_g 0.0245732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_643_369#_c_634_n 0.0015302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_643_369#_c_635_n 0.00125494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_643_369#_c_622_n 0.00356071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_643_369#_c_623_n 0.0105554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_643_369#_c_624_n 0.00220675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_643_369#_c_625_n 0.00453649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_643_369#_c_640_n 0.0058776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_643_369#_c_641_n 3.73476e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_643_369#_c_642_n 0.00752647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_643_369#_c_643_n 0.00213153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_643_369#_c_644_n 0.0321882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_643_369#_c_645_n 0.00192244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_809_369#_c_909_n 0.0244169f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_173 VPB N_A_809_369#_c_910_n 0.0174418f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_174 VPB N_A_809_369#_M1044_g 0.0159123f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_175 VPB N_A_809_369#_c_912_n 0.0374421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_809_369#_M1034_g 0.0213555f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.53
cc_177 VPB N_A_809_369#_c_914_n 0.0283508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_809_369#_c_915_n 0.00487948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_809_369#_c_916_n 0.00948235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_809_369#_c_904_n 0.00121793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_809_369#_c_905_n 3.90977e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_809_369#_c_906_n 0.0030446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_809_369#_c_907_n 0.0169522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1129_21#_M1040_g 0.0216766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1129_21#_c_1085_n 0.00176545f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_186 VPB N_A_1129_21#_c_1086_n 0.0377265f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_187 VPB N_A_1129_21#_c_1087_n 0.00566683f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.53
cc_188 VPB N_A_1129_21#_c_1088_n 7.28078e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1129_21#_c_1083_n 0.0167848f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_997_413#_M1005_g 0.0487068f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_191 VPB N_A_997_413#_M1011_g 0.0264872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_997_413#_c_1187_n 0.0126708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_997_413#_c_1177_n 0.00574591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_997_413#_c_1178_n 0.00210306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_997_413#_c_1179_n 0.00940441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_997_413#_c_1180_n 0.0035338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_997_413#_c_1181_n 0.00131078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_997_413#_c_1182_n 0.00600964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_SET_B_M1030_g 0.0241724f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_200 VPB N_SET_B_M1042_g 0.00836198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_SET_B_c_1321_n 0.00547376f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_202 VPB N_SET_B_c_1325_n 0.0429653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_SET_B_c_1326_n 0.0110097f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_204 VPB N_SET_B_c_1327_n 0.00810406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_SET_B_c_1328_n 0.015762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_SET_B_c_1329_n 0.0139047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_SET_B_c_1330_n 0.00495266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_SET_B_c_1331_n 0.00566661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_SET_B_c_1332_n 0.0044368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_SET_B_c_1333_n 0.0278673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_SET_B_c_1334_n 0.00907209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_SET_B_c_1335_n 0.00833156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_1781_295#_M1006_g 0.0347737f $X=-0.19 $Y=1.305 $X2=0.315
+ $Y2=1.695
cc_214 VPB N_A_1781_295#_c_1464_n 0.0272831f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.695
cc_215 VPB N_A_1781_295#_c_1465_n 0.00635875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_1781_295#_c_1456_n 0.010639f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_217 VPB N_A_1781_295#_c_1459_n 0.00702928f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.53
cc_218 VPB N_A_1781_295#_c_1468_n 8.64549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_1781_295#_c_1469_n 0.0187552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1597_329#_M1015_g 0.0295641f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_221 VPB N_A_1597_329#_c_1562_n 0.0248059f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_222 VPB N_A_1597_329#_M1016_g 0.0207967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1597_329#_c_1566_n 0.00277454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1597_329#_c_1567_n 0.00164223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1597_329#_c_1577_n 0.00807823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1597_329#_c_1578_n 0.00461389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1597_329#_c_1579_n 0.0057934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1597_329#_c_1580_n 0.00240039f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_1597_329#_c_1581_n 5.71433e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_A_1597_329#_c_1582_n 0.00171978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_1597_329#_c_1583_n 0.0341616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_1597_329#_c_1584_n 0.0168553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_2227_47#_M1003_g 0.0193752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_2227_47#_M1024_g 0.0183907f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_235 VPB N_A_2227_47#_M1028_g 0.0183913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_2227_47#_M1045_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_A_2227_47#_c_1729_n 0.0112012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_2227_47#_c_1722_n 0.00194757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_A_2227_47#_c_1724_n 0.0160627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_27_369#_c_1810_n 0.0170416f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_241 VPB N_A_27_369#_c_1811_n 0.00117506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_A_27_369#_c_1812_n 0.00939815f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_243 VPB N_A_27_369#_c_1813_n 0.00262476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1852_n 0.00242115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1853_n 0.00888562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1854_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1855_n 0.00500806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1856_n 0.00488885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1857_n 0.0024119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1858_n 0.00359948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1859_n 0.0113268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1860_n 0.0485139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1861_n 0.0459023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1862_n 0.00564769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1863_n 0.0271668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1864_n 0.00631397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1865_n 0.0182605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1866_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1867_n 0.0143786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1868_n 0.0161129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1869_n 0.0507059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1870_n 0.016761f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1871_n 0.0257651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1872_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1873_n 0.00391805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1874_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1875_n 0.0133604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1876_n 0.0199681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1877_n 0.0192332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1878_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1879_n 0.0055597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1851_n 0.0681155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_A_181_47#_c_2066_n 0.00388703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_A_181_47#_c_2067_n 0.00300946f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_275 VPB N_A_181_47#_c_2062_n 0.00201708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_A_181_47#_c_2069_n 0.0248372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_A_181_47#_c_2070_n 0.00312327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_A_181_47#_c_2065_n 0.00329791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_A_181_47#_c_2072_n 0.00436874f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB Q 0.00153701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 N_SCD_c_283_n N_SCE_M1012_g 0.00583208f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_282 N_SCD_c_284_n N_SCE_M1012_g 0.0484084f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_283 SCD N_SCE_M1012_g 2.56735e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_284 N_SCD_c_283_n N_SCE_c_317_n 0.0200842f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_285 SCD N_SCE_c_317_n 3.421e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_286 N_SCD_c_287_n N_SCE_M1002_g 0.00453523f $X=0.315 $Y=1.62 $X2=0 $Y2=0
cc_287 N_SCD_c_289_n N_SCE_M1002_g 0.0327721f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_288 SCD N_SCE_M1002_g 2.04234e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_289 N_SCD_c_283_n SCE 0.00799654f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_290 N_SCD_c_289_n SCE 0.00146655f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_291 SCD SCE 0.0593537f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_292 SCD N_SCE_c_340_n 0.00158165f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_293 N_SCD_c_288_n N_A_27_369#_c_1811_n 0.014189f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_294 N_SCD_c_283_n N_A_27_369#_c_1812_n 5.05332e-19 $X=0.315 $Y=1.325 $X2=0
+ $Y2=0
cc_295 N_SCD_c_289_n N_A_27_369#_c_1812_n 0.00316572f $X=0.47 $Y=1.695 $X2=0
+ $Y2=0
cc_296 SCD N_A_27_369#_c_1812_n 0.0226954f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_297 N_SCD_c_288_n N_A_27_369#_c_1818_n 4.39242e-19 $X=0.47 $Y=1.77 $X2=0
+ $Y2=0
cc_298 N_SCD_c_288_n N_VPWR_c_1852_n 0.00863247f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_299 N_SCD_c_288_n N_VPWR_c_1867_n 0.00346207f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_300 N_SCD_c_288_n N_VPWR_c_1851_n 0.00509645f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_301 N_SCD_c_284_n N_A_181_47#_c_2073_n 2.6495e-19 $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_302 N_SCD_c_283_n N_VGND_c_2268_n 0.00480402f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_303 N_SCD_c_284_n N_VGND_c_2268_n 0.0218413f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_304 SCD N_VGND_c_2268_n 0.0221354f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_305 SCD N_VGND_c_2275_n 9.88088e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_306 N_SCE_M1012_g N_D_c_424_n 0.0160455f $X=0.83 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_307 N_SCE_c_317_n N_D_M1004_g 0.0911662f $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_308 SCE N_D_M1004_g 6.11571e-19 $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_309 N_SCE_M1012_g D 0.00302957f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_310 N_SCE_c_317_n D 0.00293745f $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_311 SCE D 0.0531526f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_312 N_SCE_c_320_n D 0.023169f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_313 N_SCE_c_340_n D 0.00219522f $X=0.835 $Y=1.19 $X2=0 $Y2=0
cc_314 N_SCE_M1012_g N_D_c_427_n 0.0194304f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_315 SCE N_D_c_427_n 3.39482e-19 $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_316 N_SCE_c_320_n N_D_c_427_n 0.00134139f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_317 N_SCE_c_320_n N_A_319_21#_c_466_n 0.00255736f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_318 N_SCE_M1026_g N_A_319_21#_c_467_n 0.00659955f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_319 N_SCE_M1013_g N_A_319_21#_c_467_n 0.00270542f $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_320 N_SCE_c_320_n N_A_319_21#_c_467_n 0.0170338f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_321 N_SCE_c_356_p N_A_319_21#_c_467_n 6.89964e-19 $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_322 N_SCE_c_321_n N_A_319_21#_c_467_n 0.00247217f $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_SCE_c_322_n N_A_319_21#_c_467_n 0.0398183f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_324 N_SCE_c_320_n N_A_319_21#_c_468_n 0.00396034f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_325 N_SCE_c_321_n N_A_319_21#_c_468_n 0.0212905f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_326 N_SCE_c_322_n N_A_319_21#_c_468_n 7.06022e-19 $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_SCE_M1013_g N_A_319_21#_c_469_n 0.00531082f $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_328 N_SCE_c_320_n N_A_319_21#_c_469_n 0.00905152f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_329 N_SCE_c_356_p N_A_319_21#_c_469_n 0.00104259f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_330 N_SCE_c_321_n N_A_319_21#_c_469_n 0.002964f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_331 N_SCE_c_322_n N_A_319_21#_c_469_n 0.00979853f $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_SCE_M1013_g N_A_319_21#_c_470_n 0.00284252f $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_333 N_SCE_M1026_g N_A_319_21#_c_476_n 0.00209962f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_334 N_SCE_c_321_n N_A_319_21#_c_476_n 4.82439e-19 $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_335 N_SCE_c_322_n N_A_319_21#_c_476_n 0.0105043f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_336 N_SCE_M1013_g N_CLK_c_542_n 0.00166043f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_337 N_SCE_M1013_g CLK 0.00584669f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_338 N_SCE_M1026_g CLK 0.00891234f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_339 N_SCE_M1026_g CLK 0.00218466f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_340 N_SCE_c_356_p CLK 0.0017785f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_341 N_SCE_c_321_n CLK 0.00323603f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_342 N_SCE_c_322_n CLK 0.0351412f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_343 N_SCE_M1026_g N_CLK_c_545_n 0.00124122f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_344 N_SCE_c_321_n N_CLK_c_545_n 0.00327928f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_345 N_SCE_c_322_n N_CLK_c_545_n 3.62704e-19 $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_346 N_SCE_c_321_n N_CLK_c_546_n 0.00166043f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_347 N_SCE_M1026_g N_A_643_369#_c_646_n 0.00345048f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_348 N_SCE_M1013_g N_A_643_369#_c_619_n 0.00346504f $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_349 N_SCE_M1026_g N_A_643_369#_c_635_n 0.00127534f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_350 N_SCE_M1013_g N_A_643_369#_c_621_n 5.16475e-19 $X=2.64 $Y=0.445 $X2=0
+ $Y2=0
cc_351 N_SCE_c_317_n N_A_27_369#_c_1811_n 7.65221e-19 $X=0.89 $Y=1.415 $X2=0
+ $Y2=0
cc_352 N_SCE_M1002_g N_A_27_369#_c_1811_n 0.0123242f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_353 SCE N_A_27_369#_c_1811_n 0.0185939f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_354 N_SCE_c_320_n N_A_27_369#_c_1811_n 0.00666807f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_355 N_SCE_c_340_n N_A_27_369#_c_1811_n 0.00141465f $X=0.835 $Y=1.19 $X2=0
+ $Y2=0
cc_356 N_SCE_M1002_g N_A_27_369#_c_1818_n 0.00487221f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_357 N_SCE_M1002_g N_A_27_369#_c_1825_n 0.00389743f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_358 N_SCE_M1002_g N_VPWR_c_1852_n 0.00292936f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_359 N_SCE_M1026_g N_VPWR_c_1853_n 0.00501988f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_360 N_SCE_M1002_g N_VPWR_c_1861_n 0.00428647f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_361 N_SCE_M1026_g N_VPWR_c_1861_n 0.00585385f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_362 N_SCE_M1002_g N_VPWR_c_1851_n 0.00564895f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_363 N_SCE_M1026_g N_VPWR_c_1851_n 0.0132032f $X=2.61 $Y=2.165 $X2=0 $Y2=0
cc_364 N_SCE_M1012_g N_A_181_47#_c_2073_n 0.00497883f $X=0.83 $Y=0.445 $X2=0
+ $Y2=0
cc_365 N_SCE_c_317_n N_A_181_47#_c_2073_n 9.02625e-19 $X=0.89 $Y=1.415 $X2=0
+ $Y2=0
cc_366 N_SCE_c_320_n N_A_181_47#_c_2073_n 0.00870107f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_367 N_SCE_c_320_n N_A_181_47#_c_2077_n 0.00434157f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_368 N_SCE_c_320_n N_A_181_47#_c_2063_n 0.00452657f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_369 N_SCE_M1026_g N_A_181_47#_c_2069_n 0.00616318f $X=2.61 $Y=2.165 $X2=0
+ $Y2=0
cc_370 N_SCE_c_320_n N_A_181_47#_c_2069_n 0.0490896f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_371 N_SCE_c_356_p N_A_181_47#_c_2069_n 0.0249445f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_372 N_SCE_c_321_n N_A_181_47#_c_2069_n 4.55029e-19 $X=2.535 $Y=1.16 $X2=0
+ $Y2=0
cc_373 N_SCE_c_322_n N_A_181_47#_c_2069_n 0.017172f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_374 N_SCE_c_320_n N_A_181_47#_c_2070_n 0.0258361f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_375 N_SCE_c_320_n N_A_181_47#_c_2065_n 0.0179698f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_376 N_SCE_M1013_g N_VGND_c_2250_n 0.00193415f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_377 N_SCE_c_320_n N_VGND_c_2250_n 0.00127321f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_378 N_SCE_M1013_g N_VGND_c_2251_n 0.00958993f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_379 N_SCE_c_322_n N_VGND_c_2251_n 2.63385e-19 $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_380 N_SCE_M1012_g N_VGND_c_2258_n 0.005323f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_381 N_SCE_M1013_g N_VGND_c_2262_n 0.00486043f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_382 N_SCE_M1012_g N_VGND_c_2268_n 0.00412734f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_383 N_SCE_c_317_n N_VGND_c_2268_n 3.91104e-19 $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_384 SCE N_VGND_c_2268_n 0.0111408f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_385 N_SCE_c_340_n N_VGND_c_2268_n 6.88562e-19 $X=0.835 $Y=1.19 $X2=0 $Y2=0
cc_386 N_SCE_M1012_g N_VGND_c_2275_n 0.00728858f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_387 N_SCE_M1013_g N_VGND_c_2275_n 0.00965187f $X=2.64 $Y=0.445 $X2=0 $Y2=0
cc_388 SCE N_VGND_c_2275_n 0.00510613f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_389 N_D_c_424_n N_A_319_21#_M1031_g 0.0310205f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_390 D N_A_319_21#_M1031_g 3.21313e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_391 N_D_c_427_n N_A_319_21#_M1031_g 0.020121f $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_392 N_D_M1004_g N_A_319_21#_c_466_n 0.056689f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_393 D N_A_319_21#_c_466_n 0.00150183f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_394 D N_A_27_369#_c_1811_n 0.00629694f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_395 N_D_M1004_g N_A_27_369#_c_1813_n 0.012106f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_396 D N_A_27_369#_c_1813_n 0.00435308f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_397 N_D_M1004_g N_VPWR_c_1861_n 0.00357877f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_398 N_D_M1004_g N_VPWR_c_1851_n 0.00515774f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_399 N_D_c_424_n N_A_181_47#_c_2073_n 0.0121647f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_400 D N_A_181_47#_c_2073_n 0.0192899f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_401 N_D_c_427_n N_A_181_47#_c_2073_n 2.99729e-19 $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_402 N_D_M1004_g N_A_181_47#_c_2077_n 0.00326172f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_403 D N_A_181_47#_c_2077_n 0.00267197f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_404 N_D_c_424_n N_A_181_47#_c_2063_n 0.00357781f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_405 D N_A_181_47#_c_2063_n 0.00301423f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_406 N_D_c_427_n N_A_181_47#_c_2063_n 3.93323e-19 $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_407 D N_A_181_47#_c_2070_n 0.00763475f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_408 N_D_M1004_g N_A_181_47#_c_2065_n 0.00514875f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_409 D N_A_181_47#_c_2065_n 0.0638647f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_410 N_D_c_427_n N_A_181_47#_c_2065_n 0.00166259f $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_411 N_D_c_424_n N_VGND_c_2258_n 0.00357877f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_412 N_D_c_424_n N_VGND_c_2275_n 0.00528062f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_413 N_A_319_21#_c_469_n CLK 0.00859062f $X=2.39 $Y=0.715 $X2=0 $Y2=0
cc_414 N_A_319_21#_c_476_n CLK 0.00581744f $X=2.4 $Y=1.99 $X2=0 $Y2=0
cc_415 N_A_319_21#_c_476_n N_A_27_369#_M1001_d 0.00519628f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_416 N_A_319_21#_M1001_g N_A_27_369#_c_1813_n 0.00914137f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_417 N_A_319_21#_c_475_n N_A_27_369#_c_1813_n 0.0148151f $X=2.395 $Y=1.927
+ $X2=0 $Y2=0
cc_418 N_A_319_21#_c_476_n N_A_27_369#_c_1813_n 0.0132953f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_419 N_A_319_21#_M1001_g N_VPWR_c_1861_n 0.00357877f $X=1.67 $Y=2.165 $X2=0
+ $Y2=0
cc_420 N_A_319_21#_c_475_n N_VPWR_c_1861_n 0.0154197f $X=2.395 $Y=1.927 $X2=0
+ $Y2=0
cc_421 N_A_319_21#_c_476_n N_VPWR_c_1861_n 0.00432835f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_422 N_A_319_21#_M1026_s N_VPWR_c_1851_n 0.00261392f $X=2.275 $Y=1.845 $X2=0
+ $Y2=0
cc_423 N_A_319_21#_M1001_g N_VPWR_c_1851_n 0.00657948f $X=1.67 $Y=2.165 $X2=0
+ $Y2=0
cc_424 N_A_319_21#_c_475_n N_VPWR_c_1851_n 0.00941222f $X=2.395 $Y=1.927 $X2=0
+ $Y2=0
cc_425 N_A_319_21#_c_476_n N_VPWR_c_1851_n 0.00699224f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_426 N_A_319_21#_M1001_g N_A_181_47#_c_2077_n 0.00536988f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_427 N_A_319_21#_c_476_n N_A_181_47#_c_2077_n 0.0199612f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_428 N_A_319_21#_M1031_g N_A_181_47#_c_2063_n 0.0158472f $X=1.67 $Y=0.445
+ $X2=0 $Y2=0
cc_429 N_A_319_21#_c_469_n N_A_181_47#_c_2063_n 0.00724643f $X=2.39 $Y=0.715
+ $X2=0 $Y2=0
cc_430 N_A_319_21#_c_470_n N_A_181_47#_c_2063_n 0.00506574f $X=2.43 $Y=0.44
+ $X2=0 $Y2=0
cc_431 N_A_319_21#_c_467_n N_A_181_47#_c_2069_n 0.0169458f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_432 N_A_319_21#_c_468_n N_A_181_47#_c_2069_n 0.00172463f $X=1.95 $Y=1.16
+ $X2=0 $Y2=0
cc_433 N_A_319_21#_c_476_n N_A_181_47#_c_2069_n 0.0111897f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_434 N_A_319_21#_M1001_g N_A_181_47#_c_2070_n 0.00423017f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_435 N_A_319_21#_c_467_n N_A_181_47#_c_2070_n 0.0027962f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_436 N_A_319_21#_M1031_g N_A_181_47#_c_2065_n 0.00370215f $X=1.67 $Y=0.445
+ $X2=0 $Y2=0
cc_437 N_A_319_21#_M1001_g N_A_181_47#_c_2065_n 0.0103628f $X=1.67 $Y=2.165
+ $X2=0 $Y2=0
cc_438 N_A_319_21#_c_466_n N_A_181_47#_c_2065_n 0.0084262f $X=1.67 $Y=1.16 $X2=0
+ $Y2=0
cc_439 N_A_319_21#_c_467_n N_A_181_47#_c_2065_n 0.0614598f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_440 N_A_319_21#_c_469_n N_A_181_47#_c_2065_n 0.00798473f $X=2.39 $Y=0.715
+ $X2=0 $Y2=0
cc_441 N_A_319_21#_c_476_n N_A_181_47#_c_2065_n 0.00599428f $X=2.4 $Y=1.99 $X2=0
+ $Y2=0
cc_442 N_A_319_21#_M1031_g N_VGND_c_2250_n 0.005626f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_443 N_A_319_21#_c_468_n N_VGND_c_2250_n 0.00128608f $X=1.95 $Y=1.16 $X2=0
+ $Y2=0
cc_444 N_A_319_21#_c_469_n N_VGND_c_2250_n 0.0174596f $X=2.39 $Y=0.715 $X2=0
+ $Y2=0
cc_445 N_A_319_21#_c_470_n N_VGND_c_2250_n 0.0233255f $X=2.43 $Y=0.44 $X2=0
+ $Y2=0
cc_446 N_A_319_21#_M1031_g N_VGND_c_2258_n 0.00464258f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_447 N_A_319_21#_c_469_n N_VGND_c_2262_n 0.00268684f $X=2.39 $Y=0.715 $X2=0
+ $Y2=0
cc_448 N_A_319_21#_c_470_n N_VGND_c_2262_n 0.0173307f $X=2.43 $Y=0.44 $X2=0
+ $Y2=0
cc_449 N_A_319_21#_M1013_s N_VGND_c_2275_n 0.0036554f $X=2.305 $Y=0.235 $X2=0
+ $Y2=0
cc_450 N_A_319_21#_M1031_g N_VGND_c_2275_n 0.00862073f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_451 N_A_319_21#_c_469_n N_VGND_c_2275_n 0.00551711f $X=2.39 $Y=0.715 $X2=0
+ $Y2=0
cc_452 N_A_319_21#_c_470_n N_VGND_c_2275_n 0.00983733f $X=2.43 $Y=0.44 $X2=0
+ $Y2=0
cc_453 N_CLK_c_547_n N_A_643_369#_M1029_g 0.00719527f $X=3.52 $Y=1.62 $X2=0
+ $Y2=0
cc_454 N_CLK_c_548_n N_A_643_369#_M1029_g 0.0304072f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_455 CLK N_A_643_369#_M1029_g 2.61881e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_456 N_CLK_c_541_n N_A_643_369#_c_614_n 0.0138105f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_457 N_CLK_c_542_n N_A_643_369#_c_618_n 0.00767217f $X=3.58 $Y=0.805 $X2=0
+ $Y2=0
cc_458 N_CLK_c_541_n N_A_643_369#_c_619_n 0.00270983f $X=3.58 $Y=0.73 $X2=0
+ $Y2=0
cc_459 N_CLK_c_548_n N_A_643_369#_c_634_n 0.0140471f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_460 CLK N_A_643_369#_c_634_n 0.00782756f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_461 N_CLK_c_548_n N_A_643_369#_c_635_n 3.1659e-19 $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_462 CLK N_A_643_369#_c_635_n 0.0108188f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_463 CLK N_A_643_369#_c_635_n 0.0113567f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_464 N_CLK_c_545_n N_A_643_369#_c_635_n 5.89316e-19 $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_465 N_CLK_c_541_n N_A_643_369#_c_620_n 0.00390588f $X=3.58 $Y=0.73 $X2=0
+ $Y2=0
cc_466 N_CLK_c_542_n N_A_643_369#_c_620_n 0.00637134f $X=3.58 $Y=0.805 $X2=0
+ $Y2=0
cc_467 CLK N_A_643_369#_c_620_n 0.00797093f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_468 N_CLK_c_546_n N_A_643_369#_c_620_n 0.00151794f $X=3.43 $Y=1.09 $X2=0
+ $Y2=0
cc_469 N_CLK_c_542_n N_A_643_369#_c_621_n 0.00352145f $X=3.58 $Y=0.805 $X2=0
+ $Y2=0
cc_470 CLK N_A_643_369#_c_621_n 0.0136403f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_471 CLK N_A_643_369#_c_621_n 0.0161115f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_472 N_CLK_c_545_n N_A_643_369#_c_621_n 8.54762e-19 $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_473 N_CLK_c_546_n N_A_643_369#_c_621_n 5.61645e-19 $X=3.43 $Y=1.09 $X2=0
+ $Y2=0
cc_474 N_CLK_c_548_n N_A_643_369#_c_622_n 0.0025963f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_475 CLK N_A_643_369#_c_622_n 0.0052596f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_476 CLK N_A_643_369#_c_622_n 0.0064932f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_477 CLK N_A_643_369#_c_622_n 0.0439523f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_478 N_CLK_c_546_n N_A_643_369#_c_622_n 0.0037422f $X=3.43 $Y=1.09 $X2=0 $Y2=0
cc_479 CLK N_A_643_369#_c_623_n 3.7897e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_480 N_CLK_c_545_n N_A_643_369#_c_623_n 0.0213743f $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_481 N_CLK_c_546_n N_A_643_369#_c_630_n 0.0064798f $X=3.43 $Y=1.09 $X2=0 $Y2=0
cc_482 CLK N_VPWR_M1026_d 0.00205142f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_483 N_CLK_c_548_n N_VPWR_c_1853_n 0.00394857f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_484 CLK N_VPWR_c_1853_n 0.00606401f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_485 N_CLK_c_548_n N_VPWR_c_1854_n 0.00836773f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_486 N_CLK_c_548_n N_VPWR_c_1868_n 0.00348948f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_487 CLK N_VPWR_c_1868_n 0.00148905f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_488 N_CLK_c_548_n N_VPWR_c_1851_n 0.00553267f $X=3.52 $Y=1.77 $X2=0 $Y2=0
cc_489 CLK N_VPWR_c_1851_n 0.00297482f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_490 N_CLK_c_547_n N_A_181_47#_c_2069_n 0.00100904f $X=3.52 $Y=1.62 $X2=0
+ $Y2=0
cc_491 N_CLK_c_548_n N_A_181_47#_c_2069_n 0.00182678f $X=3.52 $Y=1.77 $X2=0
+ $Y2=0
cc_492 CLK N_A_181_47#_c_2069_n 5.20642e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_493 CLK N_A_181_47#_c_2069_n 0.00387206f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_494 CLK N_A_181_47#_c_2069_n 0.0427426f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_495 N_CLK_c_541_n N_VGND_c_2251_n 0.00224354f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_496 CLK N_VGND_c_2251_n 0.0163599f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_497 N_CLK_c_541_n N_VGND_c_2252_n 0.00767804f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_498 N_CLK_c_541_n N_VGND_c_2263_n 0.00348405f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_499 N_CLK_c_542_n N_VGND_c_2263_n 2.82692e-19 $X=3.58 $Y=0.805 $X2=0 $Y2=0
cc_500 N_CLK_c_541_n N_VGND_c_2275_n 0.00552264f $X=3.58 $Y=0.73 $X2=0 $Y2=0
cc_501 CLK N_VGND_c_2275_n 7.78553e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_502 N_A_643_369#_c_640_n N_A_809_369#_M1029_d 0.00106464f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_503 N_A_643_369#_c_641_n N_A_809_369#_M1029_d 4.96569e-19 $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_504 N_A_643_369#_M1029_g N_A_809_369#_c_909_n 0.0121191f $X=3.97 $Y=2.165
+ $X2=0 $Y2=0
cc_505 N_A_643_369#_c_640_n N_A_809_369#_c_909_n 0.00114519f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_506 N_A_643_369#_c_644_n N_A_809_369#_c_909_n 0.0032436f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_507 N_A_643_369#_c_644_n N_A_809_369#_c_899_n 0.0085606f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_508 N_A_643_369#_c_645_n N_A_809_369#_c_899_n 2.0638e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_509 N_A_643_369#_c_616_n N_A_809_369#_M1021_g 0.0193318f $X=4.94 $Y=0.73
+ $X2=0 $Y2=0
cc_510 N_A_643_369#_M1017_g N_A_809_369#_M1044_g 0.0141749f $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_511 N_A_643_369#_M1033_g N_A_809_369#_M1044_g 0.0173162f $X=9 $Y=0.445 $X2=0
+ $Y2=0
cc_512 N_A_643_369#_c_624_n N_A_809_369#_M1044_g 0.00869456f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_513 N_A_643_369#_c_625_n N_A_809_369#_M1044_g 0.0206167f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_514 N_A_643_369#_c_626_n N_A_809_369#_M1044_g 0.0157656f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_515 N_A_643_369#_c_628_n N_A_809_369#_M1044_g 0.00142299f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_516 N_A_643_369#_c_629_n N_A_809_369#_M1044_g 0.0109721f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_517 N_A_643_369#_M1017_g N_A_809_369#_c_912_n 0.00409586f $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_518 N_A_643_369#_c_626_n N_A_809_369#_c_912_n 0.00124923f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_519 N_A_643_369#_c_696_p N_A_809_369#_c_912_n 0.00205153f $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_520 N_A_643_369#_M1017_g N_A_809_369#_M1034_g 0.0125619f $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_521 N_A_643_369#_c_696_p N_A_809_369#_M1034_g 0.00121481f $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_522 N_A_643_369#_M1038_g N_A_809_369#_c_914_n 0.0161622f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_523 N_A_643_369#_c_640_n N_A_809_369#_c_914_n 0.00565079f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_524 N_A_643_369#_c_643_n N_A_809_369#_c_914_n 7.24988e-19 $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_525 N_A_643_369#_c_644_n N_A_809_369#_c_914_n 0.00461659f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_526 N_A_643_369#_c_645_n N_A_809_369#_c_914_n 5.74415e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_527 N_A_643_369#_c_640_n N_A_809_369#_c_915_n 0.00228522f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_528 N_A_643_369#_M1029_g N_A_809_369#_c_916_n 0.00920763f $X=3.97 $Y=2.165
+ $X2=0 $Y2=0
cc_529 N_A_643_369#_c_706_p N_A_809_369#_c_916_n 0.0115657f $X=3.865 $Y=1.83
+ $X2=0 $Y2=0
cc_530 N_A_643_369#_c_640_n N_A_809_369#_c_916_n 0.0191192f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_531 N_A_643_369#_c_641_n N_A_809_369#_c_916_n 0.00278251f $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_532 N_A_643_369#_c_615_n N_A_809_369#_c_902_n 0.00100605f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_533 N_A_643_369#_c_624_n N_A_809_369#_c_902_n 0.023168f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_534 N_A_643_369#_c_625_n N_A_809_369#_c_902_n 0.00288312f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_535 N_A_643_369#_c_626_n N_A_809_369#_c_902_n 0.0116627f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_536 N_A_643_369#_c_640_n N_A_809_369#_c_902_n 0.0075219f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_537 N_A_643_369#_c_642_n N_A_809_369#_c_902_n 0.047224f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_538 N_A_643_369#_c_643_n N_A_809_369#_c_902_n 0.0126603f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_539 N_A_643_369#_c_645_n N_A_809_369#_c_902_n 6.70475e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_540 N_A_643_369#_c_615_n N_A_809_369#_c_903_n 0.00234075f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_541 N_A_643_369#_c_622_n N_A_809_369#_c_903_n 0.00138833f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_542 N_A_643_369#_c_615_n N_A_809_369#_c_904_n 0.00183262f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_543 N_A_643_369#_c_623_n N_A_809_369#_c_904_n 0.0031868f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_544 N_A_643_369#_c_624_n N_A_809_369#_c_905_n 0.00209286f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_545 N_A_643_369#_c_626_n N_A_809_369#_c_905_n 0.00487486f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_546 N_A_643_369#_c_628_n N_A_809_369#_c_905_n 0.00614212f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_547 N_A_643_369#_c_629_n N_A_809_369#_c_905_n 0.00367564f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_548 N_A_643_369#_M1017_g N_A_809_369#_c_906_n 6.25086e-19 $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_549 N_A_643_369#_c_624_n N_A_809_369#_c_906_n 0.0254561f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_550 N_A_643_369#_c_625_n N_A_809_369#_c_906_n 4.15885e-19 $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_551 N_A_643_369#_c_626_n N_A_809_369#_c_906_n 0.0149273f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_552 N_A_643_369#_c_628_n N_A_809_369#_c_906_n 0.0116275f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_553 N_A_643_369#_c_629_n N_A_809_369#_c_906_n 0.00117508f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_554 N_A_643_369#_c_696_p N_A_809_369#_c_906_n 0.0125472f $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_555 N_A_643_369#_c_615_n N_A_809_369#_c_907_n 0.0487935f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_556 N_A_643_369#_c_622_n N_A_809_369#_c_907_n 3.00848e-19 $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_557 N_A_643_369#_c_623_n N_A_809_369#_c_907_n 0.0203131f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_558 N_A_643_369#_c_614_n N_A_809_369#_c_908_n 0.00458005f $X=4 $Y=0.73 $X2=0
+ $Y2=0
cc_559 N_A_643_369#_c_615_n N_A_809_369#_c_908_n 0.0132045f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_560 N_A_643_369#_c_620_n N_A_809_369#_c_908_n 0.0129402f $X=3.735 $Y=0.8
+ $X2=0 $Y2=0
cc_561 N_A_643_369#_c_622_n N_A_809_369#_c_908_n 0.0686527f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_562 N_A_643_369#_c_630_n N_A_809_369#_c_908_n 0.0031868f $X=3.917 $Y=1.09
+ $X2=0 $Y2=0
cc_563 N_A_643_369#_M1038_g N_A_1129_21#_M1040_g 0.0211742f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_564 N_A_643_369#_c_642_n N_A_1129_21#_M1040_g 0.00306453f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_565 N_A_643_369#_c_642_n N_A_1129_21#_c_1085_n 0.0108654f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_566 N_A_643_369#_c_642_n N_A_1129_21#_c_1086_n 0.00401276f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_567 N_A_643_369#_c_644_n N_A_1129_21#_c_1086_n 0.0130435f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_568 N_A_643_369#_c_696_p N_A_1129_21#_c_1087_n 8.15517e-19 $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_569 N_A_643_369#_c_642_n N_A_1129_21#_c_1087_n 0.0251481f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_570 N_A_643_369#_c_642_n N_A_1129_21#_c_1088_n 0.00322176f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_571 N_A_643_369#_c_642_n N_A_997_413#_M1005_g 0.00379884f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_572 N_A_643_369#_M1017_g N_A_997_413#_M1011_g 0.0521194f $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_573 N_A_643_369#_c_624_n N_A_997_413#_M1011_g 0.0025506f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_574 N_A_643_369#_c_696_p N_A_997_413#_M1011_g 0.0141577f $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_575 N_A_643_369#_c_752_p N_A_997_413#_M1011_g 0.00166615f $X=7.645 $Y=1.87
+ $X2=0 $Y2=0
cc_576 N_A_643_369#_c_615_n N_A_997_413#_c_1176_n 0.0042049f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_577 N_A_643_369#_c_616_n N_A_997_413#_c_1176_n 0.00613402f $X=4.94 $Y=0.73
+ $X2=0 $Y2=0
cc_578 N_A_643_369#_M1038_g N_A_997_413#_c_1201_n 0.0121756f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_579 N_A_643_369#_c_640_n N_A_997_413#_c_1201_n 0.00362812f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_580 N_A_643_369#_c_642_n N_A_997_413#_c_1201_n 0.00492445f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_581 N_A_643_369#_c_643_n N_A_997_413#_c_1201_n 0.00506476f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_582 N_A_643_369#_c_644_n N_A_997_413#_c_1201_n 9.46198e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_583 N_A_643_369#_c_645_n N_A_997_413#_c_1201_n 0.0108411f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_584 N_A_643_369#_M1038_g N_A_997_413#_c_1187_n 0.00392912f $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_585 N_A_643_369#_c_642_n N_A_997_413#_c_1187_n 0.0149262f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_586 N_A_643_369#_c_643_n N_A_997_413#_c_1187_n 0.00307458f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_587 N_A_643_369#_c_644_n N_A_997_413#_c_1187_n 0.00212617f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_588 N_A_643_369#_c_645_n N_A_997_413#_c_1187_n 0.0263544f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_589 N_A_643_369#_c_640_n N_A_997_413#_c_1177_n 0.00396196f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_590 N_A_643_369#_c_642_n N_A_997_413#_c_1177_n 0.00354029f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_591 N_A_643_369#_c_643_n N_A_997_413#_c_1177_n 0.0032583f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_592 N_A_643_369#_c_644_n N_A_997_413#_c_1177_n 0.00293864f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_593 N_A_643_369#_c_645_n N_A_997_413#_c_1177_n 0.014754f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_594 N_A_643_369#_c_624_n N_A_997_413#_c_1178_n 0.0270221f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_595 N_A_643_369#_c_625_n N_A_997_413#_c_1178_n 0.00191823f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_596 N_A_643_369#_c_696_p N_A_997_413#_c_1178_n 0.00984522f $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_597 N_A_643_369#_c_642_n N_A_997_413#_c_1178_n 0.00128054f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_598 N_A_643_369#_c_642_n N_A_997_413#_c_1180_n 0.0077952f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_599 N_A_643_369#_c_624_n N_A_997_413#_c_1182_n 3.87262e-19 $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_600 N_A_643_369#_c_625_n N_A_997_413#_c_1182_n 0.0521194f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_601 N_A_643_369#_c_696_p N_A_997_413#_c_1182_n 0.00160602f $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_602 N_A_643_369#_c_624_n N_A_997_413#_c_1184_n 0.00223303f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_603 N_A_643_369#_c_627_n N_A_997_413#_c_1184_n 0.00403072f $X=8.135 $Y=0.812
+ $X2=0 $Y2=0
cc_604 N_A_643_369#_c_642_n N_SET_B_M1030_g 0.00452095f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_605 N_A_643_369#_M1017_g N_SET_B_c_1329_n 0.00161248f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_606 N_A_643_369#_c_624_n N_SET_B_c_1329_n 0.0216722f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_607 N_A_643_369#_c_626_n N_SET_B_c_1329_n 0.00356101f $X=8.82 $Y=0.812 $X2=0
+ $Y2=0
cc_608 N_A_643_369#_c_628_n N_SET_B_c_1329_n 0.00179525f $X=8.94 $Y=1.09 $X2=0
+ $Y2=0
cc_609 N_A_643_369#_c_629_n N_SET_B_c_1329_n 3.78285e-19 $X=8.94 $Y=1.09 $X2=0
+ $Y2=0
cc_610 N_A_643_369#_c_696_p N_SET_B_c_1329_n 0.0121308f $X=7.885 $Y=1.812 $X2=0
+ $Y2=0
cc_611 N_A_643_369#_c_642_n N_SET_B_c_1329_n 0.0499417f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_612 N_A_643_369#_c_752_p N_SET_B_c_1329_n 0.0261637f $X=7.645 $Y=1.87 $X2=0
+ $Y2=0
cc_613 N_A_643_369#_c_642_n N_SET_B_c_1330_n 0.0265307f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_614 N_A_643_369#_c_628_n N_SET_B_c_1331_n 0.00630037f $X=8.94 $Y=1.09 $X2=0
+ $Y2=0
cc_615 N_A_643_369#_c_628_n N_SET_B_c_1332_n 0.0155825f $X=8.94 $Y=1.09 $X2=0
+ $Y2=0
cc_616 N_A_643_369#_c_629_n N_SET_B_c_1332_n 6.03712e-19 $X=8.94 $Y=1.09 $X2=0
+ $Y2=0
cc_617 N_A_643_369#_c_696_p N_SET_B_c_1333_n 0.00427048f $X=7.885 $Y=1.812 $X2=0
+ $Y2=0
cc_618 N_A_643_369#_c_642_n N_SET_B_c_1333_n 0.00390363f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_619 N_A_643_369#_c_696_p N_SET_B_c_1334_n 0.00821773f $X=7.885 $Y=1.812 $X2=0
+ $Y2=0
cc_620 N_A_643_369#_c_642_n N_SET_B_c_1334_n 0.00855439f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_621 N_A_643_369#_c_629_n N_A_1781_295#_c_1465_n 0.0104506f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_622 N_A_643_369#_M1033_g N_A_1781_295#_M1035_g 0.0362711f $X=9 $Y=0.445 $X2=0
+ $Y2=0
cc_623 N_A_643_369#_c_626_n N_A_1781_295#_M1035_g 0.00188431f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_624 N_A_643_369#_M1033_g N_A_1781_295#_c_1457_n 3.86539e-19 $X=9 $Y=0.445
+ $X2=0 $Y2=0
cc_625 N_A_643_369#_c_626_n N_A_1781_295#_c_1457_n 0.00343189f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_626 N_A_643_369#_c_628_n N_A_1781_295#_c_1457_n 0.0180302f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_627 N_A_643_369#_c_628_n N_A_1781_295#_c_1458_n 0.00202933f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_628 N_A_643_369#_c_629_n N_A_1781_295#_c_1458_n 0.0362711f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_629 N_A_643_369#_c_628_n N_A_1781_295#_c_1468_n 0.00398684f $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_630 N_A_643_369#_c_626_n N_A_1597_329#_M1044_d 0.00212707f $X=8.82 $Y=0.812
+ $X2=-0.19 $Y2=-0.24
cc_631 N_A_643_369#_c_624_n N_A_1597_329#_M1017_d 2.5336e-19 $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_632 N_A_643_369#_c_696_p N_A_1597_329#_M1017_d 0.00547966f $X=7.885 $Y=1.812
+ $X2=0 $Y2=0
cc_633 N_A_643_369#_M1017_g N_A_1597_329#_c_1588_n 0.00138656f $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_634 N_A_643_369#_M1033_g N_A_1597_329#_c_1589_n 0.0142183f $X=9 $Y=0.445
+ $X2=0 $Y2=0
cc_635 N_A_643_369#_c_626_n N_A_1597_329#_c_1589_n 0.0389425f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_636 N_A_643_369#_c_629_n N_A_1597_329#_c_1589_n 4.18621e-19 $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_637 N_A_643_369#_c_626_n N_A_1597_329#_c_1568_n 0.00224983f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_638 N_A_643_369#_c_626_n N_A_1597_329#_c_1569_n 0.00266946f $X=8.82 $Y=0.812
+ $X2=0 $Y2=0
cc_639 N_A_643_369#_c_628_n N_A_1597_329#_c_1580_n 7.54131e-19 $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_640 N_A_643_369#_c_629_n N_A_1597_329#_c_1580_n 3.84956e-19 $X=8.94 $Y=1.09
+ $X2=0 $Y2=0
cc_641 N_A_643_369#_c_634_n N_VPWR_M1036_d 6.64995e-19 $X=3.735 $Y=1.915 $X2=0
+ $Y2=0
cc_642 N_A_643_369#_c_706_p N_VPWR_M1036_d 0.00137413f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_643 N_A_643_369#_c_696_p N_VPWR_M1030_d 0.00884603f $X=7.885 $Y=1.812 $X2=0
+ $Y2=0
cc_644 N_A_643_369#_c_646_n N_VPWR_c_1853_n 0.0102695f $X=3.34 $Y=2.16 $X2=0
+ $Y2=0
cc_645 N_A_643_369#_M1029_g N_VPWR_c_1854_n 0.00819473f $X=3.97 $Y=2.165 $X2=0
+ $Y2=0
cc_646 N_A_643_369#_c_634_n N_VPWR_c_1854_n 0.00397675f $X=3.735 $Y=1.915 $X2=0
+ $Y2=0
cc_647 N_A_643_369#_c_706_p N_VPWR_c_1854_n 0.00628707f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_648 N_A_643_369#_c_641_n N_VPWR_c_1854_n 8.45658e-19 $X=4.055 $Y=1.87 $X2=0
+ $Y2=0
cc_649 N_A_643_369#_c_646_n N_VPWR_c_1868_n 0.00593494f $X=3.34 $Y=2.16 $X2=0
+ $Y2=0
cc_650 N_A_643_369#_c_634_n N_VPWR_c_1868_n 0.0020032f $X=3.735 $Y=1.915 $X2=0
+ $Y2=0
cc_651 N_A_643_369#_M1029_g N_VPWR_c_1869_n 0.0039838f $X=3.97 $Y=2.165 $X2=0
+ $Y2=0
cc_652 N_A_643_369#_M1038_g N_VPWR_c_1869_n 0.00357877f $X=5.33 $Y=2.275 $X2=0
+ $Y2=0
cc_653 N_A_643_369#_c_706_p N_VPWR_c_1869_n 0.00102589f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_654 N_A_643_369#_c_642_n N_VPWR_c_1875_n 0.00139085f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_655 N_A_643_369#_M1017_g N_VPWR_c_1877_n 0.0199583f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_656 N_A_643_369#_c_696_p N_VPWR_c_1877_n 0.0428613f $X=7.885 $Y=1.812 $X2=0
+ $Y2=0
cc_657 N_A_643_369#_c_642_n N_VPWR_c_1877_n 0.00782266f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_658 N_A_643_369#_c_752_p N_VPWR_c_1877_n 0.00338024f $X=7.645 $Y=1.87 $X2=0
+ $Y2=0
cc_659 N_A_643_369#_M1036_s N_VPWR_c_1851_n 0.00387904f $X=3.215 $Y=1.845 $X2=0
+ $Y2=0
cc_660 N_A_643_369#_M1029_g N_VPWR_c_1851_n 0.00530391f $X=3.97 $Y=2.165 $X2=0
+ $Y2=0
cc_661 N_A_643_369#_M1038_g N_VPWR_c_1851_n 0.00539327f $X=5.33 $Y=2.275 $X2=0
+ $Y2=0
cc_662 N_A_643_369#_c_646_n N_VPWR_c_1851_n 0.00591039f $X=3.34 $Y=2.16 $X2=0
+ $Y2=0
cc_663 N_A_643_369#_c_634_n N_VPWR_c_1851_n 0.00457428f $X=3.735 $Y=1.915 $X2=0
+ $Y2=0
cc_664 N_A_643_369#_c_706_p N_VPWR_c_1851_n 0.00152919f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_665 N_A_643_369#_c_696_p N_VPWR_c_1851_n 0.00668331f $X=7.885 $Y=1.812 $X2=0
+ $Y2=0
cc_666 N_A_643_369#_c_640_n N_VPWR_c_1851_n 0.0529901f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_667 N_A_643_369#_c_641_n N_VPWR_c_1851_n 0.0139738f $X=4.055 $Y=1.87 $X2=0
+ $Y2=0
cc_668 N_A_643_369#_c_642_n N_VPWR_c_1851_n 0.0935903f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_669 N_A_643_369#_c_643_n N_VPWR_c_1851_n 0.0156394f $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_670 N_A_643_369#_c_752_p N_VPWR_c_1851_n 0.0143849f $X=7.645 $Y=1.87 $X2=0
+ $Y2=0
cc_671 N_A_643_369#_c_615_n N_A_181_47#_c_2061_n 0.00755734f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_672 N_A_643_369#_c_616_n N_A_181_47#_c_2061_n 0.00248143f $X=4.94 $Y=0.73
+ $X2=0 $Y2=0
cc_673 N_A_643_369#_c_640_n N_A_181_47#_c_2066_n 6.0342e-19 $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_674 N_A_643_369#_c_644_n N_A_181_47#_c_2066_n 2.97118e-19 $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_675 N_A_643_369#_c_645_n N_A_181_47#_c_2066_n 0.00145104f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_676 N_A_643_369#_M1038_g N_A_181_47#_c_2067_n 2.14497e-19 $X=5.33 $Y=2.275
+ $X2=0 $Y2=0
cc_677 N_A_643_369#_c_640_n N_A_181_47#_c_2067_n 0.016219f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_678 N_A_643_369#_c_643_n N_A_181_47#_c_2067_n 0.00279803f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_679 N_A_643_369#_c_644_n N_A_181_47#_c_2067_n 0.00239106f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_680 N_A_643_369#_c_645_n N_A_181_47#_c_2067_n 0.0106345f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_681 N_A_643_369#_c_615_n N_A_181_47#_c_2064_n 0.00896128f $X=4.865 $Y=0.805
+ $X2=0 $Y2=0
cc_682 N_A_643_369#_M1029_g N_A_181_47#_c_2069_n 0.00390687f $X=3.97 $Y=2.165
+ $X2=0 $Y2=0
cc_683 N_A_643_369#_c_618_n N_A_181_47#_c_2069_n 0.00230404f $X=3.992 $Y=0.805
+ $X2=0 $Y2=0
cc_684 N_A_643_369#_c_634_n N_A_181_47#_c_2069_n 0.00799158f $X=3.735 $Y=1.915
+ $X2=0 $Y2=0
cc_685 N_A_643_369#_c_635_n N_A_181_47#_c_2069_n 0.00136429f $X=3.425 $Y=1.915
+ $X2=0 $Y2=0
cc_686 N_A_643_369#_c_620_n N_A_181_47#_c_2069_n 0.00559677f $X=3.735 $Y=0.8
+ $X2=0 $Y2=0
cc_687 N_A_643_369#_c_621_n N_A_181_47#_c_2069_n 7.07979e-19 $X=3.455 $Y=0.8
+ $X2=0 $Y2=0
cc_688 N_A_643_369#_c_622_n N_A_181_47#_c_2069_n 0.0217647f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_689 N_A_643_369#_c_623_n N_A_181_47#_c_2069_n 4.51301e-19 $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_690 N_A_643_369#_c_640_n N_A_181_47#_c_2069_n 0.0490885f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_691 N_A_643_369#_c_641_n N_A_181_47#_c_2069_n 0.0254571f $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_692 N_A_643_369#_c_640_n N_A_181_47#_c_2072_n 0.0264737f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_693 N_A_643_369#_c_644_n N_A_181_47#_c_2072_n 0.00127036f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_694 N_A_643_369#_c_645_n N_A_181_47#_c_2072_n 0.00208921f $X=5.33 $Y=1.74
+ $X2=0 $Y2=0
cc_695 N_A_643_369#_c_696_p A_1525_329# 0.00168642f $X=7.885 $Y=1.812 $X2=-0.19
+ $Y2=-0.24
cc_696 N_A_643_369#_c_752_p A_1525_329# 0.00159132f $X=7.645 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_697 N_A_643_369#_c_619_n N_VGND_c_2251_n 0.0239406f $X=3.37 $Y=0.44 $X2=0
+ $Y2=0
cc_698 N_A_643_369#_c_614_n N_VGND_c_2252_n 0.00919432f $X=4 $Y=0.73 $X2=0 $Y2=0
cc_699 N_A_643_369#_c_620_n N_VGND_c_2252_n 0.0223223f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_700 N_A_643_369#_c_623_n N_VGND_c_2252_n 4.22312e-19 $X=3.91 $Y=1.255 $X2=0
+ $Y2=0
cc_701 N_A_643_369#_c_619_n N_VGND_c_2263_n 0.0125902f $X=3.37 $Y=0.44 $X2=0
+ $Y2=0
cc_702 N_A_643_369#_c_620_n N_VGND_c_2263_n 0.00240298f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_703 N_A_643_369#_c_614_n N_VGND_c_2264_n 0.00427781f $X=4 $Y=0.73 $X2=0 $Y2=0
cc_704 N_A_643_369#_c_615_n N_VGND_c_2264_n 0.00382237f $X=4.865 $Y=0.805 $X2=0
+ $Y2=0
cc_705 N_A_643_369#_c_616_n N_VGND_c_2264_n 0.00564131f $X=4.94 $Y=0.73 $X2=0
+ $Y2=0
cc_706 N_A_643_369#_c_620_n N_VGND_c_2264_n 5.94794e-19 $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_707 N_A_643_369#_M1033_g N_VGND_c_2265_n 0.00362032f $X=9 $Y=0.445 $X2=0
+ $Y2=0
cc_708 N_A_643_369#_c_626_n N_VGND_c_2265_n 0.00429175f $X=8.82 $Y=0.812 $X2=0
+ $Y2=0
cc_709 N_A_643_369#_c_627_n N_VGND_c_2265_n 0.00405482f $X=8.135 $Y=0.812 $X2=0
+ $Y2=0
cc_710 N_A_643_369#_c_627_n N_VGND_c_2272_n 0.00757355f $X=8.135 $Y=0.812 $X2=0
+ $Y2=0
cc_711 N_A_643_369#_M1000_s N_VGND_c_2275_n 0.00323692f $X=3.245 $Y=0.235 $X2=0
+ $Y2=0
cc_712 N_A_643_369#_c_614_n N_VGND_c_2275_n 0.00792209f $X=4 $Y=0.73 $X2=0 $Y2=0
cc_713 N_A_643_369#_c_615_n N_VGND_c_2275_n 0.00372099f $X=4.865 $Y=0.805 $X2=0
+ $Y2=0
cc_714 N_A_643_369#_c_616_n N_VGND_c_2275_n 0.0115324f $X=4.94 $Y=0.73 $X2=0
+ $Y2=0
cc_715 N_A_643_369#_M1033_g N_VGND_c_2275_n 0.00557586f $X=9 $Y=0.445 $X2=0
+ $Y2=0
cc_716 N_A_643_369#_c_619_n N_VGND_c_2275_n 0.00703355f $X=3.37 $Y=0.44 $X2=0
+ $Y2=0
cc_717 N_A_643_369#_c_620_n N_VGND_c_2275_n 0.0062796f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_718 N_A_643_369#_c_626_n N_VGND_c_2275_n 0.00863847f $X=8.82 $Y=0.812 $X2=0
+ $Y2=0
cc_719 N_A_643_369#_c_627_n N_VGND_c_2275_n 0.00706476f $X=8.135 $Y=0.812 $X2=0
+ $Y2=0
cc_720 N_A_643_369#_c_626_n A_1514_47# 0.00233778f $X=8.82 $Y=0.812 $X2=-0.19
+ $Y2=-0.24
cc_721 N_A_643_369#_c_627_n A_1514_47# 0.00819269f $X=8.135 $Y=0.812 $X2=-0.19
+ $Y2=-0.24
cc_722 N_A_809_369#_M1021_g N_A_1129_21#_M1023_g 0.0598207f $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_723 N_A_809_369#_c_902_n N_A_1129_21#_c_1085_n 5.84337e-19 $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_724 N_A_809_369#_c_902_n N_A_1129_21#_c_1079_n 0.00911256f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_725 N_A_809_369#_M1021_g N_A_1129_21#_c_1081_n 4.79914e-19 $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_726 N_A_809_369#_c_902_n N_A_1129_21#_c_1081_n 0.00859525f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_727 N_A_809_369#_c_902_n N_A_1129_21#_c_1082_n 0.00455149f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_728 N_A_809_369#_M1021_g N_A_1129_21#_c_1083_n 0.00652836f $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_729 N_A_809_369#_c_902_n N_A_1129_21#_c_1083_n 0.00266737f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_730 N_A_809_369#_c_899_n N_A_997_413#_c_1176_n 0.0138219f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_731 N_A_809_369#_M1021_g N_A_997_413#_c_1176_n 0.0212478f $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_732 N_A_809_369#_c_902_n N_A_997_413#_c_1176_n 0.0327595f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_733 N_A_809_369#_c_899_n N_A_997_413#_c_1177_n 0.00618953f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_734 N_A_809_369#_c_902_n N_A_997_413#_c_1177_n 0.0242139f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_735 N_A_809_369#_c_907_n N_A_997_413#_c_1177_n 3.67923e-19 $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_736 N_A_809_369#_c_902_n N_A_997_413#_c_1178_n 0.048307f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_737 N_A_809_369#_c_902_n N_A_997_413#_c_1179_n 0.00146532f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_738 N_A_809_369#_c_902_n N_A_997_413#_c_1180_n 0.0174294f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_739 N_A_809_369#_c_902_n N_A_997_413#_c_1181_n 0.0111401f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_740 N_A_809_369#_M1044_g N_SET_B_c_1329_n 0.00175794f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_741 N_A_809_369#_c_912_n N_SET_B_c_1329_n 0.00264635f $X=8.54 $Y=1.905 $X2=0
+ $Y2=0
cc_742 N_A_809_369#_c_902_n N_SET_B_c_1329_n 0.121254f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_743 N_A_809_369#_c_905_n N_SET_B_c_1329_n 0.0256417f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_744 N_A_809_369#_c_906_n N_SET_B_c_1329_n 0.014244f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_745 N_A_809_369#_c_902_n N_SET_B_c_1330_n 0.0264445f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_746 N_A_809_369#_c_912_n N_SET_B_c_1331_n 6.80967e-19 $X=8.54 $Y=1.905 $X2=0
+ $Y2=0
cc_747 N_A_809_369#_c_906_n N_SET_B_c_1331_n 0.00267262f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_748 N_A_809_369#_M1044_g N_SET_B_c_1332_n 3.92661e-19 $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_749 N_A_809_369#_c_912_n N_SET_B_c_1332_n 8.48728e-19 $X=8.54 $Y=1.905 $X2=0
+ $Y2=0
cc_750 N_A_809_369#_c_906_n N_SET_B_c_1332_n 0.0160216f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_751 N_A_809_369#_c_902_n N_SET_B_c_1334_n 9.31754e-19 $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_752 N_A_809_369#_M1034_g N_A_1781_295#_M1006_g 0.0304162f $X=8.54 $Y=2.275
+ $X2=0 $Y2=0
cc_753 N_A_809_369#_c_906_n N_A_1781_295#_M1006_g 0.00103116f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_754 N_A_809_369#_M1044_g N_A_1781_295#_c_1465_n 0.00238845f $X=8.39 $Y=0.555
+ $X2=0 $Y2=0
cc_755 N_A_809_369#_c_912_n N_A_1781_295#_c_1465_n 0.020974f $X=8.54 $Y=1.905
+ $X2=0 $Y2=0
cc_756 N_A_809_369#_c_906_n N_A_1781_295#_c_1465_n 4.76657e-19 $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_757 N_A_809_369#_c_905_n N_A_1781_295#_c_1456_n 9.56757e-19 $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_758 N_A_809_369#_c_906_n N_A_1781_295#_c_1456_n 0.00282361f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_759 N_A_809_369#_c_905_n N_A_1781_295#_c_1468_n 0.00122442f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_760 N_A_809_369#_c_906_n N_A_1781_295#_c_1468_n 0.0024305f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_761 N_A_809_369#_c_912_n N_A_1597_329#_c_1588_n 0.00488486f $X=8.54 $Y=1.905
+ $X2=0 $Y2=0
cc_762 N_A_809_369#_M1034_g N_A_1597_329#_c_1588_n 0.0113397f $X=8.54 $Y=2.275
+ $X2=0 $Y2=0
cc_763 N_A_809_369#_c_906_n N_A_1597_329#_c_1588_n 0.0108833f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_764 N_A_809_369#_M1034_g N_A_1597_329#_c_1580_n 0.00469548f $X=8.54 $Y=2.275
+ $X2=0 $Y2=0
cc_765 N_A_809_369#_c_906_n N_A_1597_329#_c_1580_n 7.30124e-19 $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_766 N_A_809_369#_M1034_g N_VPWR_c_1863_n 0.00358923f $X=8.54 $Y=2.275 $X2=0
+ $Y2=0
cc_767 N_A_809_369#_c_910_n N_VPWR_c_1869_n 0.00585385f $X=4.91 $Y=1.99 $X2=0
+ $Y2=0
cc_768 N_A_809_369#_c_914_n N_VPWR_c_1869_n 0.00216624f $X=4.91 $Y=1.915 $X2=0
+ $Y2=0
cc_769 N_A_809_369#_c_915_n N_VPWR_c_1869_n 0.023872f $X=4.18 $Y=2.3 $X2=0 $Y2=0
cc_770 N_A_809_369#_M1034_g N_VPWR_c_1877_n 0.00159206f $X=8.54 $Y=2.275 $X2=0
+ $Y2=0
cc_771 N_A_809_369#_M1029_d N_VPWR_c_1851_n 0.00210742f $X=4.045 $Y=1.845 $X2=0
+ $Y2=0
cc_772 N_A_809_369#_c_910_n N_VPWR_c_1851_n 0.00769758f $X=4.91 $Y=1.99 $X2=0
+ $Y2=0
cc_773 N_A_809_369#_M1034_g N_VPWR_c_1851_n 0.0057638f $X=8.54 $Y=2.275 $X2=0
+ $Y2=0
cc_774 N_A_809_369#_c_914_n N_VPWR_c_1851_n 0.00143264f $X=4.91 $Y=1.915 $X2=0
+ $Y2=0
cc_775 N_A_809_369#_c_915_n N_VPWR_c_1851_n 0.00624504f $X=4.18 $Y=2.3 $X2=0
+ $Y2=0
cc_776 N_A_809_369#_c_1036_p N_A_181_47#_c_2061_n 0.0256294f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_777 N_A_809_369#_c_909_n N_A_181_47#_c_2066_n 0.00538723f $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_778 N_A_809_369#_c_899_n N_A_181_47#_c_2066_n 0.0014889f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_779 N_A_809_369#_c_914_n N_A_181_47#_c_2066_n 0.00150693f $X=4.91 $Y=1.915
+ $X2=0 $Y2=0
cc_780 N_A_809_369#_c_916_n N_A_181_47#_c_2066_n 0.00936332f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_781 N_A_809_369#_c_902_n N_A_181_47#_c_2066_n 8.95626e-19 $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_782 N_A_809_369#_c_909_n N_A_181_47#_c_2067_n 0.00448337f $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_783 N_A_809_369#_c_910_n N_A_181_47#_c_2067_n 0.0039304f $X=4.91 $Y=1.99
+ $X2=0 $Y2=0
cc_784 N_A_809_369#_c_914_n N_A_181_47#_c_2067_n 0.0125452f $X=4.91 $Y=1.915
+ $X2=0 $Y2=0
cc_785 N_A_809_369#_c_916_n N_A_181_47#_c_2067_n 0.0631002f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_786 N_A_809_369#_c_909_n N_A_181_47#_c_2062_n 6.71081e-19 $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_787 N_A_809_369#_c_899_n N_A_181_47#_c_2062_n 0.00723713f $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_788 N_A_809_369#_c_916_n N_A_181_47#_c_2062_n 0.00124944f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_789 N_A_809_369#_c_902_n N_A_181_47#_c_2062_n 0.0120122f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_790 N_A_809_369#_c_903_n N_A_181_47#_c_2062_n 0.00235599f $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_791 N_A_809_369#_c_904_n N_A_181_47#_c_2062_n 0.0217629f $X=4.37 $Y=1.19
+ $X2=0 $Y2=0
cc_792 N_A_809_369#_c_907_n N_A_181_47#_c_2062_n 0.00624074f $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_793 N_A_809_369#_c_908_n N_A_181_47#_c_2062_n 0.00789495f $X=4.327 $Y=1.09
+ $X2=0 $Y2=0
cc_794 N_A_809_369#_M1021_g N_A_181_47#_c_2064_n 8.04362e-19 $X=5.36 $Y=0.445
+ $X2=0 $Y2=0
cc_795 N_A_809_369#_c_902_n N_A_181_47#_c_2064_n 0.00605448f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_796 N_A_809_369#_c_903_n N_A_181_47#_c_2064_n 5.00901e-19 $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_797 N_A_809_369#_c_907_n N_A_181_47#_c_2064_n 0.00356774f $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_798 N_A_809_369#_c_908_n N_A_181_47#_c_2064_n 0.0256294f $X=4.327 $Y=1.09
+ $X2=0 $Y2=0
cc_799 N_A_809_369#_c_909_n N_A_181_47#_c_2069_n 0.00307634f $X=4.615 $Y=1.84
+ $X2=0 $Y2=0
cc_800 N_A_809_369#_c_916_n N_A_181_47#_c_2069_n 0.0163681f $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_801 N_A_809_369#_c_902_n N_A_181_47#_c_2069_n 0.0135911f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_802 N_A_809_369#_c_903_n N_A_181_47#_c_2069_n 0.0254082f $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_803 N_A_809_369#_c_904_n N_A_181_47#_c_2069_n 0.0014472f $X=4.37 $Y=1.19
+ $X2=0 $Y2=0
cc_804 N_A_809_369#_c_907_n N_A_181_47#_c_2069_n 8.3882e-19 $X=4.69 $Y=1.255
+ $X2=0 $Y2=0
cc_805 N_A_809_369#_c_899_n N_A_181_47#_c_2072_n 4.09059e-19 $X=5.285 $Y=1.165
+ $X2=0 $Y2=0
cc_806 N_A_809_369#_c_914_n N_A_181_47#_c_2072_n 4.12766e-19 $X=4.91 $Y=1.915
+ $X2=0 $Y2=0
cc_807 N_A_809_369#_c_916_n N_A_181_47#_c_2072_n 5.70177e-19 $X=4.267 $Y=2.135
+ $X2=0 $Y2=0
cc_808 N_A_809_369#_c_902_n N_A_181_47#_c_2072_n 0.0264737f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_809 N_A_809_369#_M1021_g N_VGND_c_2264_n 0.00592053f $X=5.36 $Y=0.445 $X2=0
+ $Y2=0
cc_810 N_A_809_369#_c_1036_p N_VGND_c_2264_n 0.0143008f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_811 N_A_809_369#_M1044_g N_VGND_c_2265_n 0.00437171f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_812 N_A_809_369#_M1044_g N_VGND_c_2272_n 0.0148051f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_813 N_A_809_369#_c_902_n N_VGND_c_2272_n 0.00606746f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_814 N_A_809_369#_M1039_d N_VGND_c_2275_n 0.00382094f $X=4.075 $Y=0.235 $X2=0
+ $Y2=0
cc_815 N_A_809_369#_M1021_g N_VGND_c_2275_n 0.00511765f $X=5.36 $Y=0.445 $X2=0
+ $Y2=0
cc_816 N_A_809_369#_M1044_g N_VGND_c_2275_n 0.00784322f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_817 N_A_809_369#_c_1036_p N_VGND_c_2275_n 0.00798371f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_818 N_A_1129_21#_M1040_g N_A_997_413#_M1005_g 0.011154f $X=5.84 $Y=2.275
+ $X2=0 $Y2=0
cc_819 N_A_1129_21#_c_1085_n N_A_997_413#_M1005_g 0.00217932f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_820 N_A_1129_21#_c_1086_n N_A_997_413#_M1005_g 0.0167577f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_821 N_A_1129_21#_c_1087_n N_A_997_413#_M1005_g 0.0130957f $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_822 N_A_1129_21#_c_1083_n N_A_997_413#_M1005_g 0.00524709f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_823 N_A_1129_21#_c_1079_n N_A_997_413#_c_1174_n 0.00169799f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_824 N_A_1129_21#_M1023_g N_A_997_413#_c_1175_n 8.48075e-19 $X=5.72 $Y=0.445
+ $X2=0 $Y2=0
cc_825 N_A_1129_21#_c_1079_n N_A_997_413#_c_1175_n 0.00789989f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_826 N_A_1129_21#_c_1081_n N_A_997_413#_c_1175_n 0.00106627f $X=5.81 $Y=0.72
+ $X2=0 $Y2=0
cc_827 N_A_1129_21#_c_1082_n N_A_997_413#_c_1175_n 0.00775546f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_828 N_A_1129_21#_M1023_g N_A_997_413#_c_1176_n 0.00369174f $X=5.72 $Y=0.445
+ $X2=0 $Y2=0
cc_829 N_A_1129_21#_c_1081_n N_A_997_413#_c_1176_n 0.0259255f $X=5.81 $Y=0.72
+ $X2=0 $Y2=0
cc_830 N_A_1129_21#_c_1083_n N_A_997_413#_c_1176_n 0.00259391f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_831 N_A_1129_21#_c_1085_n N_A_997_413#_c_1187_n 0.0251699f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_832 N_A_1129_21#_c_1088_n N_A_997_413#_c_1187_n 0.010676f $X=6.095 $Y=2.02
+ $X2=0 $Y2=0
cc_833 N_A_1129_21#_c_1083_n N_A_997_413#_c_1187_n 0.0119128f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_834 N_A_1129_21#_c_1081_n N_A_997_413#_c_1177_n 0.00585658f $X=5.81 $Y=0.72
+ $X2=0 $Y2=0
cc_835 N_A_1129_21#_c_1082_n N_A_997_413#_c_1177_n 0.00298561f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_836 N_A_1129_21#_c_1087_n N_A_997_413#_c_1178_n 0.00198283f $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_837 N_A_1129_21#_c_1079_n N_A_997_413#_c_1179_n 0.00227132f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_838 N_A_1129_21#_c_1087_n N_A_997_413#_c_1179_n 6.97279e-19 $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_839 N_A_1129_21#_c_1083_n N_A_997_413#_c_1179_n 0.0114262f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_840 N_A_1129_21#_c_1085_n N_A_997_413#_c_1180_n 0.0109804f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_841 N_A_1129_21#_c_1086_n N_A_997_413#_c_1180_n 0.00260846f $X=6.01 $Y=1.74
+ $X2=0 $Y2=0
cc_842 N_A_1129_21#_c_1079_n N_A_997_413#_c_1180_n 0.00808722f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_843 N_A_1129_21#_c_1087_n N_A_997_413#_c_1180_n 0.00696445f $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_844 N_A_1129_21#_c_1081_n N_A_997_413#_c_1180_n 0.0109475f $X=5.81 $Y=0.72
+ $X2=0 $Y2=0
cc_845 N_A_1129_21#_c_1082_n N_A_997_413#_c_1180_n 7.94205e-19 $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_846 N_A_1129_21#_c_1083_n N_A_997_413#_c_1180_n 0.0129003f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_847 N_A_1129_21#_c_1079_n N_A_997_413#_c_1181_n 0.0178097f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_848 N_A_1129_21#_c_1081_n N_A_997_413#_c_1181_n 0.00200868f $X=5.81 $Y=0.72
+ $X2=0 $Y2=0
cc_849 N_A_1129_21#_c_1082_n N_A_997_413#_c_1181_n 0.00156611f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_850 N_A_1129_21#_c_1083_n N_A_997_413#_c_1181_n 0.00171161f $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_851 N_A_1129_21#_c_1083_n N_A_997_413#_c_1183_n 5.49747e-19 $X=5.955 $Y=1.575
+ $X2=0 $Y2=0
cc_852 N_A_1129_21#_c_1087_n N_SET_B_M1030_g 0.00493354f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_853 N_A_1129_21#_c_1085_n N_SET_B_c_1330_n 0.00168184f $X=6.01 $Y=1.74 $X2=0
+ $Y2=0
cc_854 N_A_1129_21#_c_1087_n N_SET_B_c_1330_n 3.32046e-19 $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_855 N_A_1129_21#_c_1087_n N_SET_B_c_1333_n 0.00107555f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_856 N_A_1129_21#_c_1085_n N_SET_B_c_1334_n 0.00504977f $X=6.01 $Y=1.74 $X2=0
+ $Y2=0
cc_857 N_A_1129_21#_c_1087_n N_SET_B_c_1334_n 0.0122653f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_858 N_A_1129_21#_c_1087_n N_VPWR_M1040_d 0.00281587f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_859 N_A_1129_21#_c_1088_n N_VPWR_M1040_d 0.00142005f $X=6.095 $Y=2.02 $X2=0
+ $Y2=0
cc_860 N_A_1129_21#_M1040_g N_VPWR_c_1869_n 0.00585385f $X=5.84 $Y=2.275 $X2=0
+ $Y2=0
cc_861 N_A_1129_21#_M1040_g N_VPWR_c_1875_n 0.00335682f $X=5.84 $Y=2.275 $X2=0
+ $Y2=0
cc_862 N_A_1129_21#_c_1086_n N_VPWR_c_1875_n 7.77116e-19 $X=6.01 $Y=1.74 $X2=0
+ $Y2=0
cc_863 N_A_1129_21#_c_1087_n N_VPWR_c_1875_n 0.0164669f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_864 N_A_1129_21#_c_1088_n N_VPWR_c_1875_n 0.00947355f $X=6.095 $Y=2.02 $X2=0
+ $Y2=0
cc_865 N_A_1129_21#_c_1087_n N_VPWR_c_1876_n 0.00399899f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_866 N_A_1129_21#_c_1154_p N_VPWR_c_1876_n 0.0132089f $X=6.715 $Y=2.285 $X2=0
+ $Y2=0
cc_867 N_A_1129_21#_M1005_d N_VPWR_c_1851_n 0.00275725f $X=6.555 $Y=2.065 $X2=0
+ $Y2=0
cc_868 N_A_1129_21#_M1040_g N_VPWR_c_1851_n 0.00693532f $X=5.84 $Y=2.275 $X2=0
+ $Y2=0
cc_869 N_A_1129_21#_c_1087_n N_VPWR_c_1851_n 0.00374474f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_870 N_A_1129_21#_c_1088_n N_VPWR_c_1851_n 7.82982e-19 $X=6.095 $Y=2.02 $X2=0
+ $Y2=0
cc_871 N_A_1129_21#_c_1154_p N_VPWR_c_1851_n 0.00381852f $X=6.715 $Y=2.285 $X2=0
+ $Y2=0
cc_872 N_A_1129_21#_c_1079_n N_VGND_M1023_d 8.64202e-19 $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_873 N_A_1129_21#_c_1081_n N_VGND_M1023_d 0.00132848f $X=5.81 $Y=0.72 $X2=0
+ $Y2=0
cc_874 N_A_1129_21#_M1023_g N_VGND_c_2264_n 0.013328f $X=5.72 $Y=0.445 $X2=0
+ $Y2=0
cc_875 N_A_1129_21#_c_1079_n N_VGND_c_2264_n 0.00919218f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_876 N_A_1129_21#_c_1080_n N_VGND_c_2264_n 0.0163221f $X=6.45 $Y=0.51 $X2=0
+ $Y2=0
cc_877 N_A_1129_21#_c_1081_n N_VGND_c_2264_n 0.021134f $X=5.81 $Y=0.72 $X2=0
+ $Y2=0
cc_878 N_A_1129_21#_c_1082_n N_VGND_c_2264_n 8.18098e-19 $X=5.81 $Y=0.93 $X2=0
+ $Y2=0
cc_879 N_A_1129_21#_c_1079_n N_VGND_c_2271_n 0.00346394f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_880 N_A_1129_21#_c_1080_n N_VGND_c_2271_n 0.0170207f $X=6.45 $Y=0.51 $X2=0
+ $Y2=0
cc_881 N_A_1129_21#_c_1079_n N_VGND_c_2272_n 0.0135163f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_882 N_A_1129_21#_M1008_s N_VGND_c_2275_n 0.00268769f $X=6.325 $Y=0.235 $X2=0
+ $Y2=0
cc_883 N_A_1129_21#_c_1079_n N_VGND_c_2275_n 0.00594673f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_884 N_A_1129_21#_c_1080_n N_VGND_c_2275_n 0.00949852f $X=6.45 $Y=0.51 $X2=0
+ $Y2=0
cc_885 N_A_1129_21#_c_1081_n N_VGND_c_2275_n 0.00150511f $X=5.81 $Y=0.72 $X2=0
+ $Y2=0
cc_886 N_A_997_413#_M1005_g N_SET_B_M1030_g 0.0138848f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_887 N_A_997_413#_c_1174_n N_SET_B_M1043_g 0.0503064f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_888 N_A_997_413#_c_1178_n N_SET_B_M1043_g 0.0112575f $X=7.355 $Y=1.125 $X2=0
+ $Y2=0
cc_889 N_A_997_413#_c_1182_n N_SET_B_M1043_g 0.0213587f $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_890 N_A_997_413#_c_1183_n N_SET_B_M1043_g 0.0104446f $X=6.39 $Y=1.095 $X2=0
+ $Y2=0
cc_891 N_A_997_413#_c_1184_n N_SET_B_M1043_g 0.0223803f $X=7.465 $Y=0.995 $X2=0
+ $Y2=0
cc_892 N_A_997_413#_M1011_g N_SET_B_c_1321_n 0.00155652f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_893 N_A_997_413#_c_1178_n N_SET_B_c_1321_n 0.0063144f $X=7.355 $Y=1.125 $X2=0
+ $Y2=0
cc_894 N_A_997_413#_c_1179_n N_SET_B_c_1321_n 0.00545541f $X=6.39 $Y=1.23 $X2=0
+ $Y2=0
cc_895 N_A_997_413#_c_1181_n N_SET_B_c_1321_n 6.1772e-19 $X=6.475 $Y=1.185 $X2=0
+ $Y2=0
cc_896 N_A_997_413#_M1011_g N_SET_B_c_1329_n 0.00453798f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_897 N_A_997_413#_c_1178_n N_SET_B_c_1329_n 0.00989598f $X=7.355 $Y=1.125
+ $X2=0 $Y2=0
cc_898 N_A_997_413#_c_1182_n N_SET_B_c_1329_n 7.77586e-19 $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_899 N_A_997_413#_M1005_g N_SET_B_c_1330_n 0.00451637f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_900 N_A_997_413#_c_1178_n N_SET_B_c_1330_n 0.00232629f $X=7.355 $Y=1.125
+ $X2=0 $Y2=0
cc_901 N_A_997_413#_M1005_g N_SET_B_c_1333_n 0.0200627f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_902 N_A_997_413#_c_1178_n N_SET_B_c_1333_n 7.95701e-19 $X=7.355 $Y=1.125
+ $X2=0 $Y2=0
cc_903 N_A_997_413#_M1005_g N_SET_B_c_1334_n 0.00489625f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_904 N_A_997_413#_M1011_g N_SET_B_c_1334_n 0.00360395f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_905 N_A_997_413#_c_1178_n N_SET_B_c_1334_n 0.0278918f $X=7.355 $Y=1.125 $X2=0
+ $Y2=0
cc_906 N_A_997_413#_M1005_g N_SET_B_c_1335_n 0.00545541f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_907 N_A_997_413#_M1011_g N_SET_B_c_1335_n 0.0293466f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_908 N_A_997_413#_c_1201_n N_VPWR_c_1869_n 0.042644f $X=5.585 $Y=2.3 $X2=0
+ $Y2=0
cc_909 N_A_997_413#_M1005_g N_VPWR_c_1875_n 0.00604582f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_910 N_A_997_413#_M1005_g N_VPWR_c_1876_n 0.00422112f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_911 N_A_997_413#_M1011_g N_VPWR_c_1877_n 0.0234385f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_912 N_A_997_413#_M1007_d N_VPWR_c_1851_n 0.00212626f $X=4.985 $Y=2.065 $X2=0
+ $Y2=0
cc_913 N_A_997_413#_M1005_g N_VPWR_c_1851_n 0.00619761f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_914 N_A_997_413#_c_1201_n N_VPWR_c_1851_n 0.0122201f $X=5.585 $Y=2.3 $X2=0
+ $Y2=0
cc_915 N_A_997_413#_c_1176_n N_A_181_47#_c_2061_n 0.0591375f $X=5.15 $Y=0.42
+ $X2=0 $Y2=0
cc_916 N_A_997_413#_c_1187_n N_A_181_47#_c_2066_n 0.00197049f $X=5.67 $Y=2.135
+ $X2=0 $Y2=0
cc_917 N_A_997_413#_c_1177_n N_A_181_47#_c_2062_n 0.0111326f $X=5.755 $Y=1.31
+ $X2=0 $Y2=0
cc_918 N_A_997_413#_c_1187_n N_A_181_47#_c_2072_n 0.00424021f $X=5.67 $Y=2.135
+ $X2=0 $Y2=0
cc_919 N_A_997_413#_c_1201_n A_1081_413# 0.0063224f $X=5.585 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_920 N_A_997_413#_c_1187_n A_1081_413# 0.0012628f $X=5.67 $Y=2.135 $X2=-0.19
+ $Y2=-0.24
cc_921 N_A_997_413#_c_1174_n N_VGND_c_2264_n 0.00201299f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_922 N_A_997_413#_c_1176_n N_VGND_c_2264_n 0.0262729f $X=5.15 $Y=0.42 $X2=0
+ $Y2=0
cc_923 N_A_997_413#_c_1174_n N_VGND_c_2271_n 0.0046653f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_924 N_A_997_413#_c_1175_n N_VGND_c_2271_n 0.00120334f $X=6.66 $Y=0.805 $X2=0
+ $Y2=0
cc_925 N_A_997_413#_c_1174_n N_VGND_c_2272_n 0.0137178f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_926 N_A_997_413#_c_1175_n N_VGND_c_2272_n 0.00215939f $X=6.66 $Y=0.805 $X2=0
+ $Y2=0
cc_927 N_A_997_413#_c_1178_n N_VGND_c_2272_n 0.0750884f $X=7.355 $Y=1.125 $X2=0
+ $Y2=0
cc_928 N_A_997_413#_c_1182_n N_VGND_c_2272_n 7.09663e-19 $X=7.44 $Y=1.16 $X2=0
+ $Y2=0
cc_929 N_A_997_413#_c_1184_n N_VGND_c_2272_n 0.0317395f $X=7.465 $Y=0.995 $X2=0
+ $Y2=0
cc_930 N_A_997_413#_M1020_d N_VGND_c_2275_n 0.00215201f $X=5.015 $Y=0.235 $X2=0
+ $Y2=0
cc_931 N_A_997_413#_c_1174_n N_VGND_c_2275_n 0.00929621f $X=6.66 $Y=0.73 $X2=0
+ $Y2=0
cc_932 N_A_997_413#_c_1175_n N_VGND_c_2275_n 0.00120242f $X=6.66 $Y=0.805 $X2=0
+ $Y2=0
cc_933 N_A_997_413#_c_1176_n N_VGND_c_2275_n 0.0159733f $X=5.15 $Y=0.42 $X2=0
+ $Y2=0
cc_934 N_SET_B_c_1325_n N_A_1781_295#_M1006_g 0.014668f $X=9.715 $Y=1.985 $X2=0
+ $Y2=0
cc_935 N_SET_B_c_1327_n N_A_1781_295#_M1006_g 2.95112e-19 $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_936 N_SET_B_c_1328_n N_A_1781_295#_M1006_g 0.00434236f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_937 N_SET_B_c_1332_n N_A_1781_295#_M1006_g 0.0047394f $X=9.025 $Y=1.53 $X2=0
+ $Y2=0
cc_938 N_SET_B_c_1327_n N_A_1781_295#_c_1464_n 0.0159041f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_939 N_SET_B_c_1328_n N_A_1781_295#_c_1464_n 0.005442f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_940 N_SET_B_c_1331_n N_A_1781_295#_c_1464_n 0.00168581f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_941 N_SET_B_c_1332_n N_A_1781_295#_c_1464_n 0.00484506f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_942 N_SET_B_c_1332_n N_A_1781_295#_c_1465_n 0.00336779f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_943 N_SET_B_M1042_g N_A_1781_295#_M1035_g 0.027178f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_944 N_SET_B_M1042_g N_A_1781_295#_c_1456_n 0.0106852f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_945 N_SET_B_c_1326_n N_A_1781_295#_c_1456_n 0.005442f $X=9.78 $Y=1.6 $X2=0
+ $Y2=0
cc_946 N_SET_B_c_1331_n N_A_1781_295#_c_1456_n 0.00153181f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_947 N_SET_B_c_1332_n N_A_1781_295#_c_1456_n 0.00158925f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_948 N_SET_B_M1042_g N_A_1781_295#_c_1457_n 0.00143395f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_949 N_SET_B_M1042_g N_A_1781_295#_c_1458_n 0.0205597f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_950 N_SET_B_c_1325_n N_A_1781_295#_c_1458_n 4.53409e-19 $X=9.715 $Y=1.985
+ $X2=0 $Y2=0
cc_951 N_SET_B_c_1327_n N_A_1781_295#_c_1458_n 4.53365e-19 $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_952 N_SET_B_M1042_g N_A_1781_295#_c_1459_n 0.0109095f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_953 N_SET_B_c_1326_n N_A_1781_295#_c_1459_n 0.00326242f $X=9.78 $Y=1.6 $X2=0
+ $Y2=0
cc_954 N_SET_B_c_1327_n N_A_1781_295#_c_1459_n 0.028507f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_955 N_SET_B_c_1327_n N_A_1781_295#_c_1468_n 0.0157183f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_956 N_SET_B_c_1328_n N_A_1597_329#_M1015_g 0.0026354f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_957 N_SET_B_M1042_g N_A_1597_329#_c_1564_n 0.0177927f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_958 N_SET_B_M1042_g N_A_1597_329#_c_1565_n 0.0130002f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_959 N_SET_B_c_1326_n N_A_1597_329#_c_1566_n 0.0177927f $X=9.78 $Y=1.6 $X2=0
+ $Y2=0
cc_960 N_SET_B_c_1329_n N_A_1597_329#_c_1588_n 0.0147002f $X=8.88 $Y=1.53 $X2=0
+ $Y2=0
cc_961 N_SET_B_M1042_g N_A_1597_329#_c_1589_n 0.010118f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_962 N_SET_B_c_1325_n N_A_1597_329#_c_1577_n 0.00952217f $X=9.715 $Y=1.985
+ $X2=0 $Y2=0
cc_963 N_SET_B_c_1327_n N_A_1597_329#_c_1577_n 0.038857f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_964 N_SET_B_c_1331_n N_A_1597_329#_c_1577_n 0.00107674f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_965 N_SET_B_c_1332_n N_A_1597_329#_c_1577_n 0.0100658f $X=9.025 $Y=1.53 $X2=0
+ $Y2=0
cc_966 N_SET_B_c_1325_n N_A_1597_329#_c_1578_n 0.0056593f $X=9.715 $Y=1.985
+ $X2=0 $Y2=0
cc_967 N_SET_B_M1042_g N_A_1597_329#_c_1568_n 0.00810025f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_968 N_SET_B_M1042_g N_A_1597_329#_c_1569_n 0.00619235f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_969 N_SET_B_M1042_g N_A_1597_329#_c_1570_n 0.00290265f $X=9.84 $Y=0.445 $X2=0
+ $Y2=0
cc_970 N_SET_B_c_1325_n N_A_1597_329#_c_1580_n 4.4972e-19 $X=9.715 $Y=1.985
+ $X2=0 $Y2=0
cc_971 N_SET_B_c_1329_n N_A_1597_329#_c_1580_n 0.00169667f $X=8.88 $Y=1.53 $X2=0
+ $Y2=0
cc_972 N_SET_B_c_1331_n N_A_1597_329#_c_1580_n 6.9852e-19 $X=9.025 $Y=1.53 $X2=0
+ $Y2=0
cc_973 N_SET_B_c_1332_n N_A_1597_329#_c_1580_n 0.00798024f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_974 N_SET_B_c_1325_n N_A_1597_329#_c_1581_n 0.0143973f $X=9.715 $Y=1.985
+ $X2=0 $Y2=0
cc_975 N_SET_B_c_1327_n N_A_1597_329#_c_1581_n 0.0216774f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_976 N_SET_B_c_1325_n N_A_1597_329#_c_1582_n 2.01999e-19 $X=9.715 $Y=1.985
+ $X2=0 $Y2=0
cc_977 N_SET_B_c_1327_n N_A_1597_329#_c_1582_n 0.00856603f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_978 N_SET_B_c_1328_n N_A_1597_329#_c_1582_n 0.00258524f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_979 N_SET_B_c_1326_n N_A_1597_329#_c_1583_n 0.0151566f $X=9.78 $Y=1.6 $X2=0
+ $Y2=0
cc_980 N_SET_B_c_1327_n N_A_1597_329#_c_1583_n 0.00215089f $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_981 N_SET_B_c_1327_n N_A_1597_329#_c_1584_n 2.24875e-19 $X=9.78 $Y=1.63 $X2=0
+ $Y2=0
cc_982 N_SET_B_c_1325_n N_VPWR_c_1855_n 0.00193129f $X=9.715 $Y=1.985 $X2=0
+ $Y2=0
cc_983 N_SET_B_c_1325_n N_VPWR_c_1856_n 0.00155122f $X=9.715 $Y=1.985 $X2=0
+ $Y2=0
cc_984 N_SET_B_c_1325_n N_VPWR_c_1870_n 0.00484982f $X=9.715 $Y=1.985 $X2=0
+ $Y2=0
cc_985 N_SET_B_M1030_g N_VPWR_c_1876_n 0.00585385f $X=6.97 $Y=2.275 $X2=0 $Y2=0
cc_986 N_SET_B_M1030_g N_VPWR_c_1877_n 0.00385005f $X=6.97 $Y=2.275 $X2=0 $Y2=0
cc_987 N_SET_B_c_1329_n N_VPWR_c_1877_n 9.98887e-19 $X=8.88 $Y=1.53 $X2=0 $Y2=0
cc_988 N_SET_B_M1030_g N_VPWR_c_1851_n 0.00672875f $X=6.97 $Y=2.275 $X2=0 $Y2=0
cc_989 N_SET_B_c_1325_n N_VPWR_c_1851_n 0.00743094f $X=9.715 $Y=1.985 $X2=0
+ $Y2=0
cc_990 N_SET_B_c_1333_n N_VPWR_c_1851_n 4.0446e-19 $X=6.9 $Y=1.68 $X2=0 $Y2=0
cc_991 N_SET_B_M1042_g N_VGND_c_2253_n 0.00503921f $X=9.84 $Y=0.445 $X2=0 $Y2=0
cc_992 N_SET_B_M1042_g N_VGND_c_2265_n 0.00369278f $X=9.84 $Y=0.445 $X2=0 $Y2=0
cc_993 N_SET_B_M1043_g N_VGND_c_2272_n 0.0259455f $X=7.02 $Y=0.445 $X2=0 $Y2=0
cc_994 N_SET_B_c_1321_n N_VGND_c_2272_n 2.2914e-19 $X=6.995 $Y=1.365 $X2=0 $Y2=0
cc_995 N_SET_B_M1042_g N_VGND_c_2275_n 0.00584149f $X=9.84 $Y=0.445 $X2=0 $Y2=0
cc_996 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1562_n 0.00134819f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_997 N_A_1781_295#_c_1462_n N_A_1597_329#_c_1562_n 0.0170978f $X=10.785
+ $Y=1.28 $X2=0 $Y2=0
cc_998 N_A_1781_295#_c_1460_n N_A_1597_329#_M1009_g 7.3983e-19 $X=10.8 $Y=1.195
+ $X2=0 $Y2=0
cc_999 N_A_1781_295#_c_1461_n N_A_1597_329#_M1009_g 0.00103278f $X=10.74 $Y=0.42
+ $X2=0 $Y2=0
cc_1000 N_A_1781_295#_c_1460_n N_A_1597_329#_c_1564_n 0.0015106f $X=10.8
+ $Y=1.195 $X2=0 $Y2=0
cc_1001 N_A_1781_295#_c_1460_n N_A_1597_329#_c_1565_n 0.00692101f $X=10.8
+ $Y=1.195 $X2=0 $Y2=0
cc_1002 N_A_1781_295#_c_1461_n N_A_1597_329#_c_1565_n 0.00753262f $X=10.74
+ $Y=0.42 $X2=0 $Y2=0
cc_1003 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1566_n 0.00781309f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1004 N_A_1781_295#_c_1461_n N_A_1597_329#_c_1566_n 6.04442e-19 $X=10.74
+ $Y=0.42 $X2=0 $Y2=0
cc_1005 N_A_1781_295#_M1006_g N_A_1597_329#_c_1588_n 5.40489e-19 $X=8.98
+ $Y=2.275 $X2=0 $Y2=0
cc_1006 N_A_1781_295#_M1035_g N_A_1597_329#_c_1589_n 0.0150662f $X=9.36 $Y=0.445
+ $X2=0 $Y2=0
cc_1007 N_A_1781_295#_c_1457_n N_A_1597_329#_c_1589_n 0.00772929f $X=9.42
+ $Y=1.02 $X2=0 $Y2=0
cc_1008 N_A_1781_295#_c_1458_n N_A_1597_329#_c_1589_n 0.00105093f $X=9.42
+ $Y=1.02 $X2=0 $Y2=0
cc_1009 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1589_n 0.00516419f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1010 N_A_1781_295#_M1006_g N_A_1597_329#_c_1577_n 0.00670763f $X=8.98
+ $Y=2.275 $X2=0 $Y2=0
cc_1011 N_A_1781_295#_c_1464_n N_A_1597_329#_c_1577_n 0.00206452f $X=9.285
+ $Y=1.55 $X2=0 $Y2=0
cc_1012 N_A_1781_295#_M1006_g N_A_1597_329#_c_1578_n 5.4779e-19 $X=8.98 $Y=2.275
+ $X2=0 $Y2=0
cc_1013 N_A_1781_295#_M1035_g N_A_1597_329#_c_1568_n 0.00215102f $X=9.36
+ $Y=0.445 $X2=0 $Y2=0
cc_1014 N_A_1781_295#_c_1461_n N_A_1597_329#_c_1568_n 0.00100359f $X=10.74
+ $Y=0.42 $X2=0 $Y2=0
cc_1015 N_A_1781_295#_M1035_g N_A_1597_329#_c_1569_n 7.49727e-19 $X=9.36
+ $Y=0.445 $X2=0 $Y2=0
cc_1016 N_A_1781_295#_c_1457_n N_A_1597_329#_c_1569_n 0.0125386f $X=9.42 $Y=1.02
+ $X2=0 $Y2=0
cc_1017 N_A_1781_295#_c_1458_n N_A_1597_329#_c_1569_n 0.00101557f $X=9.42
+ $Y=1.02 $X2=0 $Y2=0
cc_1018 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1569_n 0.0150084f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1019 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1570_n 0.0426229f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1020 N_A_1781_295#_c_1460_n N_A_1597_329#_c_1570_n 0.0196589f $X=10.8
+ $Y=1.195 $X2=0 $Y2=0
cc_1021 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1571_n 0.00428401f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1022 N_A_1781_295#_c_1460_n N_A_1597_329#_c_1571_n 0.00662579f $X=10.8
+ $Y=1.195 $X2=0 $Y2=0
cc_1023 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1579_n 0.00649166f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1024 N_A_1781_295#_M1006_g N_A_1597_329#_c_1580_n 0.0144696f $X=8.98 $Y=2.275
+ $X2=0 $Y2=0
cc_1025 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1581_n 7.5421e-19 $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1026 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1582_n 0.0185636f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1027 N_A_1781_295#_c_1469_n N_A_1597_329#_c_1582_n 0.0356427f $X=10.74
+ $Y=2.285 $X2=0 $Y2=0
cc_1028 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1583_n 0.00132138f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1029 N_A_1781_295#_c_1459_n N_A_1597_329#_c_1584_n 0.0103214f $X=10.655
+ $Y=1.28 $X2=0 $Y2=0
cc_1030 N_A_1781_295#_c_1469_n N_A_1597_329#_c_1584_n 0.0229243f $X=10.74
+ $Y=2.285 $X2=0 $Y2=0
cc_1031 N_A_1781_295#_c_1461_n N_A_2227_47#_c_1721_n 0.0596011f $X=10.74 $Y=0.42
+ $X2=0 $Y2=0
cc_1032 N_A_1781_295#_c_1469_n N_A_2227_47#_c_1729_n 0.0883079f $X=10.74
+ $Y=2.285 $X2=0 $Y2=0
cc_1033 N_A_1781_295#_c_1462_n N_A_2227_47#_c_1729_n 0.0031876f $X=10.785
+ $Y=1.28 $X2=0 $Y2=0
cc_1034 N_A_1781_295#_c_1460_n N_A_2227_47#_c_1723_n 0.0172076f $X=10.8 $Y=1.195
+ $X2=0 $Y2=0
cc_1035 N_A_1781_295#_c_1462_n N_A_2227_47#_c_1723_n 0.0110951f $X=10.785
+ $Y=1.28 $X2=0 $Y2=0
cc_1036 N_A_1781_295#_M1006_g N_VPWR_c_1855_n 0.00540847f $X=8.98 $Y=2.275 $X2=0
+ $Y2=0
cc_1037 N_A_1781_295#_M1006_g N_VPWR_c_1863_n 0.00390259f $X=8.98 $Y=2.275 $X2=0
+ $Y2=0
cc_1038 N_A_1781_295#_c_1469_n N_VPWR_c_1871_n 0.018001f $X=10.74 $Y=2.285 $X2=0
+ $Y2=0
cc_1039 N_A_1781_295#_M1015_d N_VPWR_c_1851_n 0.00382897f $X=10.605 $Y=2.065
+ $X2=0 $Y2=0
cc_1040 N_A_1781_295#_M1006_g N_VPWR_c_1851_n 0.00606164f $X=8.98 $Y=2.275 $X2=0
+ $Y2=0
cc_1041 N_A_1781_295#_c_1469_n N_VPWR_c_1851_n 0.00993603f $X=10.74 $Y=2.285
+ $X2=0 $Y2=0
cc_1042 N_A_1781_295#_c_1461_n N_VGND_c_2253_n 0.0187962f $X=10.74 $Y=0.42 $X2=0
+ $Y2=0
cc_1043 N_A_1781_295#_M1035_g N_VGND_c_2265_n 0.00362032f $X=9.36 $Y=0.445 $X2=0
+ $Y2=0
cc_1044 N_A_1781_295#_c_1461_n N_VGND_c_2266_n 0.0234496f $X=10.74 $Y=0.42 $X2=0
+ $Y2=0
cc_1045 N_A_1781_295#_M1010_d N_VGND_c_2275_n 0.00537869f $X=10.485 $Y=0.235
+ $X2=0 $Y2=0
cc_1046 N_A_1781_295#_M1035_g N_VGND_c_2275_n 0.0053092f $X=9.36 $Y=0.445 $X2=0
+ $Y2=0
cc_1047 N_A_1781_295#_c_1461_n N_VGND_c_2275_n 0.0129422f $X=10.74 $Y=0.42 $X2=0
+ $Y2=0
cc_1048 N_A_1597_329#_M1009_g N_A_2227_47#_c_1717_n 0.00910136f $X=11.47 $Y=0.56
+ $X2=0 $Y2=0
cc_1049 N_A_1597_329#_c_1567_n N_A_2227_47#_M1003_g 0.0110183f $X=11.47 $Y=1.28
+ $X2=0 $Y2=0
cc_1050 N_A_1597_329#_M1009_g N_A_2227_47#_c_1721_n 0.0095769f $X=11.47 $Y=0.56
+ $X2=0 $Y2=0
cc_1051 N_A_1597_329#_c_1562_n N_A_2227_47#_c_1729_n 0.00689943f $X=11.395
+ $Y=1.28 $X2=0 $Y2=0
cc_1052 N_A_1597_329#_M1016_g N_A_2227_47#_c_1729_n 0.0105932f $X=11.47 $Y=1.985
+ $X2=0 $Y2=0
cc_1053 N_A_1597_329#_c_1584_n N_A_2227_47#_c_1729_n 0.00154523f $X=10.38
+ $Y=1.555 $X2=0 $Y2=0
cc_1054 N_A_1597_329#_c_1562_n N_A_2227_47#_c_1722_n 0.00283006f $X=11.395
+ $Y=1.28 $X2=0 $Y2=0
cc_1055 N_A_1597_329#_M1009_g N_A_2227_47#_c_1722_n 0.0152048f $X=11.47 $Y=0.56
+ $X2=0 $Y2=0
cc_1056 N_A_1597_329#_c_1567_n N_A_2227_47#_c_1722_n 0.00895869f $X=11.47
+ $Y=1.28 $X2=0 $Y2=0
cc_1057 N_A_1597_329#_c_1562_n N_A_2227_47#_c_1723_n 0.009972f $X=11.395 $Y=1.28
+ $X2=0 $Y2=0
cc_1058 N_A_1597_329#_c_1571_n N_A_2227_47#_c_1723_n 2.95153e-19 $X=10.35
+ $Y=0.93 $X2=0 $Y2=0
cc_1059 N_A_1597_329#_M1009_g N_A_2227_47#_c_1724_n 0.021471f $X=11.47 $Y=0.56
+ $X2=0 $Y2=0
cc_1060 N_A_1597_329#_c_1582_n N_VPWR_M1015_s 0.00274492f $X=10.32 $Y=1.69 $X2=0
+ $Y2=0
cc_1061 N_A_1597_329#_c_1577_n N_VPWR_c_1855_n 0.0242002f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1062 N_A_1597_329#_c_1580_n N_VPWR_c_1855_n 0.0166484f $X=8.905 $Y=1.98 $X2=0
+ $Y2=0
cc_1063 N_A_1597_329#_M1015_g N_VPWR_c_1856_n 0.00966829f $X=10.53 $Y=2.275
+ $X2=0 $Y2=0
cc_1064 N_A_1597_329#_c_1578_n N_VPWR_c_1856_n 0.0164574f $X=9.8 $Y=2.285 $X2=0
+ $Y2=0
cc_1065 N_A_1597_329#_c_1582_n N_VPWR_c_1856_n 0.0244903f $X=10.32 $Y=1.69 $X2=0
+ $Y2=0
cc_1066 N_A_1597_329#_c_1583_n N_VPWR_c_1856_n 0.00123619f $X=10.32 $Y=1.69
+ $X2=0 $Y2=0
cc_1067 N_A_1597_329#_M1016_g N_VPWR_c_1857_n 0.0167405f $X=11.47 $Y=1.985 $X2=0
+ $Y2=0
cc_1068 N_A_1597_329#_c_1588_n N_VPWR_c_1863_n 0.0371085f $X=8.82 $Y=2.292 $X2=0
+ $Y2=0
cc_1069 N_A_1597_329#_c_1577_n N_VPWR_c_1863_n 0.00284657f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1070 N_A_1597_329#_c_1580_n N_VPWR_c_1863_n 0.00925064f $X=8.905 $Y=1.98
+ $X2=0 $Y2=0
cc_1071 N_A_1597_329#_c_1577_n N_VPWR_c_1870_n 0.00268845f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1072 N_A_1597_329#_c_1578_n N_VPWR_c_1870_n 0.0174202f $X=9.8 $Y=2.285 $X2=0
+ $Y2=0
cc_1073 N_A_1597_329#_c_1579_n N_VPWR_c_1870_n 0.00331215f $X=10.155 $Y=1.98
+ $X2=0 $Y2=0
cc_1074 N_A_1597_329#_M1015_g N_VPWR_c_1871_n 0.0046653f $X=10.53 $Y=2.275 $X2=0
+ $Y2=0
cc_1075 N_A_1597_329#_M1016_g N_VPWR_c_1871_n 0.0046653f $X=11.47 $Y=1.985 $X2=0
+ $Y2=0
cc_1076 N_A_1597_329#_M1017_d N_VPWR_c_1851_n 0.00601652f $X=7.985 $Y=1.645
+ $X2=0 $Y2=0
cc_1077 N_A_1597_329#_M1025_d N_VPWR_c_1851_n 0.00209863f $X=9.665 $Y=2.065
+ $X2=0 $Y2=0
cc_1078 N_A_1597_329#_M1015_g N_VPWR_c_1851_n 0.00929867f $X=10.53 $Y=2.275
+ $X2=0 $Y2=0
cc_1079 N_A_1597_329#_M1016_g N_VPWR_c_1851_n 0.00921786f $X=11.47 $Y=1.985
+ $X2=0 $Y2=0
cc_1080 N_A_1597_329#_c_1588_n N_VPWR_c_1851_n 0.0231897f $X=8.82 $Y=2.292 $X2=0
+ $Y2=0
cc_1081 N_A_1597_329#_c_1577_n N_VPWR_c_1851_n 0.00983239f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1082 N_A_1597_329#_c_1578_n N_VPWR_c_1851_n 0.0114315f $X=9.8 $Y=2.285 $X2=0
+ $Y2=0
cc_1083 N_A_1597_329#_c_1579_n N_VPWR_c_1851_n 0.00529433f $X=10.155 $Y=1.98
+ $X2=0 $Y2=0
cc_1084 N_A_1597_329#_c_1580_n N_VPWR_c_1851_n 0.00603799f $X=8.905 $Y=1.98
+ $X2=0 $Y2=0
cc_1085 N_A_1597_329#_c_1582_n N_VPWR_c_1851_n 0.00152519f $X=10.32 $Y=1.69
+ $X2=0 $Y2=0
cc_1086 N_A_1597_329#_c_1588_n A_1723_413# 0.00493444f $X=8.82 $Y=2.292
+ $X2=-0.19 $Y2=-0.24
cc_1087 N_A_1597_329#_c_1580_n A_1723_413# 0.00180472f $X=8.905 $Y=1.98
+ $X2=-0.19 $Y2=-0.24
cc_1088 N_A_1597_329#_c_1564_n N_VGND_c_2253_n 0.00298286f $X=10.35 $Y=0.9 $X2=0
+ $Y2=0
cc_1089 N_A_1597_329#_c_1565_n N_VGND_c_2253_n 0.00962162f $X=10.35 $Y=0.765
+ $X2=0 $Y2=0
cc_1090 N_A_1597_329#_c_1589_n N_VGND_c_2253_n 0.0188589f $X=9.71 $Y=0.41 $X2=0
+ $Y2=0
cc_1091 N_A_1597_329#_c_1570_n N_VGND_c_2253_n 0.0126026f $X=10.35 $Y=0.93 $X2=0
+ $Y2=0
cc_1092 N_A_1597_329#_M1009_g N_VGND_c_2254_n 0.0123425f $X=11.47 $Y=0.56 $X2=0
+ $Y2=0
cc_1093 N_A_1597_329#_c_1589_n N_VGND_c_2265_n 0.0745808f $X=9.71 $Y=0.41 $X2=0
+ $Y2=0
cc_1094 N_A_1597_329#_M1009_g N_VGND_c_2266_n 0.0046653f $X=11.47 $Y=0.56 $X2=0
+ $Y2=0
cc_1095 N_A_1597_329#_c_1565_n N_VGND_c_2266_n 0.0046653f $X=10.35 $Y=0.765
+ $X2=0 $Y2=0
cc_1096 N_A_1597_329#_M1044_d N_VGND_c_2275_n 0.00371781f $X=8.465 $Y=0.235
+ $X2=0 $Y2=0
cc_1097 N_A_1597_329#_M1009_g N_VGND_c_2275_n 0.00921786f $X=11.47 $Y=0.56 $X2=0
+ $Y2=0
cc_1098 N_A_1597_329#_c_1565_n N_VGND_c_2275_n 0.00566354f $X=10.35 $Y=0.765
+ $X2=0 $Y2=0
cc_1099 N_A_1597_329#_c_1589_n N_VGND_c_2275_n 0.0518412f $X=9.71 $Y=0.41 $X2=0
+ $Y2=0
cc_1100 N_A_1597_329#_c_1570_n N_VGND_c_2275_n 0.0132422f $X=10.35 $Y=0.93 $X2=0
+ $Y2=0
cc_1101 N_A_1597_329#_c_1589_n A_1815_47# 0.00482916f $X=9.71 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1102 N_A_1597_329#_c_1589_n A_1887_47# 0.00620261f $X=9.71 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1103 N_A_2227_47#_M1003_g N_VPWR_c_1857_n 0.00185392f $X=11.945 $Y=1.985
+ $X2=0 $Y2=0
cc_1104 N_A_2227_47#_c_1722_n N_VPWR_c_1857_n 0.0248205f $X=11.89 $Y=1.16 $X2=0
+ $Y2=0
cc_1105 N_A_2227_47#_c_1724_n N_VPWR_c_1857_n 0.00248507f $X=13.255 $Y=1.16
+ $X2=0 $Y2=0
cc_1106 N_A_2227_47#_M1024_g N_VPWR_c_1858_n 0.00402871f $X=12.365 $Y=1.985
+ $X2=0 $Y2=0
cc_1107 N_A_2227_47#_M1028_g N_VPWR_c_1858_n 0.00153851f $X=12.835 $Y=1.985
+ $X2=0 $Y2=0
cc_1108 N_A_2227_47#_c_1724_n N_VPWR_c_1858_n 0.00300514f $X=13.255 $Y=1.16
+ $X2=0 $Y2=0
cc_1109 N_A_2227_47#_M1045_g N_VPWR_c_1860_n 0.00325148f $X=13.255 $Y=1.985
+ $X2=0 $Y2=0
cc_1110 N_A_2227_47#_M1003_g N_VPWR_c_1865_n 0.00583607f $X=11.945 $Y=1.985
+ $X2=0 $Y2=0
cc_1111 N_A_2227_47#_M1024_g N_VPWR_c_1865_n 0.004671f $X=12.365 $Y=1.985 $X2=0
+ $Y2=0
cc_1112 N_A_2227_47#_c_1729_n N_VPWR_c_1871_n 0.018001f $X=11.26 $Y=1.955 $X2=0
+ $Y2=0
cc_1113 N_A_2227_47#_M1028_g N_VPWR_c_1872_n 0.00541359f $X=12.835 $Y=1.985
+ $X2=0 $Y2=0
cc_1114 N_A_2227_47#_M1045_g N_VPWR_c_1872_n 0.00541359f $X=13.255 $Y=1.985
+ $X2=0 $Y2=0
cc_1115 N_A_2227_47#_M1016_s N_VPWR_c_1851_n 0.00382897f $X=11.135 $Y=1.485
+ $X2=0 $Y2=0
cc_1116 N_A_2227_47#_M1003_g N_VPWR_c_1851_n 0.010591f $X=11.945 $Y=1.985 $X2=0
+ $Y2=0
cc_1117 N_A_2227_47#_M1024_g N_VPWR_c_1851_n 0.00793368f $X=12.365 $Y=1.985
+ $X2=0 $Y2=0
cc_1118 N_A_2227_47#_M1028_g N_VPWR_c_1851_n 0.00962851f $X=12.835 $Y=1.985
+ $X2=0 $Y2=0
cc_1119 N_A_2227_47#_M1045_g N_VPWR_c_1851_n 0.0105203f $X=13.255 $Y=1.985 $X2=0
+ $Y2=0
cc_1120 N_A_2227_47#_c_1729_n N_VPWR_c_1851_n 0.00993603f $X=11.26 $Y=1.955
+ $X2=0 $Y2=0
cc_1121 N_A_2227_47#_c_1718_n N_Q_c_2209_n 4.88119e-19 $X=12.365 $Y=0.995 $X2=0
+ $Y2=0
cc_1122 N_A_2227_47#_c_1719_n N_Q_c_2209_n 0.0100463f $X=12.835 $Y=0.995 $X2=0
+ $Y2=0
cc_1123 N_A_2227_47#_c_1720_n N_Q_c_2209_n 0.0131951f $X=13.255 $Y=0.995 $X2=0
+ $Y2=0
cc_1124 N_A_2227_47#_c_1724_n N_Q_c_2209_n 0.00789313f $X=13.255 $Y=1.16 $X2=0
+ $Y2=0
cc_1125 N_A_2227_47#_M1024_g N_Q_c_2213_n 7.32109e-19 $X=12.365 $Y=1.985 $X2=0
+ $Y2=0
cc_1126 N_A_2227_47#_M1028_g N_Q_c_2213_n 0.0152626f $X=12.835 $Y=1.985 $X2=0
+ $Y2=0
cc_1127 N_A_2227_47#_M1045_g N_Q_c_2213_n 0.0201414f $X=13.255 $Y=1.985 $X2=0
+ $Y2=0
cc_1128 N_A_2227_47#_c_1724_n N_Q_c_2216_n 0.0469367f $X=13.255 $Y=1.16 $X2=0
+ $Y2=0
cc_1129 N_A_2227_47#_c_1724_n N_Q_c_2217_n 0.0226865f $X=13.255 $Y=1.16 $X2=0
+ $Y2=0
cc_1130 N_A_2227_47#_c_1718_n Q 0.00383491f $X=12.365 $Y=0.995 $X2=0 $Y2=0
cc_1131 N_A_2227_47#_c_1724_n Q 0.00103509f $X=13.255 $Y=1.16 $X2=0 $Y2=0
cc_1132 N_A_2227_47#_c_1722_n Q 0.0227711f $X=11.89 $Y=1.16 $X2=0 $Y2=0
cc_1133 N_A_2227_47#_c_1724_n Q 0.0108353f $X=13.255 $Y=1.16 $X2=0 $Y2=0
cc_1134 N_A_2227_47#_M1003_g Q 0.0038601f $X=11.945 $Y=1.985 $X2=0 $Y2=0
cc_1135 N_A_2227_47#_M1024_g Q 0.00471923f $X=12.365 $Y=1.985 $X2=0 $Y2=0
cc_1136 N_A_2227_47#_M1028_g Q 8.13158e-19 $X=12.835 $Y=1.985 $X2=0 $Y2=0
cc_1137 N_A_2227_47#_M1024_g Q 0.0156806f $X=12.365 $Y=1.985 $X2=0 $Y2=0
cc_1138 N_A_2227_47#_c_1718_n N_Q_c_2226_n 0.00628523f $X=12.365 $Y=0.995 $X2=0
+ $Y2=0
cc_1139 N_A_2227_47#_c_1719_n N_Q_c_2226_n 5.39143e-19 $X=12.835 $Y=0.995 $X2=0
+ $Y2=0
cc_1140 N_A_2227_47#_c_1717_n Q 0.00387953f $X=11.945 $Y=0.995 $X2=0 $Y2=0
cc_1141 N_A_2227_47#_c_1718_n Q 0.00430017f $X=12.365 $Y=0.995 $X2=0 $Y2=0
cc_1142 N_A_2227_47#_c_1722_n Q 0.00454727f $X=11.89 $Y=1.16 $X2=0 $Y2=0
cc_1143 N_A_2227_47#_c_1724_n Q 0.00477356f $X=13.255 $Y=1.16 $X2=0 $Y2=0
cc_1144 N_A_2227_47#_M1024_g Q 0.00383491f $X=12.365 $Y=1.985 $X2=0 $Y2=0
cc_1145 N_A_2227_47#_c_1724_n Q 0.00105578f $X=13.255 $Y=1.16 $X2=0 $Y2=0
cc_1146 N_A_2227_47#_c_1717_n N_VGND_c_2254_n 0.00185392f $X=11.945 $Y=0.995
+ $X2=0 $Y2=0
cc_1147 N_A_2227_47#_c_1722_n N_VGND_c_2254_n 0.0248205f $X=11.89 $Y=1.16 $X2=0
+ $Y2=0
cc_1148 N_A_2227_47#_c_1724_n N_VGND_c_2254_n 0.00248507f $X=13.255 $Y=1.16
+ $X2=0 $Y2=0
cc_1149 N_A_2227_47#_c_1718_n N_VGND_c_2255_n 0.00319678f $X=12.365 $Y=0.995
+ $X2=0 $Y2=0
cc_1150 N_A_2227_47#_c_1719_n N_VGND_c_2255_n 0.00153851f $X=12.835 $Y=0.995
+ $X2=0 $Y2=0
cc_1151 N_A_2227_47#_c_1724_n N_VGND_c_2255_n 0.00323182f $X=13.255 $Y=1.16
+ $X2=0 $Y2=0
cc_1152 N_A_2227_47#_c_1720_n N_VGND_c_2257_n 0.00325148f $X=13.255 $Y=0.995
+ $X2=0 $Y2=0
cc_1153 N_A_2227_47#_c_1717_n N_VGND_c_2260_n 0.00583607f $X=11.945 $Y=0.995
+ $X2=0 $Y2=0
cc_1154 N_A_2227_47#_c_1718_n N_VGND_c_2260_n 0.00467644f $X=12.365 $Y=0.995
+ $X2=0 $Y2=0
cc_1155 N_A_2227_47#_c_1721_n N_VGND_c_2266_n 0.018001f $X=11.26 $Y=0.425 $X2=0
+ $Y2=0
cc_1156 N_A_2227_47#_c_1719_n N_VGND_c_2267_n 0.00541359f $X=12.835 $Y=0.995
+ $X2=0 $Y2=0
cc_1157 N_A_2227_47#_c_1720_n N_VGND_c_2267_n 0.00541359f $X=13.255 $Y=0.995
+ $X2=0 $Y2=0
cc_1158 N_A_2227_47#_M1009_s N_VGND_c_2275_n 0.00382897f $X=11.135 $Y=0.235
+ $X2=0 $Y2=0
cc_1159 N_A_2227_47#_c_1717_n N_VGND_c_2275_n 0.0106371f $X=11.945 $Y=0.995
+ $X2=0 $Y2=0
cc_1160 N_A_2227_47#_c_1718_n N_VGND_c_2275_n 0.00794368f $X=12.365 $Y=0.995
+ $X2=0 $Y2=0
cc_1161 N_A_2227_47#_c_1719_n N_VGND_c_2275_n 0.00962851f $X=12.835 $Y=0.995
+ $X2=0 $Y2=0
cc_1162 N_A_2227_47#_c_1720_n N_VGND_c_2275_n 0.0105203f $X=13.255 $Y=0.995
+ $X2=0 $Y2=0
cc_1163 N_A_2227_47#_c_1721_n N_VGND_c_2275_n 0.00993603f $X=11.26 $Y=0.425
+ $X2=0 $Y2=0
cc_1164 N_A_27_369#_c_1811_n N_VPWR_M1018_d 0.00303015f $X=0.955 $Y=1.935
+ $X2=-0.19 $Y2=1.305
cc_1165 N_A_27_369#_c_1811_n N_VPWR_c_1852_n 0.0142338f $X=0.955 $Y=1.935 $X2=0
+ $Y2=0
cc_1166 N_A_27_369#_c_1811_n N_VPWR_c_1861_n 0.00224471f $X=0.955 $Y=1.935 $X2=0
+ $Y2=0
cc_1167 N_A_27_369#_c_1825_n N_VPWR_c_1861_n 0.00965331f $X=1.125 $Y=2.36 $X2=0
+ $Y2=0
cc_1168 N_A_27_369#_c_1813_n N_VPWR_c_1861_n 0.0521802f $X=1.88 $Y=2.34 $X2=0
+ $Y2=0
cc_1169 N_A_27_369#_c_1810_n N_VPWR_c_1867_n 0.0178803f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1170 N_A_27_369#_c_1811_n N_VPWR_c_1867_n 0.00212534f $X=0.955 $Y=1.935 $X2=0
+ $Y2=0
cc_1171 N_A_27_369#_M1018_s N_VPWR_c_1851_n 0.00231948f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_1172 N_A_27_369#_M1001_d N_VPWR_c_1851_n 0.00209344f $X=1.745 $Y=1.845 $X2=0
+ $Y2=0
cc_1173 N_A_27_369#_c_1810_n N_VPWR_c_1851_n 0.00991202f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1174 N_A_27_369#_c_1811_n N_VPWR_c_1851_n 0.0089533f $X=0.955 $Y=1.935 $X2=0
+ $Y2=0
cc_1175 N_A_27_369#_c_1825_n N_VPWR_c_1851_n 0.00648546f $X=1.125 $Y=2.36 $X2=0
+ $Y2=0
cc_1176 N_A_27_369#_c_1813_n N_VPWR_c_1851_n 0.0329812f $X=1.88 $Y=2.34 $X2=0
+ $Y2=0
cc_1177 N_A_27_369#_c_1811_n A_193_369# 0.00140409f $X=0.955 $Y=1.935 $X2=-0.19
+ $Y2=1.305
cc_1178 N_A_27_369#_c_1825_n A_193_369# 9.36188e-19 $X=1.125 $Y=2.36 $X2=-0.19
+ $Y2=1.305
cc_1179 N_A_27_369#_c_1813_n N_A_181_47#_M1004_d 0.00313816f $X=1.88 $Y=2.34
+ $X2=0 $Y2=0
cc_1180 N_A_27_369#_c_1813_n N_A_181_47#_c_2077_n 0.0195387f $X=1.88 $Y=2.34
+ $X2=0 $Y2=0
cc_1181 N_A_27_369#_c_1813_n N_A_181_47#_c_2070_n 0.00156994f $X=1.88 $Y=2.34
+ $X2=0 $Y2=0
cc_1182 N_VPWR_c_1851_n A_193_369# 0.00168632f $X=13.57 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1183 N_VPWR_c_1851_n N_A_181_47#_M1004_d 0.00216833f $X=13.57 $Y=2.72 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1851_n N_A_181_47#_M1007_s 0.00197307f $X=13.57 $Y=2.72 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1869_n N_A_181_47#_c_2067_n 0.0132015f $X=5.945 $Y=2.72 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1851_n N_A_181_47#_c_2067_n 0.00390749f $X=13.57 $Y=2.72 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1853_n N_A_181_47#_c_2069_n 0.00784985f $X=2.82 $Y=2.34 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1851_n A_1081_413# 0.00244888f $X=13.57 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1189 N_VPWR_c_1877_n A_1525_329# 9.61034e-19 $X=8.015 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1190 N_VPWR_c_1851_n A_1723_413# 0.00232248f $X=13.57 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1191 N_VPWR_c_1851_n N_Q_M1003_d 0.00285153f $X=13.57 $Y=2.72 $X2=0 $Y2=0
cc_1192 N_VPWR_c_1851_n N_Q_M1028_d 0.00215201f $X=13.57 $Y=2.72 $X2=0 $Y2=0
cc_1193 N_VPWR_c_1872_n N_Q_c_2213_n 0.0189039f $X=13.38 $Y=2.72 $X2=0 $Y2=0
cc_1194 N_VPWR_c_1851_n N_Q_c_2213_n 0.0122217f $X=13.57 $Y=2.72 $X2=0 $Y2=0
cc_1195 N_VPWR_c_1858_n N_Q_c_2216_n 0.0134126f $X=12.625 $Y=1.66 $X2=0 $Y2=0
cc_1196 N_VPWR_c_1865_n Q 0.0179105f $X=12.54 $Y=2.72 $X2=0 $Y2=0
cc_1197 N_VPWR_c_1851_n Q 0.0121049f $X=13.57 $Y=2.72 $X2=0 $Y2=0
cc_1198 N_VPWR_c_1858_n Q 0.0704764f $X=12.625 $Y=1.66 $X2=0 $Y2=0
cc_1199 N_VPWR_c_1860_n N_VGND_c_2257_n 0.011741f $X=13.465 $Y=1.66 $X2=0 $Y2=0
cc_1200 N_A_181_47#_c_2063_n N_VGND_c_2250_n 0.0207323f $X=1.6 $Y=0.805 $X2=0
+ $Y2=0
cc_1201 N_A_181_47#_c_2073_n N_VGND_c_2258_n 0.0281961f $X=1.38 $Y=0.425 $X2=0
+ $Y2=0
cc_1202 N_A_181_47#_c_2063_n N_VGND_c_2258_n 0.0160536f $X=1.6 $Y=0.805 $X2=0
+ $Y2=0
cc_1203 N_A_181_47#_c_2061_n N_VGND_c_2264_n 0.0220997f $X=4.73 $Y=0.42 $X2=0
+ $Y2=0
cc_1204 N_A_181_47#_M1012_d N_VGND_c_2275_n 0.00215227f $X=0.905 $Y=0.235 $X2=0
+ $Y2=0
cc_1205 N_A_181_47#_M1020_s N_VGND_c_2275_n 0.00330824f $X=4.605 $Y=0.235 $X2=0
+ $Y2=0
cc_1206 N_A_181_47#_c_2073_n N_VGND_c_2275_n 0.0183005f $X=1.38 $Y=0.425 $X2=0
+ $Y2=0
cc_1207 N_A_181_47#_c_2061_n N_VGND_c_2275_n 0.0124358f $X=4.73 $Y=0.42 $X2=0
+ $Y2=0
cc_1208 N_A_181_47#_c_2063_n N_VGND_c_2275_n 0.0109812f $X=1.6 $Y=0.805 $X2=0
+ $Y2=0
cc_1209 N_A_181_47#_c_2063_n A_265_47# 0.00396213f $X=1.6 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_1210 N_Q_c_2216_n N_VGND_c_2255_n 0.0134124f $X=12.88 $Y=1.19 $X2=0 $Y2=0
cc_1211 N_Q_c_2226_n N_VGND_c_2255_n 0.044839f $X=12.155 $Y=0.44 $X2=0 $Y2=0
cc_1212 N_Q_c_2226_n N_VGND_c_2260_n 0.0173391f $X=12.155 $Y=0.44 $X2=0 $Y2=0
cc_1213 N_Q_c_2209_n N_VGND_c_2267_n 0.0189039f $X=13.045 $Y=0.36 $X2=0 $Y2=0
cc_1214 N_Q_M1022_d N_VGND_c_2275_n 0.00290484f $X=12.02 $Y=0.235 $X2=0 $Y2=0
cc_1215 N_Q_M1032_d N_VGND_c_2275_n 0.00215201f $X=12.91 $Y=0.235 $X2=0 $Y2=0
cc_1216 N_Q_c_2209_n N_VGND_c_2275_n 0.0122217f $X=13.045 $Y=0.36 $X2=0 $Y2=0
cc_1217 N_Q_c_2226_n N_VGND_c_2275_n 0.0121108f $X=12.155 $Y=0.44 $X2=0 $Y2=0
cc_1218 N_VGND_c_2268_n A_109_47# 9.17637e-19 $X=0.23 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1219 N_VGND_c_2275_n A_109_47# 7.33531e-19 $X=13.57 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1220 N_VGND_c_2275_n A_265_47# 0.00216812f $X=13.57 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1221 N_VGND_c_2275_n A_1087_47# 0.00726675f $X=13.57 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1222 N_VGND_c_2272_n A_1514_47# 0.0113551f $X=7.715 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1223 N_VGND_c_2275_n A_1514_47# 0.0128754f $X=13.57 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1224 N_VGND_c_2275_n A_1815_47# 0.00169327f $X=13.57 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1225 N_VGND_c_2275_n A_1887_47# 0.00266073f $X=13.57 $Y=0 $X2=-0.19 $Y2=-0.24

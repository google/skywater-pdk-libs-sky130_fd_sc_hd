* File: sky130_fd_sc_hd__dlrtp_1.spice
* Created: Thu Aug 27 14:17:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlrtp_1.spice.pex"
.subckt sky130_fd_sc_hd__dlrtp_1  VNB VPB GATE D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_GATE_M1019_g N_A_27_47#_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_193_47#_M1010_d N_A_27_47#_M1010_g N_VGND_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_D_M1003_g N_A_299_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1006 A_465_47# N_A_299_47#_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07665 AS=0.0567 PD=0.785 PS=0.69 NRD=36.42 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_560_425#_M1007_d N_A_193_47#_M1007_g A_465_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.07665 PD=0.7 PS=0.785 NRD=0 NRS=36.42 M=1 R=2.8
+ SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 A_654_47# N_A_27_47#_M1015_g N_A_560_425#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.05985 AS=0.0588 PD=0.705 PS=0.7 NRD=24.996 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_711_21#_M1016_g A_654_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.05985 PD=1.36 PS=0.705 NRD=0 NRS=24.996 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_929_47# N_A_560_425#_M1005_g N_A_711_21#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10725 AS=0.169 PD=0.98 PS=1.82 NRD=20.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_RESET_B_M1008_g A_929_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.10725 PD=0.96 PS=0.98 NRD=6.456 NRS=20.304 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_Q_M1017_d N_A_711_21#_M1017_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10075 PD=1.82 PS=0.96 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VPWR_M1009_d N_GATE_M1009_g N_A_27_47#_M1009_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_VPWR_M1014_d N_D_M1014_g N_A_299_47#_M1014_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1012 A_465_369# N_A_299_47#_M1012_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.11968 AS=0.0864 PD=1.2352 PS=0.91 NRD=40.6214 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75002 A=0.096 P=1.58 MULT=1
MM1004 N_A_560_425#_M1004_d N_A_27_47#_M1004_g A_465_369# VPB PHIGHVT L=0.15
+ W=0.36 AD=0.0666 AS=0.06732 PD=0.73 PS=0.6948 NRD=19.1484 NRS=72.2202 M=1
+ R=2.4 SA=75001.1 SB=75003 A=0.054 P=1.02 MULT=1
MM1001 A_664_425# N_A_193_47#_M1001_g N_A_560_425#_M1004_d VPB PHIGHVT L=0.15
+ W=0.36 AD=0.0758769 AS=0.0666 PD=0.770769 PS=0.73 NRD=85.2222 NRS=30.0819 M=1
+ R=2.4 SA=75001.6 SB=75002.4 A=0.054 P=1.02 MULT=1
MM1018 N_VPWR_M1018_d N_A_711_21#_M1018_g A_664_425# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.118665 AS=0.0885231 PD=0.952394 PS=0.899231 NRD=0 NRS=73.0476 M=1 R=2.8
+ SA=75001.9 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 N_A_711_21#_M1002_d N_A_560_425#_M1002_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.165 AS=0.282535 PD=1.33 PS=2.26761 NRD=5.8903 NRS=0 M=1
+ R=6.66667 SA=75001.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_RESET_B_M1013_g N_A_711_21#_M1002_d VPB PHIGHVT L=0.15
+ W=1 AD=0.155 AS=0.165 PD=1.31 PS=1.33 NRD=6.8753 NRS=3.9203 M=1 R=6.66667
+ SA=75001.7 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_Q_M1011_d N_A_711_21#_M1011_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.155 PD=2.52 PS=1.31 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_134 VPB 0 2.44684e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dlrtp_1.spice.SKY130_FD_SC_HD__DLRTP_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__and4bb_2.spice
* Created: Thu Aug 27 14:09:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and4bb_2.spice.pex"
.subckt sky130_fd_sc_hd__and4bb_2  VNB VPB A_N C D B_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B_N	B_N
* D	D
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1013_d N_A_174_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.08775 PD=1.18458 PS=0.92 NRD=9.228 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_174_21#_M1015_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 A_476_47# N_A_27_47#_M1010_g N_A_174_21#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1011 A_548_47# N_A_505_280#_M1011_g A_476_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=27.852 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 A_639_47# N_C_M1009_g A_548_47# VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.06405 PD=0.69 PS=0.725 NRD=22.848 NRS=27.852 M=1 R=2.8 SA=75001
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_D_M1004_g A_639_47# VNB NSHORT L=0.15 W=0.42 AD=0.0924
+ AS=0.0567 PD=0.86 PS=0.69 NRD=47.136 NRS=22.848 M=1 R=2.8 SA=75001.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_505_280#_M1008_d N_B_N_M1008_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0924 PD=1.36 PS=0.86 NRD=0 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_27_47#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0832606 AS=0.1092 PD=0.783803 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.8 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1005_d N_A_174_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.198239 AS=0.135 PD=1.8662 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75000.4 SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_174_21#_M1001_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.465845 AS=0.135 PD=2.40141 PS=1.27 NRD=14.7553 NRS=0 M=1 R=6.66667
+ SA=75000.8 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_174_21#_M1002_d N_A_27_47#_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0672 AS=0.195655 PD=0.74 PS=1.00859 NRD=21.0987 NRS=4.6886 M=1
+ R=2.8 SA=75001.9 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_505_280#_M1012_g N_A_174_21#_M1002_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_174_21#_M1006_d N_C_M1006_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.0588 PD=0.69 PS=0.7 NRD=0 NRS=2.3443 M=1 R=2.8 SA=75002.8
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_D_M1014_g N_A_174_21#_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0924 AS=0.0567 PD=0.86 PS=0.69 NRD=77.3816 NRS=0 M=1 R=2.8 SA=75003.3
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_505_280#_M1007_d N_B_N_M1007_g N_VPWR_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0924 PD=1.36 PS=0.86 NRD=0 NRS=0 M=1 R=2.8 SA=75003.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hd__and4bb_2.spice.SKY130_FD_SC_HD__AND4BB_2.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__and4bb_2.pex.spice
* Created: Thu Aug 27 14:09:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4BB_2%A_N 3 7 9 10 17
c27 7 0 1.57019e-19 $X=0.47 $Y=2.275
r28 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r29 9 10 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.16 $X2=0.24
+ $Y2=1.53
r30 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r31 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r32 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.275
r33 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r34 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%A_174_21# 1 2 3 10 12 15 17 19 22 26 27 29
+ 30 33 36 39 41 42 45 48
r105 53 55 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.945 $Y=1.16
+ $X2=1.365 $Y2=1.16
r106 50 52 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.32 $Y=2 $X2=2.48
+ $Y2=2
r107 47 48 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.095 $Y=0.72
+ $X2=2.32 $Y2=0.72
r108 43 45 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.33 $Y=2.085
+ $X2=3.33 $Y2=2.3
r109 42 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=2 $X2=2.48
+ $Y2=2
r110 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=2
+ $X2=3.33 $Y2=2.085
r111 41 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.245 $Y=2
+ $X2=2.565 $Y2=2
r112 37 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=2.085
+ $X2=2.48 $Y2=2
r113 37 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.48 $Y=2.085
+ $X2=2.48 $Y2=2.3
r114 36 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=1.915
+ $X2=2.32 $Y2=2
r115 35 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=0.805
+ $X2=2.32 $Y2=0.72
r116 35 36 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=2.32 $Y=0.805
+ $X2=2.32 $Y2=1.915
r117 31 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.635
+ $X2=2.095 $Y2=0.72
r118 31 33 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.095 $Y=0.635
+ $X2=2.095 $Y2=0.42
r119 29 47 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=0.72
+ $X2=2.095 $Y2=0.72
r120 29 30 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.01 $Y=0.72
+ $X2=1.585 $Y2=0.72
r121 27 55 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.5 $Y=1.16
+ $X2=1.365 $Y2=1.16
r122 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.16 $X2=1.5 $Y2=1.16
r123 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.5 $Y=0.805
+ $X2=1.585 $Y2=0.72
r124 24 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.5 $Y=0.805
+ $X2=1.5 $Y2=1.16
r125 20 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.16
r126 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.365 $Y=1.325
+ $X2=1.365 $Y2=1.985
r127 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=1.16
r128 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=0.56
r129 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.325
+ $X2=0.945 $Y2=1.16
r130 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.945 $Y=1.325
+ $X2=0.945 $Y2=1.985
r131 10 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=1.16
r132 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.56
r133 3 45 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=2.065 $X2=3.33 $Y2=2.3
r134 2 39 600 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=2.065 $X2=2.48 $Y2=2.3
r135 1 33 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.095 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%A_27_47# 1 2 7 9 11 13 16 20 23 24 25 27 30
+ 38
r91 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=1.16 $X2=1.98 $Y2=1.16
r92 35 38 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.84 $Y=1.16
+ $X2=1.98 $Y2=1.16
r93 32 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.26 $Y=1.97
+ $X2=0.585 $Y2=1.97
r94 28 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.26 $Y=0.72
+ $X2=0.585 $Y2=0.72
r95 26 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.16
r96 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.885
r97 25 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.97
+ $X2=0.585 $Y2=1.97
r98 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.755 $Y=1.97
+ $X2=1.84 $Y2=1.885
r99 24 25 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=1.755 $Y=1.97
+ $X2=0.67 $Y2=1.97
r100 23 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=1.885
+ $X2=0.585 $Y2=1.97
r101 22 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=0.805
+ $X2=0.585 $Y2=0.72
r102 22 23 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=0.585 $Y=0.805
+ $X2=0.585 $Y2=1.885
r103 18 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.055
+ $X2=0.26 $Y2=1.97
r104 18 20 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.26 $Y=2.055
+ $X2=0.26 $Y2=2.3
r105 14 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.72
r106 14 16 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.42
r107 11 39 69.2658 $w=4.45e-07 $l=5.17581e-07 $layer=POLY_cond $X=2.305 $Y=0.73
+ $X2=2.112 $Y2=1.16
r108 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.305 $Y=0.73
+ $X2=2.305 $Y2=0.445
r109 7 39 40.5624 $w=4.45e-07 $l=2.12238e-07 $layer=POLY_cond $X=2.22 $Y=1.325
+ $X2=2.112 $Y2=1.16
r110 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.22 $Y=1.325
+ $X2=2.22 $Y2=2.275
r111 2 20 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r112 1 16 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%A_505_280# 1 2 9 13 15 18 19 20 23 26 28 29
+ 36 38
c72 28 0 1.43093e-19 $X=2.66 $Y=1.565
c73 20 0 1.25206e-19 $X=3.755 $Y=2
r74 34 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.34 $Y=0.42 $X2=4.43
+ $Y2=0.42
r75 29 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.565
+ $X2=2.66 $Y2=1.73
r76 29 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.565
+ $X2=2.66 $Y2=1.4
r77 28 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.66 $Y=1.565
+ $X2=2.66 $Y2=1.66
r78 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.565 $X2=2.66 $Y2=1.565
r79 26 38 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=4.43 $Y=1.915
+ $X2=4.385 $Y2=2
r80 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=0.585
+ $X2=4.43 $Y2=0.42
r81 25 26 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=4.43 $Y=0.585
+ $X2=4.43 $Y2=1.915
r82 21 38 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.385 $Y=2.085
+ $X2=4.385 $Y2=2
r83 21 23 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=4.385 $Y=2.085
+ $X2=4.385 $Y2=2.3
r84 19 38 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.255 $Y=2 $X2=4.385
+ $Y2=2
r85 19 20 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.255 $Y=2 $X2=3.755
+ $Y2=2
r86 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=1.915
+ $X2=3.755 $Y2=2
r87 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.67 $Y=1.745
+ $X2=3.67 $Y2=1.915
r88 16 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=1.66
+ $X2=2.66 $Y2=1.66
r89 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.585 $Y=1.66
+ $X2=3.67 $Y2=1.745
r90 15 16 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.585 $Y=1.66
+ $X2=2.745 $Y2=1.66
r91 13 41 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.69 $Y=2.275
+ $X2=2.69 $Y2=1.73
r92 9 40 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=2.665 $Y=0.445
+ $X2=2.665 $Y2=1.4
r93 2 23 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=2.065 $X2=4.34 $Y2=2.3
r94 1 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.235 $X2=4.34 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%C 3 6 8 9 10 15 17
c40 8 0 1.27131e-19 $X=2.995 $Y=0.51
c41 6 0 1.25206e-19 $X=3.12 $Y=2.275
r42 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.94
+ $X2=3.09 $Y2=1.105
r43 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.94
+ $X2=3.09 $Y2=0.775
r44 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=0.94 $X2=3.09 $Y2=0.94
r45 10 16 10.8721 $w=2.63e-07 $l=2.5e-07 $layer=LI1_cond $X=3.042 $Y=1.19
+ $X2=3.042 $Y2=0.94
r46 9 16 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=3.042 $Y=0.85 $X2=3.042
+ $Y2=0.94
r47 8 9 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=3.042 $Y=0.51
+ $X2=3.042 $Y2=0.85
r48 6 18 599.936 $w=1.5e-07 $l=1.17e-06 $layer=POLY_cond $X=3.12 $Y=2.275
+ $X2=3.12 $Y2=1.105
r49 3 17 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.12 $Y=0.445 $X2=3.12
+ $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%D 3 7 9 10 11 16
c44 9 0 1.43093e-19 $X=3.455 $Y=0.51
r45 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.24
+ $X2=3.57 $Y2=1.405
r46 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.24
+ $X2=3.57 $Y2=1.075
r47 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.24 $X2=3.57 $Y2=1.24
r48 11 17 1.88925 $w=3.03e-07 $l=5e-08 $layer=LI1_cond $X=3.502 $Y=1.19
+ $X2=3.502 $Y2=1.24
r49 10 11 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=3.502 $Y=0.85
+ $X2=3.502 $Y2=1.19
r50 9 10 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=3.502 $Y=0.51
+ $X2=3.502 $Y2=0.85
r51 7 19 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.54 $Y=2.275
+ $X2=3.54 $Y2=1.405
r52 3 18 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.54 $Y=0.445
+ $X2=3.54 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%B_N 3 6 8 9 13 15
r36 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=0.93
+ $X2=4.09 $Y2=1.095
r37 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=0.93
+ $X2=4.09 $Y2=0.765
r38 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=0.93 $X2=4.09 $Y2=0.93
r39 9 14 8.56101 $w=3.48e-07 $l=2.6e-07 $layer=LI1_cond $X=4 $Y=1.19 $X2=4
+ $Y2=0.93
r40 8 14 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=4 $Y=0.85 $X2=4
+ $Y2=0.93
r41 6 16 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=4.13 $Y=2.275
+ $X2=4.13 $Y2=1.095
r42 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.13 $Y=0.445
+ $X2=4.13 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%VPWR 1 2 3 4 15 19 23 25 27 37 42 49 50 53
+ 57 61 63 66
r79 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r80 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 59 61 8.20096 $w=5.48e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=2.53 $X2=2.16
+ $Y2=2.53
r82 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r83 56 59 1.63102 $w=5.48e-07 $l=7.5e-08 $layer=LI1_cond $X=1.995 $Y=2.53
+ $X2=2.07 $Y2=2.53
r84 56 57 17.2259 $w=5.48e-07 $l=5.05e-07 $layer=LI1_cond $X=1.995 $Y=2.53
+ $X2=1.49 $Y2=2.53
r85 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r87 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r88 47 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=3.92 $Y2=2.72
r89 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=4.37 $Y2=2.72
r90 46 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r91 46 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r92 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r93 43 63 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=2.905 $Y2=2.72
r94 43 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=3.45 $Y2=2.72
r95 42 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.92 $Y2=2.72
r96 42 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.45 $Y2=2.72
r97 41 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r98 41 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r99 40 61 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.53 $Y=2.72 $X2=2.16
+ $Y2=2.72
r100 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r101 37 63 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.735 $Y=2.72
+ $X2=2.905 $Y2=2.72
r102 37 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.735 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 36 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r104 36 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 35 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=1.49 $Y2=2.72
r106 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r107 33 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r108 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r109 27 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r110 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r111 25 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r112 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r113 21 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.92 $Y2=2.72
r114 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.92 $Y2=2.34
r115 17 63 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=2.635
+ $X2=2.905 $Y2=2.72
r116 17 19 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.905 $Y=2.635
+ $X2=2.905 $Y2=2.34
r117 13 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r118 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r119 4 23 600 $w=1.7e-07 $l=4.20595e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=2.065 $X2=3.92 $Y2=2.34
r120 3 19 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=2.065 $X2=2.9 $Y2=2.34
r121 2 56 300 $w=1.7e-07 $l=1.09798e-06 $layer=licon1_PDIFF $count=2 $X=1.44
+ $Y=1.485 $X2=1.995 $Y2=2.34
r122 1 15 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%X 1 2 7 8 9 16 24
c22 9 0 1.57019e-19 $X=1.07 $Y=1.445
r23 24 26 0.768295 $w=2.23e-07 $l=1.5e-08 $layer=LI1_cond $X=1.127 $Y=1.53
+ $X2=1.127 $Y2=1.545
r24 9 26 2.39662 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.155 $Y=1.58
+ $X2=1.155 $Y2=1.545
r25 9 24 1.79269 $w=2.23e-07 $l=3.5e-08 $layer=LI1_cond $X=1.127 $Y=1.495
+ $X2=1.127 $Y2=1.53
r26 8 9 15.622 $w=2.23e-07 $l=3.05e-07 $layer=LI1_cond $X=1.127 $Y=1.19
+ $X2=1.127 $Y2=1.495
r27 7 8 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.19
r28 7 16 22.0245 $w=2.23e-07 $l=4.3e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.42
r29 2 9 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.485 $X2=1.155 $Y2=1.63
r30 1 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_2%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
c76 20 0 1.27131e-19 $X=3.92 $Y=0.42
r77 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r78 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r79 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r80 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r81 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r82 39 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=3.96
+ $Y2=0
r83 39 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.37
+ $Y2=0
r84 38 52 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r85 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r86 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r87 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.575
+ $Y2=0
r88 35 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=2.07
+ $Y2=0
r89 34 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.835 $Y=0 $X2=3.96
+ $Y2=0
r90 34 37 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=3.835 $Y=0 $X2=2.07
+ $Y2=0
r91 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r92 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r93 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r94 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r95 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r96 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.575
+ $Y2=0
r97 29 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.15
+ $Y2=0
r98 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r99 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r100 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r101 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r102 18 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0
r103 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0.42
r104 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0
r105 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0.38
r106 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r107 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r108 3 20 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.235 $X2=3.92 $Y2=0.42
r109 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.575 $Y2=0.38
r110 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__nor4_1.spice
* Created: Thu Aug 27 14:32:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor4_1.pex.spice"
.subckt sky130_fd_sc_hd__nor4_1  VNB VPB D C B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_D_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.118625 AS=0.169 PD=1.015 PS=1.82 NRD=16.608 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_C_M1003_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.118625 PD=0.925 PS=1.015 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.089375 PD=0.92 PS=0.925 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1005 A_109_297# N_D_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.13 AS=0.26
+ PD=1.26 PS=2.52 NRD=14.7553 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.5 A=0.15
+ P=2.3 MULT=1
MM1004 A_191_297# N_C_M1004_g A_109_297# VPB PHIGHVT L=0.15 W=1 AD=0.19 AS=0.13
+ PD=1.38 PS=1.26 NRD=26.5753 NRS=14.7553 M=1 R=6.66667 SA=75000.6 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1000 A_297_297# N_B_M1000_g A_191_297# VPB PHIGHVT L=0.15 W=1 AD=0.135 AS=0.19
+ PD=1.27 PS=1.38 NRD=15.7403 NRS=26.5753 M=1 R=6.66667 SA=75001.1 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_297_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75001.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__nor4_1.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.065000 1.720000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985000 0.305000 7.320000 0.730000 ;
        RECT 6.985000 0.730000 8.655000 0.900000 ;
        RECT 6.985000 1.465000 8.655000 1.635000 ;
        RECT 6.985000 1.635000 7.320000 2.395000 ;
        RECT 7.840000 0.305000 8.175000 0.730000 ;
        RECT 7.840000 1.635000 8.170000 2.395000 ;
        RECT 8.410000 0.900000 8.655000 1.465000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.740000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.455000  0.085000 1.705000 0.545000 ;
        RECT 3.400000  0.085000 3.770000 0.585000 ;
        RECT 5.625000  0.085000 5.795000 0.615000 ;
        RECT 6.625000  0.085000 6.795000 0.565000 ;
        RECT 7.495000  0.085000 7.665000 0.560000 ;
        RECT 8.345000  0.085000 8.515000 0.560000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.740000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.440000 2.175000 1.705000 2.635000 ;
        RECT 3.610000 1.835000 3.780000 2.635000 ;
        RECT 5.490000 2.135000 5.705000 2.635000 ;
        RECT 6.625000 1.855000 6.805000 2.635000 ;
        RECT 7.500000 1.805000 7.670000 2.635000 ;
        RECT 8.340000 1.805000 8.510000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.840000 0.805000 ;
      RECT 0.175000 1.795000 0.840000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.610000 0.805000 0.840000 1.795000 ;
      RECT 1.015000 0.345000 1.240000 2.465000 ;
      RECT 1.890000 0.365000 2.220000 0.535000 ;
      RECT 1.890000 0.535000 2.060000 2.065000 ;
      RECT 1.890000 2.065000 2.125000 2.440000 ;
      RECT 2.230000 0.705000 2.810000 1.035000 ;
      RECT 2.230000 1.035000 2.470000 1.905000 ;
      RECT 2.370000 2.190000 3.440000 2.360000 ;
      RECT 2.400000 0.365000 3.150000 0.535000 ;
      RECT 2.660000 1.655000 3.100000 2.010000 ;
      RECT 2.980000 0.535000 3.150000 1.315000 ;
      RECT 2.980000 1.315000 3.780000 1.485000 ;
      RECT 3.270000 1.485000 3.780000 1.575000 ;
      RECT 3.270000 1.575000 3.440000 2.190000 ;
      RECT 3.320000 0.765000 4.120000 1.065000 ;
      RECT 3.320000 1.065000 3.490000 1.095000 ;
      RECT 3.610000 1.245000 3.780000 1.315000 ;
      RECT 3.950000 0.365000 4.410000 0.535000 ;
      RECT 3.950000 0.535000 4.120000 0.765000 ;
      RECT 3.950000 1.065000 4.120000 2.135000 ;
      RECT 3.950000 2.135000 4.200000 2.465000 ;
      RECT 4.290000 0.705000 4.840000 1.035000 ;
      RECT 4.290000 1.245000 4.480000 1.965000 ;
      RECT 4.425000 2.165000 5.310000 2.335000 ;
      RECT 4.640000 0.365000 5.310000 0.535000 ;
      RECT 4.650000 1.035000 4.840000 1.575000 ;
      RECT 4.650000 1.575000 4.970000 1.905000 ;
      RECT 5.140000 0.535000 5.310000 1.075000 ;
      RECT 5.140000 1.075000 6.230000 1.245000 ;
      RECT 5.140000 1.245000 5.310000 2.165000 ;
      RECT 5.480000 1.500000 6.590000 1.670000 ;
      RECT 5.480000 1.670000 6.340000 1.830000 ;
      RECT 6.090000 0.295000 6.450000 0.735000 ;
      RECT 6.090000 0.735000 6.590000 0.905000 ;
      RECT 6.170000 1.830000 6.340000 2.455000 ;
      RECT 6.420000 0.905000 6.590000 1.075000 ;
      RECT 6.420000 1.075000 8.240000 1.245000 ;
      RECT 6.420000 1.245000 6.590000 1.500000 ;
    LAYER mcon ;
      RECT 0.610000 1.785000 0.780000 1.955000 ;
      RECT 1.070000 0.765000 1.240000 0.935000 ;
      RECT 2.470000 0.765000 2.640000 0.935000 ;
      RECT 2.930000 1.785000 3.100000 1.955000 ;
      RECT 4.310000 0.765000 4.480000 0.935000 ;
      RECT 4.310000 1.785000 4.480000 1.955000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 4.540000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 4.540000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.410000 0.735000 2.700000 0.780000 ;
      RECT 2.410000 0.920000 2.700000 0.965000 ;
      RECT 2.870000 1.755000 3.160000 1.800000 ;
      RECT 2.870000 1.940000 3.160000 1.985000 ;
      RECT 4.250000 0.735000 4.540000 0.780000 ;
      RECT 4.250000 0.920000 4.540000 0.965000 ;
      RECT 4.250000 1.755000 4.540000 1.800000 ;
      RECT 4.250000 1.940000 4.540000 1.985000 ;
  END
END sky130_fd_sc_hd__dfxtp_4

* File: sky130_fd_sc_hd__a311oi_4.pxi.spice
* Created: Thu Aug 27 14:04:28 2020
* 
x_PM_SKY130_FD_SC_HD__A311OI_4%A3 N_A3_c_107_n N_A3_M1015_g N_A3_M1004_g
+ N_A3_c_108_n N_A3_M1021_g N_A3_M1007_g N_A3_c_109_n N_A3_M1026_g N_A3_M1027_g
+ N_A3_c_110_n N_A3_M1039_g N_A3_M1037_g A3 A3 A3 A3 N_A3_c_111_n
+ PM_SKY130_FD_SC_HD__A311OI_4%A3
x_PM_SKY130_FD_SC_HD__A311OI_4%A2 N_A2_c_177_n N_A2_M1022_g N_A2_M1001_g
+ N_A2_c_178_n N_A2_M1028_g N_A2_M1008_g N_A2_c_179_n N_A2_M1034_g N_A2_M1031_g
+ N_A2_c_180_n N_A2_M1035_g N_A2_M1038_g A2 A2 A2 A2 N_A2_c_182_n
+ PM_SKY130_FD_SC_HD__A311OI_4%A2
x_PM_SKY130_FD_SC_HD__A311OI_4%A1 N_A1_M1003_g N_A1_M1012_g N_A1_c_248_n
+ N_A1_M1013_g N_A1_M1017_g N_A1_c_249_n N_A1_M1016_g N_A1_M1025_g N_A1_c_250_n
+ N_A1_M1023_g N_A1_c_251_n N_A1_M1029_g A1 A1 A1 A1 N_A1_c_252_n
+ PM_SKY130_FD_SC_HD__A311OI_4%A1
x_PM_SKY130_FD_SC_HD__A311OI_4%B1 N_B1_c_316_n N_B1_M1010_g N_B1_M1002_g
+ N_B1_c_317_n N_B1_M1014_g N_B1_M1005_g N_B1_c_318_n N_B1_M1019_g N_B1_M1009_g
+ N_B1_c_319_n N_B1_M1024_g N_B1_M1032_g B1 B1 B1 N_B1_c_320_n N_B1_c_321_n
+ PM_SKY130_FD_SC_HD__A311OI_4%B1
x_PM_SKY130_FD_SC_HD__A311OI_4%C1 N_C1_c_386_n N_C1_M1011_g N_C1_M1000_g
+ N_C1_c_387_n N_C1_M1018_g N_C1_M1006_g N_C1_c_388_n N_C1_M1030_g N_C1_M1020_g
+ N_C1_c_389_n N_C1_M1033_g N_C1_M1036_g C1 C1 C1 C1 N_C1_c_390_n
+ PM_SKY130_FD_SC_HD__A311OI_4%C1
x_PM_SKY130_FD_SC_HD__A311OI_4%VPWR N_VPWR_M1004_s N_VPWR_M1007_s N_VPWR_M1037_s
+ N_VPWR_M1008_s N_VPWR_M1038_s N_VPWR_M1012_d N_VPWR_M1025_d N_VPWR_c_461_n
+ N_VPWR_c_462_n N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n N_VPWR_c_466_n
+ N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n
+ N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n VPWR
+ N_VPWR_c_476_n N_VPWR_c_477_n N_VPWR_c_478_n N_VPWR_c_460_n N_VPWR_c_480_n
+ N_VPWR_c_481_n N_VPWR_c_482_n PM_SKY130_FD_SC_HD__A311OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A311OI_4%A_109_297# N_A_109_297#_M1004_d
+ N_A_109_297#_M1027_d N_A_109_297#_M1001_d N_A_109_297#_M1031_d
+ N_A_109_297#_M1003_s N_A_109_297#_M1017_s N_A_109_297#_M1002_d
+ N_A_109_297#_M1009_d N_A_109_297#_c_647_n N_A_109_297#_c_598_n
+ N_A_109_297#_c_602_n N_A_109_297#_c_651_n N_A_109_297#_c_604_n
+ N_A_109_297#_c_655_n N_A_109_297#_c_610_n N_A_109_297#_c_659_n
+ N_A_109_297#_c_614_n N_A_109_297#_c_663_n N_A_109_297#_c_622_n
+ N_A_109_297#_c_667_n N_A_109_297#_c_597_n N_A_109_297#_c_606_n
+ N_A_109_297#_c_616_n N_A_109_297#_c_618_n N_A_109_297#_c_629_n
+ PM_SKY130_FD_SC_HD__A311OI_4%A_109_297#
x_PM_SKY130_FD_SC_HD__A311OI_4%A_1139_297# N_A_1139_297#_M1002_s
+ N_A_1139_297#_M1005_s N_A_1139_297#_M1032_s N_A_1139_297#_M1006_d
+ N_A_1139_297#_M1036_d N_A_1139_297#_c_679_n N_A_1139_297#_c_680_n
+ N_A_1139_297#_c_681_n PM_SKY130_FD_SC_HD__A311OI_4%A_1139_297#
x_PM_SKY130_FD_SC_HD__A311OI_4%Y N_Y_M1013_s N_Y_M1016_s N_Y_M1029_s N_Y_M1014_s
+ N_Y_M1024_s N_Y_M1018_s N_Y_M1033_s N_Y_M1000_s N_Y_M1020_s N_Y_c_720_n
+ N_Y_c_802_p N_Y_c_733_n N_Y_c_742_n N_Y_c_743_n N_Y_c_747_n N_Y_c_749_n
+ N_Y_c_805_p N_Y_c_753_n N_Y_c_808_p N_Y_c_737_n N_Y_c_739_n N_Y_c_762_n
+ N_Y_c_764_n Y Y Y Y Y Y PM_SKY130_FD_SC_HD__A311OI_4%Y
x_PM_SKY130_FD_SC_HD__A311OI_4%A_27_47# N_A_27_47#_M1015_d N_A_27_47#_M1021_d
+ N_A_27_47#_M1039_d N_A_27_47#_M1028_s N_A_27_47#_M1035_s N_A_27_47#_c_856_p
+ N_A_27_47#_c_831_n N_A_27_47#_c_835_n N_A_27_47#_c_859_p N_A_27_47#_c_837_n
+ N_A_27_47#_c_862_p N_A_27_47#_c_830_n N_A_27_47#_c_841_n N_A_27_47#_c_849_n
+ PM_SKY130_FD_SC_HD__A311OI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__A311OI_4%VGND N_VGND_M1015_s N_VGND_M1026_s N_VGND_M1010_d
+ N_VGND_M1019_d N_VGND_M1011_d N_VGND_M1030_d N_VGND_c_880_n N_VGND_c_881_n
+ N_VGND_c_882_n N_VGND_c_883_n N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n
+ VGND N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n
+ N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n N_VGND_c_895_n
+ N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n N_VGND_c_899_n
+ PM_SKY130_FD_SC_HD__A311OI_4%VGND
x_PM_SKY130_FD_SC_HD__A311OI_4%A_445_47# N_A_445_47#_M1022_d N_A_445_47#_M1034_d
+ N_A_445_47#_M1013_d N_A_445_47#_M1023_d N_A_445_47#_c_1030_n
+ PM_SKY130_FD_SC_HD__A311OI_4%A_445_47#
cc_1 VNB N_A3_c_107_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A3_c_108_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A3_c_109_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A3_c_110_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A3_c_111_n 0.0941763f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_6 VNB N_A2_c_177_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_7 VNB N_A2_c_178_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_8 VNB N_A2_c_179_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_9 VNB N_A2_c_180_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_10 VNB A2 0.00613911f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_11 VNB N_A2_c_182_n 0.0609554f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_12 VNB N_A1_c_248_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_13 VNB N_A1_c_249_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_14 VNB N_A1_c_250_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_15 VNB N_A1_c_251_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_16 VNB N_A1_c_252_n 0.094602f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.16
cc_17 VNB N_B1_c_316_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_18 VNB N_B1_c_317_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_19 VNB N_B1_c_318_n 0.0157734f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_20 VNB N_B1_c_319_n 0.0176599f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_21 VNB N_B1_c_320_n 0.00205078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_B1_c_321_n 0.0677119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_C1_c_386_n 0.0176711f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_24 VNB N_C1_c_387_n 0.0157752f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_25 VNB N_C1_c_388_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_26 VNB N_C1_c_389_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_27 VNB N_C1_c_390_n 0.0963992f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.16
cc_28 VNB N_VPWR_c_460_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_720_n 0.00209549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB Y 0.0111366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_830_n 0.00248013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_880_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_881_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_34 VNB N_VGND_c_882_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_35 VNB N_VGND_c_883_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_884_n 0.0169862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_885_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_38 VNB N_VGND_c_886_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_39 VNB N_VGND_c_887_n 0.0151407f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_40 VNB N_VGND_c_888_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_41 VNB N_VGND_c_889_n 0.102905f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.16
cc_42 VNB N_VGND_c_890_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_891_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_892_n 0.0151407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_893_n 0.452945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_894_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_895_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_896_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_897_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_898_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_899_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_445_47#_c_1030_n 0.00650014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_A3_M1004_g 0.02509f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_54 VPB N_A3_M1007_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_55 VPB N_A3_M1027_g 0.0182793f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_56 VPB N_A3_M1037_g 0.0185651f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_57 VPB N_A3_c_111_n 0.0188402f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_58 VPB N_A2_M1001_g 0.0185651f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_59 VPB N_A2_M1008_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_60 VPB N_A2_M1031_g 0.0182793f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_61 VPB N_A2_M1038_g 0.0185651f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_62 VPB A2 0.00216082f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_63 VPB N_A2_c_182_n 0.0100051f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_64 VPB N_A1_M1003_g 0.01753f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_65 VPB N_A1_M1012_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A1_M1017_g 0.0172788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A1_M1025_g 0.0208795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A1_c_252_n 0.0335064f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_69 VPB N_B1_M1002_g 0.0223275f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_70 VPB N_B1_M1005_g 0.0171325f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_71 VPB N_B1_M1009_g 0.0178141f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_72 VPB N_B1_M1032_g 0.0207779f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_73 VPB N_B1_c_320_n 0.00504128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B1_c_321_n 0.0136011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_C1_M1000_g 0.0208084f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_76 VPB N_C1_M1006_g 0.0185023f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_77 VPB N_C1_M1020_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_78 VPB N_C1_M1036_g 0.0259842f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_79 VPB N_C1_c_390_n 0.0217476f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_80 VPB N_VPWR_c_461_n 0.0103102f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_81 VPB N_VPWR_c_462_n 0.0386297f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_82 VPB N_VPWR_c_463_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_83 VPB N_VPWR_c_464_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_465_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_85 VPB N_VPWR_c_466_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_86 VPB N_VPWR_c_467_n 0.0124915f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_87 VPB N_VPWR_c_468_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_469_n 0.00551074f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_89 VPB N_VPWR_c_470_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_471_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_91 VPB N_VPWR_c_472_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_473_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_474_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_475_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_476_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_477_n 0.0117278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_478_n 0.100841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_460_n 0.0471986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_480_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_481_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_482_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_109_297#_c_597_n 0.00842332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_1139_297#_c_679_n 0.00218948f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_104 VPB N_A_1139_297#_c_680_n 0.00747916f $X=-0.19 $Y=1.305 $X2=1.73
+ $Y2=1.985
cc_105 VPB N_A_1139_297#_c_681_n 0.0166149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB Y 0.00519606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 N_A3_c_110_n N_A2_c_177_n 0.0234661f $X=1.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_108 N_A3_M1037_g N_A2_M1001_g 0.0234661f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_109 A3 A2 0.0258519f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_110 N_A3_c_111_n A2 0.00289706f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_111 A3 N_A2_c_182_n 2.92893e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_112 N_A3_c_111_n N_A2_c_182_n 0.0234661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A3_M1004_g N_VPWR_c_462_n 0.0149251f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A3_M1007_g N_VPWR_c_462_n 7.5193e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_115 A3 N_VPWR_c_462_n 0.0166542f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_116 N_A3_c_111_n N_VPWR_c_462_n 0.00632846f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A3_M1004_g N_VPWR_c_463_n 6.0901e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A3_M1007_g N_VPWR_c_463_n 0.0102874f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A3_M1027_g N_VPWR_c_463_n 0.0102874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A3_M1037_g N_VPWR_c_463_n 6.0901e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A3_M1027_g N_VPWR_c_464_n 6.0901e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A3_M1037_g N_VPWR_c_464_n 0.0102535f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A3_M1027_g N_VPWR_c_470_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A3_M1037_g N_VPWR_c_470_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A3_M1004_g N_VPWR_c_476_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A3_M1007_g N_VPWR_c_476_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A3_M1004_g N_VPWR_c_460_n 0.00789179f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A3_M1007_g N_VPWR_c_460_n 0.00789179f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A3_M1027_g N_VPWR_c_460_n 0.00789179f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A3_M1037_g N_VPWR_c_460_n 0.00789179f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A3_M1007_g N_A_109_297#_c_598_n 0.0136764f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A3_M1027_g N_A_109_297#_c_598_n 0.0141087f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_133 A3 N_A_109_297#_c_598_n 0.0409723f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A3_c_111_n N_A_109_297#_c_598_n 0.00201785f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_135 A3 N_A_109_297#_c_602_n 0.0134105f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A3_c_111_n N_A_109_297#_c_602_n 0.00209661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A3_M1037_g N_A_109_297#_c_604_n 0.0162466f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_138 A3 N_A_109_297#_c_604_n 0.00758912f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_139 A3 N_A_109_297#_c_606_n 0.0134105f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A3_c_111_n N_A_109_297#_c_606_n 0.00209661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A3_c_107_n N_A_27_47#_c_831_n 0.0127817f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A3_c_108_n N_A_27_47#_c_831_n 0.0115294f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_143 A3 N_A_27_47#_c_831_n 0.0375135f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A3_c_111_n N_A_27_47#_c_831_n 0.0019918f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_145 A3 N_A_27_47#_c_835_n 0.0123848f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A3_c_111_n N_A_27_47#_c_835_n 0.00386661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A3_c_109_n N_A_27_47#_c_837_n 0.0115735f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A3_c_110_n N_A_27_47#_c_837_n 0.0136104f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_149 A3 N_A_27_47#_c_837_n 0.0312246f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A3_c_111_n N_A_27_47#_c_837_n 0.0019918f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_151 A3 N_A_27_47#_c_841_n 0.0121035f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A3_c_111_n N_A_27_47#_c_841_n 0.00205824f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A3_c_107_n N_VGND_c_880_n 0.00834749f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A3_c_108_n N_VGND_c_880_n 0.00664421f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A3_c_109_n N_VGND_c_880_n 5.08801e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A3_c_108_n N_VGND_c_881_n 5.08801e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A3_c_109_n N_VGND_c_881_n 0.00664421f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A3_c_110_n N_VGND_c_881_n 0.00784221f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A3_c_107_n N_VGND_c_887_n 0.00339367f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A3_c_108_n N_VGND_c_888_n 0.00339367f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A3_c_109_n N_VGND_c_888_n 0.00339367f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A3_c_110_n N_VGND_c_889_n 0.00339367f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A3_c_107_n N_VGND_c_893_n 0.00489827f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A3_c_108_n N_VGND_c_893_n 0.00394406f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A3_c_109_n N_VGND_c_893_n 0.00394406f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A3_c_110_n N_VGND_c_893_n 0.00397127f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_M1038_g N_A1_M1003_g 0.0226383f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_168 A2 A1 0.021551f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A2_c_182_n A1 3.44632e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_170 A2 N_A1_c_252_n 0.00276779f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A2_c_182_n N_A1_c_252_n 0.0226383f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A2_M1001_g N_VPWR_c_464_n 0.0102535f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A2_M1008_g N_VPWR_c_464_n 6.0901e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A2_M1001_g N_VPWR_c_465_n 6.0901e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A2_M1008_g N_VPWR_c_465_n 0.0102874f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A2_M1031_g N_VPWR_c_465_n 0.0102874f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M1038_g N_VPWR_c_465_n 6.0901e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_M1031_g N_VPWR_c_466_n 6.0901e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_M1038_g N_VPWR_c_466_n 0.0102535f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_VPWR_c_472_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A2_M1008_g N_VPWR_c_472_n 0.0046653f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A2_M1031_g N_VPWR_c_474_n 0.0046653f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A2_M1038_g N_VPWR_c_474_n 0.0046653f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A2_M1001_g N_VPWR_c_460_n 0.00789179f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A2_M1008_g N_VPWR_c_460_n 0.00789179f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A2_M1031_g N_VPWR_c_460_n 0.00789179f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A2_M1038_g N_VPWR_c_460_n 0.00789179f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A2_M1001_g N_A_109_297#_c_604_n 0.0141087f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_189 A2 N_A_109_297#_c_604_n 0.0214312f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_190 N_A2_M1008_g N_A_109_297#_c_610_n 0.0141528f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A2_M1031_g N_A_109_297#_c_610_n 0.0141528f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_192 A2 N_A_109_297#_c_610_n 0.0409723f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_193 N_A2_c_182_n N_A_109_297#_c_610_n 0.00201785f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A2_M1038_g N_A_109_297#_c_614_n 0.0141087f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_195 A2 N_A_109_297#_c_614_n 0.0155848f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_196 A2 N_A_109_297#_c_616_n 0.0134105f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_197 N_A2_c_182_n N_A_109_297#_c_616_n 0.00209661f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_198 A2 N_A_109_297#_c_618_n 0.0134105f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A2_c_182_n N_A_109_297#_c_618_n 0.00209661f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A2_c_177_n N_A_27_47#_c_830_n 0.011544f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A2_c_178_n N_A_27_47#_c_830_n 0.00847802f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A2_c_179_n N_A_27_47#_c_830_n 0.00847802f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A2_c_180_n N_A_27_47#_c_830_n 0.00847802f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_204 A2 N_A_27_47#_c_830_n 0.0872482f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_205 N_A2_c_182_n N_A_27_47#_c_830_n 0.00597539f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_206 A2 N_A_27_47#_c_849_n 0.00680018f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_207 N_A2_c_177_n N_VGND_c_881_n 0.00116167f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A2_c_177_n N_VGND_c_889_n 0.00413298f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A2_c_178_n N_VGND_c_889_n 0.00366111f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A2_c_179_n N_VGND_c_889_n 0.00366111f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A2_c_180_n N_VGND_c_889_n 0.00366111f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A2_c_177_n N_VGND_c_893_n 0.00570263f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A2_c_178_n N_VGND_c_893_n 0.00524008f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A2_c_179_n N_VGND_c_893_n 0.00524008f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A2_c_180_n N_VGND_c_893_n 0.00661716f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A2_c_177_n N_A_445_47#_c_1030_n 0.00245853f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A2_c_178_n N_A_445_47#_c_1030_n 0.00789149f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A2_c_179_n N_A_445_47#_c_1030_n 0.00789149f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A2_c_180_n N_A_445_47#_c_1030_n 0.00999448f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A1_c_251_n N_B1_c_316_n 0.0257108f $X=5.61 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_221 A1 N_B1_c_320_n 0.02034f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_222 N_A1_c_252_n N_B1_c_320_n 0.0187421f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_223 N_A1_c_252_n N_B1_c_321_n 0.0216032f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_224 N_A1_M1003_g N_VPWR_c_466_n 0.0102535f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A1_M1012_g N_VPWR_c_466_n 6.0901e-19 $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A1_M1003_g N_VPWR_c_467_n 0.0046653f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A1_M1012_g N_VPWR_c_467_n 0.0046653f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A1_M1003_g N_VPWR_c_468_n 6.0901e-19 $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A1_M1012_g N_VPWR_c_468_n 0.0102874f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A1_M1017_g N_VPWR_c_468_n 0.010268f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_M1025_g N_VPWR_c_468_n 5.59199e-19 $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A1_M1017_g N_VPWR_c_469_n 5.08801e-19 $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_M1025_g N_VPWR_c_469_n 0.00774571f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A1_M1017_g N_VPWR_c_477_n 0.0046653f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A1_M1025_g N_VPWR_c_477_n 0.00339367f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A1_M1003_g N_VPWR_c_460_n 0.00789179f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A1_M1012_g N_VPWR_c_460_n 0.00789179f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A1_M1017_g N_VPWR_c_460_n 0.00789179f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A1_M1025_g N_VPWR_c_460_n 0.00394406f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A1_M1003_g N_A_109_297#_c_614_n 0.0155129f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_241 A1 N_A_109_297#_c_614_n 0.00901737f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_242 N_A1_M1012_g N_A_109_297#_c_622_n 0.0141087f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A1_M1017_g N_A_109_297#_c_622_n 0.0136764f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_244 A1 N_A_109_297#_c_622_n 0.0543828f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_245 N_A1_c_252_n N_A_109_297#_c_622_n 0.00493857f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_246 N_A1_M1025_g N_A_109_297#_c_597_n 0.0135496f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_247 A1 N_A_109_297#_c_597_n 0.0107554f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_248 N_A1_c_252_n N_A_109_297#_c_597_n 0.0111383f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_249 A1 N_A_109_297#_c_629_n 0.0134105f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_250 N_A1_c_252_n N_A_109_297#_c_629_n 0.00217288f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_251 N_A1_c_248_n N_Y_c_720_n 0.00847802f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_249_n N_Y_c_720_n 0.00847802f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_250_n N_Y_c_720_n 0.00847802f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_251_n N_Y_c_720_n 0.0132923f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_255 A1 N_Y_c_720_n 0.0853445f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_256 N_A1_c_252_n N_Y_c_720_n 0.0143752f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_257 N_A1_c_252_n N_A_27_47#_c_830_n 0.00121861f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_258 N_A1_c_251_n N_VGND_c_882_n 0.0018398f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_c_248_n N_VGND_c_889_n 0.00366111f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A1_c_249_n N_VGND_c_889_n 0.00366111f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A1_c_250_n N_VGND_c_889_n 0.00366111f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A1_c_251_n N_VGND_c_889_n 0.00413298f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A1_c_248_n N_VGND_c_893_n 0.00661716f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A1_c_249_n N_VGND_c_893_n 0.00524008f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A1_c_250_n N_VGND_c_893_n 0.00524008f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A1_c_251_n N_VGND_c_893_n 0.00574665f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A1_c_248_n N_A_445_47#_c_1030_n 0.00999448f $X=4.35 $Y=0.995 $X2=0
+ $Y2=0
cc_268 N_A1_c_249_n N_A_445_47#_c_1030_n 0.00789149f $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A1_c_250_n N_A_445_47#_c_1030_n 0.00789149f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A1_c_251_n N_A_445_47#_c_1030_n 0.00363095f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_271 A1 N_A_445_47#_c_1030_n 0.00542351f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_272 N_A1_c_252_n N_A_445_47#_c_1030_n 0.00423751f $X=5.19 $Y=1.17 $X2=0 $Y2=0
cc_273 N_B1_c_319_n N_C1_c_386_n 0.013756f $X=7.29 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_274 N_B1_M1032_g N_C1_M1000_g 0.013756f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B1_c_321_n N_C1_c_390_n 0.013756f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B1_M1002_g N_VPWR_c_469_n 0.00294182f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B1_M1002_g N_VPWR_c_478_n 0.00366111f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B1_M1005_g N_VPWR_c_478_n 0.00366111f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B1_M1009_g N_VPWR_c_478_n 0.00366111f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B1_M1032_g N_VPWR_c_478_n 0.00366111f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B1_M1002_g N_VPWR_c_460_n 0.00656615f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_282 N_B1_M1005_g N_VPWR_c_460_n 0.00524008f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_283 N_B1_M1009_g N_VPWR_c_460_n 0.00524008f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B1_M1032_g N_VPWR_c_460_n 0.00571579f $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_285 N_B1_c_320_n N_A_109_297#_M1002_d 0.00219451f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B1_M1002_g N_A_109_297#_c_597_n 0.0111157f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_287 N_B1_M1005_g N_A_109_297#_c_597_n 0.00901269f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_B1_M1009_g N_A_109_297#_c_597_n 0.0113392f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_289 N_B1_M1032_g N_A_109_297#_c_597_n 0.00487813f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_B1_c_320_n N_A_109_297#_c_597_n 0.0477267f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_291 N_B1_c_321_n N_A_109_297#_c_597_n 0.00295878f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B1_c_320_n N_A_1139_297#_M1002_s 0.00340475f $X=6.77 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_293 N_B1_c_320_n N_A_1139_297#_M1005_s 0.00219451f $X=6.77 $Y=1.16 $X2=0
+ $Y2=0
cc_294 N_B1_M1002_g N_A_1139_297#_c_679_n 0.00789149f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_B1_M1005_g N_A_1139_297#_c_679_n 0.00789149f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_B1_M1009_g N_A_1139_297#_c_679_n 0.00789149f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_B1_M1032_g N_A_1139_297#_c_679_n 0.0115259f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_B1_c_316_n N_Y_c_720_n 0.00957617f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B1_c_317_n N_Y_c_720_n 0.0115735f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B1_c_320_n N_Y_c_720_n 0.0554268f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_301 N_B1_c_321_n N_Y_c_720_n 0.0031865f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_302 N_B1_c_318_n N_Y_c_733_n 0.0142491f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B1_c_319_n N_Y_c_733_n 0.0170066f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_304 N_B1_c_320_n N_Y_c_733_n 0.00603295f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_305 N_B1_c_321_n N_Y_c_733_n 0.00330881f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_306 N_B1_c_320_n N_Y_c_737_n 0.0127201f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_307 N_B1_c_321_n N_Y_c_737_n 0.00205824f $X=7.29 $Y=1.16 $X2=0 $Y2=0
cc_308 N_B1_M1032_g N_Y_c_739_n 5.48211e-19 $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_309 N_B1_c_319_n Y 0.015829f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B1_c_320_n Y 0.0186894f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_311 N_B1_c_316_n N_VGND_c_882_n 0.0093418f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_312 N_B1_c_317_n N_VGND_c_882_n 0.00664421f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B1_c_318_n N_VGND_c_882_n 5.08801e-19 $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B1_c_317_n N_VGND_c_883_n 5.08801e-19 $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_315 N_B1_c_318_n N_VGND_c_883_n 0.00664421f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B1_c_319_n N_VGND_c_883_n 0.00796297f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B1_c_319_n N_VGND_c_884_n 0.00339367f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_319_n N_VGND_c_885_n 8.8473e-19 $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_319 N_B1_c_316_n N_VGND_c_889_n 0.00339367f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_320 N_B1_c_317_n N_VGND_c_890_n 0.00339367f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_321 N_B1_c_318_n N_VGND_c_890_n 0.00339367f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B1_c_316_n N_VGND_c_893_n 0.00401529f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B1_c_317_n N_VGND_c_893_n 0.00394406f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_324 N_B1_c_318_n N_VGND_c_893_n 0.00394406f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_325 N_B1_c_319_n N_VGND_c_893_n 0.00441977f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B1_c_316_n N_A_445_47#_c_1030_n 4.913e-19 $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_327 N_C1_M1000_g N_VPWR_c_478_n 0.00366111f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_328 N_C1_M1006_g N_VPWR_c_478_n 0.00366111f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_329 N_C1_M1020_g N_VPWR_c_478_n 0.00366111f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_330 N_C1_M1036_g N_VPWR_c_478_n 0.00366111f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_331 N_C1_M1000_g N_VPWR_c_460_n 0.00577307f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_332 N_C1_M1006_g N_VPWR_c_460_n 0.00524008f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_333 N_C1_M1020_g N_VPWR_c_460_n 0.00524008f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_334 N_C1_M1036_g N_VPWR_c_460_n 0.00619429f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_335 N_C1_M1000_g N_A_109_297#_c_597_n 4.8914e-19 $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_336 N_C1_M1000_g N_A_1139_297#_c_679_n 0.0122896f $X=7.93 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_C1_M1006_g N_A_1139_297#_c_679_n 0.00931965f $X=8.35 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_C1_M1020_g N_A_1139_297#_c_679_n 0.00931965f $X=8.77 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_C1_M1036_g N_A_1139_297#_c_679_n 0.0115553f $X=9.19 $Y=1.985 $X2=0
+ $Y2=0
cc_340 C1 N_A_1139_297#_c_681_n 0.00732571f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_341 N_C1_c_390_n N_A_1139_297#_c_681_n 0.00451952f $X=9.415 $Y=1.16 $X2=0
+ $Y2=0
cc_342 N_C1_c_386_n N_Y_c_742_n 0.00514161f $X=7.93 $Y=0.995 $X2=0 $Y2=0
cc_343 N_C1_c_386_n N_Y_c_743_n 0.0149256f $X=7.93 $Y=0.995 $X2=0 $Y2=0
cc_344 N_C1_c_387_n N_Y_c_743_n 0.0115735f $X=8.35 $Y=0.995 $X2=0 $Y2=0
cc_345 C1 N_Y_c_743_n 0.0305713f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_346 N_C1_c_390_n N_Y_c_743_n 0.0019918f $X=9.415 $Y=1.16 $X2=0 $Y2=0
cc_347 N_C1_M1000_g N_Y_c_747_n 0.0108927f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_348 C1 N_Y_c_747_n 0.00229682f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_349 N_C1_M1006_g N_Y_c_749_n 0.00876469f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_350 N_C1_M1020_g N_Y_c_749_n 0.00876469f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_351 C1 N_Y_c_749_n 0.0268173f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_352 N_C1_c_390_n N_Y_c_749_n 0.00195183f $X=9.415 $Y=1.16 $X2=0 $Y2=0
cc_353 N_C1_c_388_n N_Y_c_753_n 0.0115294f $X=8.77 $Y=0.995 $X2=0 $Y2=0
cc_354 N_C1_c_389_n N_Y_c_753_n 0.0127817f $X=9.19 $Y=0.995 $X2=0 $Y2=0
cc_355 C1 N_Y_c_753_n 0.0498983f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_356 N_C1_c_390_n N_Y_c_753_n 0.0058584f $X=9.415 $Y=1.16 $X2=0 $Y2=0
cc_357 N_C1_M1000_g N_Y_c_739_n 0.0071106f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_358 N_C1_M1006_g N_Y_c_739_n 0.00800641f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_359 N_C1_M1020_g N_Y_c_739_n 0.00108523f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_360 C1 N_Y_c_739_n 0.0186506f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_361 N_C1_c_390_n N_Y_c_739_n 0.00204168f $X=9.415 $Y=1.16 $X2=0 $Y2=0
cc_362 C1 N_Y_c_762_n 0.0121035f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_363 N_C1_c_390_n N_Y_c_762_n 0.00205824f $X=9.415 $Y=1.16 $X2=0 $Y2=0
cc_364 N_C1_M1006_g N_Y_c_764_n 0.00108523f $X=8.35 $Y=1.985 $X2=0 $Y2=0
cc_365 N_C1_M1020_g N_Y_c_764_n 0.00774392f $X=8.77 $Y=1.985 $X2=0 $Y2=0
cc_366 N_C1_M1036_g N_Y_c_764_n 0.0168837f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_367 C1 N_Y_c_764_n 0.0176184f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_368 N_C1_c_390_n N_Y_c_764_n 0.00202223f $X=9.415 $Y=1.16 $X2=0 $Y2=0
cc_369 N_C1_M1000_g Y 0.00291124f $X=7.93 $Y=1.985 $X2=0 $Y2=0
cc_370 N_C1_c_390_n Y 0.00737944f $X=9.415 $Y=1.16 $X2=0 $Y2=0
cc_371 N_C1_c_386_n Y 0.00737944f $X=7.93 $Y=0.995 $X2=0 $Y2=0
cc_372 C1 Y 0.0242824f $X=9.34 $Y=1.105 $X2=0 $Y2=0
cc_373 N_C1_c_386_n N_VGND_c_883_n 8.88674e-19 $X=7.93 $Y=0.995 $X2=0 $Y2=0
cc_374 N_C1_c_386_n N_VGND_c_884_n 0.00339367f $X=7.93 $Y=0.995 $X2=0 $Y2=0
cc_375 N_C1_c_386_n N_VGND_c_885_n 0.00904556f $X=7.93 $Y=0.995 $X2=0 $Y2=0
cc_376 N_C1_c_387_n N_VGND_c_885_n 0.00664421f $X=8.35 $Y=0.995 $X2=0 $Y2=0
cc_377 N_C1_c_388_n N_VGND_c_885_n 5.08801e-19 $X=8.77 $Y=0.995 $X2=0 $Y2=0
cc_378 N_C1_c_387_n N_VGND_c_886_n 5.08801e-19 $X=8.35 $Y=0.995 $X2=0 $Y2=0
cc_379 N_C1_c_388_n N_VGND_c_886_n 0.00664421f $X=8.77 $Y=0.995 $X2=0 $Y2=0
cc_380 N_C1_c_389_n N_VGND_c_886_n 0.00834749f $X=9.19 $Y=0.995 $X2=0 $Y2=0
cc_381 N_C1_c_387_n N_VGND_c_891_n 0.00339367f $X=8.35 $Y=0.995 $X2=0 $Y2=0
cc_382 N_C1_c_388_n N_VGND_c_891_n 0.00339367f $X=8.77 $Y=0.995 $X2=0 $Y2=0
cc_383 N_C1_c_389_n N_VGND_c_892_n 0.00339367f $X=9.19 $Y=0.995 $X2=0 $Y2=0
cc_384 N_C1_c_386_n N_VGND_c_893_n 0.00448104f $X=7.93 $Y=0.995 $X2=0 $Y2=0
cc_385 N_C1_c_387_n N_VGND_c_893_n 0.00394406f $X=8.35 $Y=0.995 $X2=0 $Y2=0
cc_386 N_C1_c_388_n N_VGND_c_893_n 0.00394406f $X=8.77 $Y=0.995 $X2=0 $Y2=0
cc_387 N_C1_c_389_n N_VGND_c_893_n 0.00489827f $X=9.19 $Y=0.995 $X2=0 $Y2=0
cc_388 N_VPWR_c_460_n N_A_109_297#_M1004_d 0.00562358f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_389 N_VPWR_c_460_n N_A_109_297#_M1027_d 0.00562358f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_460_n N_A_109_297#_M1001_d 0.00562358f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_460_n N_A_109_297#_M1031_d 0.00562358f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_460_n N_A_109_297#_M1003_s 0.00562358f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_460_n N_A_109_297#_M1017_s 0.00405853f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_460_n N_A_109_297#_M1002_d 0.00219239f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_460_n N_A_109_297#_M1009_d 0.00219239f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_476_n N_A_109_297#_c_647_n 0.0113958f $X=0.935 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_460_n N_A_109_297#_c_647_n 0.00646998f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_398 N_VPWR_M1007_s N_A_109_297#_c_598_n 0.00342716f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_463_n N_A_109_297#_c_598_n 0.0127176f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_400 N_VPWR_c_470_n N_A_109_297#_c_651_n 0.0113958f $X=1.775 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_460_n N_A_109_297#_c_651_n 0.00646998f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_M1037_s N_A_109_297#_c_604_n 0.00564044f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_464_n N_A_109_297#_c_604_n 0.0127176f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_404 N_VPWR_c_472_n N_A_109_297#_c_655_n 0.0113958f $X=2.615 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_460_n N_A_109_297#_c_655_n 0.00646998f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_M1008_s N_A_109_297#_c_610_n 0.00342716f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_465_n N_A_109_297#_c_610_n 0.0127176f $X=2.78 $Y=2 $X2=0 $Y2=0
cc_408 N_VPWR_c_474_n N_A_109_297#_c_659_n 0.0113958f $X=3.455 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_460_n N_A_109_297#_c_659_n 0.00646998f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_M1038_s N_A_109_297#_c_614_n 0.0077029f $X=3.485 $Y=1.485 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_466_n N_A_109_297#_c_614_n 0.0127176f $X=3.62 $Y=2 $X2=0 $Y2=0
cc_412 N_VPWR_c_467_n N_A_109_297#_c_663_n 0.0113958f $X=4.295 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_460_n N_A_109_297#_c_663_n 0.00646998f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_M1012_d N_A_109_297#_c_622_n 0.0034223f $X=4.325 $Y=1.485 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_468_n N_A_109_297#_c_622_n 0.0127176f $X=4.46 $Y=2 $X2=0 $Y2=0
cc_416 N_VPWR_c_477_n N_A_109_297#_c_667_n 0.0113958f $X=5.135 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_460_n N_A_109_297#_c_667_n 0.00646998f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_M1025_d N_A_109_297#_c_597_n 0.00626492f $X=5.165 $Y=1.485 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_469_n N_A_109_297#_c_597_n 0.0206068f $X=5.3 $Y=2.34 $X2=0 $Y2=0
cc_420 N_VPWR_c_477_n N_A_109_297#_c_597_n 0.00243651f $X=5.135 $Y=2.72 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_478_n N_A_109_297#_c_597_n 0.00346265f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_460_n N_A_109_297#_c_597_n 0.013968f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_423 N_VPWR_c_460_n N_A_1139_297#_M1002_s 0.00211652f $X=9.43 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_424 N_VPWR_c_460_n N_A_1139_297#_M1005_s 0.00217615f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_460_n N_A_1139_297#_M1032_s 0.00399252f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_460_n N_A_1139_297#_M1006_d 0.00217615f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_460_n N_A_1139_297#_M1036_d 0.00211581f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_469_n N_A_1139_297#_c_679_n 0.0137364f $X=5.3 $Y=2.34 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_478_n N_A_1139_297#_c_679_n 0.163054f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_460_n N_A_1139_297#_c_679_n 0.126943f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_478_n N_A_1139_297#_c_680_n 0.0136988f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_460_n N_A_1139_297#_c_680_n 0.00939829f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_460_n N_Y_M1000_s 0.00219239f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_434 N_VPWR_c_460_n N_Y_M1020_s 0.00219239f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_435 N_A_109_297#_c_597_n N_A_1139_297#_M1002_s 0.00552234f $X=7.08 $Y=2
+ $X2=-0.19 $Y2=1.305
cc_436 N_A_109_297#_c_597_n N_A_1139_297#_M1005_s 0.00357959f $X=7.08 $Y=2 $X2=0
+ $Y2=0
cc_437 N_A_109_297#_M1002_d N_A_1139_297#_c_679_n 0.00325828f $X=6.105 $Y=1.485
+ $X2=0 $Y2=0
cc_438 N_A_109_297#_M1009_d N_A_1139_297#_c_679_n 0.00325828f $X=6.945 $Y=1.485
+ $X2=0 $Y2=0
cc_439 N_A_109_297#_c_597_n N_A_1139_297#_c_679_n 0.0797617f $X=7.08 $Y=2 $X2=0
+ $Y2=0
cc_440 N_A_1139_297#_c_679_n N_Y_M1000_s 0.00325424f $X=9.315 $Y=2.34 $X2=0
+ $Y2=0
cc_441 N_A_1139_297#_c_679_n N_Y_M1020_s 0.00325424f $X=9.315 $Y=2.34 $X2=0
+ $Y2=0
cc_442 N_A_1139_297#_M1032_s N_Y_c_747_n 0.00402452f $X=7.365 $Y=1.485 $X2=0
+ $Y2=0
cc_443 N_A_1139_297#_c_679_n N_Y_c_747_n 0.00507861f $X=9.315 $Y=2.34 $X2=0
+ $Y2=0
cc_444 N_A_1139_297#_M1006_d N_Y_c_749_n 0.00457143f $X=8.425 $Y=1.485 $X2=0
+ $Y2=0
cc_445 N_A_1139_297#_c_679_n N_Y_c_749_n 0.011054f $X=9.315 $Y=2.34 $X2=0 $Y2=0
cc_446 N_A_1139_297#_c_679_n N_Y_c_739_n 0.0158292f $X=9.315 $Y=2.34 $X2=0 $Y2=0
cc_447 N_A_1139_297#_c_679_n N_Y_c_764_n 0.0157959f $X=9.315 $Y=2.34 $X2=0 $Y2=0
cc_448 N_A_1139_297#_M1032_s Y 0.0129123f $X=7.365 $Y=1.485 $X2=0 $Y2=0
cc_449 N_A_1139_297#_c_679_n Y 0.0156553f $X=9.315 $Y=2.34 $X2=0 $Y2=0
cc_450 N_A_1139_297#_M1032_s Y 0.00148304f $X=7.365 $Y=1.485 $X2=0 $Y2=0
cc_451 N_Y_c_720_n N_A_27_47#_c_830_n 0.0145425f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_452 N_Y_c_720_n N_VGND_M1010_d 0.00312394f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_453 N_Y_c_733_n N_VGND_M1019_d 0.00517199f $X=7.415 $Y=0.72 $X2=0 $Y2=0
cc_454 N_Y_c_743_n N_VGND_M1011_d 0.00312394f $X=8.475 $Y=0.72 $X2=0 $Y2=0
cc_455 N_Y_c_753_n N_VGND_M1030_d 0.00312394f $X=9.315 $Y=0.72 $X2=0 $Y2=0
cc_456 N_Y_c_720_n N_VGND_c_882_n 0.0159625f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_457 N_Y_c_733_n N_VGND_c_883_n 0.0159625f $X=7.415 $Y=0.72 $X2=0 $Y2=0
cc_458 N_Y_c_733_n N_VGND_c_884_n 0.00244309f $X=7.415 $Y=0.72 $X2=0 $Y2=0
cc_459 N_Y_c_742_n N_VGND_c_884_n 0.0116048f $X=7.5 $Y=0.42 $X2=0 $Y2=0
cc_460 N_Y_c_743_n N_VGND_c_884_n 0.00360658f $X=8.475 $Y=0.72 $X2=0 $Y2=0
cc_461 Y N_VGND_c_884_n 0.00289856f $X=7.53 $Y=0.765 $X2=0 $Y2=0
cc_462 N_Y_c_742_n N_VGND_c_885_n 0.00817611f $X=7.5 $Y=0.42 $X2=0 $Y2=0
cc_463 N_Y_c_743_n N_VGND_c_885_n 0.0159625f $X=8.475 $Y=0.72 $X2=0 $Y2=0
cc_464 N_Y_c_753_n N_VGND_c_886_n 0.0159625f $X=9.315 $Y=0.72 $X2=0 $Y2=0
cc_465 N_Y_c_720_n N_VGND_c_889_n 0.00775032f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_466 N_Y_c_720_n N_VGND_c_890_n 0.00244309f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_467 N_Y_c_802_p N_VGND_c_890_n 0.0112274f $X=6.66 $Y=0.42 $X2=0 $Y2=0
cc_468 N_Y_c_733_n N_VGND_c_890_n 0.00244309f $X=7.415 $Y=0.72 $X2=0 $Y2=0
cc_469 N_Y_c_743_n N_VGND_c_891_n 0.00244309f $X=8.475 $Y=0.72 $X2=0 $Y2=0
cc_470 N_Y_c_805_p N_VGND_c_891_n 0.0112274f $X=8.56 $Y=0.42 $X2=0 $Y2=0
cc_471 N_Y_c_753_n N_VGND_c_891_n 0.00244309f $X=9.315 $Y=0.72 $X2=0 $Y2=0
cc_472 N_Y_c_753_n N_VGND_c_892_n 0.00244309f $X=9.315 $Y=0.72 $X2=0 $Y2=0
cc_473 N_Y_c_808_p N_VGND_c_892_n 0.01143f $X=9.4 $Y=0.42 $X2=0 $Y2=0
cc_474 N_Y_M1013_s N_VGND_c_893_n 0.00212464f $X=4.015 $Y=0.235 $X2=0 $Y2=0
cc_475 N_Y_M1016_s N_VGND_c_893_n 0.00219239f $X=4.845 $Y=0.235 $X2=0 $Y2=0
cc_476 N_Y_M1029_s N_VGND_c_893_n 0.00315309f $X=5.685 $Y=0.235 $X2=0 $Y2=0
cc_477 N_Y_M1014_s N_VGND_c_893_n 0.00249348f $X=6.525 $Y=0.235 $X2=0 $Y2=0
cc_478 N_Y_M1024_s N_VGND_c_893_n 0.00509403f $X=7.365 $Y=0.235 $X2=0 $Y2=0
cc_479 N_Y_M1018_s N_VGND_c_893_n 0.00249348f $X=8.425 $Y=0.235 $X2=0 $Y2=0
cc_480 N_Y_M1033_s N_VGND_c_893_n 0.00368727f $X=9.265 $Y=0.235 $X2=0 $Y2=0
cc_481 N_Y_c_720_n N_VGND_c_893_n 0.0218108f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_482 N_Y_c_802_p N_VGND_c_893_n 0.00643448f $X=6.66 $Y=0.42 $X2=0 $Y2=0
cc_483 N_Y_c_733_n N_VGND_c_893_n 0.00984256f $X=7.415 $Y=0.72 $X2=0 $Y2=0
cc_484 N_Y_c_742_n N_VGND_c_893_n 0.00646998f $X=7.5 $Y=0.42 $X2=0 $Y2=0
cc_485 N_Y_c_743_n N_VGND_c_893_n 0.0118672f $X=8.475 $Y=0.72 $X2=0 $Y2=0
cc_486 N_Y_c_805_p N_VGND_c_893_n 0.00643448f $X=8.56 $Y=0.42 $X2=0 $Y2=0
cc_487 N_Y_c_753_n N_VGND_c_893_n 0.00984256f $X=9.315 $Y=0.72 $X2=0 $Y2=0
cc_488 N_Y_c_808_p N_VGND_c_893_n 0.00643448f $X=9.4 $Y=0.42 $X2=0 $Y2=0
cc_489 Y N_VGND_c_893_n 0.00451323f $X=7.53 $Y=0.765 $X2=0 $Y2=0
cc_490 N_Y_c_720_n N_A_445_47#_M1013_d 0.00312766f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_491 N_Y_c_720_n N_A_445_47#_M1023_d 0.00409235f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_492 N_Y_M1013_s N_A_445_47#_c_1030_n 0.00476093f $X=4.015 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_Y_M1016_s N_A_445_47#_c_1030_n 0.00315945f $X=4.845 $Y=0.235 $X2=0
+ $Y2=0
cc_494 N_Y_c_720_n N_A_445_47#_c_1030_n 0.0797583f $X=6.575 $Y=0.72 $X2=0 $Y2=0
cc_495 N_A_27_47#_c_831_n N_VGND_M1015_s 0.00312394f $X=1.015 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_496 N_A_27_47#_c_837_n N_VGND_M1026_s 0.00312394f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_831_n N_VGND_c_880_n 0.0159625f $X=1.015 $Y=0.72 $X2=0 $Y2=0
cc_498 N_A_27_47#_c_837_n N_VGND_c_881_n 0.0159625f $X=1.855 $Y=0.72 $X2=0 $Y2=0
cc_499 N_A_27_47#_c_856_p N_VGND_c_887_n 0.01143f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_500 N_A_27_47#_c_831_n N_VGND_c_887_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_c_831_n N_VGND_c_888_n 0.00244309f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_c_859_p N_VGND_c_888_n 0.0112274f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_503 N_A_27_47#_c_837_n N_VGND_c_888_n 0.00244309f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_c_837_n N_VGND_c_889_n 0.00244309f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_c_862_p N_VGND_c_889_n 0.0112274f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_506 N_A_27_47#_c_830_n N_VGND_c_889_n 0.00245287f $X=3.62 $Y=0.72 $X2=0 $Y2=0
cc_507 N_A_27_47#_M1015_d N_VGND_c_893_n 0.00368727f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_M1021_d N_VGND_c_893_n 0.00249348f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_M1039_d N_VGND_c_893_n 0.00249348f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_M1028_s N_VGND_c_893_n 0.00219239f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_M1035_s N_VGND_c_893_n 0.00212464f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_512 N_A_27_47#_c_856_p N_VGND_c_893_n 0.00643448f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_513 N_A_27_47#_c_831_n N_VGND_c_893_n 0.00984256f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_859_p N_VGND_c_893_n 0.00643448f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_515 N_A_27_47#_c_837_n N_VGND_c_893_n 0.00984256f $X=1.855 $Y=0.72 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_c_862_p N_VGND_c_893_n 0.00643448f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_517 N_A_27_47#_c_830_n N_VGND_c_893_n 0.00707809f $X=3.62 $Y=0.72 $X2=0 $Y2=0
cc_518 N_A_27_47#_c_830_n N_A_445_47#_M1022_d 0.00312766f $X=3.62 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_519 N_A_27_47#_c_830_n N_A_445_47#_M1034_d 0.00312766f $X=3.62 $Y=0.72 $X2=0
+ $Y2=0
cc_520 N_A_27_47#_M1028_s N_A_445_47#_c_1030_n 0.00315945f $X=2.645 $Y=0.235
+ $X2=0 $Y2=0
cc_521 N_A_27_47#_M1035_s N_A_445_47#_c_1030_n 0.00498385f $X=3.485 $Y=0.235
+ $X2=0 $Y2=0
cc_522 N_A_27_47#_c_830_n N_A_445_47#_c_1030_n 0.0797583f $X=3.62 $Y=0.72 $X2=0
+ $Y2=0
cc_523 N_VGND_c_893_n N_A_445_47#_M1022_d 0.00217615f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_524 N_VGND_c_893_n N_A_445_47#_M1034_d 0.00217615f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_893_n N_A_445_47#_M1013_d 0.00217615f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_893_n N_A_445_47#_M1023_d 0.00217615f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_882_n N_A_445_47#_c_1030_n 0.00545039f $X=6.24 $Y=0.38 $X2=0
+ $Y2=0
cc_528 N_VGND_c_889_n N_A_445_47#_c_1030_n 0.151358f $X=6.075 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_893_n N_A_445_47#_c_1030_n 0.117456f $X=9.43 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__xor2_1.spice
* Created: Tue Sep  1 19:33:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__xor2_1.pex.spice"
.subckt sky130_fd_sc_hd__xor2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1005 N_A_35_297#_M1005_d N_B_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_M1008_g N_A_35_297#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1000 A_285_47# N_A_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001 SB=75001.6
+ A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_B_M1003_g A_285_47# VNB NSHORT L=0.15 W=0.65 AD=0.25025
+ AS=0.08775 PD=1.42 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75001.4 SB=75001.2
+ A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A_35_297#_M1001_g N_X_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.208 AS=0.25025 PD=1.94 PS=1.42 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 A_117_297# N_B_M1009_g N_A_35_297#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_117_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75000.6 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1004 N_A_285_297#_M1004_d N_A_M1004_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g N_A_285_297#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_35_297#_M1007_g N_A_285_297#_M1007_s VPB PHIGHVT L=0.15
+ W=1 AD=0.3 AS=0.26 PD=2.6 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__xor2_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o41a_4.spice.pex
* Created: Thu Aug 27 14:41:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O41A_4%A_79_21# 1 2 3 12 16 20 24 28 32 36 40 42 50
+ 52 56 60 68 75
c126 60 0 8.97448e-20 $X=2.88 $Y=0.72
r127 72 73 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r128 64 65 13.3588 $w=3.79e-07 $l=4.15e-07 $layer=LI1_cond $X=2.43 $Y=0.77
+ $X2=2.43 $Y2=1.185
r129 58 64 2.72394 $w=2.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.665 $Y=0.77
+ $X2=2.43 $Y2=0.77
r130 58 60 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.665 $Y=0.77
+ $X2=2.88 $Y2=0.77
r131 57 65 11.1055 $w=3.79e-07 $l=3.45e-07 $layer=LI1_cond $X=2.43 $Y=1.53
+ $X2=2.43 $Y2=1.185
r132 56 68 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=1.53
+ $X2=3.7 $Y2=1.53
r133 56 57 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.575 $Y=1.53
+ $X2=2.545 $Y2=1.53
r134 52 54 22.3903 $w=3.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.37 $Y=1.66
+ $X2=2.37 $Y2=2.34
r135 50 57 2.82783 $w=3.79e-07 $l=1.11018e-07 $layer=LI1_cond $X=2.37 $Y=1.615
+ $X2=2.43 $Y2=1.53
r136 50 52 1.48171 $w=3.48e-07 $l=4.5e-08 $layer=LI1_cond $X=2.37 $Y=1.615
+ $X2=2.37 $Y2=1.66
r137 49 75 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=1.525 $Y=1.16
+ $X2=1.73 $Y2=1.16
r138 49 73 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=1.525 $Y=1.16
+ $X2=1.31 $Y2=1.16
r139 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.16 $X2=1.525 $Y2=1.16
r140 45 72 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=0.68 $Y=1.16
+ $X2=0.89 $Y2=1.16
r141 45 69 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=0.68 $Y=1.16
+ $X2=0.47 $Y2=1.16
r142 44 48 44.2643 $w=2.18e-07 $l=8.45e-07 $layer=LI1_cond $X=0.68 $Y=1.185
+ $X2=1.525 $Y2=1.185
r143 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=1.16 $X2=0.68 $Y2=1.16
r144 42 65 3.91961 $w=2.2e-07 $l=2.35e-07 $layer=LI1_cond $X=2.195 $Y=1.185
+ $X2=2.43 $Y2=1.185
r145 42 48 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=2.195 $Y=1.185
+ $X2=1.525 $Y2=1.185
r146 38 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r147 38 40 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r148 34 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r149 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r150 30 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r151 30 32 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r152 26 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r153 26 28 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r154 22 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r155 22 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r156 18 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.16
r157 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r158 14 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r159 14 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.985
r160 10 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r161 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
r162 3 68 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=3.605
+ $Y=1.485 $X2=3.74 $Y2=1.61
r163 2 54 400 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.38 $Y2=2.34
r164 2 52 400 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.38 $Y2=1.66
r165 1 60 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%B1 3 5 6 9 13 17 19 26
r51 24 26 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=3 $Y=1.16 $X2=3.09
+ $Y2=1.16
r52 22 24 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.67 $Y=1.16 $X2=3
+ $Y2=1.16
r53 21 22 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=2.59 $Y=1.16 $X2=2.67
+ $Y2=1.16
r54 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=1.16
+ $X2=3 $Y2=1.16
r55 15 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=1.16
r56 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=0.56
r57 11 22 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=1.16
r58 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=0.56
r59 7 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.59 $Y=1.295
+ $X2=2.59 $Y2=1.16
r60 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.59 $Y=1.295 $X2=2.59
+ $Y2=1.985
r61 5 21 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.515 $Y=1.16 $X2=2.59
+ $Y2=1.16
r62 5 6 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.515 $Y=1.16
+ $X2=2.225 $Y2=1.16
r63 1 6 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.225 $Y2=1.16
r64 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295 $X2=2.15
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A4 3 7 11 15 17 18 26
c51 7 0 6.70685e-20 $X=3.53 $Y=1.985
c52 3 0 8.97448e-20 $X=3.53 $Y=0.56
r53 24 26 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=3.74 $Y=1.16
+ $X2=3.95 $Y2=1.16
r54 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.16 $X2=3.74 $Y2=1.16
r55 21 24 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=3.53 $Y=1.16
+ $X2=3.74 $Y2=1.16
r56 18 25 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=3.955 $Y=1.175
+ $X2=3.74 $Y2=1.175
r57 17 25 13.5864 $w=1.98e-07 $l=2.45e-07 $layer=LI1_cond $X=3.495 $Y=1.175
+ $X2=3.74 $Y2=1.175
r58 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.95 $Y=1.295
+ $X2=3.95 $Y2=1.16
r59 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.95 $Y=1.295
+ $X2=3.95 $Y2=1.985
r60 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.95 $Y=1.025
+ $X2=3.95 $Y2=1.16
r61 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.95 $Y=1.025
+ $X2=3.95 $Y2=0.56
r62 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.53 $Y=1.295
+ $X2=3.53 $Y2=1.16
r63 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.53 $Y=1.295 $X2=3.53
+ $Y2=1.985
r64 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.53 $Y=1.025
+ $X2=3.53 $Y2=1.16
r65 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.53 $Y=1.025
+ $X2=3.53 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A3 3 7 11 15 17 18 26
r48 24 26 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.58 $Y=1.16
+ $X2=4.79 $Y2=1.16
r49 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.58
+ $Y=1.16 $X2=4.58 $Y2=1.16
r50 21 24 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.37 $Y=1.16
+ $X2=4.58 $Y2=1.16
r51 18 25 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=4.875 $Y=1.175
+ $X2=4.58 $Y2=1.175
r52 17 25 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=1.175
+ $X2=4.58 $Y2=1.175
r53 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.79 $Y=1.295
+ $X2=4.79 $Y2=1.16
r54 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.79 $Y=1.295
+ $X2=4.79 $Y2=1.985
r55 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.79 $Y=1.025
+ $X2=4.79 $Y2=1.16
r56 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.79 $Y=1.025
+ $X2=4.79 $Y2=0.56
r57 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.37 $Y=1.295
+ $X2=4.37 $Y2=1.16
r58 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.37 $Y=1.295 $X2=4.37
+ $Y2=1.985
r59 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.37 $Y=1.025
+ $X2=4.37 $Y2=1.16
r60 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.37 $Y=1.025
+ $X2=4.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A2 3 7 11 15 17 18 19 20 24 33
c54 33 0 1.92379e-19 $X=6.19 $Y=1.16
c55 17 0 1.14128e-19 $X=5.305 $Y=1.16
r56 31 33 9.99782 $w=2.7e-07 $l=4.5e-08 $layer=POLY_cond $X=6.145 $Y=1.16
+ $X2=6.19 $Y2=1.16
r57 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.145
+ $Y=1.16 $X2=6.145 $Y2=1.16
r58 29 31 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=5.99 $Y=1.16
+ $X2=6.145 $Y2=1.16
r59 28 29 48.8782 $w=2.7e-07 $l=2.2e-07 $layer=POLY_cond $X=5.77 $Y=1.16
+ $X2=5.99 $Y2=1.16
r60 24 28 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.695 $Y=1.16
+ $X2=5.77 $Y2=1.16
r61 24 26 84.426 $w=2.7e-07 $l=3.8e-07 $layer=POLY_cond $X=5.695 $Y=1.16
+ $X2=5.315 $Y2=1.16
r62 20 32 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=6.275 $Y=1.175
+ $X2=6.145 $Y2=1.175
r63 19 32 18.3 $w=1.98e-07 $l=3.3e-07 $layer=LI1_cond $X=5.815 $Y=1.175
+ $X2=6.145 $Y2=1.175
r64 18 19 27.7273 $w=1.98e-07 $l=5e-07 $layer=LI1_cond $X=5.315 $Y=1.175
+ $X2=5.815 $Y2=1.175
r65 18 26 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.315
+ $Y=1.16 $X2=5.315 $Y2=1.16
r66 17 26 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=5.305 $Y=1.16
+ $X2=5.315 $Y2=1.16
r67 13 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.19 $Y=1.295
+ $X2=6.19 $Y2=1.16
r68 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.19 $Y=1.295
+ $X2=6.19 $Y2=1.985
r69 9 29 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.99 $Y=1.025
+ $X2=5.99 $Y2=1.16
r70 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.99 $Y=1.025
+ $X2=5.99 $Y2=0.56
r71 5 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.77 $Y=1.295
+ $X2=5.77 $Y2=1.16
r72 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.77 $Y=1.295 $X2=5.77
+ $Y2=1.985
r73 1 17 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=5.23 $Y=1.025
+ $X2=5.305 $Y2=1.16
r74 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.23 $Y=1.025
+ $X2=5.23 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A1 3 7 11 15 17 21 22 23 28 38
c42 23 0 1.92379e-19 $X=7.55 $Y=1.105
r43 29 38 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=7.315 $Y=1.175
+ $X2=7.615 $Y2=1.175
r44 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.315
+ $Y=1.16 $X2=7.315 $Y2=1.16
r45 23 38 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=7.635 $Y=1.175
+ $X2=7.615 $Y2=1.175
r46 22 29 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=7.195 $Y=1.175
+ $X2=7.315 $Y2=1.175
r47 21 22 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.735 $Y=1.175
+ $X2=7.195 $Y2=1.175
r48 18 20 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.61 $Y=1.16 $X2=7.03
+ $Y2=1.16
r49 17 28 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=7.105 $Y=1.16
+ $X2=7.315 $Y2=1.16
r50 17 20 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=7.105 $Y=1.16
+ $X2=7.03 $Y2=1.16
r51 13 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.03 $Y=1.295
+ $X2=7.03 $Y2=1.16
r52 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.03 $Y=1.295
+ $X2=7.03 $Y2=1.985
r53 9 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.03 $Y=1.025
+ $X2=7.03 $Y2=1.16
r54 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.03 $Y=1.025
+ $X2=7.03 $Y2=0.56
r55 5 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.61 $Y=1.295
+ $X2=6.61 $Y2=1.16
r56 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.61 $Y=1.295 $X2=6.61
+ $Y2=1.985
r57 1 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.61 $Y=1.025
+ $X2=6.61 $Y2=1.16
r58 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.61 $Y=1.025
+ $X2=6.61 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%VPWR 1 2 3 4 5 16 18 22 26 32 36 39 40 42 43
+ 45 46 47 59 65 66 72
r100 72 73 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r101 66 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r102 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r103 63 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.985 $Y=2.72
+ $X2=6.82 $Y2=2.72
r104 63 65 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.985 $Y=2.72
+ $X2=7.59 $Y2=2.72
r105 62 73 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=6.67 $Y2=2.72
r106 61 62 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r107 59 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.655 $Y=2.72
+ $X2=6.82 $Y2=2.72
r108 59 61 239.107 $w=1.68e-07 $l=3.665e-06 $layer=LI1_cond $X=6.655 $Y=2.72
+ $X2=2.99 $Y2=2.72
r109 58 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r110 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r111 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r113 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 49 69 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r116 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 47 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 47 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r119 45 57 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.715 $Y=2.72
+ $X2=2.84 $Y2=2.72
r121 44 61 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=2.99 $Y2=2.72
r122 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=2.84 $Y2=2.72
r123 42 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r124 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.94 $Y2=2.72
r125 41 57 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.53 $Y2=2.72
r126 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.94 $Y2=2.72
r127 39 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r128 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r129 38 54 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r130 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r131 34 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=2.635
+ $X2=6.82 $Y2=2.72
r132 34 36 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=6.82 $Y=2.635
+ $X2=6.82 $Y2=1.95
r133 30 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=2.635
+ $X2=2.84 $Y2=2.72
r134 30 32 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.84 $Y=2.635
+ $X2=2.84 $Y2=2
r135 26 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.94 $Y=1.66
+ $X2=1.94 $Y2=2.34
r136 24 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r137 24 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.34
r138 20 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r139 20 22 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r140 16 69 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r141 16 18 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2
r142 5 36 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=6.685
+ $Y=1.485 $X2=6.82 $Y2=1.95
r143 4 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=2
r144 3 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.34
r145 3 26 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.66
r146 2 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r147 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%X 1 2 3 4 15 19 21 22 23 24 27 29 31 35 36 37
r67 37 59 24.6773 $w=1.98e-07 $l=4.45e-07 $layer=LI1_cond $X=0.235 $Y=1.565
+ $X2=0.68 $Y2=1.565
r68 37 44 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=0.235 $Y=1.565
+ $X2=0.215 $Y2=1.565
r69 37 44 0.443247 $w=2.58e-07 $l=1e-08 $layer=LI1_cond $X=0.215 $Y=1.455
+ $X2=0.215 $Y2=1.465
r70 36 37 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=0.215 $Y=1.19
+ $X2=0.215 $Y2=1.455
r71 35 43 1.16746 $w=1.88e-07 $l=2e-08 $layer=LI1_cond $X=0.235 $Y=0.81
+ $X2=0.215 $Y2=0.81
r72 35 36 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=0.215 $Y=0.92
+ $X2=0.215 $Y2=1.19
r73 35 43 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.215 $Y=0.92
+ $X2=0.215 $Y2=0.905
r74 29 34 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=1.52 $Y=1.665 $X2=1.52
+ $Y2=1.565
r75 29 31 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r76 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=0.715
+ $X2=1.52 $Y2=0.38
r77 24 59 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.565
+ $X2=0.68 $Y2=1.565
r78 23 34 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.565
+ $X2=1.52 $Y2=1.565
r79 23 24 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.565
+ $X2=0.845 $Y2=1.565
r80 21 25 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.355 $Y=0.81
+ $X2=1.52 $Y2=0.715
r81 21 22 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=0.81
+ $X2=0.845 $Y2=0.81
r82 19 59 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=2.34
+ $X2=0.68 $Y2=1.665
r83 13 22 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.81
+ $X2=0.845 $Y2=0.81
r84 13 35 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=0.68 $Y=0.81
+ $X2=0.235 $Y2=0.81
r85 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.715
+ $X2=0.68 $Y2=0.38
r86 4 34 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r87 4 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r88 3 59 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r89 3 19 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r90 2 27 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r91 1 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A_639_297# 1 2 3 12 14 15 16 19 20 27
c49 20 0 1.18248e-19 $X=4.835 $Y=1.53
c50 16 0 6.70685e-20 $X=4.16 $Y=1.615
r51 21 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=1.53
+ $X2=4.16 $Y2=1.53
r52 20 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=1.53 $X2=5
+ $Y2=1.53
r53 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.835 $Y=1.53
+ $X2=4.325 $Y2=1.53
r54 17 19 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=4.16 $Y=2.295
+ $X2=4.16 $Y2=2.29
r55 16 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.615 $X2=4.16
+ $Y2=1.53
r56 16 19 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.16 $Y=1.615
+ $X2=4.16 $Y2=2.29
r57 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.995 $Y=2.38
+ $X2=4.16 $Y2=2.295
r58 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.995 $Y=2.38
+ $X2=3.405 $Y2=2.38
r59 10 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.27 $Y=2.295
+ $X2=3.405 $Y2=2.38
r60 10 12 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.27 $Y=2.295
+ $X2=3.27 $Y2=2
r61 3 27 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5 $Y2=1.61
r62 2 25 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.485 $X2=4.16 $Y2=1.61
r63 2 19 400 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.485 $X2=4.16 $Y2=2.29
r64 1 12 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=3.195
+ $Y=1.485 $X2=3.32 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A_889_297# 1 2 9 11 12 15
r21 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=5.98 $Y=2.295
+ $X2=5.98 $Y2=1.95
r22 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.815 $Y=2.38
+ $X2=5.98 $Y2=2.295
r23 11 12 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=5.815 $Y=2.38
+ $X2=4.665 $Y2=2.38
r24 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.58 $Y=2.295
+ $X2=4.665 $Y2=2.38
r25 7 9 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.58 $Y=2.295 $X2=4.58
+ $Y2=1.95
r26 2 15 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.845
+ $Y=1.485 $X2=5.98 $Y2=1.95
r27 1 9 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.445
+ $Y=1.485 $X2=4.58 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A_1083_297# 1 2 3 12 16 18 20 22 25 27
r40 20 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=1.615 $X2=7.43
+ $Y2=1.53
r41 20 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.43 $Y=1.615
+ $X2=7.43 $Y2=2.29
r42 19 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=1.53 $X2=6.4
+ $Y2=1.53
r43 18 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=1.53
+ $X2=7.43 $Y2=1.53
r44 18 19 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.265 $Y=1.53
+ $X2=6.485 $Y2=1.53
r45 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=1.615 $X2=6.4
+ $Y2=1.53
r46 14 16 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.4 $Y=1.615
+ $X2=6.4 $Y2=2.29
r47 13 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.645 $Y=1.53
+ $X2=5.52 $Y2=1.53
r48 12 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.315 $Y=1.53 $X2=6.4
+ $Y2=1.53
r49 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.315 $Y=1.53
+ $X2=5.645 $Y2=1.53
r50 3 29 400 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=1 $X=7.105
+ $Y=1.485 $X2=7.43 $Y2=1.61
r51 3 22 400 $w=1.7e-07 $l=9.53756e-07 $layer=licon1_PDIFF $count=1 $X=7.105
+ $Y=1.485 $X2=7.43 $Y2=2.29
r52 2 27 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=6.265
+ $Y=1.485 $X2=6.4 $Y2=1.61
r53 2 16 400 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=6.265
+ $Y=1.485 $X2=6.4 $Y2=2.29
r54 1 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.415
+ $Y=1.485 $X2=5.56 $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 47 48
+ 50 51 53 54 56 57 58 64 84 85 91 96 99
r125 98 99 9.78215 $w=6.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.78 $Y=0.23
+ $X2=5.915 $Y2=0.23
r126 94 98 0.569561 $w=6.28e-07 $l=3e-08 $layer=LI1_cond $X=5.75 $Y=0.23
+ $X2=5.78 $Y2=0.23
r127 94 96 15.6676 $w=6.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.75 $Y=0.23
+ $X2=5.305 $Y2=0.23
r128 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r129 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r130 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r131 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r132 82 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=5.75
+ $Y2=0
r133 81 99 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=5.915 $Y2=0
r134 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r135 78 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r136 77 96 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.29 $Y=0 $X2=5.305
+ $Y2=0
r137 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r138 74 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r139 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r140 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r141 71 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.07 $Y2=0
r142 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r143 68 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=1.98
+ $Y2=0
r144 68 70 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=2.105 $Y=0
+ $X2=3.45 $Y2=0
r145 67 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r146 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r147 64 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.98
+ $Y2=0
r148 64 66 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r149 63 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r150 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r151 60 88 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r152 60 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r153 58 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r154 58 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r155 56 81 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.685 $Y=0 $X2=6.67
+ $Y2=0
r156 56 57 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.685 $Y=0 $X2=6.82
+ $Y2=0
r157 55 84 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.955 $Y=0
+ $X2=7.59 $Y2=0
r158 55 57 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.955 $Y=0 $X2=6.82
+ $Y2=0
r159 53 73 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.37
+ $Y2=0
r160 53 54 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.58
+ $Y2=0
r161 52 77 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=5.29 $Y2=0
r162 52 54 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.58
+ $Y2=0
r163 50 70 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.655 $Y=0
+ $X2=3.45 $Y2=0
r164 50 51 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.765
+ $Y2=0
r165 49 73 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.875 $Y=0
+ $X2=4.37 $Y2=0
r166 49 51 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.765
+ $Y2=0
r167 47 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r168 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r169 46 66 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r170 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r171 42 57 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=0.085
+ $X2=6.82 $Y2=0
r172 42 44 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.82 $Y=0.085
+ $X2=6.82 $Y2=0.38
r173 38 54 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r174 38 40 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.38
r175 34 51 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0.085
+ $X2=3.765 $Y2=0
r176 34 36 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.765 $Y=0.085
+ $X2=3.765 $Y2=0.38
r177 30 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r178 30 32 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.38
r179 26 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r180 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r181 22 88 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r182 22 24 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.38
r183 7 44 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.685
+ $Y=0.235 $X2=6.82 $Y2=0.38
r184 6 98 91 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_NDIFF $count=2 $X=5.305
+ $Y=0.235 $X2=5.78 $Y2=0.38
r185 5 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.58 $Y2=0.38
r186 4 36 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.235 $X2=3.74 $Y2=0.38
r187 3 32 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r188 2 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r189 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O41A_4%A_467_47# 1 2 3 4 5 6 19 23 26 27 28 31 33 37
+ 39 43 45 49 53 54 55
c101 39 0 1.14128e-19 $X=6.24 $Y=0.82
c102 33 0 1.18248e-19 $X=4.915 $Y=0.82
r103 47 49 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=7.43 $Y=0.735
+ $X2=7.43 $Y2=0.42
r104 46 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=0.82
+ $X2=6.325 $Y2=0.82
r105 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.265 $Y=0.82
+ $X2=7.43 $Y2=0.735
r106 45 46 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=7.265 $Y=0.82
+ $X2=6.41 $Y2=0.82
r107 41 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=0.735
+ $X2=6.325 $Y2=0.82
r108 41 43 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.325 $Y=0.735
+ $X2=6.325 $Y2=0.42
r109 40 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=0.82 $X2=5
+ $Y2=0.82
r110 39 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=0.82
+ $X2=6.325 $Y2=0.82
r111 39 40 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=6.24 $Y=0.82
+ $X2=5.085 $Y2=0.82
r112 35 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.735 $X2=5
+ $Y2=0.82
r113 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5 $Y=0.735 $X2=5
+ $Y2=0.42
r114 34 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.82
+ $X2=4.16 $Y2=0.82
r115 33 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0.82 $X2=5
+ $Y2=0.82
r116 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.915 $Y=0.82
+ $X2=4.245 $Y2=0.82
r117 29 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=0.735
+ $X2=4.16 $Y2=0.82
r118 29 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.16 $Y=0.735
+ $X2=4.16 $Y2=0.42
r119 27 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=0.82
+ $X2=4.16 $Y2=0.82
r120 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.075 $Y=0.82
+ $X2=3.485 $Y2=0.82
r121 24 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.36 $Y=0.735
+ $X2=3.485 $Y2=0.82
r122 24 26 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.36 $Y=0.735
+ $X2=3.36 $Y2=0.72
r123 23 52 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.36 $Y=0.465
+ $X2=3.36 $Y2=0.36
r124 23 26 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.36 $Y=0.465
+ $X2=3.36 $Y2=0.72
r125 19 52 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=0.36
+ $X2=3.36 $Y2=0.36
r126 19 21 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=3.235 $Y=0.36
+ $X2=2.46 $Y2=0.36
r127 6 49 91 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=2 $X=7.105
+ $Y=0.235 $X2=7.43 $Y2=0.42
r128 5 43 91 $w=1.7e-07 $l=3.40147e-07 $layer=licon1_NDIFF $count=2 $X=6.065
+ $Y=0.235 $X2=6.325 $Y2=0.42
r129 4 37 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.865
+ $Y=0.235 $X2=5 $Y2=0.42
r130 3 31 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.025
+ $Y=0.235 $X2=4.16 $Y2=0.42
r131 2 52 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.32 $Y2=0.38
r132 2 26 182 $w=1.7e-07 $l=5.57136e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.32 $Y2=0.72
r133 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__nor2b_4.spice
* Created: Thu Aug 27 14:31:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor2b_4.spice.pex"
.subckt sky130_fd_sc_hd__nor2b_4  VNB VPB A B_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B_N	B_N
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1002_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1008_d N_A_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1009_s N_A_419_21#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_419_21#_M1010_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1010_d N_A_419_21#_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_A_419_21#_M1016_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B_N_M1003_g N_A_419_21#_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.182 PD=1.84 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1001_d N_A_M1012_g N_A_27_297#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_27_297#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1014_d N_A_M1017_g N_A_27_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_A_27_297#_M1017_s N_A_419_21#_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1006 N_A_27_297#_M1006_d N_A_419_21#_M1006_g N_Y_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1007 N_A_27_297#_M1006_d N_A_419_21#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1015 N_A_27_297#_M1015_d N_A_419_21#_M1015_g N_Y_M1007_s VPB PHIGHVT L=0.15
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_B_N_M1011_g N_A_419_21#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.27 PD=2.56 PS=2.54 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=8.7312 P=14.09
c_46 VNB 0 1.68547e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__nor2b_4.spice.SKY130_FD_SC_HD__NOR2B_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_2.spice
* Created: Tue Sep  1 19:11:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_clkinvkapwr_2.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_2  VNB VPB A Y KAPWR VGND VPWR
* 
* VGND	VGND
* KAPWR	KAPWR
* Y	Y
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1004 N_Y_M1002_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1092 PD=0.7 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1000 N_KAPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1001 N_KAPWR_M1000_d N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MM1003 N_KAPWR_M1003_d N_A_M1003_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX5_noxref VNB VPB NWDIODE A=3.5631 P=7.65
*
.include "sky130_fd_sc_hd__lpflow_clkinvkapwr_2.pxi.spice"
*
.ends
*
*

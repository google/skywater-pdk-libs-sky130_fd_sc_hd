* File: sky130_fd_sc_hd__a22o_1.spice
* Created: Tue Sep  1 18:53:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a22o_1.pex.spice"
.subckt sky130_fd_sc_hd__a22o_1  VNB VPB B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1008 A_109_47# N_B2_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65 AD=0.07475
+ AS=0.169 PD=0.88 PS=1.82 NRD=11.076 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_297#_M1001_d N_B1_M1001_g A_109_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.07475 PD=1.82 PS=0.88 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 A_373_47# N_A1_M1006_g N_A_27_297#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.169 PD=1 PS=1.82 NRD=22.152 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_373_47# VNB NSHORT L=0.15 W=0.65 AD=0.10075
+ AS=0.11375 PD=0.96 PS=1 NRD=6.456 NRS=22.152 M=1 R=4.33333 SA=75000.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_27_297#_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10075 PD=1.82 PS=0.96 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_109_297#_M1004_d N_B2_M1004_g N_A_27_297#_M1004_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_27_297#_M1002_d N_B1_M1002_g N_A_109_297#_M1004_d VPB PHIGHVT L=0.15
+ W=1 AD=0.25285 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_109_297#_M1000_d N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.2529 PD=1.32 PS=2.52 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_109_297#_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.16 PD=1.31 PS=1.32 NRD=6.8753 NRS=6.8753 M=1 R=6.66667
+ SA=75000.6 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1009_d N_A_27_297#_M1009_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.155 PD=2.52 PS=1.31 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a22o_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__macro_sparecell.spice
* Created: Thu Aug 27 14:27:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__macro_sparecell.spice.pex"
.subckt sky130_fd_sc_hd__macro_sparecell  VNB VPB LO VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* LO	LO
* VPB	VPB
* VNB	VNB
MXsky130_fd_sc_hd__inv_2_1/M1001
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1001_g
+ N_VGND_Xsky130_fd_sc_hd__inv_2_1/M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__inv_2_1/M1003
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1003_g
+ N_VGND_Xsky130_fd_sc_hd__inv_2_1/M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1001
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1001_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1001_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.5
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1002
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1001_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1002_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75001
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1003
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1003_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1003_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1004
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1003_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1004_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_1/M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1003
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1003_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1003_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1003_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1004
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1004_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1004_g
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1003_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1002
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1004_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1002_g
+ N_VGND_Xsky130_fd_sc_hd__nand2_2_1/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1007
+ N_XSKY130_FD_SC_HD__NAND2_2_1/A_27_47#_Xsky130_fd_sc_hd__nand2_2_1/M1007_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1007_g
+ N_VGND_Xsky130_fd_sc_hd__nand2_2_1/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1002
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1002_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1002_g
+ N_VGND_Xsky130_fd_sc_hd__nand2_2_0/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.4
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1007
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1007_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1007_g
+ N_VGND_Xsky130_fd_sc_hd__nand2_2_0/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75001
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1003
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1007_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1003_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1003_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1004
+ N_XSKY130_FD_SC_HD__NAND2_2_0/A_27_47#_Xsky130_fd_sc_hd__nand2_2_0/M1004_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1004_g
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1003_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1001
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1001_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1001_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.4
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1002
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1001_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1002_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75001
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1003
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1003_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1003_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1004
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1003_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1004_g
+ N_VGND_Xsky130_fd_sc_hd__nor2_2_0/M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__inv_2_0/M1001
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1001_g
+ N_VGND_Xsky130_fd_sc_hd__inv_2_0/M1001_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__inv_2_0/M1003
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1001_d
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1003_g
+ N_VGND_Xsky130_fd_sc_hd__inv_2_0/M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MXsky130_fd_sc_hd__inv_2_1/M1000 N_VPWR_Xsky130_fd_sc_hd__inv_2_1/M1000_d
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__inv_2_1/M1002 N_VPWR_Xsky130_fd_sc_hd__inv_2_1/M1002_d
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__inv_2_1/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_1/Y_Xsky130_fd_sc_hd__inv_2_1/M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1005
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1005_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1005_g
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1006
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1006_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1006_g
+ N_SKY130_FD_SC_HD__INV_2_1/A_Xsky130_fd_sc_hd__nor2_2_1/M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1000 N_VPWR_Xsky130_fd_sc_hd__nor2_2_1/M1000_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1000_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1006_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75000.6 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_1/M1007 N_VPWR_Xsky130_fd_sc_hd__nor2_2_1/M1000_d
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nor2_2_1/M1007_g
+ N_XSKY130_FD_SC_HD__NOR2_2_1/A_27_297#_Xsky130_fd_sc_hd__nor2_2_1/M1007_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1000
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1000_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1000_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.4 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1001
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1000_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1001_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1005
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1005_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1005_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_1/M1006
+ N_SKY130_FD_SC_HD__NOR2_2_1/B_Xsky130_fd_sc_hd__nand2_2_1/M1005_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_1/M1006_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_1/M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75000.2 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1000
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1000_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1000_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.4 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1001
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1000_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1001_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1005
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1005_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1005_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nand2_2_0/M1006
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nand2_2_0/M1005_d
+ N_LO_Xsky130_fd_sc_hd__nand2_2_0/M1006_g
+ N_VPWR_Xsky130_fd_sc_hd__nand2_2_0/M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75000.2 A=0.15
+ P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1000 N_VPWR_Xsky130_fd_sc_hd__nor2_2_0/M1000_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1000_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1000_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1007 N_VPWR_Xsky130_fd_sc_hd__nor2_2_0/M1000_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1007_g
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1007_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1005
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1007_s
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75000.6 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__nor2_2_0/M1006
+ N_XSKY130_FD_SC_HD__NOR2_2_0/A_27_297#_Xsky130_fd_sc_hd__nor2_2_0/M1006_d
+ N_SKY130_FD_SC_HD__NOR2_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1006_g
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__nor2_2_0/M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__inv_2_0/M1000 N_VPWR_Xsky130_fd_sc_hd__inv_2_0/M1000_d
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1000_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MXsky130_fd_sc_hd__inv_2_0/M1002 N_VPWR_Xsky130_fd_sc_hd__inv_2_0/M1002_d
+ N_SKY130_FD_SC_HD__INV_2_0/A_Xsky130_fd_sc_hd__inv_2_0/M1002_g
+ N_SKY130_FD_SC_HD__INV_2_0/Y_Xsky130_fd_sc_hd__inv_2_0/M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=22.0206 P=30.65
rXsky130_fd_sc_hd__conb_1_0/R1 SKY130_FD_SC_HD__CONB_1_0/HI
+ N_VPWR_Xsky130_fd_sc_hd__conb_1_0/R1_neg SHORT 0.01 M=1
rXsky130_fd_sc_hd__conb_1_0/R0 N_VGND_Xsky130_fd_sc_hd__conb_1_0/R0_pos
+ N_LO_Xsky130_fd_sc_hd__conb_1_0/R0_neg SHORT 0.01 M=1
c_130 VNB 0 1.32973e-19 $X=0.145 $Y=-0.085
c_238 VPB 0 3.3186e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__macro_sparecell.spice.SKY130_FD_SC_HD__MACRO_SPARECELL.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_1.pxi.spice
* Created: Thu Aug 27 14:23:54 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%A N_A_M1000_g N_A_M1002_g N_A_M1001_g
+ A A A N_A_c_24_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%KAPWR N_KAPWR_M1000_d N_KAPWR_M1001_d
+ N_KAPWR_c_53_n N_KAPWR_c_54_n KAPWR N_KAPWR_c_55_n N_KAPWR_c_56_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%Y N_Y_M1002_s N_Y_M1000_s N_Y_c_78_n
+ N_Y_c_80_n Y Y PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%Y
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%VGND N_VGND_M1002_d N_VGND_c_105_n
+ N_VGND_c_106_n VGND N_VGND_c_107_n N_VGND_c_108_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%VPWR VPWR N_VPWR_c_121_n
+ N_VPWR_c_120_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_1%VPWR
cc_1 VNB N_A_M1002_g 0.0411839f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=0.445
cc_2 VNB A 0.0444627f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_3 VNB N_A_c_24_n 0.0756236f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_4 VNB N_Y_c_78_n 0.00128525f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.345
cc_5 VNB Y 0.0346199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_VGND_c_105_n 0.0103648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_VGND_c_106_n 0.0193127f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=0.445
cc_8 VNB N_VGND_c_107_n 0.0294553f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=2.065
cc_9 VNB N_VGND_c_108_n 0.114657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VPWR_c_120_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.345
cc_11 VPB N_A_M1000_g 0.037104f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.065
cc_12 VPB N_A_M1001_g 0.037104f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=2.065
cc_13 VPB A 0.00366f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.425
cc_14 VPB N_A_c_24_n 0.0176333f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.16
cc_15 VPB N_KAPWR_c_53_n 0.00876329f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=0.445
cc_16 VPB N_KAPWR_c_54_n 0.00876329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_17 VPB N_KAPWR_c_55_n 0.0273169f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_18 VPB N_KAPWR_c_56_n 0.0276178f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_19 VPB N_Y_c_80_n 0.00609894f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.425
cc_20 VPB N_VPWR_c_121_n 0.039878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_120_n 0.0418774f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.345
cc_22 N_A_M1000_g N_KAPWR_c_53_n 0.00580645f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_23 N_A_M1001_g N_KAPWR_c_53_n 0.00580645f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_24 N_A_M1000_g N_KAPWR_c_55_n 0.0118305f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_25 A N_KAPWR_c_55_n 0.0123519f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_26 N_A_c_24_n N_KAPWR_c_55_n 0.00307083f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_27 N_A_M1001_g N_KAPWR_c_56_n 0.0110392f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_28 N_A_M1002_g N_Y_c_78_n 0.0135245f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_29 A N_Y_c_78_n 0.0220349f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_30 N_A_M1000_g N_Y_c_80_n 0.00771009f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_31 N_A_M1001_g N_Y_c_80_n 0.00771009f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_32 A N_Y_c_80_n 0.00166044f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_33 N_A_c_24_n N_Y_c_80_n 0.00655811f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_34 N_A_M1002_g Y 0.0145962f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_35 A Y 0.0307235f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_36 N_A_c_24_n Y 0.0382611f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_37 N_A_M1002_g N_VGND_c_106_n 0.00453359f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_38 N_A_M1002_g N_VGND_c_107_n 0.00426974f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_39 A N_VGND_c_107_n 0.00966373f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_40 N_A_M1002_g N_VGND_c_108_n 0.00816786f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_41 A N_VGND_c_108_n 0.00857725f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_42 N_A_M1000_g N_VPWR_c_121_n 0.00541359f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_43 N_A_M1001_g N_VPWR_c_121_n 0.00541359f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_44 N_A_M1000_g N_VPWR_c_120_n 0.00600702f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_45 N_A_M1001_g N_VPWR_c_120_n 0.0060257f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_46 N_KAPWR_c_53_n N_Y_M1000_s 0.00424434f $X=0.995 $Y=2.24 $X2=0 $Y2=0
cc_47 N_KAPWR_c_53_n N_Y_c_80_n 0.018737f $X=0.995 $Y=2.24 $X2=0 $Y2=0
cc_48 N_KAPWR_c_54_n N_Y_c_80_n 4.06353e-19 $X=0.385 $Y=2.24 $X2=0 $Y2=0
cc_49 N_KAPWR_c_55_n N_Y_c_80_n 0.0325469f $X=0.26 $Y=1.83 $X2=0 $Y2=0
cc_50 N_KAPWR_c_56_n N_Y_c_80_n 0.0327379f $X=1.1 $Y=1.83 $X2=0 $Y2=0
cc_51 N_KAPWR_c_56_n Y 0.0167148f $X=1.1 $Y=1.83 $X2=0 $Y2=0
cc_52 N_KAPWR_c_53_n N_VPWR_c_121_n 0.00217232f $X=0.995 $Y=2.24 $X2=0 $Y2=0
cc_53 N_KAPWR_c_54_n N_VPWR_c_121_n 3.1468e-19 $X=0.385 $Y=2.24 $X2=0 $Y2=0
cc_54 N_KAPWR_c_55_n N_VPWR_c_121_n 0.0217551f $X=0.26 $Y=1.83 $X2=0 $Y2=0
cc_55 N_KAPWR_c_56_n N_VPWR_c_121_n 0.0231615f $X=1.1 $Y=1.83 $X2=0 $Y2=0
cc_56 N_KAPWR_M1000_d N_VPWR_c_120_n 0.0010704f $X=0.135 $Y=1.645 $X2=0 $Y2=0
cc_57 N_KAPWR_M1001_d N_VPWR_c_120_n 0.00115538f $X=0.965 $Y=1.645 $X2=0 $Y2=0
cc_58 N_KAPWR_c_54_n N_VPWR_c_120_n 0.127401f $X=0.385 $Y=2.24 $X2=0 $Y2=0
cc_59 N_KAPWR_c_55_n N_VPWR_c_120_n 0.00308845f $X=0.26 $Y=1.83 $X2=0 $Y2=0
cc_60 N_KAPWR_c_56_n N_VPWR_c_120_n 0.00327408f $X=1.1 $Y=1.83 $X2=0 $Y2=0
cc_61 Y N_VGND_c_106_n 0.0245139f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_62 N_Y_c_78_n N_VGND_c_107_n 0.0153589f $X=0.675 $Y=0.435 $X2=0 $Y2=0
cc_63 Y N_VGND_c_107_n 0.00239287f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_64 N_Y_M1002_s N_VGND_c_108_n 0.00351653f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_65 N_Y_c_78_n N_VGND_c_108_n 0.00934584f $X=0.675 $Y=0.435 $X2=0 $Y2=0
cc_66 Y N_VGND_c_108_n 0.00508538f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_67 N_Y_c_80_n N_VPWR_c_121_n 0.0113958f $X=0.68 $Y=1.83 $X2=0 $Y2=0
cc_68 N_Y_M1000_s N_VPWR_c_120_n 0.00149677f $X=0.545 $Y=1.645 $X2=0 $Y2=0
cc_69 N_Y_c_80_n N_VPWR_c_120_n 0.00155926f $X=0.68 $Y=1.83 $X2=0 $Y2=0

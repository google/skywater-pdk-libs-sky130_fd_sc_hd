* File: sky130_fd_sc_hd__a211oi_4.spice
* Created: Thu Aug 27 13:59:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a211oi_4.pex.spice"
.subckt sky130_fd_sc_hd__a211oi_4  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_109_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75006.6 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A2_M1018_g N_A_109_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75006.2 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1018_d N_A2_M1025_g N_A_109_47#_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75005.8 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_A1_M1013_g N_A_109_47#_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1013_d N_A1_M1014_g N_A_109_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1020_d N_A1_M1020_g N_A_109_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1024 N_Y_M1020_d N_A1_M1024_g N_A_109_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1030 N_VGND_M1030_d N_A2_M1030_g N_A_109_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.08775 PD=0.985 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1002_d N_B1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.091 PD=0.985 PS=0.93 NRD=7.38 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1023_d N_B1_M1023_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.091 PD=0.925 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1023_d N_C1_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.08775 PD=0.925 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1021 N_Y_M1021_d N_C1_M1021_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1027 N_Y_M1021_d N_C1_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1031 N_Y_M1031_d N_C1_M1031_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.08775 PD=0.93 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75006.1 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1026 N_Y_M1031_d N_B1_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.1885 PD=0.93 PS=1.88 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75006.6 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM16_noxref N_VPWR_M16_noxref_d N_A2_M16_noxref_g N_noxref_7_M16_noxref_s VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75006.6 A=0.15 P=2.3 MULT=1
MM17_noxref N_noxref_7_M17_noxref_d N_A2_M17_noxref_g N_VPWR_M16_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75006.2 A=0.15 P=2.3 MULT=1
MM18_noxref N_VPWR_M18_noxref_d N_A2_M18_noxref_g N_noxref_7_M17_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75005.8 A=0.15 P=2.3 MULT=1
MM19_noxref N_noxref_7_M19_noxref_d N_A1_M19_noxref_g N_VPWR_M18_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.4 SB=75005.3 A=0.15 P=2.3 MULT=1
MM20_noxref N_VPWR_M20_noxref_d N_A1_M20_noxref_g N_noxref_7_M19_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75004.9 A=0.15 P=2.3 MULT=1
MM21_noxref N_noxref_7_M21_noxref_d N_A1_M21_noxref_g N_VPWR_M20_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75004.5 A=0.15 P=2.3 MULT=1
MM22_noxref N_VPWR_M22_noxref_d N_A1_M22_noxref_g N_noxref_7_M21_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.7 SB=75004.1 A=0.15 P=2.3 MULT=1
MM23_noxref N_noxref_7_M23_noxref_d N_A2_M23_noxref_g N_VPWR_M22_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.1 SB=75003.7 A=0.15 P=2.3 MULT=1
MM24_noxref N_noxref_9_M24_noxref_d N_B1_M24_noxref_g N_noxref_7_M23_noxref_d
+ VPB PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1
+ R=6.66667 SA=75003.5 SB=75003.2 A=0.15 P=2.3 MULT=1
MM25_noxref N_noxref_7_M25_noxref_d N_B1_M25_noxref_g N_noxref_9_M24_noxref_d
+ VPB PHIGHVT L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1
+ R=6.66667 SA=75004 SB=75002.8 A=0.15 P=2.3 MULT=1
MM26_noxref noxref_10 N_B1_M26_noxref_g N_noxref_7_M25_noxref_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.135 PD=1.3 PS=1.27 NRD=18.6953 NRS=0 M=1 R=6.66667
+ SA=75004.4 SB=75002.4 A=0.15 P=2.3 MULT=1
MM27_noxref N_Y_M27_noxref_d N_C1_M27_noxref_g noxref_10 VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=18.6953 M=1 R=6.66667 SA=75004.8
+ SB=75002 A=0.15 P=2.3 MULT=1
MM28_noxref N_noxref_9_M28_noxref_d N_C1_M28_noxref_g N_Y_M27_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75005.3 SB=75001.5 A=0.15 P=2.3 MULT=1
MM29_noxref N_Y_M29_noxref_d N_C1_M29_noxref_g N_noxref_9_M28_noxref_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=3.9203 NRS=0 M=1
+ R=6.66667 SA=75005.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM30_noxref noxref_12 N_C1_M30_noxref_g N_Y_M29_noxref_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.15 PD=1.31 PS=1.3 NRD=19.6803 NRS=0 M=1 R=6.66667 SA=75006.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM31_noxref N_noxref_7_M31_noxref_d N_B1_M31_noxref_g noxref_12 VPB PHIGHVT
+ L=0.15 W=1 AD=0.26 AS=0.155 PD=2.52 PS=1.31 NRD=0 NRS=19.6803 M=1 R=6.66667
+ SA=75006.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=12.4227 P=18.69
*
.include "sky130_fd_sc_hd__a211oi_4.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_204_309# VPB phighvt w=940000u l=150000u
+  ad=1.3263e+12p pd=1.231e+07u as=2.3452e+12p ps=2.234e+07u
M1001 Z A a_204_309# VPB phighvt w=1e+06u l=150000u
+  ad=1.08e+12p pd=1.016e+07u as=0p ps=0u
M1002 a_215_47# A Z VNB nshort w=650000u l=150000u
+  ad=1.61525e+12p pd=1.667e+07u as=7.02e+11p ps=7.36e+06u
M1003 Z A a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Z A a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_204_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_204_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z A a_204_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_215_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.71e+11p ps=9.18e+06u
M1009 VGND a_27_47# a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR TE_B a_204_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_215_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_47# a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR TE_B a_204_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_27_47# a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_215_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_204_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_27_47# a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_215_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_204_309# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_204_309# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_215_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Z A a_204_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR TE_B a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1024 a_204_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Z A a_204_309# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_204_309# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_215_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR TE_B a_204_309# VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_204_309# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND TE_B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1031 Z A a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_215_47# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Z A a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

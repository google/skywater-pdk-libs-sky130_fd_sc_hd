* NGSPICE file created from sky130_fd_sc_hd__and2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
M1000 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.7e+11p pd=5.14e+06u as=1.2115e+12p ps=1.051e+07u
M1001 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_33_199# A_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=3.64e+11p pd=3.72e+06u as=6.685e+11p ps=6.01e+06u
M1004 a_33_199# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 VPWR a_27_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# a_33_199# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.43e+11p ps=1.74e+06u
M1012 a_109_47# a_33_199# a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1013 VPWR a_27_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__o21a_1.spice
* Created: Thu Aug 27 14:35:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21a_1.pex.spice"
.subckt sky130_fd_sc_hd__o21a_1  VNB VPB B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_79_21#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_297_47#_M1001_d N_B1_M1001_g N_A_79_21#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10075 AS=0.169 PD=0.96 PS=1.82 NRD=6.456 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_297_47#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10075 PD=0.92 PS=0.96 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1003 N_A_297_47#_M1003_d N_A1_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_79_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3275 AS=0.28 PD=1.655 PS=2.56 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1002 N_A_79_21#_M1002_d N_B1_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.3275 PD=1.39 PS=1.655 NRD=13.7703 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1004 A_382_297# N_A2_M1004_g N_A_79_21#_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.195 PD=1.305 PS=1.39 NRD=19.1878 NRS=7.8603 M=1 R=6.66667
+ SA=75001.5 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_382_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.1525 PD=2.52 PS=1.305 NRD=0 NRS=19.1878 M=1 R=6.66667 SA=75002 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
c_51 VPB 0 5.84632e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__o21a_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__maj3_2.pex.spice
* Created: Tue Sep  1 19:14:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MAJ3_2%C 3 7 11 15 18 20 21 22 28 29 33 40 46 48
c85 33 0 1.13272e-19 $X=2.58 $Y=1.52
r86 40 48 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=2.54 $Y=1.54 $X2=2.53
+ $Y2=1.54
r87 33 36 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.58 $Y=1.52
+ $X2=2.58 $Y2=1.655
r88 33 35 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.58 $Y=1.52
+ $X2=2.58 $Y2=1.385
r89 28 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r90 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r91 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r92 21 48 1.75171 $w=2.48e-07 $l=3.8e-08 $layer=LI1_cond $X=2.492 $Y=1.54
+ $X2=2.53 $Y2=1.54
r93 21 46 4.73668 $w=2.48e-07 $l=7.7e-08 $layer=LI1_cond $X=2.492 $Y=1.54
+ $X2=2.415 $Y2=1.54
r94 21 22 18.8079 $w=2.48e-07 $l=4.08e-07 $layer=LI1_cond $X=2.577 $Y=1.54
+ $X2=2.985 $Y2=1.54
r95 21 40 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=2.577 $Y=1.54
+ $X2=2.54 $Y2=1.54
r96 21 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.52 $X2=2.58 $Y2=1.52
r97 20 29 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.6 $Y=1.19 $X2=0.6
+ $Y2=1.16
r98 19 20 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.6 $Y=1.495
+ $X2=0.6 $Y2=1.19
r99 18 19 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.775 $Y=1.58
+ $X2=0.6 $Y2=1.495
r100 18 46 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=0.775 $Y=1.58
+ $X2=2.415 $Y2=1.58
r101 15 36 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.49 $Y=2.165
+ $X2=2.49 $Y2=1.655
r102 11 35 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.49 $Y=0.445 $X2=2.49
+ $Y2=1.385
r103 7 31 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.57 $Y=2.165
+ $X2=0.57 $Y2=1.325
r104 3 30 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.57 $Y=0.445
+ $X2=0.57 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_2%A 3 7 11 15 17 18 26
c45 26 0 1.85037e-19 $X=1.35 $Y=1.16
r46 24 26 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.14 $Y=1.16
+ $X2=1.35 $Y2=1.16
r47 21 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.93 $Y=1.16
+ $X2=1.14 $Y2=1.16
r48 17 18 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.14 $Y=1.16
+ $X2=1.61 $Y2=1.16
r49 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.16 $X2=1.14 $Y2=1.16
r50 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=1.16
r51 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=2.165
r52 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=1.16
r53 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.35 $Y=0.995
+ $X2=1.35 $Y2=0.445
r54 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.16
r55 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.93 $Y=1.325 $X2=0.93
+ $Y2=2.165
r56 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.16
r57 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.93 $Y=0.995 $X2=0.93
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_2%B 3 7 11 15 17 24
c43 17 0 1.85037e-19 $X=2.07 $Y=1.19
r44 22 24 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.95 $Y=1.16 $X2=2.13
+ $Y2=1.16
r45 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.16 $X2=1.95 $Y2=1.16
r46 19 22 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.71 $Y=1.16
+ $X2=1.95 $Y2=1.16
r47 17 23 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.07 $Y=1.16 $X2=1.95
+ $Y2=1.16
r48 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.325
+ $X2=2.13 $Y2=1.16
r49 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.13 $Y=1.325
+ $X2=2.13 $Y2=2.165
r50 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=0.995
+ $X2=2.13 $Y2=1.16
r51 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.13 $Y=0.995
+ $X2=2.13 $Y2=0.445
r52 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.325
+ $X2=1.71 $Y2=1.16
r53 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.71 $Y=1.325 $X2=1.71
+ $Y2=2.165
r54 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=0.995
+ $X2=1.71 $Y2=1.16
r55 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.71 $Y=0.995 $X2=1.71
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_2%A_47_47# 1 2 3 4 15 19 23 27 31 33 37 41 44
+ 46 50 51 55 57 61 67
c141 67 0 6.84111e-20 $X=3.66 $Y=1.16
r142 66 67 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.24 $Y=1.16
+ $X2=3.66 $Y2=1.16
r143 62 66 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=3.11 $Y=1.16
+ $X2=3.24 $Y2=1.16
r144 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.16 $X2=3.11 $Y2=1.16
r145 58 61 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.015 $Y=1.16
+ $X2=3.11 $Y2=1.16
r146 50 53 1.8054 $w=5.28e-07 $l=8e-08 $layer=LI1_cond $X=0.35 $Y=1.92 $X2=0.35
+ $Y2=2
r147 50 51 7.89897 $w=5.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.92
+ $X2=0.35 $Y2=1.835
r148 49 51 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.835
r149 48 49 6.73996 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=0.74
+ $X2=0.305 $Y2=0.825
r150 46 48 7.72661 $w=4.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.305 $Y=0.445
+ $X2=0.305 $Y2=0.74
r151 44 58 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=1.075
+ $X2=3.015 $Y2=1.16
r152 43 44 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=3.015 $Y=0.825
+ $X2=3.015 $Y2=1.075
r153 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=0.74
+ $X2=1.92 $Y2=0.74
r154 41 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.925 $Y=0.74
+ $X2=3.015 $Y2=0.825
r155 41 42 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.925 $Y=0.74
+ $X2=2.085 $Y2=0.74
r156 35 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=0.655
+ $X2=1.92 $Y2=0.74
r157 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.92 $Y=0.655
+ $X2=1.92 $Y2=0.36
r158 34 50 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=0.615 $Y=1.92
+ $X2=0.35 $Y2=1.92
r159 33 57 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=1.92
+ $X2=1.92 $Y2=1.92
r160 33 34 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=1.755 $Y=1.92
+ $X2=0.615 $Y2=1.92
r161 32 48 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=0.74
+ $X2=0.305 $Y2=0.74
r162 31 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=0.74
+ $X2=1.92 $Y2=0.74
r163 31 32 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=1.755 $Y=0.74
+ $X2=0.525 $Y2=0.74
r164 25 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.66 $Y=1.295
+ $X2=3.66 $Y2=1.16
r165 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.66 $Y=1.295
+ $X2=3.66 $Y2=1.985
r166 21 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.66 $Y=1.025
+ $X2=3.66 $Y2=1.16
r167 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.66 $Y=1.025
+ $X2=3.66 $Y2=0.56
r168 17 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.24 $Y=1.295
+ $X2=3.24 $Y2=1.16
r169 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.24 $Y=1.295
+ $X2=3.24 $Y2=1.985
r170 13 66 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.24 $Y=1.025
+ $X2=3.24 $Y2=1.16
r171 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.24 $Y=1.025
+ $X2=3.24 $Y2=0.56
r172 4 57 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.785
+ $Y=1.845 $X2=1.92 $Y2=2
r173 3 53 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.235
+ $Y=1.845 $X2=0.36 $Y2=2
r174 2 37 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.235 $X2=1.92 $Y2=0.36
r175 1 46 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.235 $X2=0.36 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_2%VPWR 1 2 3 12 16 18 20 25 26 27 29 41 46 50
r60 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r64 41 49 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.962 $Y2=2.72
r65 41 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 40 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r68 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 36 39 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.14 $Y2=2.72
r73 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 32 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=1.14 $Y2=2.72
r77 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 27 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 25 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.535 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 25 26 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.535 $Y=2.72
+ $X2=2.697 $Y2=2.72
r81 24 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.86 $Y=2.72 $X2=3.45
+ $Y2=2.72
r82 24 26 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=2.86 $Y=2.72
+ $X2=2.697 $Y2=2.72
r83 20 23 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.92 $Y=1.66
+ $X2=3.92 $Y2=2.34
r84 18 49 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.962 $Y2=2.72
r85 18 23 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.92 $Y2=2.34
r86 14 26 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.697 $Y=2.635
+ $X2=2.697 $Y2=2.72
r87 14 16 22.517 $w=3.23e-07 $l=6.35e-07 $layer=LI1_cond $X=2.697 $Y=2.635
+ $X2=2.697 $Y2=2
r88 10 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.72
r89 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.34
r90 3 23 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.735
+ $Y=1.485 $X2=3.87 $Y2=2.34
r91 3 20 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.735
+ $Y=1.485 $X2=3.87 $Y2=1.66
r92 2 16 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.565
+ $Y=1.845 $X2=2.7 $Y2=2
r93 1 12 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.845 $X2=1.14 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_2%X 1 2 9 11 16 17 18 21
c33 9 0 1.13272e-19 $X=3.45 $Y=1.66
r34 18 21 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.45 $Y=0.51
+ $X2=3.45 $Y2=0.4
r35 16 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.53 $Y=0.905
+ $X2=3.53 $Y2=1.495
r36 15 18 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.45 $Y=0.74
+ $X2=3.45 $Y2=0.51
r37 15 16 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=0.74
+ $X2=3.45 $Y2=0.905
r38 9 17 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=1.66
+ $X2=3.45 $Y2=1.495
r39 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.45 $Y=1.66 $X2=3.45
+ $Y2=2.34
r40 2 11 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.485 $X2=3.45 $Y2=2.34
r41 2 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.485 $X2=3.45 $Y2=1.66
r42 1 21 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.315
+ $Y=0.235 $X2=3.45 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_2%VGND 1 2 3 12 16 18 20 23 24 25 27 39 44 48
c61 16 0 6.84111e-20 $X=2.8 $Y=0.38
r62 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r63 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r64 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r65 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r66 39 47 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.962
+ $Y2=0
r67 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.45
+ $Y2=0
r68 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r69 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r70 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r71 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r72 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r73 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r75 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.61
+ $Y2=0
r76 30 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r77 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r78 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r79 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.69
+ $Y2=0
r80 25 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r81 23 37 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.53
+ $Y2=0
r82 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.8
+ $Y2=0
r83 22 41 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=3.45
+ $Y2=0
r84 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.8
+ $Y2=0
r85 18 47 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.92 $Y=0.085
+ $X2=3.962 $Y2=0
r86 18 20 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.92 $Y=0.085
+ $X2=3.92 $Y2=0.4
r87 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r88 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.38
r89 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r90 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.36
r91 3 20 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.735
+ $Y=0.235 $X2=3.87 $Y2=0.4
r92 2 16 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.235 $X2=2.8 $Y2=0.38
r93 1 12 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.14 $Y2=0.36
.ends


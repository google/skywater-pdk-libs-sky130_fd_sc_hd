* File: sky130_fd_sc_hd__dlxtp_1.pxi.spice
* Created: Tue Sep  1 19:06:25 2020
* 
x_PM_SKY130_FD_SC_HD__DLXTP_1%GATE N_GATE_c_132_n N_GATE_c_127_n N_GATE_M1016_g
+ N_GATE_c_133_n N_GATE_M1011_g N_GATE_c_128_n N_GATE_c_134_n GATE GATE
+ N_GATE_c_130_n N_GATE_c_131_n PM_SKY130_FD_SC_HD__DLXTP_1%GATE
x_PM_SKY130_FD_SC_HD__DLXTP_1%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1012_g N_A_27_47#_M1000_g N_A_27_47#_M1004_g N_A_27_47#_c_171_n
+ N_A_27_47#_c_172_n N_A_27_47#_M1007_g N_A_27_47#_c_183_n N_A_27_47#_c_307_p
+ N_A_27_47#_c_174_n N_A_27_47#_c_175_n N_A_27_47#_c_184_n N_A_27_47#_c_185_n
+ N_A_27_47#_c_176_n N_A_27_47#_c_177_n N_A_27_47#_c_187_n N_A_27_47#_c_188_n
+ N_A_27_47#_c_189_n N_A_27_47#_c_190_n N_A_27_47#_c_191_n N_A_27_47#_c_192_n
+ N_A_27_47#_c_178_n PM_SKY130_FD_SC_HD__DLXTP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLXTP_1%D N_D_M1005_g N_D_M1014_g D N_D_c_318_n
+ N_D_c_319_n PM_SKY130_FD_SC_HD__DLXTP_1%D
x_PM_SKY130_FD_SC_HD__DLXTP_1%A_299_47# N_A_299_47#_M1005_s N_A_299_47#_M1014_s
+ N_A_299_47#_M1010_g N_A_299_47#_M1013_g N_A_299_47#_c_364_n
+ N_A_299_47#_c_357_n N_A_299_47#_c_365_n N_A_299_47#_c_366_n
+ N_A_299_47#_c_358_n N_A_299_47#_c_359_n N_A_299_47#_c_360_n
+ N_A_299_47#_c_361_n N_A_299_47#_c_362_n PM_SKY130_FD_SC_HD__DLXTP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__DLXTP_1%A_193_47# N_A_193_47#_M1012_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1015_g N_A_193_47#_M1002_g N_A_193_47#_c_439_n
+ N_A_193_47#_c_446_n N_A_193_47#_c_440_n N_A_193_47#_c_441_n
+ N_A_193_47#_c_447_n N_A_193_47#_c_448_n N_A_193_47#_c_449_n
+ N_A_193_47#_c_450_n N_A_193_47#_c_442_n N_A_193_47#_c_451_n
+ N_A_193_47#_c_452_n N_A_193_47#_c_443_n PM_SKY130_FD_SC_HD__DLXTP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLXTP_1%A_713_21# N_A_713_21#_M1008_s N_A_713_21#_M1001_s
+ N_A_713_21#_M1006_g N_A_713_21#_M1009_g N_A_713_21#_M1017_g
+ N_A_713_21#_M1003_g N_A_713_21#_c_571_n N_A_713_21#_c_572_n
+ N_A_713_21#_c_611_p N_A_713_21#_c_564_n N_A_713_21#_c_573_n
+ N_A_713_21#_c_565_n N_A_713_21#_c_566_n N_A_713_21#_c_591_p
+ N_A_713_21#_c_587_p N_A_713_21#_c_593_p N_A_713_21#_c_567_n
+ PM_SKY130_FD_SC_HD__DLXTP_1%A_713_21#
x_PM_SKY130_FD_SC_HD__DLXTP_1%A_560_47# N_A_560_47#_M1015_d N_A_560_47#_M1004_d
+ N_A_560_47#_c_640_n N_A_560_47#_M1008_g N_A_560_47#_M1001_g
+ N_A_560_47#_c_641_n N_A_560_47#_c_642_n N_A_560_47#_c_651_n
+ N_A_560_47#_c_652_n N_A_560_47#_c_643_n N_A_560_47#_c_649_n
+ N_A_560_47#_c_644_n N_A_560_47#_c_645_n PM_SKY130_FD_SC_HD__DLXTP_1%A_560_47#
x_PM_SKY130_FD_SC_HD__DLXTP_1%VPWR N_VPWR_M1011_d N_VPWR_M1014_d N_VPWR_M1009_d
+ N_VPWR_M1001_d N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_726_n N_VPWR_c_727_n
+ N_VPWR_c_728_n N_VPWR_c_729_n N_VPWR_c_730_n N_VPWR_c_731_n VPWR
+ N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_723_n N_VPWR_c_736_n
+ N_VPWR_c_737_n PM_SKY130_FD_SC_HD__DLXTP_1%VPWR
x_PM_SKY130_FD_SC_HD__DLXTP_1%Q N_Q_M1017_d N_Q_M1003_d Q Q Q Q N_Q_c_816_n
+ PM_SKY130_FD_SC_HD__DLXTP_1%Q
x_PM_SKY130_FD_SC_HD__DLXTP_1%VGND N_VGND_M1016_d N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_M1008_d N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n
+ N_VGND_c_834_n N_VGND_c_835_n VGND N_VGND_c_836_n N_VGND_c_837_n
+ N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n
+ N_VGND_c_843_n PM_SKY130_FD_SC_HD__DLXTP_1%VGND
cc_1 VNB N_GATE_c_127_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_c_128_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE 0.0153903f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_c_130_n 0.0210048f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_c_131_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1012_g 0.0397896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_171_n 0.0132134f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_c_172_n 0.00481939f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_9 VNB N_A_27_47#_M1007_g 0.0454581f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_10 VNB N_A_27_47#_c_174_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_175_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_176_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_177_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_178_n 0.0230671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_D_M1005_g 0.025905f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_16 VNB N_D_M1014_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_17 VNB N_D_c_318_n 0.00407935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_18 VNB N_D_c_319_n 0.0421785f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_19 VNB N_A_299_47#_M1013_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_299_47#_c_357_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_299_47#_c_358_n 0.00497129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_359_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_23 VNB N_A_299_47#_c_360_n 0.00265154f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_24 VNB N_A_299_47#_c_361_n 0.0272829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_299_47#_c_362_n 0.0166781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_c_439_n 0.0140955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_440_n 0.0280162f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_28 VNB N_A_193_47#_c_441_n 0.00381134f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_29 VNB N_A_193_47#_c_442_n 0.0176526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_443_n 0.00466868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_713_21#_M1006_g 0.0508363f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_32 VNB N_A_713_21#_c_564_n 0.00253778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_713_21#_c_565_n 0.00316203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_713_21#_c_566_n 0.0247079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_713_21#_c_567_n 0.0196499f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_560_47#_c_640_n 0.0195151f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_37 VNB N_A_560_47#_c_641_n 0.0441682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_560_47#_c_642_n 0.00807186f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_39 VNB N_A_560_47#_c_643_n 0.00754924f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_40 VNB N_A_560_47#_c_644_n 0.0034004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_560_47#_c_645_n 0.00905941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_723_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB Q 0.0131477f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_44 VNB N_Q_c_816_n 0.0251065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_830_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_46 VNB N_VGND_c_831_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_47 VNB N_VGND_c_832_n 0.00714112f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_48 VNB N_VGND_c_833_n 0.00491327f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_49 VNB N_VGND_c_834_n 0.0200635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_835_n 0.00394313f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.53
cc_51 VNB N_VGND_c_836_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_837_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_838_n 0.0394571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_839_n 0.0199269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_840_n 0.29854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_841_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_842_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_843_n 0.00507544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VPB N_GATE_c_132_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_60 VPB N_GATE_c_133_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_61 VPB N_GATE_c_134_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_62 VPB GATE 0.0153801f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_63 VPB N_GATE_c_130_n 0.0106763f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_64 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_65 VPB N_A_27_47#_M1004_g 0.0300163f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_66 VPB N_A_27_47#_c_171_n 0.0172363f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_67 VPB N_A_27_47#_c_172_n 0.00940865f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_68 VPB N_A_27_47#_c_183_n 0.0121148f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_69 VPB N_A_27_47#_c_184_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_185_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_176_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_187_n 0.0224566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_188_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_189_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_190_n 0.00344459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_191_n 0.00529835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_192_n 0.00947367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_178_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_D_M1014_g 0.0462501f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_80 VPB N_D_c_318_n 0.00235013f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_81 VPB N_A_299_47#_M1013_g 0.036646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_299_47#_c_364_n 0.00712099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_299_47#_c_365_n 0.00409088f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_84 VPB N_A_299_47#_c_366_n 0.00290124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_299_47#_c_359_n 0.00355393f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_86 VPB N_A_193_47#_M1002_g 0.020263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_193_47#_c_439_n 0.00804665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_193_47#_c_446_n 0.00293933f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_89 VPB N_A_193_47#_c_447_n 0.00873764f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.19
cc_90 VPB N_A_193_47#_c_448_n 0.00238602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_193_47#_c_449_n 0.00711634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_193_47#_c_450_n 0.00239593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_193_47#_c_451_n 0.0270871f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_193_47#_c_452_n 0.00849735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_193_47#_c_443_n 0.00250944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_713_21#_M1006_g 0.0154265f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_97 VPB N_A_713_21#_M1009_g 0.0258593f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_98 VPB N_A_713_21#_M1003_g 0.022522f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_99 VPB N_A_713_21#_c_571_n 0.00551022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_713_21#_c_572_n 0.0473509f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_101 VPB N_A_713_21#_c_573_n 0.00370604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_713_21#_c_565_n 0.00305444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_713_21#_c_566_n 0.00673586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_560_47#_M1001_g 0.0223351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_560_47#_c_641_n 0.0150381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_560_47#_c_642_n 5.11268e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_107 VPB N_A_560_47#_c_649_n 0.00530349f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_108 VPB N_A_560_47#_c_644_n 0.00210101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_724_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_110 VPB N_VPWR_c_725_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_111 VPB N_VPWR_c_726_n 0.00470153f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_112 VPB N_VPWR_c_727_n 0.00491327f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_113 VPB N_VPWR_c_728_n 0.0395284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_729_n 0.00324376f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.53
cc_115 VPB N_VPWR_c_730_n 0.021856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_731_n 0.00391723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_732_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_733_n 0.0295132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_734_n 0.0192621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_723_n 0.0594177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_736_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_737_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB Q 0.00545527f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_124 VPB Q 0.0250272f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_125 VPB N_Q_c_816_n 0.0158513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 N_GATE_c_127_n N_A_27_47#_M1012_g 0.0187834f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_127 N_GATE_c_131_n N_A_27_47#_M1012_g 0.00419721f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_128 N_GATE_c_134_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_129 N_GATE_c_130_n N_A_27_47#_M1000_g 0.00527139f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_130 N_GATE_c_127_n N_A_27_47#_c_174_n 0.00663556f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_131 N_GATE_c_128_n N_A_27_47#_c_174_n 0.0105293f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_132 N_GATE_c_128_n N_A_27_47#_c_175_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_133 GATE N_A_27_47#_c_175_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_134 N_GATE_c_130_n N_A_27_47#_c_175_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_135 N_GATE_c_133_n N_A_27_47#_c_184_n 0.0135489f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_136 N_GATE_c_134_n N_A_27_47#_c_184_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_137 N_GATE_c_133_n N_A_27_47#_c_185_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_138 N_GATE_c_134_n N_A_27_47#_c_185_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_139 GATE N_A_27_47#_c_185_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_140 N_GATE_c_130_n N_A_27_47#_c_185_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_141 N_GATE_c_130_n N_A_27_47#_c_176_n 0.00319349f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_142 N_GATE_c_128_n N_A_27_47#_c_177_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_143 GATE N_A_27_47#_c_177_n 0.0288278f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_144 N_GATE_c_131_n N_A_27_47#_c_177_n 0.00151818f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_145 N_GATE_c_132_n N_A_27_47#_c_188_n 0.0033897f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_146 N_GATE_c_134_n N_A_27_47#_c_188_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_147 GATE N_A_27_47#_c_188_n 0.00653562f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_148 N_GATE_c_132_n N_A_27_47#_c_189_n 7.602e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_149 N_GATE_c_134_n N_A_27_47#_c_189_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_150 GATE N_A_27_47#_c_178_n 9.06856e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_151 N_GATE_c_130_n N_A_27_47#_c_178_n 0.0165768f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_152 N_GATE_c_133_n N_VPWR_c_724_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_153 N_GATE_c_133_n N_VPWR_c_732_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_154 N_GATE_c_133_n N_VPWR_c_723_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_155 N_GATE_c_127_n N_VGND_c_830_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_156 N_GATE_c_127_n N_VGND_c_836_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_157 N_GATE_c_128_n N_VGND_c_836_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_158 N_GATE_c_127_n N_VGND_c_840_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_187_n N_D_M1014_g 0.00583826f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_187_n N_D_c_318_n 0.0087134f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_161 N_A_27_47#_M1012_g N_D_c_319_n 0.00520956f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_27_47#_M1004_g N_A_299_47#_M1013_g 0.0360425f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_172_n N_A_299_47#_M1013_g 0.0248435f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_187_n N_A_299_47#_M1013_g 0.00493352f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_190_n N_A_299_47#_M1013_g 0.00140912f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_191_n N_A_299_47#_M1013_g 0.00239179f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_187_n N_A_299_47#_c_365_n 0.0116439f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_190_n N_A_299_47#_c_365_n 0.00130924f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_191_n N_A_299_47#_c_365_n 0.00675603f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_187_n N_A_299_47#_c_366_n 0.0115067f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_187_n N_A_299_47#_c_358_n 0.00675641f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_187_n N_A_299_47#_c_359_n 0.0108494f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_190_n N_A_299_47#_c_359_n 0.00124596f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_191_n N_A_299_47#_c_359_n 0.00570493f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_187_n N_A_299_47#_c_361_n 0.00107604f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1004_g N_A_193_47#_M1002_g 0.0197558f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_M1012_g N_A_193_47#_c_439_n 0.00779983f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_174_n N_A_193_47#_c_439_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_176_n N_A_193_47#_c_439_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_177_n N_A_193_47#_c_439_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_187_n N_A_193_47#_c_439_n 0.0184539f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_188_n N_A_193_47#_c_439_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_189_n N_A_193_47#_c_439_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_184_n N_A_193_47#_c_446_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_187_n N_A_193_47#_c_446_n 0.00195186f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_178_n N_A_193_47#_c_446_n 0.00779983f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_172_n N_A_193_47#_c_440_n 0.0197851f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1007_g N_A_193_47#_c_440_n 0.0192857f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_191_n N_A_193_47#_c_440_n 5.32999e-19 $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_171_n N_A_193_47#_c_441_n 7.03475e-19 $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_172_n N_A_193_47#_c_441_n 0.00136018f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1007_g N_A_193_47#_c_441_n 0.00256371f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_191_n N_A_193_47#_c_441_n 0.00180905f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1004_g N_A_193_47#_c_447_n 0.00738725f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_195 N_A_27_47#_c_171_n N_A_193_47#_c_447_n 0.00118095f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_183_n N_A_193_47#_c_447_n 0.00190431f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_187_n N_A_193_47#_c_447_n 0.0871075f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_190_n N_A_193_47#_c_447_n 0.0266027f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_191_n N_A_193_47#_c_447_n 0.00879307f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_M1000_g N_A_193_47#_c_448_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_184_n N_A_193_47#_c_448_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_187_n N_A_193_47#_c_448_n 0.0259095f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_189_n N_A_193_47#_c_448_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_M1000_g N_A_193_47#_c_449_n 0.00779983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_M1004_g N_A_193_47#_c_450_n 0.00144777f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_206 N_A_27_47#_c_171_n N_A_193_47#_c_450_n 0.00114785f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1007_g N_A_193_47#_c_442_n 0.0155884f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_M1004_g N_A_193_47#_c_451_n 0.0114263f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_171_n N_A_193_47#_c_451_n 0.0184478f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_183_n N_A_193_47#_c_451_n 0.00489663f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_M1004_g N_A_193_47#_c_452_n 0.00476768f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_212 N_A_27_47#_c_171_n N_A_193_47#_c_452_n 0.00413065f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_183_n N_A_193_47#_c_452_n 0.0026326f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_171_n N_A_193_47#_c_443_n 0.0127486f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_M1007_g N_A_193_47#_c_443_n 0.00492704f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_190_n N_A_193_47#_c_443_n 0.00148697f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_191_n N_A_193_47#_c_443_n 0.0232128f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_192_n N_A_193_47#_c_443_n 0.0026326f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_M1007_g N_A_713_21#_M1006_g 0.0546091f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1004_g N_A_560_47#_c_651_n 0.00377685f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_221 N_A_27_47#_M1007_g N_A_560_47#_c_652_n 0.0123233f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_M1007_g N_A_560_47#_c_643_n 0.00527917f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_171_n N_A_560_47#_c_649_n 6.38593e-19 $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_M1007_g N_A_560_47#_c_645_n 0.00328462f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_184_n N_VPWR_M1011_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_226 N_A_27_47#_M1000_g N_VPWR_c_724_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_184_n N_VPWR_c_724_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_185_n N_VPWR_c_724_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_188_n N_VPWR_c_724_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_230 N_A_27_47#_M1004_g N_VPWR_c_725_n 0.0040344f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_187_n N_VPWR_c_725_n 0.0019389f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_232 N_A_27_47#_M1004_g N_VPWR_c_728_n 0.0054153f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_184_n N_VPWR_c_732_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_185_n N_VPWR_c_732_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_235 N_A_27_47#_M1000_g N_VPWR_c_733_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_M1000_g N_VPWR_c_723_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1004_g N_VPWR_c_723_n 0.00634589f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_184_n N_VPWR_c_723_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_185_n N_VPWR_c_723_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_174_n N_VGND_M1016_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_241 N_A_27_47#_M1012_g N_VGND_c_830_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_174_n N_VGND_c_830_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_176_n N_VGND_c_830_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_178_n N_VGND_c_830_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_M1007_g N_VGND_c_832_n 0.00181257f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_307_p N_VGND_c_836_n 0.00713694f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_174_n N_VGND_c_836_n 0.00243651f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_248 N_A_27_47#_M1012_g N_VGND_c_837_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_249 N_A_27_47#_M1007_g N_VGND_c_838_n 0.0037981f $X=3.22 $Y=0.415 $X2=0 $Y2=0
cc_250 N_A_27_47#_M1016_s N_VGND_c_840_n 0.003754f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_251 N_A_27_47#_M1012_g N_VGND_c_840_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1007_g N_VGND_c_840_n 0.00557956f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_307_p N_VGND_c_840_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_174_n N_VGND_c_840_n 0.00549708f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_255 N_D_c_319_n N_A_299_47#_M1013_g 0.03863f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_256 N_D_M1014_g N_A_299_47#_c_364_n 0.012851f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_257 N_D_M1005_g N_A_299_47#_c_357_n 0.0144498f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_258 N_D_c_318_n N_A_299_47#_c_357_n 0.00627239f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_259 N_D_c_319_n N_A_299_47#_c_357_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_260 N_D_M1014_g N_A_299_47#_c_365_n 0.00794545f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_261 N_D_M1014_g N_A_299_47#_c_366_n 0.00412429f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_262 N_D_c_318_n N_A_299_47#_c_366_n 0.0229667f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_263 N_D_c_319_n N_A_299_47#_c_366_n 0.00131849f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_264 N_D_M1005_g N_A_299_47#_c_358_n 0.00563568f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_265 N_D_c_318_n N_A_299_47#_c_358_n 0.0107593f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_266 N_D_c_318_n N_A_299_47#_c_359_n 0.0164827f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_267 N_D_c_319_n N_A_299_47#_c_359_n 0.00552652f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_268 N_D_M1005_g N_A_299_47#_c_360_n 0.00120855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_269 N_D_c_318_n N_A_299_47#_c_360_n 0.0138491f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_270 N_D_c_319_n N_A_299_47#_c_360_n 0.0042466f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_271 N_D_M1005_g N_A_299_47#_c_361_n 0.0197208f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_272 N_D_M1005_g N_A_299_47#_c_362_n 0.015283f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_273 N_D_M1005_g N_A_193_47#_c_439_n 0.00203374f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_274 N_D_M1014_g N_A_193_47#_c_439_n 0.00459933f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_275 N_D_c_318_n N_A_193_47#_c_439_n 0.0209974f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_276 N_D_c_319_n N_A_193_47#_c_439_n 0.00256393f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_277 N_D_M1014_g N_A_193_47#_c_446_n 0.00134564f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_278 N_D_M1014_g N_A_193_47#_c_447_n 0.00294239f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_279 N_D_M1014_g N_VPWR_c_725_n 0.00304701f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_280 N_D_M1014_g N_VPWR_c_733_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_281 N_D_M1014_g N_VPWR_c_723_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_282 N_D_M1005_g N_VGND_c_831_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_283 N_D_M1005_g N_VGND_c_837_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_284 N_D_M1005_g N_VGND_c_840_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_285 N_D_c_319_n N_VGND_c_840_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_286 N_A_299_47#_c_364_n N_A_193_47#_c_439_n 0.0010921f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_287 N_A_299_47#_c_366_n N_A_193_47#_c_439_n 0.00859001f $X=1.785 $Y=1.58
+ $X2=0 $Y2=0
cc_288 N_A_299_47#_c_360_n N_A_193_47#_c_439_n 0.0191833f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_289 N_A_299_47#_c_364_n N_A_193_47#_c_446_n 0.0471072f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_290 N_A_299_47#_c_358_n N_A_193_47#_c_440_n 9.5712e-19 $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_291 N_A_299_47#_c_361_n N_A_193_47#_c_440_n 0.0126737f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_292 N_A_299_47#_c_358_n N_A_193_47#_c_441_n 0.012908f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_293 N_A_299_47#_c_361_n N_A_193_47#_c_441_n 9.1294e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_294 N_A_299_47#_M1013_g N_A_193_47#_c_447_n 0.00364042f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_295 N_A_299_47#_c_364_n N_A_193_47#_c_447_n 0.022748f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_296 N_A_299_47#_c_365_n N_A_193_47#_c_447_n 0.00551435f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_297 N_A_299_47#_c_364_n N_A_193_47#_c_448_n 0.00273055f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_298 N_A_299_47#_c_362_n N_A_193_47#_c_442_n 0.0262132f $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_299 N_A_299_47#_M1013_g N_A_193_47#_c_443_n 0.00370009f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_300 N_A_299_47#_c_358_n N_A_193_47#_c_443_n 0.00178567f $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_301 N_A_299_47#_c_361_n N_A_193_47#_c_443_n 9.9633e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_302 N_A_299_47#_M1013_g N_A_560_47#_c_651_n 4.99236e-19 $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_303 N_A_299_47#_M1013_g N_VPWR_c_725_n 0.0234565f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_304 N_A_299_47#_c_364_n N_VPWR_c_725_n 0.0232987f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_305 N_A_299_47#_c_365_n N_VPWR_c_725_n 0.013562f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_306 N_A_299_47#_M1013_g N_VPWR_c_728_n 0.00212864f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_307 N_A_299_47#_c_364_n N_VPWR_c_733_n 0.0159418f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_308 N_A_299_47#_M1014_s N_VPWR_c_723_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_309 N_A_299_47#_M1013_g N_VPWR_c_723_n 0.00261509f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_310 N_A_299_47#_c_364_n N_VPWR_c_723_n 0.00576627f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_311 N_A_299_47#_c_358_n N_VGND_M1005_d 0.00156939f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_312 N_A_299_47#_c_357_n N_VGND_c_831_n 0.00259081f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_313 N_A_299_47#_c_358_n N_VGND_c_831_n 0.0141976f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_314 N_A_299_47#_c_362_n N_VGND_c_831_n 0.0094968f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_315 N_A_299_47#_c_357_n N_VGND_c_837_n 0.00255672f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_316 N_A_299_47#_c_360_n N_VGND_c_837_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_317 N_A_299_47#_c_361_n N_VGND_c_838_n 9.84895e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_318 N_A_299_47#_c_362_n N_VGND_c_838_n 0.0046653f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_319 N_A_299_47#_M1005_s N_VGND_c_840_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_320 N_A_299_47#_c_357_n N_VGND_c_840_n 0.00473142f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_321 N_A_299_47#_c_358_n N_VGND_c_840_n 0.00552372f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_322 N_A_299_47#_c_360_n N_VGND_c_840_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_323 N_A_299_47#_c_361_n N_VGND_c_840_n 0.00117722f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_324 N_A_299_47#_c_362_n N_VGND_c_840_n 0.00440683f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_325 N_A_193_47#_c_443_n N_A_713_21#_M1006_g 9.87052e-19 $X=3.095 $Y=1.575
+ $X2=0 $Y2=0
cc_326 N_A_193_47#_M1002_g N_A_713_21#_M1009_g 0.0253509f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_327 N_A_193_47#_c_452_n N_A_713_21#_M1009_g 3.29084e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_328 N_A_193_47#_c_451_n N_A_713_21#_c_572_n 0.0157438f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_329 N_A_193_47#_c_452_n N_A_713_21#_c_572_n 3.93081e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_330 N_A_193_47#_M1002_g N_A_560_47#_c_651_n 0.00872591f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_331 N_A_193_47#_c_447_n N_A_560_47#_c_651_n 0.00241909f $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_332 N_A_193_47#_c_450_n N_A_560_47#_c_651_n 0.00255896f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_333 N_A_193_47#_c_451_n N_A_560_47#_c_651_n 0.00219621f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_334 N_A_193_47#_c_452_n N_A_560_47#_c_651_n 0.0133551f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_335 N_A_193_47#_c_440_n N_A_560_47#_c_652_n 0.00209266f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_336 N_A_193_47#_c_441_n N_A_560_47#_c_652_n 0.0177949f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_337 N_A_193_47#_c_441_n N_A_560_47#_c_643_n 0.0184898f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_338 N_A_193_47#_M1002_g N_A_560_47#_c_649_n 0.00559487f $X=3.145 $Y=2.275
+ $X2=0 $Y2=0
cc_339 N_A_193_47#_c_450_n N_A_560_47#_c_649_n 0.00130177f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_340 N_A_193_47#_c_451_n N_A_560_47#_c_649_n 0.00171665f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_341 N_A_193_47#_c_452_n N_A_560_47#_c_649_n 0.0309805f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_342 N_A_193_47#_c_443_n N_A_560_47#_c_649_n 0.0113314f $X=3.095 $Y=1.575
+ $X2=0 $Y2=0
cc_343 N_A_193_47#_c_441_n N_A_560_47#_c_645_n 0.0027819f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_344 N_A_193_47#_c_451_n N_A_560_47#_c_645_n 4.91178e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_345 N_A_193_47#_c_443_n N_A_560_47#_c_645_n 0.0167533f $X=3.095 $Y=1.575
+ $X2=0 $Y2=0
cc_346 N_A_193_47#_c_447_n N_VPWR_M1014_d 6.81311e-19 $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_347 N_A_193_47#_c_449_n N_VPWR_c_724_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_348 N_A_193_47#_c_447_n N_VPWR_c_725_n 0.0184727f $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_349 N_A_193_47#_c_450_n N_VPWR_c_725_n 9.60836e-19 $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_350 N_A_193_47#_c_452_n N_VPWR_c_725_n 0.0021853f $X=3.18 $Y=1.74 $X2=0 $Y2=0
cc_351 N_A_193_47#_M1002_g N_VPWR_c_728_n 0.00366111f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_352 N_A_193_47#_c_449_n N_VPWR_c_733_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_353 N_A_193_47#_M1002_g N_VPWR_c_723_n 0.00541284f $X=3.145 $Y=2.275 $X2=0
+ $Y2=0
cc_354 N_A_193_47#_c_447_n N_VPWR_c_723_n 0.0750686f $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_355 N_A_193_47#_c_448_n N_VPWR_c_723_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_356 N_A_193_47#_c_449_n N_VPWR_c_723_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_357 N_A_193_47#_c_450_n N_VPWR_c_723_n 0.0147399f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_358 N_A_193_47#_c_447_n A_465_369# 0.00387108f $X=2.87 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_359 N_A_193_47#_c_442_n N_VGND_c_831_n 0.00184485f $X=2.792 $Y=0.705 $X2=0
+ $Y2=0
cc_360 N_A_193_47#_c_439_n N_VGND_c_837_n 0.00732874f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_361 N_A_193_47#_c_440_n N_VGND_c_838_n 6.62516e-19 $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_362 N_A_193_47#_c_441_n N_VGND_c_838_n 0.00182549f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_363 N_A_193_47#_c_442_n N_VGND_c_838_n 0.00500228f $X=2.792 $Y=0.705 $X2=0
+ $Y2=0
cc_364 N_A_193_47#_M1012_d N_VGND_c_840_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_365 N_A_193_47#_c_439_n N_VGND_c_840_n 0.00616598f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_366 N_A_193_47#_c_440_n N_VGND_c_840_n 9.75233e-19 $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_367 N_A_193_47#_c_441_n N_VGND_c_840_n 0.00344069f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_368 N_A_193_47#_c_442_n N_VGND_c_840_n 0.00848363f $X=2.792 $Y=0.705 $X2=0
+ $Y2=0
cc_369 N_A_713_21#_c_564_n N_A_560_47#_c_640_n 0.00671379f $X=4.43 $Y=0.995
+ $X2=0 $Y2=0
cc_370 N_A_713_21#_c_567_n N_A_560_47#_c_640_n 0.0210784f $X=5.01 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A_713_21#_M1003_g N_A_560_47#_M1001_g 0.0224331f $X=5.025 $Y=1.985
+ $X2=0 $Y2=0
cc_372 N_A_713_21#_c_572_n N_A_560_47#_M1001_g 0.00407044f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_373 N_A_713_21#_c_573_n N_A_560_47#_M1001_g 0.00755466f $X=4.43 $Y=1.535
+ $X2=0 $Y2=0
cc_374 N_A_713_21#_c_587_p N_A_560_47#_M1001_g 8.96335e-19 $X=4.38 $Y=1.755
+ $X2=0 $Y2=0
cc_375 N_A_713_21#_M1006_g N_A_560_47#_c_641_n 0.0181721f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_376 N_A_713_21#_c_571_n N_A_560_47#_c_641_n 0.00755072f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_377 N_A_713_21#_c_572_n N_A_560_47#_c_641_n 0.00639877f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_378 N_A_713_21#_c_591_p N_A_560_47#_c_641_n 0.00182108f $X=4.38 $Y=0.58 $X2=0
+ $Y2=0
cc_379 N_A_713_21#_c_587_p N_A_560_47#_c_641_n 0.00212837f $X=4.38 $Y=1.755
+ $X2=0 $Y2=0
cc_380 N_A_713_21#_c_593_p N_A_560_47#_c_641_n 0.017901f $X=4.43 $Y=1.16 $X2=0
+ $Y2=0
cc_381 N_A_713_21#_c_565_n N_A_560_47#_c_642_n 0.0218426f $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_382 N_A_713_21#_c_566_n N_A_560_47#_c_642_n 0.0214946f $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_383 N_A_713_21#_M1009_g N_A_560_47#_c_651_n 0.00475392f $X=3.64 $Y=2.275
+ $X2=0 $Y2=0
cc_384 N_A_713_21#_M1006_g N_A_560_47#_c_652_n 0.00147432f $X=3.64 $Y=0.415
+ $X2=0 $Y2=0
cc_385 N_A_713_21#_M1006_g N_A_560_47#_c_643_n 0.0107407f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_386 N_A_713_21#_M1006_g N_A_560_47#_c_649_n 0.0114592f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_387 N_A_713_21#_M1009_g N_A_560_47#_c_649_n 0.015786f $X=3.64 $Y=2.275 $X2=0
+ $Y2=0
cc_388 N_A_713_21#_c_571_n N_A_560_47#_c_649_n 0.0192517f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_389 N_A_713_21#_c_572_n N_A_560_47#_c_649_n 0.00911775f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_390 N_A_713_21#_M1006_g N_A_560_47#_c_644_n 0.0164414f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_391 N_A_713_21#_c_571_n N_A_560_47#_c_644_n 0.0221958f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_392 N_A_713_21#_c_572_n N_A_560_47#_c_644_n 0.00776367f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_393 N_A_713_21#_c_593_p N_A_560_47#_c_644_n 0.0277655f $X=4.43 $Y=1.16 $X2=0
+ $Y2=0
cc_394 N_A_713_21#_M1006_g N_A_560_47#_c_645_n 0.0059144f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_395 N_A_713_21#_M1009_g N_VPWR_c_726_n 0.00622935f $X=3.64 $Y=2.275 $X2=0
+ $Y2=0
cc_396 N_A_713_21#_c_571_n N_VPWR_c_726_n 0.00562825f $X=4.295 $Y=1.7 $X2=0
+ $Y2=0
cc_397 N_A_713_21#_c_572_n N_VPWR_c_726_n 0.00481721f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_398 N_A_713_21#_c_611_p N_VPWR_c_726_n 0.013068f $X=4.38 $Y=2.27 $X2=0 $Y2=0
cc_399 N_A_713_21#_M1003_g N_VPWR_c_727_n 0.00366919f $X=5.025 $Y=1.985 $X2=0
+ $Y2=0
cc_400 N_A_713_21#_c_565_n N_VPWR_c_727_n 0.0123213f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_401 N_A_713_21#_c_566_n N_VPWR_c_727_n 5.14689e-19 $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_402 N_A_713_21#_M1009_g N_VPWR_c_728_n 0.00526858f $X=3.64 $Y=2.275 $X2=0
+ $Y2=0
cc_403 N_A_713_21#_c_611_p N_VPWR_c_730_n 0.0112378f $X=4.38 $Y=2.27 $X2=0 $Y2=0
cc_404 N_A_713_21#_M1003_g N_VPWR_c_734_n 0.00585385f $X=5.025 $Y=1.985 $X2=0
+ $Y2=0
cc_405 N_A_713_21#_M1001_s N_VPWR_c_723_n 0.0023739f $X=4.255 $Y=1.485 $X2=0
+ $Y2=0
cc_406 N_A_713_21#_M1009_g N_VPWR_c_723_n 0.010697f $X=3.64 $Y=2.275 $X2=0 $Y2=0
cc_407 N_A_713_21#_M1003_g N_VPWR_c_723_n 0.0115783f $X=5.025 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_A_713_21#_c_571_n N_VPWR_c_723_n 0.0125784f $X=4.295 $Y=1.7 $X2=0 $Y2=0
cc_409 N_A_713_21#_c_572_n N_VPWR_c_723_n 0.00394376f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_410 N_A_713_21#_c_611_p N_VPWR_c_723_n 0.00827281f $X=4.38 $Y=2.27 $X2=0
+ $Y2=0
cc_411 N_A_713_21#_M1003_g N_Q_c_816_n 0.00948536f $X=5.025 $Y=1.985 $X2=0 $Y2=0
cc_412 N_A_713_21#_c_565_n N_Q_c_816_n 0.0262108f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_413 N_A_713_21#_c_566_n N_Q_c_816_n 0.00755993f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_414 N_A_713_21#_c_567_n N_Q_c_816_n 0.00686745f $X=5.01 $Y=0.995 $X2=0 $Y2=0
cc_415 N_A_713_21#_M1006_g N_VGND_c_832_n 0.0111886f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_416 N_A_713_21#_c_591_p N_VGND_c_832_n 0.00639259f $X=4.38 $Y=0.58 $X2=0
+ $Y2=0
cc_417 N_A_713_21#_c_565_n N_VGND_c_833_n 0.0111962f $X=5.01 $Y=1.16 $X2=0 $Y2=0
cc_418 N_A_713_21#_c_566_n N_VGND_c_833_n 5.02062e-19 $X=5.01 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A_713_21#_c_567_n N_VGND_c_833_n 0.0032775f $X=5.01 $Y=0.995 $X2=0
+ $Y2=0
cc_420 N_A_713_21#_c_591_p N_VGND_c_834_n 0.00650283f $X=4.38 $Y=0.58 $X2=0
+ $Y2=0
cc_421 N_A_713_21#_M1006_g N_VGND_c_838_n 0.0046653f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_422 N_A_713_21#_c_567_n N_VGND_c_839_n 0.00585385f $X=5.01 $Y=0.995 $X2=0
+ $Y2=0
cc_423 N_A_713_21#_M1008_s N_VGND_c_840_n 0.00370868f $X=4.255 $Y=0.235 $X2=0
+ $Y2=0
cc_424 N_A_713_21#_M1006_g N_VGND_c_840_n 0.00799591f $X=3.64 $Y=0.415 $X2=0
+ $Y2=0
cc_425 N_A_713_21#_c_591_p N_VGND_c_840_n 0.00761394f $X=4.38 $Y=0.58 $X2=0
+ $Y2=0
cc_426 N_A_713_21#_c_567_n N_VGND_c_840_n 0.0117699f $X=5.01 $Y=0.995 $X2=0
+ $Y2=0
cc_427 N_A_560_47#_c_651_n N_VPWR_c_725_n 0.00552787f $X=3.435 $Y=2.34 $X2=0
+ $Y2=0
cc_428 N_A_560_47#_M1001_g N_VPWR_c_726_n 0.00310876f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_429 N_A_560_47#_c_651_n N_VPWR_c_726_n 0.0133617f $X=3.435 $Y=2.34 $X2=0
+ $Y2=0
cc_430 N_A_560_47#_c_649_n N_VPWR_c_726_n 0.00839059f $X=3.52 $Y=2.255 $X2=0
+ $Y2=0
cc_431 N_A_560_47#_M1001_g N_VPWR_c_727_n 0.00381684f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_432 N_A_560_47#_c_651_n N_VPWR_c_728_n 0.0373288f $X=3.435 $Y=2.34 $X2=0
+ $Y2=0
cc_433 N_A_560_47#_M1001_g N_VPWR_c_730_n 0.00585385f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_434 N_A_560_47#_M1004_d N_VPWR_c_723_n 0.00173952f $X=2.8 $Y=2.065 $X2=0
+ $Y2=0
cc_435 N_A_560_47#_M1001_g N_VPWR_c_723_n 0.0120037f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_436 N_A_560_47#_c_651_n N_VPWR_c_723_n 0.0218494f $X=3.435 $Y=2.34 $X2=0
+ $Y2=0
cc_437 N_A_560_47#_c_651_n A_644_413# 0.00670962f $X=3.435 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_438 N_A_560_47#_c_649_n A_644_413# 0.00226411f $X=3.52 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_439 N_A_560_47#_c_640_n N_VGND_c_832_n 0.00662174f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_440 N_A_560_47#_c_641_n N_VGND_c_832_n 0.00112595f $X=4.515 $Y=1.16 $X2=0
+ $Y2=0
cc_441 N_A_560_47#_c_652_n N_VGND_c_832_n 0.0127315f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_442 N_A_560_47#_c_644_n N_VGND_c_832_n 0.0121132f $X=4.09 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A_560_47#_c_640_n N_VGND_c_833_n 0.00340873f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_444 N_A_560_47#_c_640_n N_VGND_c_834_n 0.00585385f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_445 N_A_560_47#_c_652_n N_VGND_c_838_n 0.0228359f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_446 N_A_560_47#_M1015_d N_VGND_c_840_n 0.00310043f $X=2.8 $Y=0.235 $X2=0
+ $Y2=0
cc_447 N_A_560_47#_c_640_n N_VGND_c_840_n 0.0120818f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_448 N_A_560_47#_c_652_n N_VGND_c_840_n 0.022423f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_449 N_A_560_47#_c_652_n A_659_47# 0.00347857f $X=3.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_450 N_A_560_47#_c_643_n A_659_47# 7.28282e-19 $X=3.415 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_451 N_VPWR_c_723_n A_465_369# 0.00469197f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_452 N_VPWR_c_723_n A_644_413# 0.00280095f $X=5.29 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_453 N_VPWR_c_723_n N_Q_M1003_d 0.00403684f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_454 N_VPWR_c_734_n Q 0.0185715f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_455 N_VPWR_c_723_n Q 0.0108473f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_456 Q N_VGND_c_839_n 0.00948931f $X=5.23 $Y=0.425 $X2=0 $Y2=0
cc_457 N_Q_M1017_d N_VGND_c_840_n 0.00428292f $X=5.1 $Y=0.235 $X2=0 $Y2=0
cc_458 Q N_VGND_c_840_n 0.00983854f $X=5.23 $Y=0.425 $X2=0 $Y2=0
cc_459 N_VGND_c_840_n A_465_47# 0.0123065f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24
cc_460 N_VGND_c_840_n A_659_47# 0.00451958f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__sdfxtp_2.pxi.spice
* Created: Thu Aug 27 14:47:25 2020
* 
x_PM_SKY130_FD_SC_HD__SDFXTP_2%CLK N_CLK_c_214_n N_CLK_c_218_n N_CLK_c_215_n
+ N_CLK_M1031_g N_CLK_c_219_n N_CLK_M1012_g N_CLK_c_220_n CLK CLK
+ PM_SKY130_FD_SC_HD__SDFXTP_2%CLK
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_27_47# N_A_27_47#_M1031_s N_A_27_47#_M1012_s
+ N_A_27_47#_M1018_g N_A_27_47#_M1029_g N_A_27_47#_M1028_g N_A_27_47#_c_258_n
+ N_A_27_47#_c_259_n N_A_27_47#_M1030_g N_A_27_47#_M1009_g N_A_27_47#_c_260_n
+ N_A_27_47#_M1004_g N_A_27_47#_c_493_p N_A_27_47#_c_262_n N_A_27_47#_c_263_n
+ N_A_27_47#_c_275_n N_A_27_47#_c_264_n N_A_27_47#_c_381_p N_A_27_47#_c_276_n
+ N_A_27_47#_c_277_n N_A_27_47#_c_265_n N_A_27_47#_c_278_n N_A_27_47#_c_279_n
+ N_A_27_47#_c_280_n N_A_27_47#_c_281_n N_A_27_47#_c_282_n N_A_27_47#_c_266_n
+ N_A_27_47#_c_284_n N_A_27_47#_c_285_n N_A_27_47#_c_286_n N_A_27_47#_c_267_n
+ N_A_27_47#_c_268_n PM_SKY130_FD_SC_HD__SDFXTP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%SCE N_SCE_M1024_g N_SCE_M1032_g N_SCE_c_514_n
+ N_SCE_M1014_g N_SCE_M1026_g N_SCE_c_505_n N_SCE_c_506_n N_SCE_c_517_n
+ N_SCE_c_507_n N_SCE_c_532_p N_SCE_c_508_n N_SCE_c_509_n N_SCE_c_510_n
+ N_SCE_c_511_n SCE N_SCE_c_512_n PM_SKY130_FD_SC_HD__SDFXTP_2%SCE
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_299_47# N_A_299_47#_M1032_s N_A_299_47#_M1024_s
+ N_A_299_47#_M1021_g N_A_299_47#_M1007_g N_A_299_47#_c_624_n
+ N_A_299_47#_c_631_n N_A_299_47#_c_639_n N_A_299_47#_c_625_n
+ N_A_299_47#_c_641_n N_A_299_47#_c_633_n N_A_299_47#_c_626_n
+ N_A_299_47#_c_634_n N_A_299_47#_c_627_n N_A_299_47#_c_628_n
+ N_A_299_47#_c_646_n N_A_299_47#_c_635_n N_A_299_47#_c_636_n
+ PM_SKY130_FD_SC_HD__SDFXTP_2%A_299_47#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%D N_D_M1016_g N_D_M1022_g D N_D_c_754_n
+ N_D_c_755_n PM_SKY130_FD_SC_HD__SDFXTP_2%D
x_PM_SKY130_FD_SC_HD__SDFXTP_2%SCD N_SCD_M1020_g N_SCD_M1005_g SCD SCD
+ N_SCD_c_802_n PM_SKY130_FD_SC_HD__SDFXTP_2%SCD
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_193_47# N_A_193_47#_M1018_d N_A_193_47#_M1029_d
+ N_A_193_47#_M1008_g N_A_193_47#_M1001_g N_A_193_47#_c_848_n
+ N_A_193_47#_M1003_g N_A_193_47#_M1000_g N_A_193_47#_c_849_n
+ N_A_193_47#_c_865_n N_A_193_47#_c_850_n N_A_193_47#_c_851_n
+ N_A_193_47#_c_852_n N_A_193_47#_c_867_n N_A_193_47#_c_868_n
+ N_A_193_47#_c_853_n N_A_193_47#_c_854_n N_A_193_47#_c_855_n
+ N_A_193_47#_c_989_p N_A_193_47#_c_856_n N_A_193_47#_c_857_n
+ N_A_193_47#_c_858_n N_A_193_47#_c_859_n N_A_193_47#_c_860_n
+ N_A_193_47#_c_861_n PM_SKY130_FD_SC_HD__SDFXTP_2%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_1098_183# N_A_1098_183#_M1017_d
+ N_A_1098_183#_M1025_d N_A_1098_183#_M1006_g N_A_1098_183#_M1023_g
+ N_A_1098_183#_c_1067_n N_A_1098_183#_c_1093_n N_A_1098_183#_c_1113_p
+ N_A_1098_183#_c_1094_n N_A_1098_183#_c_1068_n N_A_1098_183#_c_1069_n
+ N_A_1098_183#_c_1081_n N_A_1098_183#_c_1070_n N_A_1098_183#_c_1071_n
+ PM_SKY130_FD_SC_HD__SDFXTP_2%A_1098_183#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_939_413# N_A_939_413#_M1028_d
+ N_A_939_413#_M1008_d N_A_939_413#_c_1160_n N_A_939_413#_M1025_g
+ N_A_939_413#_c_1161_n N_A_939_413#_M1017_g N_A_939_413#_c_1162_n
+ N_A_939_413#_c_1163_n N_A_939_413#_c_1164_n N_A_939_413#_c_1178_n
+ N_A_939_413#_c_1204_n N_A_939_413#_c_1165_n N_A_939_413#_c_1170_n
+ N_A_939_413#_c_1166_n PM_SKY130_FD_SC_HD__SDFXTP_2%A_939_413#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_1526_315# N_A_1526_315#_M1015_s
+ N_A_1526_315#_M1002_s N_A_1526_315#_M1019_g N_A_1526_315#_M1027_g
+ N_A_1526_315#_c_1270_n N_A_1526_315#_M1011_g N_A_1526_315#_M1010_g
+ N_A_1526_315#_c_1271_n N_A_1526_315#_M1013_g N_A_1526_315#_M1033_g
+ N_A_1526_315#_c_1280_n N_A_1526_315#_c_1281_n N_A_1526_315#_c_1293_p
+ N_A_1526_315#_c_1272_n N_A_1526_315#_c_1282_n N_A_1526_315#_c_1273_n
+ N_A_1526_315#_c_1274_n N_A_1526_315#_c_1295_p N_A_1526_315#_c_1300_p
+ N_A_1526_315#_c_1275_n PM_SKY130_FD_SC_HD__SDFXTP_2%A_1526_315#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_1355_413# N_A_1355_413#_M1003_d
+ N_A_1355_413#_M1009_d N_A_1355_413#_c_1368_n N_A_1355_413#_M1015_g
+ N_A_1355_413#_M1002_g N_A_1355_413#_c_1369_n N_A_1355_413#_c_1370_n
+ N_A_1355_413#_c_1380_n N_A_1355_413#_c_1383_n N_A_1355_413#_c_1377_n
+ N_A_1355_413#_c_1371_n N_A_1355_413#_c_1372_n N_A_1355_413#_c_1373_n
+ PM_SKY130_FD_SC_HD__SDFXTP_2%A_1355_413#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%VPWR N_VPWR_M1012_d N_VPWR_M1024_d N_VPWR_M1005_d
+ N_VPWR_M1006_d N_VPWR_M1019_d N_VPWR_M1002_d N_VPWR_M1033_s N_VPWR_c_1457_n
+ N_VPWR_c_1458_n N_VPWR_c_1459_n N_VPWR_c_1460_n N_VPWR_c_1461_n
+ N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n N_VPWR_c_1465_n
+ N_VPWR_c_1466_n N_VPWR_c_1467_n VPWR N_VPWR_c_1468_n N_VPWR_c_1469_n
+ N_VPWR_c_1470_n N_VPWR_c_1471_n N_VPWR_c_1472_n N_VPWR_c_1473_n
+ N_VPWR_c_1474_n N_VPWR_c_1475_n N_VPWR_c_1476_n N_VPWR_c_1477_n
+ N_VPWR_c_1456_n PM_SKY130_FD_SC_HD__SDFXTP_2%VPWR
x_PM_SKY130_FD_SC_HD__SDFXTP_2%A_559_369# N_A_559_369#_M1022_d
+ N_A_559_369#_M1028_s N_A_559_369#_M1016_d N_A_559_369#_M1008_s
+ N_A_559_369#_c_1632_n N_A_559_369#_c_1644_n N_A_559_369#_c_1656_n
+ N_A_559_369#_c_1621_n N_A_559_369#_c_1628_n N_A_559_369#_c_1629_n
+ N_A_559_369#_c_1622_n N_A_559_369#_c_1623_n N_A_559_369#_c_1624_n
+ N_A_559_369#_c_1625_n N_A_559_369#_c_1626_n N_A_559_369#_c_1627_n
+ N_A_559_369#_c_1631_n PM_SKY130_FD_SC_HD__SDFXTP_2%A_559_369#
x_PM_SKY130_FD_SC_HD__SDFXTP_2%Q N_Q_M1011_s N_Q_M1010_d N_Q_c_1744_n
+ N_Q_c_1742_n Q Q Q N_Q_c_1757_n PM_SKY130_FD_SC_HD__SDFXTP_2%Q
x_PM_SKY130_FD_SC_HD__SDFXTP_2%VGND N_VGND_M1031_d N_VGND_M1032_d N_VGND_M1020_d
+ N_VGND_M1023_d N_VGND_M1027_d N_VGND_M1015_d N_VGND_M1013_d N_VGND_c_1773_n
+ N_VGND_c_1774_n N_VGND_c_1775_n N_VGND_c_1776_n N_VGND_c_1777_n
+ N_VGND_c_1778_n N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n
+ N_VGND_c_1782_n VGND N_VGND_c_1783_n N_VGND_c_1784_n N_VGND_c_1785_n
+ N_VGND_c_1786_n N_VGND_c_1787_n N_VGND_c_1788_n N_VGND_c_1789_n
+ N_VGND_c_1790_n N_VGND_c_1791_n N_VGND_c_1792_n N_VGND_c_1793_n
+ N_VGND_c_1794_n PM_SKY130_FD_SC_HD__SDFXTP_2%VGND
cc_1 VNB N_CLK_c_214_n 0.0573151f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_215_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0185843f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1018_g 0.0381832f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1028_g 0.0521093f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_6 VNB N_A_27_47#_c_258_n 0.0136466f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_7 VNB N_A_27_47#_c_259_n 0.00249911f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_8 VNB N_A_27_47#_c_260_n 0.0158261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1004_g 0.043789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_262_n 0.00319094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_263_n 0.00642096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_264_n 8.11193e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_265_n 0.00238722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_266_n 0.0228343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_267_n 0.00980165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_268_n 0.00148891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_SCE_M1032_g 0.0206182f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_18 VNB N_SCE_M1026_g 0.016865f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_19 VNB N_SCE_c_505_n 0.003249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_SCE_c_506_n 0.00457186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_507_n 0.00292878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_508_n 0.00344001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_509_n 0.00118673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_510_n 0.0272672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_SCE_c_511_n 0.00148358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_SCE_c_512_n 0.0267875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_299_47#_M1021_g 0.021613f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_28 VNB N_A_299_47#_c_624_n 0.0137655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_299_47#_c_625_n 0.00261142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_299_47#_c_626_n 0.00249039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_299_47#_c_627_n 0.00280608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_299_47#_c_628_n 0.0298276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_D_M1022_g 0.0443728f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_34 VNB N_SCD_M1020_g 0.0457816f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_35 VNB SCD 0.00498049f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_36 VNB N_SCD_c_802_n 0.0137367f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_37 VNB N_A_193_47#_c_848_n 0.0180432f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_38 VNB N_A_193_47#_c_849_n 0.00330396f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.53
cc_39 VNB N_A_193_47#_c_850_n 0.00369255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_851_n 0.00403969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_193_47#_c_852_n 0.00632811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_193_47#_c_853_n 0.0492616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_193_47#_c_854_n 0.00572932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_193_47#_c_855_n 0.0101801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_193_47#_c_856_n 0.0114368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_193_47#_c_857_n 9.18319e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_193_47#_c_858_n 0.0266741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_193_47#_c_859_n 0.005674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_193_47#_c_860_n 0.0176138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_193_47#_c_861_n 0.0285203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1098_183#_M1006_g 0.0146965f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_52 VNB N_A_1098_183#_M1023_g 0.0210316f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_53 VNB N_A_1098_183#_c_1067_n 0.00354578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1098_183#_c_1068_n 0.00364457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1098_183#_c_1069_n 0.00130441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1098_183#_c_1070_n 0.00302393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1098_183#_c_1071_n 0.0338642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_939_413#_c_1160_n 0.0118275f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.135
cc_59 VNB N_A_939_413#_c_1161_n 0.0158415f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_60 VNB N_A_939_413#_c_1162_n 0.0152351f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_61 VNB N_A_939_413#_c_1163_n 0.00913873f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_62 VNB N_A_939_413#_c_1164_n 8.51874e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_939_413#_c_1165_n 0.0118271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_939_413#_c_1166_n 0.00180949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1526_315#_M1027_g 0.0482636f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_66 VNB N_A_1526_315#_c_1270_n 0.0165357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1526_315#_c_1271_n 0.0203476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1526_315#_c_1272_n 0.00161491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1526_315#_c_1273_n 0.00425124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1526_315#_c_1274_n 0.00701384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1526_315#_c_1275_n 0.0484489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1355_413#_c_1368_n 0.0205013f $X=-0.19 $Y=-0.24 $X2=0.475
+ $Y2=2.135
cc_73 VNB N_A_1355_413#_c_1369_n 0.0393229f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.445
cc_74 VNB N_A_1355_413#_c_1370_n 0.00807254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1355_413#_c_1371_n 0.00998398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1355_413#_c_1372_n 0.00584041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1355_413#_c_1373_n 0.00344545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VPWR_c_1456_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_559_369#_c_1621_n 2.29256e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_559_369#_c_1622_n 0.0119702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_559_369#_c_1623_n 0.00220658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_559_369#_c_1624_n 0.00350881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_559_369#_c_1625_n 0.00922578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_559_369#_c_1626_n 0.00246161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_559_369#_c_1627_n 0.00182501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_Q_c_1742_n 0.00103903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1773_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1774_n 0.00278677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1775_n 0.00486519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1776_n 0.0460447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1777_n 0.0058544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1778_n 0.00237946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1779_n 0.0220776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1780_n 0.00470745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1781_n 0.0110531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1782_n 0.00922231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1783_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1784_n 0.0289225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1785_n 0.0344998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1786_n 0.0430904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1787_n 0.0192854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1788_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1789_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1790_n 0.00381885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1791_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1792_n 0.00513917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1793_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1794_n 0.484781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VPB N_CLK_c_214_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_110 VPB N_CLK_c_218_n 0.0162394f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_111 VPB N_CLK_c_219_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.74
cc_112 VPB N_CLK_c_220_n 0.0235707f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_113 VPB CLK 0.0178159f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_114 VPB N_A_27_47#_M1029_g 0.03676f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_115 VPB N_A_27_47#_c_258_n 0.0143056f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_116 VPB N_A_27_47#_c_259_n 0.0052612f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_117 VPB N_A_27_47#_M1030_g 0.0191311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_M1009_g 0.033754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_260_n 0.0211567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_275_n 0.00174908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_276_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_277_n 0.00356676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_27_47#_c_278_n 0.0575467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_47#_c_279_n 0.00148899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_27_47#_c_280_n 0.00118201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_27_47#_c_281_n 8.53245e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_47#_c_282_n 0.00543917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_266_n 0.0115869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_284_n 0.0266783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_285_n 0.00853708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_286_n 0.0106236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_267_n 0.0208929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_268_n 0.00437972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_SCE_M1024_g 0.0236916f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_135 VPB N_SCE_c_514_n 0.0160433f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_136 VPB N_SCE_M1014_g 0.0195854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_SCE_c_506_n 0.00116067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_SCE_c_517_n 0.027587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_SCE_c_512_n 0.00509208f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_299_47#_M1007_g 0.0184813f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_141 VPB N_A_299_47#_c_624_n 0.0105202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_299_47#_c_631_n 0.00406887f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_143 VPB N_A_299_47#_c_625_n 0.00416757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_299_47#_c_633_n 0.00158406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_299_47#_c_634_n 0.0018061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_299_47#_c_635_n 0.0014433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_299_47#_c_636_n 0.027856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_D_M1016_g 0.0190988f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_149 VPB N_D_M1022_g 0.003603f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.135
cc_150 VPB N_D_c_754_n 0.0270161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_D_c_755_n 0.00442173f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_152 VPB N_SCD_M1005_g 0.0337159f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.135
cc_153 VPB SCD 0.0061556f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_154 VPB N_SCD_c_802_n 0.0200872f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_155 VPB N_A_193_47#_M1008_g 0.024991f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_156 VPB N_A_193_47#_M1000_g 0.0221869f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_157 VPB N_A_193_47#_c_849_n 0.00462988f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.53
cc_158 VPB N_A_193_47#_c_865_n 0.0328226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_193_47#_c_850_n 0.00311128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_193_47#_c_867_n 0.00568481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_193_47#_c_868_n 0.0266658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_193_47#_c_856_n 0.0173127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_1098_183#_M1006_g 0.049805f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_164 VPB N_A_1098_183#_c_1070_n 0.00255179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_939_413#_M1025_g 0.0226707f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.665
cc_166 VPB N_A_939_413#_c_1163_n 0.0189969f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_167 VPB N_A_939_413#_c_1164_n 0.00681499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_939_413#_c_1170_n 0.00161138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_939_413#_c_1166_n 0.00888291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1526_315#_M1019_g 0.0253795f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_171 VPB N_A_1526_315#_M1027_g 0.0179972f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_172 VPB N_A_1526_315#_M1010_g 0.0191788f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_173 VPB N_A_1526_315#_M1033_g 0.0232394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_1526_315#_c_1280_n 0.0129293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1526_315#_c_1281_n 0.040764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1526_315#_c_1282_n 0.00235569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1526_315#_c_1273_n 0.00425124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1526_315#_c_1275_n 0.00901875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1355_413#_M1002_g 0.0237342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1355_413#_c_1369_n 0.014657f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_181 VPB N_A_1355_413#_c_1370_n 5.1131e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1355_413#_c_1377_n 0.0126839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1355_413#_c_1371_n 0.00386833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1355_413#_c_1372_n 0.0050339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1457_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1458_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1459_n 0.00470486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1460_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1461_n 0.00548955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1462_n 0.0226033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1463_n 0.00472584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1464_n 0.0110272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1465_n 0.0108407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1466_n 0.0523928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1467_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1468_n 0.0156572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1469_n 0.0255003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1470_n 0.0377079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1471_n 0.0449606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1472_n 0.0192387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1473_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1474_n 0.00436214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1475_n 0.00324297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1476_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1477_n 0.00334019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1456_n 0.062548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_559_369#_c_1628_n 0.00866343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_559_369#_c_1629_n 0.00155557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_559_369#_c_1625_n 0.0111823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_559_369#_c_1631_n 0.00872065f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_Q_c_1742_n 0.00122795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 N_CLK_c_214_n N_A_27_47#_M1018_g 0.0049062f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_213 N_CLK_c_215_n N_A_27_47#_M1018_g 0.0187731f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_214 CLK N_A_27_47#_M1018_g 3.14819e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_215 N_CLK_c_218_n N_A_27_47#_M1029_g 0.00531917f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_216 N_CLK_c_220_n N_A_27_47#_M1029_g 0.0276478f $X=0.475 $Y=1.665 $X2=0 $Y2=0
cc_217 CLK N_A_27_47#_M1029_g 5.73308e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_218 N_CLK_c_214_n N_A_27_47#_c_262_n 0.00761961f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_219 N_CLK_c_215_n N_A_27_47#_c_262_n 0.00668648f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_220 CLK N_A_27_47#_c_262_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_221 N_CLK_c_214_n N_A_27_47#_c_263_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_222 CLK N_A_27_47#_c_263_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_223 N_CLK_c_219_n N_A_27_47#_c_275_n 0.0128144f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_224 N_CLK_c_220_n N_A_27_47#_c_275_n 0.0013816f $X=0.475 $Y=1.665 $X2=0 $Y2=0
cc_225 CLK N_A_27_47#_c_275_n 0.00728212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_226 N_CLK_c_214_n N_A_27_47#_c_264_n 3.98708e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_227 CLK N_A_27_47#_c_264_n 0.0516739f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_228 N_CLK_c_214_n N_A_27_47#_c_276_n 2.90926e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_229 N_CLK_c_218_n N_A_27_47#_c_276_n 7.09762e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_230 N_CLK_c_220_n N_A_27_47#_c_276_n 0.00440146f $X=0.475 $Y=1.665 $X2=0
+ $Y2=0
cc_231 N_CLK_c_214_n N_A_27_47#_c_277_n 2.26313e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_232 N_CLK_c_219_n N_A_27_47#_c_277_n 2.17882e-19 $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_233 N_CLK_c_220_n N_A_27_47#_c_277_n 0.00358837f $X=0.475 $Y=1.665 $X2=0
+ $Y2=0
cc_234 CLK N_A_27_47#_c_277_n 0.0153364f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_235 N_CLK_c_214_n N_A_27_47#_c_265_n 0.00381855f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_236 N_CLK_c_219_n N_A_27_47#_c_279_n 0.00101286f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_237 N_CLK_c_214_n N_A_27_47#_c_266_n 0.0169285f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_238 CLK N_A_27_47#_c_266_n 0.00161876f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_239 N_CLK_c_219_n N_VPWR_c_1457_n 0.00946555f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_240 N_CLK_c_219_n N_VPWR_c_1468_n 0.00332278f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_241 N_CLK_c_219_n N_VPWR_c_1456_n 0.00485269f $X=0.475 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_215_n N_VGND_c_1773_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_243 N_CLK_c_214_n N_VGND_c_1783_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_244 N_CLK_c_215_n N_VGND_c_1783_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_245 N_CLK_c_215_n N_VGND_c_1794_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_278_n N_SCE_M1024_g 0.00322296f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_278_n N_SCE_M1014_g 0.0012424f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_278_n N_SCE_c_506_n 0.00414929f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_278_n N_SCE_c_517_n 0.00351631f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_278_n N_A_299_47#_M1007_g 7.69535e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_278_n N_A_299_47#_c_624_n 0.0120648f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_278_n N_A_299_47#_c_639_n 0.0163793f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_278_n N_A_299_47#_c_625_n 0.00921137f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_278_n N_A_299_47#_c_641_n 0.0367444f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_278_n N_A_299_47#_c_633_n 0.0113096f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1018_g N_A_299_47#_c_626_n 9.61905e-19 $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_278_n N_A_299_47#_c_634_n 0.0130054f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_278_n N_A_299_47#_c_628_n 0.00277281f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_278_n N_A_299_47#_c_646_n 0.0046527f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_278_n N_A_299_47#_c_635_n 7.81108e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_278_n N_A_299_47#_c_636_n 0.0016565f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_278_n N_D_M1016_g 0.00218294f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_278_n N_D_c_754_n 0.00308822f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_278_n N_D_c_755_n 0.00838144f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_278_n N_SCD_M1005_g 0.00187497f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_278_n SCD 0.0124672f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_278_n N_A_193_47#_M1029_d 6.81311e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_278_n N_A_193_47#_M1008_g 0.00371812f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_284_n N_A_193_47#_M1008_g 0.0144165f $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_285_n N_A_193_47#_M1008_g 9.60176e-19 $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1004_g N_A_193_47#_c_848_n 0.0144677f $X=7.345 $Y=0.415 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1009_g N_A_193_47#_M1000_g 0.0175056f $X=6.7 $Y=2.275 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_282_n N_A_193_47#_M1000_g 0.00135837f $X=6.705 $Y=1.87 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_268_n N_A_193_47#_M1000_g 5.16255e-19 $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1028_g N_A_193_47#_c_849_n 0.0077284f $X=4.625 $Y=0.415 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_258_n N_A_193_47#_c_849_n 0.00687115f $X=5.01 $Y=1.32 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_259_n N_A_193_47#_c_849_n 0.00418731f $X=4.7 $Y=1.32 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_278_n N_A_193_47#_c_849_n 0.0139192f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_281_n N_A_193_47#_c_849_n 2.1733e-19 $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_284_n N_A_193_47#_c_849_n 7.29366e-19 $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_285_n N_A_193_47#_c_849_n 0.0168958f $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_286_n N_A_193_47#_c_849_n 0.00604391f $X=5.145 $Y=1.575
+ $X2=0 $Y2=0
cc_283 N_A_27_47#_c_259_n N_A_193_47#_c_865_n 0.0162569f $X=4.7 $Y=1.32 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_278_n N_A_193_47#_c_865_n 0.00545515f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_284_n N_A_193_47#_c_865_n 0.0174998f $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_285_n N_A_193_47#_c_865_n 0.00118389f $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_260_n N_A_193_47#_c_850_n 0.0117161f $X=7.27 $Y=1.32 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1004_g N_A_193_47#_c_850_n 0.00430042f $X=7.345 $Y=0.415
+ $X2=0 $Y2=0
cc_289 N_A_27_47#_c_267_n N_A_193_47#_c_850_n 0.00402309f $X=6.695 $Y=1.32 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_268_n N_A_193_47#_c_850_n 0.0234373f $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_M1018_g N_A_193_47#_c_851_n 0.00136529f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_262_n N_A_193_47#_c_851_n 0.00442897f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1004_g N_A_193_47#_c_852_n 0.0020279f $X=7.345 $Y=0.415 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_267_n N_A_193_47#_c_852_n 0.00222109f $X=6.695 $Y=1.32 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_268_n N_A_193_47#_c_852_n 0.0119224f $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_M1009_g N_A_193_47#_c_867_n 0.00117691f $X=6.7 $Y=2.275 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_260_n N_A_193_47#_c_867_n 0.00338756f $X=7.27 $Y=1.32 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_282_n N_A_193_47#_c_867_n 0.00508223f $X=6.705 $Y=1.87 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_268_n N_A_193_47#_c_867_n 0.0245744f $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_M1009_g N_A_193_47#_c_868_n 0.0130792f $X=6.7 $Y=2.275 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_260_n N_A_193_47#_c_868_n 0.0212127f $X=7.27 $Y=1.32 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_268_n N_A_193_47#_c_868_n 6.54911e-19 $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_M1028_g N_A_193_47#_c_853_n 0.00225641f $X=4.625 $Y=0.415
+ $X2=0 $Y2=0
cc_304 N_A_27_47#_M1018_g N_A_193_47#_c_854_n 0.00662116f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_262_n N_A_193_47#_c_854_n 0.0022123f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_265_n N_A_193_47#_c_854_n 0.00516669f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_267_n N_A_193_47#_c_855_n 2.10748e-19 $X=6.695 $Y=1.32 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_M1018_g N_A_193_47#_c_856_n 0.00851768f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_262_n N_A_193_47#_c_856_n 0.0055484f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_264_n N_A_193_47#_c_856_n 0.059769f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_381_p N_A_193_47#_c_856_n 0.00826673f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_265_n N_A_193_47#_c_856_n 0.00884862f $X=0.73 $Y=0.97 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_278_n N_A_193_47#_c_856_n 0.0247251f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_279_n N_A_193_47#_c_856_n 0.00244764f $X=0.87 $Y=1.87 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_266_n N_A_193_47#_c_856_n 0.0174894f $X=0.895 $Y=1.235 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_267_n N_A_193_47#_c_857_n 9.82747e-19 $X=6.695 $Y=1.32 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_268_n N_A_193_47#_c_857_n 0.00125233f $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_M1028_g N_A_193_47#_c_858_n 0.0213105f $X=4.625 $Y=0.415 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_258_n N_A_193_47#_c_858_n 0.0174066f $X=5.01 $Y=1.32 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_284_n N_A_193_47#_c_858_n 5.43883e-19 $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_285_n N_A_193_47#_c_858_n 4.76262e-19 $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_M1028_g N_A_193_47#_c_859_n 0.0116468f $X=4.625 $Y=0.415 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_258_n N_A_193_47#_c_859_n 0.00587088f $X=5.01 $Y=1.32 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_285_n N_A_193_47#_c_859_n 0.00398178f $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1028_g N_A_193_47#_c_860_n 0.0102604f $X=4.625 $Y=0.415 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_M1004_g N_A_193_47#_c_861_n 0.0193601f $X=7.345 $Y=0.415 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_267_n N_A_193_47#_c_861_n 0.020308f $X=6.695 $Y=1.32 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_280_n N_A_1098_183#_M1025_d 0.00523078f $X=6.56 $Y=1.87
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_258_n N_A_1098_183#_M1006_g 0.0113457f $X=5.01 $Y=1.32 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_M1030_g N_A_1098_183#_M1006_g 0.0276008f $X=5.085 $Y=2.275
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_280_n N_A_1098_183#_M1006_g 0.00281129f $X=6.56 $Y=1.87
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_281_n N_A_1098_183#_M1006_g 0.00148276f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_284_n N_A_1098_183#_M1006_g 0.0206011f $X=5.145 $Y=1.74
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_285_n N_A_1098_183#_M1006_g 0.0022f $X=5.145 $Y=1.74 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_280_n N_A_1098_183#_c_1081_n 0.00261642f $X=6.56 $Y=1.87
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_M1009_g N_A_1098_183#_c_1070_n 0.00455971f $X=6.7 $Y=2.275
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_280_n N_A_1098_183#_c_1070_n 0.0193938f $X=6.56 $Y=1.87
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_282_n N_A_1098_183#_c_1070_n 0.00314501f $X=6.705 $Y=1.87
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_c_267_n N_A_1098_183#_c_1070_n 0.00225153f $X=6.695 $Y=1.32
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_268_n N_A_1098_183#_c_1070_n 0.0517078f $X=6.695 $Y=1.41
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_267_n N_A_939_413#_c_1160_n 0.0158005f $X=6.695 $Y=1.32
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_c_268_n N_A_939_413#_c_1160_n 3.03019e-19 $X=6.695 $Y=1.41
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_M1009_g N_A_939_413#_M1025_g 0.0247799f $X=6.7 $Y=2.275 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_280_n N_A_939_413#_M1025_g 0.00700233f $X=6.56 $Y=1.87 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_268_n N_A_939_413#_M1025_g 8.29633e-19 $X=6.695 $Y=1.41
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_c_280_n N_A_939_413#_c_1163_n 0.00109659f $X=6.56 $Y=1.87
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_M1030_g N_A_939_413#_c_1178_n 0.00859817f $X=5.085 $Y=2.275
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_278_n N_A_939_413#_c_1178_n 0.00697565f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_280_n N_A_939_413#_c_1178_n 0.00383646f $X=6.56 $Y=1.87
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_281_n N_A_939_413#_c_1178_n 0.00159423f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_284_n N_A_939_413#_c_1178_n 5.38487e-19 $X=5.145 $Y=1.74
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_c_285_n N_A_939_413#_c_1178_n 0.0252801f $X=5.145 $Y=1.74
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_M1028_g N_A_939_413#_c_1165_n 9.86268e-19 $X=4.625 $Y=0.415
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_258_n N_A_939_413#_c_1165_n 8.14452e-19 $X=5.01 $Y=1.32
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_M1030_g N_A_939_413#_c_1170_n 9.97608e-19 $X=5.085 $Y=2.275
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_280_n N_A_939_413#_c_1170_n 0.0183205f $X=6.56 $Y=1.87 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_281_n N_A_939_413#_c_1170_n 0.00257444f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_c_284_n N_A_939_413#_c_1170_n 7.00613e-19 $X=5.145 $Y=1.74
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_285_n N_A_939_413#_c_1170_n 0.0250151f $X=5.145 $Y=1.74
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_c_258_n N_A_939_413#_c_1166_n 0.00225879f $X=5.01 $Y=1.32
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_280_n N_A_939_413#_c_1166_n 0.0176196f $X=6.56 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_281_n N_A_939_413#_c_1166_n 0.00154209f $X=5.435 $Y=1.87
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_285_n N_A_939_413#_c_1166_n 0.00980238f $X=5.145 $Y=1.74
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_286_n N_A_939_413#_c_1166_n 4.44848e-19 $X=5.145 $Y=1.575
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_M1004_g N_A_1526_315#_M1027_g 0.0463015f $X=7.345 $Y=0.415
+ $X2=0 $Y2=0
cc_366 N_A_27_47#_M1009_g N_A_1355_413#_c_1380_n 0.00281529f $X=6.7 $Y=2.275
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_c_282_n N_A_1355_413#_c_1380_n 0.00210372f $X=6.705 $Y=1.87
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_c_268_n N_A_1355_413#_c_1380_n 0.0022468f $X=6.695 $Y=1.41
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_M1004_g N_A_1355_413#_c_1383_n 0.00800808f $X=7.345 $Y=0.415
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_282_n N_A_1355_413#_c_1377_n 0.00228172f $X=6.705 $Y=1.87
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_268_n N_A_1355_413#_c_1377_n 9.63849e-19 $X=6.695 $Y=1.41
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_M1004_g N_A_1355_413#_c_1371_n 3.1587e-19 $X=7.345 $Y=0.415
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_260_n N_A_1355_413#_c_1372_n 0.00558094f $X=7.27 $Y=1.32
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_M1004_g N_A_1355_413#_c_1372_n 0.0061466f $X=7.345 $Y=0.415
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_M1004_g N_A_1355_413#_c_1373_n 0.0110517f $X=7.345 $Y=0.415
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_381_p N_VPWR_M1012_d 6.91013e-19 $X=0.73 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_377 N_A_27_47#_c_279_n N_VPWR_M1012_d 0.00178771f $X=0.87 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_378 N_A_27_47#_c_280_n N_VPWR_M1006_d 0.00678497f $X=6.56 $Y=1.87 $X2=0 $Y2=0
cc_379 N_A_27_47#_M1029_g N_VPWR_c_1457_n 0.00937841f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_275_n N_VPWR_c_1457_n 0.0031092f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_381_p N_VPWR_c_1457_n 0.0133497f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_277_n N_VPWR_c_1457_n 0.012721f $X=0.265 $Y=1.96 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_279_n N_VPWR_c_1457_n 0.00330948f $X=0.87 $Y=1.87 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_278_n N_VPWR_c_1458_n 0.00124409f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_278_n N_VPWR_c_1459_n 8.00522e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_280_n N_VPWR_c_1460_n 0.00950843f $X=6.56 $Y=1.87 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_M1030_g N_VPWR_c_1466_n 0.0037886f $X=5.085 $Y=2.275 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_275_n N_VPWR_c_1468_n 0.0018545f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_277_n N_VPWR_c_1468_n 0.0120313f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_M1029_g N_VPWR_c_1469_n 0.00442511f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_M1009_g N_VPWR_c_1471_n 0.00430107f $X=6.7 $Y=2.275 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_268_n N_VPWR_c_1471_n 0.00157744f $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_M1029_g N_VPWR_c_1456_n 0.00534571f $X=0.895 $Y=2.135 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_M1030_g N_VPWR_c_1456_n 0.00557208f $X=5.085 $Y=2.275 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_M1009_g N_VPWR_c_1456_n 0.0057371f $X=6.7 $Y=2.275 $X2=0 $Y2=0
cc_396 N_A_27_47#_c_275_n N_VPWR_c_1456_n 0.00403677f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_277_n N_VPWR_c_1456_n 0.00646745f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_278_n N_VPWR_c_1456_n 0.199302f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_399 N_A_27_47#_c_279_n N_VPWR_c_1456_n 0.0145601f $X=0.87 $Y=1.87 $X2=0 $Y2=0
cc_400 N_A_27_47#_c_280_n N_VPWR_c_1456_n 0.0532767f $X=6.56 $Y=1.87 $X2=0 $Y2=0
cc_401 N_A_27_47#_c_281_n N_VPWR_c_1456_n 0.0146717f $X=5.435 $Y=1.87 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_282_n N_VPWR_c_1456_n 0.0159329f $X=6.705 $Y=1.87 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_268_n N_VPWR_c_1456_n 0.00100625f $X=6.695 $Y=1.41 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_278_n N_A_559_369#_c_1632_n 0.00584375f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_278_n N_A_559_369#_c_1628_n 0.0229627f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_278_n N_A_559_369#_c_1629_n 0.0102321f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_M1028_g N_A_559_369#_c_1624_n 0.0044467f $X=4.625 $Y=0.415
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_M1028_g N_A_559_369#_c_1625_n 0.00902644f $X=4.625 $Y=0.415
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_278_n N_A_559_369#_c_1625_n 0.0104876f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_M1028_g N_A_559_369#_c_1626_n 0.00178202f $X=4.625 $Y=0.415
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_M1028_g N_A_559_369#_c_1627_n 0.00164257f $X=4.625 $Y=0.415
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_278_n N_A_559_369#_c_1631_n 0.0110091f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_285_n N_A_559_369#_c_1631_n 0.00314032f $X=5.145 $Y=1.74
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_278_n A_643_369# 0.00134881f $X=5.145 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_415 N_A_27_47#_c_262_n N_VGND_M1031_d 0.00166329f $X=0.615 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_416 N_A_27_47#_M1018_g N_VGND_c_1773_n 0.0100209f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_262_n N_VGND_c_1773_n 0.0150403f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_264_n N_VGND_c_1773_n 0.00108069f $X=0.73 $Y=1.085 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_266_n N_VGND_c_1773_n 5.70216e-19 $X=0.895 $Y=1.235 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_M1028_g N_VGND_c_1775_n 0.00339332f $X=4.625 $Y=0.415 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_M1028_g N_VGND_c_1776_n 0.00431421f $X=4.625 $Y=0.415 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_M1004_g N_VGND_c_1778_n 0.00230753f $X=7.345 $Y=0.415 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_493_p N_VGND_c_1783_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_262_n N_VGND_c_1783_n 0.00243651f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_M1018_g N_VGND_c_1784_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_M1004_g N_VGND_c_1786_n 0.00379696f $X=7.345 $Y=0.415 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_M1031_s N_VGND_c_1794_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_M1018_g N_VGND_c_1794_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_M1028_g N_VGND_c_1794_n 0.00721265f $X=4.625 $Y=0.415 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_M1004_g N_VGND_c_1794_n 0.00575728f $X=7.345 $Y=0.415 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_c_493_p N_VGND_c_1794_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_c_262_n N_VGND_c_1794_n 0.00564532f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_433 N_SCE_M1032_g N_A_299_47#_M1021_g 0.0181478f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_434 N_SCE_c_506_n N_A_299_47#_M1021_g 0.00148594f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_435 N_SCE_c_507_n N_A_299_47#_M1021_g 0.0106895f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_436 N_SCE_c_512_n N_A_299_47#_M1021_g 0.00259672f $X=1.865 $Y=1.385 $X2=0
+ $Y2=0
cc_437 N_SCE_M1024_g N_A_299_47#_c_624_n 0.00433634f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_438 N_SCE_M1032_g N_A_299_47#_c_624_n 0.00718205f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_439 N_SCE_c_505_n N_A_299_47#_c_624_n 0.0110051f $X=1.847 $Y=0.83 $X2=0 $Y2=0
cc_440 N_SCE_c_506_n N_A_299_47#_c_624_n 0.0621923f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_441 N_SCE_c_517_n N_A_299_47#_c_624_n 0.00716372f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_442 N_SCE_c_532_p N_A_299_47#_c_624_n 0.0130415f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_443 N_SCE_M1024_g N_A_299_47#_c_639_n 0.0125876f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_444 N_SCE_c_506_n N_A_299_47#_c_639_n 0.0103251f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_445 N_SCE_c_517_n N_A_299_47#_c_639_n 0.00410833f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_446 N_SCE_M1024_g N_A_299_47#_c_625_n 0.00143725f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_447 N_SCE_c_514_n N_A_299_47#_c_625_n 0.00760609f $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_448 N_SCE_M1014_g N_A_299_47#_c_625_n 0.00577745f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_449 N_SCE_c_506_n N_A_299_47#_c_625_n 0.0405815f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_450 N_SCE_c_517_n N_A_299_47#_c_625_n 0.00128732f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_451 N_SCE_c_512_n N_A_299_47#_c_625_n 0.00143321f $X=1.865 $Y=1.385 $X2=0
+ $Y2=0
cc_452 N_SCE_M1014_g N_A_299_47#_c_641_n 0.00557358f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_453 N_SCE_M1032_g N_A_299_47#_c_626_n 0.00239434f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_454 N_SCE_c_532_p N_A_299_47#_c_626_n 0.00168685f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_455 N_SCE_c_517_n N_A_299_47#_c_634_n 2.83838e-19 $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_456 N_SCE_c_514_n N_A_299_47#_c_627_n 4.17098e-19 $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_457 N_SCE_c_506_n N_A_299_47#_c_627_n 0.0134087f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_458 N_SCE_c_507_n N_A_299_47#_c_627_n 0.0205375f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_459 N_SCE_c_509_n N_A_299_47#_c_627_n 0.00388622f $X=3.165 $Y=0.95 $X2=0
+ $Y2=0
cc_460 N_SCE_c_512_n N_A_299_47#_c_627_n 5.19181e-19 $X=1.865 $Y=1.385 $X2=0
+ $Y2=0
cc_461 N_SCE_c_514_n N_A_299_47#_c_628_n 0.00783615f $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_462 N_SCE_c_506_n N_A_299_47#_c_628_n 0.00158198f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_463 N_SCE_c_507_n N_A_299_47#_c_628_n 0.00319888f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_464 N_SCE_c_512_n N_A_299_47#_c_628_n 0.0174165f $X=1.865 $Y=1.385 $X2=0
+ $Y2=0
cc_465 N_SCE_M1014_g N_A_299_47#_c_646_n 0.00682561f $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_466 N_SCE_c_509_n N_A_299_47#_c_635_n 0.00959271f $X=3.165 $Y=0.95 $X2=0
+ $Y2=0
cc_467 N_SCE_c_510_n N_A_299_47#_c_635_n 3.983e-19 $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_468 N_SCE_c_509_n N_A_299_47#_c_636_n 2.12418e-19 $X=3.165 $Y=0.95 $X2=0
+ $Y2=0
cc_469 N_SCE_c_510_n N_A_299_47#_c_636_n 0.0144723f $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_470 N_SCE_M1014_g N_D_M1016_g 0.0384234f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_471 N_SCE_M1026_g N_D_M1022_g 0.013704f $X=3.225 $Y=0.445 $X2=0 $Y2=0
cc_472 N_SCE_c_508_n N_D_M1022_g 0.012647f $X=3.08 $Y=0.7 $X2=0 $Y2=0
cc_473 N_SCE_c_509_n N_D_M1022_g 0.00203037f $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_474 N_SCE_c_510_n N_D_M1022_g 0.0213831f $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_475 N_SCE_c_514_n N_D_c_754_n 0.00996826f $X=2.185 $Y=1.58 $X2=0 $Y2=0
cc_476 N_SCE_c_517_n N_D_c_754_n 0.00186998f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_477 N_SCE_c_508_n N_D_c_754_n 7.55694e-19 $X=3.08 $Y=0.7 $X2=0 $Y2=0
cc_478 N_SCE_c_511_n N_D_c_754_n 0.00125086f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_479 N_SCE_c_512_n N_D_c_754_n 3.44894e-19 $X=1.865 $Y=1.385 $X2=0 $Y2=0
cc_480 N_SCE_c_514_n N_D_c_755_n 0.0012389f $X=2.185 $Y=1.58 $X2=0 $Y2=0
cc_481 N_SCE_c_507_n N_D_c_755_n 2.69368e-19 $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_482 N_SCE_c_508_n N_D_c_755_n 0.00189539f $X=3.08 $Y=0.7 $X2=0 $Y2=0
cc_483 N_SCE_c_511_n N_D_c_755_n 0.00314298f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_484 N_SCE_M1026_g N_SCD_M1020_g 0.0569691f $X=3.225 $Y=0.445 $X2=0 $Y2=0
cc_485 N_SCE_c_509_n N_SCD_M1020_g 0.00152146f $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_486 N_SCE_c_509_n SCD 0.00395967f $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_487 N_SCE_c_510_n SCD 2.88262e-19 $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_488 N_SCE_c_514_n N_A_193_47#_c_853_n 0.00163167f $X=2.185 $Y=1.58 $X2=0
+ $Y2=0
cc_489 N_SCE_M1026_g N_A_193_47#_c_853_n 5.27825e-19 $X=3.225 $Y=0.445 $X2=0
+ $Y2=0
cc_490 N_SCE_c_505_n N_A_193_47#_c_853_n 7.64766e-19 $X=1.847 $Y=0.83 $X2=0
+ $Y2=0
cc_491 N_SCE_c_506_n N_A_193_47#_c_853_n 0.0165918f $X=1.865 $Y=1.52 $X2=0 $Y2=0
cc_492 N_SCE_c_517_n N_A_193_47#_c_853_n 0.00319402f $X=1.865 $Y=1.52 $X2=0
+ $Y2=0
cc_493 N_SCE_c_507_n N_A_193_47#_c_853_n 0.0166965f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_494 N_SCE_c_532_p N_A_193_47#_c_853_n 0.0035151f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_495 N_SCE_c_508_n N_A_193_47#_c_853_n 0.0203609f $X=3.08 $Y=0.7 $X2=0 $Y2=0
cc_496 N_SCE_c_509_n N_A_193_47#_c_853_n 0.0108868f $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_497 N_SCE_c_510_n N_A_193_47#_c_853_n 0.0037338f $X=3.165 $Y=0.95 $X2=0 $Y2=0
cc_498 N_SCE_c_511_n N_A_193_47#_c_853_n 0.00735012f $X=2.562 $Y=0.7 $X2=0 $Y2=0
cc_499 N_SCE_c_512_n N_A_193_47#_c_853_n 0.0018864f $X=1.865 $Y=1.385 $X2=0
+ $Y2=0
cc_500 N_SCE_M1024_g N_A_193_47#_c_856_n 0.00160127f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_501 N_SCE_M1024_g N_VPWR_c_1458_n 0.00869424f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_502 N_SCE_M1014_g N_VPWR_c_1458_n 0.00922894f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_503 N_SCE_M1024_g N_VPWR_c_1469_n 0.00340533f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_504 N_SCE_M1014_g N_VPWR_c_1470_n 0.00354675f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_505 N_SCE_M1024_g N_VPWR_c_1456_n 0.00515557f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_506 N_SCE_M1014_g N_VPWR_c_1456_n 0.00403915f $X=2.26 $Y=2.165 $X2=0 $Y2=0
cc_507 N_SCE_c_508_n N_A_559_369#_M1022_d 0.00218892f $X=3.08 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_508 N_SCE_M1014_g N_A_559_369#_c_1632_n 5.71884e-19 $X=2.26 $Y=2.165 $X2=0
+ $Y2=0
cc_509 N_SCE_M1026_g N_A_559_369#_c_1644_n 0.00763758f $X=3.225 $Y=0.445 $X2=0
+ $Y2=0
cc_510 N_SCE_c_508_n N_A_559_369#_c_1644_n 0.0204608f $X=3.08 $Y=0.7 $X2=0 $Y2=0
cc_511 N_SCE_c_510_n N_A_559_369#_c_1644_n 2.32966e-19 $X=3.165 $Y=0.95 $X2=0
+ $Y2=0
cc_512 N_SCE_M1026_g N_A_559_369#_c_1621_n 0.00405684f $X=3.225 $Y=0.445 $X2=0
+ $Y2=0
cc_513 N_SCE_c_508_n N_A_559_369#_c_1621_n 0.00630259f $X=3.08 $Y=0.7 $X2=0
+ $Y2=0
cc_514 N_SCE_M1026_g N_A_559_369#_c_1623_n 9.7798e-19 $X=3.225 $Y=0.445 $X2=0
+ $Y2=0
cc_515 N_SCE_c_508_n N_A_559_369#_c_1623_n 0.00793437f $X=3.08 $Y=0.7 $X2=0
+ $Y2=0
cc_516 N_SCE_c_509_n N_A_559_369#_c_1623_n 0.00554533f $X=3.165 $Y=0.95 $X2=0
+ $Y2=0
cc_517 N_SCE_c_507_n N_VGND_M1032_d 0.00245508f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_518 N_SCE_M1032_g N_VGND_c_1774_n 0.00409505f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_519 N_SCE_c_507_n N_VGND_c_1774_n 0.018541f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_520 N_SCE_M1032_g N_VGND_c_1784_n 0.00409976f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_521 N_SCE_c_532_p N_VGND_c_1784_n 0.00251644f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_522 N_SCE_M1026_g N_VGND_c_1785_n 0.00362032f $X=3.225 $Y=0.445 $X2=0 $Y2=0
cc_523 N_SCE_c_507_n N_VGND_c_1785_n 0.00259773f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_524 N_SCE_c_508_n N_VGND_c_1785_n 0.00277894f $X=3.08 $Y=0.7 $X2=0 $Y2=0
cc_525 SCE N_VGND_c_1785_n 0.00782706f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_526 N_SCE_M1032_g N_VGND_c_1794_n 0.00686433f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_527 N_SCE_M1026_g N_VGND_c_1794_n 0.00526606f $X=3.225 $Y=0.445 $X2=0 $Y2=0
cc_528 N_SCE_c_507_n N_VGND_c_1794_n 0.00308055f $X=2.475 $Y=0.7 $X2=0 $Y2=0
cc_529 N_SCE_c_532_p N_VGND_c_1794_n 0.00183549f $X=1.95 $Y=0.7 $X2=0 $Y2=0
cc_530 N_SCE_c_508_n N_VGND_c_1794_n 0.00229883f $X=3.08 $Y=0.7 $X2=0 $Y2=0
cc_531 SCE N_VGND_c_1794_n 0.00302552f $X=2.475 $Y=0.425 $X2=0 $Y2=0
cc_532 SCE A_486_47# 0.00226988f $X=2.475 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_533 N_A_299_47#_M1007_g N_D_M1016_g 0.028319f $X=3.14 $Y=2.165 $X2=0 $Y2=0
cc_534 N_A_299_47#_c_625_n N_D_M1016_g 0.00113604f $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_535 N_A_299_47#_c_641_n N_D_M1016_g 0.0118472f $X=3.075 $Y=1.967 $X2=0 $Y2=0
cc_536 N_A_299_47#_c_633_n N_D_M1016_g 0.00126571f $X=3.16 $Y=1.86 $X2=0 $Y2=0
cc_537 N_A_299_47#_M1021_g N_D_M1022_g 0.0412182f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_538 N_A_299_47#_c_625_n N_D_M1022_g 0.00515026f $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_539 N_A_299_47#_c_627_n N_D_M1022_g 6.95453e-19 $X=2.295 $Y=1.04 $X2=0 $Y2=0
cc_540 N_A_299_47#_c_628_n N_D_M1022_g 0.0168449f $X=2.295 $Y=1.04 $X2=0 $Y2=0
cc_541 N_A_299_47#_c_625_n N_D_c_754_n 6.097e-19 $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_542 N_A_299_47#_c_641_n N_D_c_754_n 0.00290918f $X=3.075 $Y=1.967 $X2=0 $Y2=0
cc_543 N_A_299_47#_c_635_n N_D_c_754_n 0.0011165f $X=3.185 $Y=1.52 $X2=0 $Y2=0
cc_544 N_A_299_47#_c_636_n N_D_c_754_n 0.0197807f $X=3.185 $Y=1.52 $X2=0 $Y2=0
cc_545 N_A_299_47#_c_625_n N_D_c_755_n 0.025415f $X=2.205 $Y=1.86 $X2=0 $Y2=0
cc_546 N_A_299_47#_c_641_n N_D_c_755_n 0.0196694f $X=3.075 $Y=1.967 $X2=0 $Y2=0
cc_547 N_A_299_47#_c_635_n N_D_c_755_n 0.0157068f $X=3.185 $Y=1.52 $X2=0 $Y2=0
cc_548 N_A_299_47#_c_636_n N_D_c_755_n 0.00104193f $X=3.185 $Y=1.52 $X2=0 $Y2=0
cc_549 N_A_299_47#_M1007_g N_SCD_M1005_g 0.0359024f $X=3.14 $Y=2.165 $X2=0 $Y2=0
cc_550 N_A_299_47#_c_641_n N_SCD_M1005_g 2.17192e-19 $X=3.075 $Y=1.967 $X2=0
+ $Y2=0
cc_551 N_A_299_47#_c_633_n N_SCD_M1005_g 0.002483f $X=3.16 $Y=1.86 $X2=0 $Y2=0
cc_552 N_A_299_47#_c_635_n SCD 0.0158825f $X=3.185 $Y=1.52 $X2=0 $Y2=0
cc_553 N_A_299_47#_c_636_n SCD 0.00104429f $X=3.185 $Y=1.52 $X2=0 $Y2=0
cc_554 N_A_299_47#_c_635_n N_SCD_c_802_n 0.00107204f $X=3.185 $Y=1.52 $X2=0
+ $Y2=0
cc_555 N_A_299_47#_c_636_n N_SCD_c_802_n 0.0194305f $X=3.185 $Y=1.52 $X2=0 $Y2=0
cc_556 N_A_299_47#_c_624_n N_A_193_47#_c_851_n 0.0978566f $X=1.52 $Y=1.86 $X2=0
+ $Y2=0
cc_557 N_A_299_47#_c_626_n N_A_193_47#_c_851_n 0.00751783f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_558 N_A_299_47#_M1021_g N_A_193_47#_c_853_n 0.00170444f $X=2.355 $Y=0.445
+ $X2=0 $Y2=0
cc_559 N_A_299_47#_c_624_n N_A_193_47#_c_853_n 0.0181188f $X=1.52 $Y=1.86 $X2=0
+ $Y2=0
cc_560 N_A_299_47#_c_626_n N_A_193_47#_c_853_n 0.00465031f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_561 N_A_299_47#_c_627_n N_A_193_47#_c_853_n 0.00858868f $X=2.295 $Y=1.04
+ $X2=0 $Y2=0
cc_562 N_A_299_47#_c_628_n N_A_193_47#_c_853_n 0.00457609f $X=2.295 $Y=1.04
+ $X2=0 $Y2=0
cc_563 N_A_299_47#_c_635_n N_A_193_47#_c_853_n 0.00166362f $X=3.185 $Y=1.52
+ $X2=0 $Y2=0
cc_564 N_A_299_47#_c_636_n N_A_193_47#_c_853_n 6.70678e-19 $X=3.185 $Y=1.52
+ $X2=0 $Y2=0
cc_565 N_A_299_47#_c_624_n N_A_193_47#_c_854_n 0.00264809f $X=1.52 $Y=1.86 $X2=0
+ $Y2=0
cc_566 N_A_299_47#_c_631_n N_A_193_47#_c_856_n 0.0272627f $X=1.625 $Y=2.175
+ $X2=0 $Y2=0
cc_567 N_A_299_47#_c_634_n N_A_193_47#_c_856_n 0.0158156f $X=1.572 $Y=1.967
+ $X2=0 $Y2=0
cc_568 N_A_299_47#_c_639_n N_VPWR_M1024_d 0.00416053f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_569 N_A_299_47#_c_639_n N_VPWR_c_1458_n 0.0128774f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_570 N_A_299_47#_c_646_n N_VPWR_c_1458_n 0.00232703f $X=2.205 $Y=1.967 $X2=0
+ $Y2=0
cc_571 N_A_299_47#_c_631_n N_VPWR_c_1469_n 0.0168466f $X=1.625 $Y=2.175 $X2=0
+ $Y2=0
cc_572 N_A_299_47#_c_639_n N_VPWR_c_1469_n 0.00240758f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_573 N_A_299_47#_M1007_g N_VPWR_c_1470_n 0.00368123f $X=3.14 $Y=2.165 $X2=0
+ $Y2=0
cc_574 N_A_299_47#_c_641_n N_VPWR_c_1470_n 0.00594978f $X=3.075 $Y=1.967 $X2=0
+ $Y2=0
cc_575 N_A_299_47#_c_646_n N_VPWR_c_1470_n 0.00138725f $X=2.205 $Y=1.967 $X2=0
+ $Y2=0
cc_576 N_A_299_47#_M1024_s N_VPWR_c_1456_n 0.00184114f $X=1.5 $Y=1.845 $X2=0
+ $Y2=0
cc_577 N_A_299_47#_M1007_g N_VPWR_c_1456_n 0.00535446f $X=3.14 $Y=2.165 $X2=0
+ $Y2=0
cc_578 N_A_299_47#_c_631_n N_VPWR_c_1456_n 0.00494372f $X=1.625 $Y=2.175 $X2=0
+ $Y2=0
cc_579 N_A_299_47#_c_639_n N_VPWR_c_1456_n 0.00247958f $X=2.12 $Y=1.967 $X2=0
+ $Y2=0
cc_580 N_A_299_47#_c_641_n N_VPWR_c_1456_n 0.00548208f $X=3.075 $Y=1.967 $X2=0
+ $Y2=0
cc_581 N_A_299_47#_c_646_n N_VPWR_c_1456_n 0.00121488f $X=2.205 $Y=1.967 $X2=0
+ $Y2=0
cc_582 N_A_299_47#_c_641_n A_467_369# 0.00527104f $X=3.075 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_583 N_A_299_47#_c_641_n N_A_559_369#_M1016_d 0.00427378f $X=3.075 $Y=1.967
+ $X2=0 $Y2=0
cc_584 N_A_299_47#_M1007_g N_A_559_369#_c_1632_n 0.00811134f $X=3.14 $Y=2.165
+ $X2=0 $Y2=0
cc_585 N_A_299_47#_c_641_n N_A_559_369#_c_1632_n 0.0265702f $X=3.075 $Y=1.967
+ $X2=0 $Y2=0
cc_586 N_A_299_47#_c_636_n N_A_559_369#_c_1632_n 0.0012413f $X=3.185 $Y=1.52
+ $X2=0 $Y2=0
cc_587 N_A_299_47#_M1007_g N_A_559_369#_c_1656_n 0.00367162f $X=3.14 $Y=2.165
+ $X2=0 $Y2=0
cc_588 N_A_299_47#_M1007_g N_A_559_369#_c_1629_n 5.41855e-19 $X=3.14 $Y=2.165
+ $X2=0 $Y2=0
cc_589 N_A_299_47#_c_641_n N_A_559_369#_c_1629_n 0.00683183f $X=3.075 $Y=1.967
+ $X2=0 $Y2=0
cc_590 N_A_299_47#_c_633_n N_A_559_369#_c_1629_n 0.00221463f $X=3.16 $Y=1.86
+ $X2=0 $Y2=0
cc_591 N_A_299_47#_c_626_n N_VGND_c_1773_n 0.002159f $X=1.64 $Y=0.36 $X2=0 $Y2=0
cc_592 N_A_299_47#_M1021_g N_VGND_c_1774_n 0.00775696f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_593 N_A_299_47#_c_626_n N_VGND_c_1784_n 0.0193961f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_594 N_A_299_47#_M1021_g N_VGND_c_1785_n 0.00351072f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_595 N_A_299_47#_M1032_s N_VGND_c_1794_n 0.00183934f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_596 N_A_299_47#_M1021_g N_VGND_c_1794_n 0.00382755f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_597 N_A_299_47#_c_626_n N_VGND_c_1794_n 0.00613328f $X=1.64 $Y=0.36 $X2=0
+ $Y2=0
cc_598 N_D_M1022_g N_SCD_M1020_g 0.00527618f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_599 N_D_M1022_g N_A_193_47#_c_853_n 0.00435792f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_600 N_D_c_754_n N_A_193_47#_c_853_n 0.00255857f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_601 N_D_c_755_n N_A_193_47#_c_853_n 0.00705029f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_602 N_D_M1016_g N_VPWR_c_1458_n 0.00181264f $X=2.72 $Y=2.165 $X2=0 $Y2=0
cc_603 N_D_M1016_g N_VPWR_c_1470_n 0.00385655f $X=2.72 $Y=2.165 $X2=0 $Y2=0
cc_604 N_D_M1016_g N_VPWR_c_1456_n 0.00546011f $X=2.72 $Y=2.165 $X2=0 $Y2=0
cc_605 N_D_M1016_g N_A_559_369#_c_1632_n 0.0061739f $X=2.72 $Y=2.165 $X2=0 $Y2=0
cc_606 N_D_M1022_g N_VGND_c_1774_n 0.00140249f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_607 N_D_M1022_g N_VGND_c_1785_n 0.00422112f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_608 N_D_M1022_g N_VGND_c_1794_n 0.0056538f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_609 N_SCD_M1020_g N_A_193_47#_c_853_n 0.00244488f $X=3.605 $Y=0.445 $X2=0
+ $Y2=0
cc_610 SCD N_A_193_47#_c_853_n 0.012926f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_611 N_SCD_M1005_g N_VPWR_c_1459_n 0.00615911f $X=3.605 $Y=2.165 $X2=0 $Y2=0
cc_612 N_SCD_M1005_g N_VPWR_c_1470_n 0.00412211f $X=3.605 $Y=2.165 $X2=0 $Y2=0
cc_613 N_SCD_M1005_g N_VPWR_c_1456_n 0.00690372f $X=3.605 $Y=2.165 $X2=0 $Y2=0
cc_614 N_SCD_M1005_g N_A_559_369#_c_1632_n 0.00494628f $X=3.605 $Y=2.165 $X2=0
+ $Y2=0
cc_615 N_SCD_M1020_g N_A_559_369#_c_1644_n 0.00444746f $X=3.605 $Y=0.445 $X2=0
+ $Y2=0
cc_616 N_SCD_M1005_g N_A_559_369#_c_1656_n 0.00680709f $X=3.605 $Y=2.165 $X2=0
+ $Y2=0
cc_617 N_SCD_M1020_g N_A_559_369#_c_1621_n 0.00632492f $X=3.605 $Y=0.445 $X2=0
+ $Y2=0
cc_618 N_SCD_M1005_g N_A_559_369#_c_1628_n 0.00857305f $X=3.605 $Y=2.165 $X2=0
+ $Y2=0
cc_619 SCD N_A_559_369#_c_1628_n 0.0307973f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_620 N_SCD_c_802_n N_A_559_369#_c_1628_n 5.47062e-19 $X=3.665 $Y=1.355 $X2=0
+ $Y2=0
cc_621 N_SCD_M1005_g N_A_559_369#_c_1629_n 0.00252323f $X=3.605 $Y=2.165 $X2=0
+ $Y2=0
cc_622 SCD N_A_559_369#_c_1629_n 0.00360851f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_623 N_SCD_M1020_g N_A_559_369#_c_1622_n 0.00825998f $X=3.605 $Y=0.445 $X2=0
+ $Y2=0
cc_624 SCD N_A_559_369#_c_1622_n 0.0302838f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_625 N_SCD_c_802_n N_A_559_369#_c_1622_n 5.22038e-19 $X=3.665 $Y=1.355 $X2=0
+ $Y2=0
cc_626 N_SCD_M1020_g N_A_559_369#_c_1623_n 0.00227426f $X=3.605 $Y=0.445 $X2=0
+ $Y2=0
cc_627 SCD N_A_559_369#_c_1623_n 0.00391935f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_628 N_SCD_M1020_g N_A_559_369#_c_1624_n 0.0021982f $X=3.605 $Y=0.445 $X2=0
+ $Y2=0
cc_629 N_SCD_M1020_g N_A_559_369#_c_1625_n 0.00402041f $X=3.605 $Y=0.445 $X2=0
+ $Y2=0
cc_630 N_SCD_M1005_g N_A_559_369#_c_1625_n 0.00422492f $X=3.605 $Y=2.165 $X2=0
+ $Y2=0
cc_631 SCD N_A_559_369#_c_1625_n 0.0469263f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_632 N_SCD_c_802_n N_A_559_369#_c_1625_n 0.00140293f $X=3.665 $Y=1.355 $X2=0
+ $Y2=0
cc_633 N_SCD_M1005_g N_A_559_369#_c_1631_n 0.00281601f $X=3.605 $Y=2.165 $X2=0
+ $Y2=0
cc_634 N_SCD_M1020_g N_VGND_c_1775_n 0.00562907f $X=3.605 $Y=0.445 $X2=0 $Y2=0
cc_635 N_SCD_M1020_g N_VGND_c_1785_n 0.00404961f $X=3.605 $Y=0.445 $X2=0 $Y2=0
cc_636 N_SCD_M1020_g N_VGND_c_1794_n 0.00665506f $X=3.605 $Y=0.445 $X2=0 $Y2=0
cc_637 N_A_193_47#_c_852_n N_A_1098_183#_M1017_d 0.00133652f $X=6.97 $Y=0.87
+ $X2=-0.19 $Y2=-0.24
cc_638 N_A_193_47#_c_855_n N_A_1098_183#_M1017_d 9.65449e-19 $X=6.57 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_639 N_A_193_47#_c_857_n N_A_1098_183#_M1017_d 6.4695e-19 $X=6.715 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_640 N_A_193_47#_c_855_n N_A_1098_183#_M1023_g 0.00208483f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_641 N_A_193_47#_c_860_n N_A_1098_183#_M1023_g 0.013781f $X=5.045 $Y=0.705
+ $X2=0 $Y2=0
cc_642 N_A_193_47#_c_855_n N_A_1098_183#_c_1067_n 0.0221014f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_643 N_A_193_47#_c_857_n N_A_1098_183#_c_1093_n 8.93965e-19 $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_644 N_A_193_47#_c_852_n N_A_1098_183#_c_1094_n 0.00716698f $X=6.97 $Y=0.87
+ $X2=0 $Y2=0
cc_645 N_A_193_47#_c_855_n N_A_1098_183#_c_1094_n 0.00363224f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_646 N_A_193_47#_c_857_n N_A_1098_183#_c_1094_n 0.00168986f $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_647 N_A_193_47#_c_855_n N_A_1098_183#_c_1068_n 0.00899288f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_648 N_A_193_47#_c_850_n N_A_1098_183#_c_1069_n 0.00114045f $X=7.065 $Y=1.575
+ $X2=0 $Y2=0
cc_649 N_A_193_47#_c_852_n N_A_1098_183#_c_1069_n 0.018732f $X=6.97 $Y=0.87
+ $X2=0 $Y2=0
cc_650 N_A_193_47#_c_855_n N_A_1098_183#_c_1069_n 0.0176435f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_651 N_A_193_47#_c_857_n N_A_1098_183#_c_1069_n 0.00185392f $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_652 N_A_193_47#_c_861_n N_A_1098_183#_c_1069_n 5.82389e-19 $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_653 N_A_193_47#_c_850_n N_A_1098_183#_c_1070_n 0.00620052f $X=7.065 $Y=1.575
+ $X2=0 $Y2=0
cc_654 N_A_193_47#_c_855_n N_A_1098_183#_c_1071_n 0.00299829f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_655 N_A_193_47#_c_858_n N_A_1098_183#_c_1071_n 0.0179412f $X=5.045 $Y=0.87
+ $X2=0 $Y2=0
cc_656 N_A_193_47#_c_850_n N_A_939_413#_c_1160_n 6.31337e-19 $X=7.065 $Y=1.575
+ $X2=0 $Y2=0
cc_657 N_A_193_47#_c_848_n N_A_939_413#_c_1161_n 0.00957285f $X=6.83 $Y=0.705
+ $X2=0 $Y2=0
cc_658 N_A_193_47#_c_852_n N_A_939_413#_c_1161_n 0.00100831f $X=6.97 $Y=0.87
+ $X2=0 $Y2=0
cc_659 N_A_193_47#_c_850_n N_A_939_413#_c_1162_n 3.37852e-19 $X=7.065 $Y=1.575
+ $X2=0 $Y2=0
cc_660 N_A_193_47#_c_861_n N_A_939_413#_c_1162_n 0.00957285f $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_661 N_A_193_47#_M1008_g N_A_939_413#_c_1178_n 0.00188835f $X=4.62 $Y=2.275
+ $X2=0 $Y2=0
cc_662 N_A_193_47#_c_849_n N_A_939_413#_c_1178_n 0.00286257f $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_663 N_A_193_47#_c_865_n N_A_939_413#_c_1178_n 6.94615e-19 $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_664 N_A_193_47#_c_855_n N_A_939_413#_c_1204_n 0.00506965f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_665 N_A_193_47#_c_989_p N_A_939_413#_c_1204_n 0.00100579f $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_666 N_A_193_47#_c_858_n N_A_939_413#_c_1204_n 0.00256542f $X=5.045 $Y=0.87
+ $X2=0 $Y2=0
cc_667 N_A_193_47#_c_859_n N_A_939_413#_c_1204_n 0.0237558f $X=5.045 $Y=0.87
+ $X2=0 $Y2=0
cc_668 N_A_193_47#_c_860_n N_A_939_413#_c_1204_n 0.00840911f $X=5.045 $Y=0.705
+ $X2=0 $Y2=0
cc_669 N_A_193_47#_c_849_n N_A_939_413#_c_1165_n 0.00981359f $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_670 N_A_193_47#_c_855_n N_A_939_413#_c_1165_n 0.0188221f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_671 N_A_193_47#_c_989_p N_A_939_413#_c_1165_n 4.66512e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_672 N_A_193_47#_c_859_n N_A_939_413#_c_1165_n 0.0239925f $X=5.045 $Y=0.87
+ $X2=0 $Y2=0
cc_673 N_A_193_47#_c_860_n N_A_939_413#_c_1165_n 0.00604394f $X=5.045 $Y=0.705
+ $X2=0 $Y2=0
cc_674 N_A_193_47#_c_849_n N_A_939_413#_c_1166_n 0.00649323f $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_675 N_A_193_47#_c_855_n N_A_939_413#_c_1166_n 0.00803733f $X=6.57 $Y=0.85
+ $X2=0 $Y2=0
cc_676 N_A_193_47#_M1000_g N_A_1526_315#_c_1281_n 0.018025f $X=7.12 $Y=2.275
+ $X2=0 $Y2=0
cc_677 N_A_193_47#_c_868_n N_A_1526_315#_c_1281_n 0.0119764f $X=7.205 $Y=1.74
+ $X2=0 $Y2=0
cc_678 N_A_193_47#_M1000_g N_A_1355_413#_c_1380_n 0.00974744f $X=7.12 $Y=2.275
+ $X2=0 $Y2=0
cc_679 N_A_193_47#_c_867_n N_A_1355_413#_c_1380_n 0.012999f $X=7.205 $Y=1.74
+ $X2=0 $Y2=0
cc_680 N_A_193_47#_c_868_n N_A_1355_413#_c_1380_n 0.00300896f $X=7.205 $Y=1.74
+ $X2=0 $Y2=0
cc_681 N_A_193_47#_c_852_n N_A_1355_413#_c_1383_n 0.0153172f $X=6.97 $Y=0.87
+ $X2=0 $Y2=0
cc_682 N_A_193_47#_c_861_n N_A_1355_413#_c_1383_n 8.54271e-19 $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_683 N_A_193_47#_M1000_g N_A_1355_413#_c_1377_n 0.0046302f $X=7.12 $Y=2.275
+ $X2=0 $Y2=0
cc_684 N_A_193_47#_c_850_n N_A_1355_413#_c_1377_n 0.00868218f $X=7.065 $Y=1.575
+ $X2=0 $Y2=0
cc_685 N_A_193_47#_c_867_n N_A_1355_413#_c_1377_n 0.0246912f $X=7.205 $Y=1.74
+ $X2=0 $Y2=0
cc_686 N_A_193_47#_c_868_n N_A_1355_413#_c_1377_n 0.00187857f $X=7.205 $Y=1.74
+ $X2=0 $Y2=0
cc_687 N_A_193_47#_c_850_n N_A_1355_413#_c_1372_n 0.0272384f $X=7.065 $Y=1.575
+ $X2=0 $Y2=0
cc_688 N_A_193_47#_c_868_n N_A_1355_413#_c_1372_n 0.00102186f $X=7.205 $Y=1.74
+ $X2=0 $Y2=0
cc_689 N_A_193_47#_c_848_n N_A_1355_413#_c_1373_n 8.96907e-19 $X=6.83 $Y=0.705
+ $X2=0 $Y2=0
cc_690 N_A_193_47#_c_852_n N_A_1355_413#_c_1373_n 0.025625f $X=6.97 $Y=0.87
+ $X2=0 $Y2=0
cc_691 N_A_193_47#_c_857_n N_A_1355_413#_c_1373_n 8.16973e-19 $X=6.715 $Y=0.85
+ $X2=0 $Y2=0
cc_692 N_A_193_47#_c_861_n N_A_1355_413#_c_1373_n 3.08898e-19 $X=6.925 $Y=0.87
+ $X2=0 $Y2=0
cc_693 N_A_193_47#_c_856_n N_VPWR_c_1457_n 0.0127357f $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_694 N_A_193_47#_c_856_n N_VPWR_c_1458_n 5.63902e-19 $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_695 N_A_193_47#_M1008_g N_VPWR_c_1459_n 0.00262954f $X=4.62 $Y=2.275 $X2=0
+ $Y2=0
cc_696 N_A_193_47#_M1008_g N_VPWR_c_1466_n 0.005785f $X=4.62 $Y=2.275 $X2=0
+ $Y2=0
cc_697 N_A_193_47#_c_856_n N_VPWR_c_1469_n 0.015988f $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_698 N_A_193_47#_M1000_g N_VPWR_c_1471_n 0.00383564f $X=7.12 $Y=2.275 $X2=0
+ $Y2=0
cc_699 N_A_193_47#_M1008_g N_VPWR_c_1456_n 0.00734982f $X=4.62 $Y=2.275 $X2=0
+ $Y2=0
cc_700 N_A_193_47#_M1000_g N_VPWR_c_1456_n 0.00579176f $X=7.12 $Y=2.275 $X2=0
+ $Y2=0
cc_701 N_A_193_47#_c_849_n N_VPWR_c_1456_n 0.00189161f $X=4.635 $Y=1.74 $X2=0
+ $Y2=0
cc_702 N_A_193_47#_c_865_n N_VPWR_c_1456_n 4.15345e-19 $X=4.635 $Y=1.74 $X2=0
+ $Y2=0
cc_703 N_A_193_47#_c_856_n N_VPWR_c_1456_n 0.00409094f $X=1.135 $Y=0.85 $X2=0
+ $Y2=0
cc_704 N_A_193_47#_c_853_n N_A_559_369#_c_1644_n 0.00536043f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_705 N_A_193_47#_c_853_n N_A_559_369#_c_1622_n 0.0220682f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_706 N_A_193_47#_c_853_n N_A_559_369#_c_1623_n 0.00970914f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_707 N_A_193_47#_c_849_n N_A_559_369#_c_1625_n 0.058581f $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_708 N_A_193_47#_c_865_n N_A_559_369#_c_1625_n 0.0052844f $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_709 N_A_193_47#_c_853_n N_A_559_369#_c_1625_n 0.0123751f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_710 N_A_193_47#_c_989_p N_A_559_369#_c_1625_n 2.43115e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_711 N_A_193_47#_c_859_n N_A_559_369#_c_1625_n 0.012499f $X=5.045 $Y=0.87
+ $X2=0 $Y2=0
cc_712 N_A_193_47#_c_853_n N_A_559_369#_c_1626_n 0.00506513f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_713 N_A_193_47#_c_859_n N_A_559_369#_c_1626_n 6.01474e-19 $X=5.045 $Y=0.87
+ $X2=0 $Y2=0
cc_714 N_A_193_47#_c_853_n N_A_559_369#_c_1627_n 0.00562077f $X=4.685 $Y=0.85
+ $X2=0 $Y2=0
cc_715 N_A_193_47#_c_989_p N_A_559_369#_c_1627_n 2.74809e-19 $X=4.975 $Y=0.85
+ $X2=0 $Y2=0
cc_716 N_A_193_47#_c_859_n N_A_559_369#_c_1627_n 0.0122359f $X=5.045 $Y=0.87
+ $X2=0 $Y2=0
cc_717 N_A_193_47#_M1008_g N_A_559_369#_c_1631_n 0.00994993f $X=4.62 $Y=2.275
+ $X2=0 $Y2=0
cc_718 N_A_193_47#_c_849_n N_A_559_369#_c_1631_n 0.00558861f $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_719 N_A_193_47#_c_865_n N_A_559_369#_c_1631_n 9.82843e-19 $X=4.635 $Y=1.74
+ $X2=0 $Y2=0
cc_720 N_A_193_47#_c_853_n N_VGND_c_1774_n 0.00117841f $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_721 N_A_193_47#_c_853_n N_VGND_c_1775_n 8.73533e-19 $X=4.685 $Y=0.85 $X2=0
+ $Y2=0
cc_722 N_A_193_47#_c_859_n N_VGND_c_1776_n 0.00254426f $X=5.045 $Y=0.87 $X2=0
+ $Y2=0
cc_723 N_A_193_47#_c_860_n N_VGND_c_1776_n 0.0037981f $X=5.045 $Y=0.705 $X2=0
+ $Y2=0
cc_724 N_A_193_47#_c_855_n N_VGND_c_1777_n 0.00197288f $X=6.57 $Y=0.85 $X2=0
+ $Y2=0
cc_725 N_A_193_47#_c_851_n N_VGND_c_1784_n 0.0100142f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_726 N_A_193_47#_c_848_n N_VGND_c_1786_n 0.00435108f $X=6.83 $Y=0.705 $X2=0
+ $Y2=0
cc_727 N_A_193_47#_c_852_n N_VGND_c_1786_n 0.00341023f $X=6.97 $Y=0.87 $X2=0
+ $Y2=0
cc_728 N_A_193_47#_c_861_n N_VGND_c_1786_n 8.04624e-19 $X=6.925 $Y=0.87 $X2=0
+ $Y2=0
cc_729 N_A_193_47#_M1018_d N_VGND_c_1794_n 0.00281453f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_730 N_A_193_47#_c_848_n N_VGND_c_1794_n 0.00623562f $X=6.83 $Y=0.705 $X2=0
+ $Y2=0
cc_731 N_A_193_47#_c_851_n N_VGND_c_1794_n 0.00380969f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_732 N_A_193_47#_c_852_n N_VGND_c_1794_n 0.00402561f $X=6.97 $Y=0.87 $X2=0
+ $Y2=0
cc_733 N_A_193_47#_c_853_n N_VGND_c_1794_n 0.1569f $X=4.685 $Y=0.85 $X2=0 $Y2=0
cc_734 N_A_193_47#_c_854_n N_VGND_c_1794_n 0.0151167f $X=1.28 $Y=0.85 $X2=0
+ $Y2=0
cc_735 N_A_193_47#_c_855_n N_VGND_c_1794_n 0.0732377f $X=6.57 $Y=0.85 $X2=0
+ $Y2=0
cc_736 N_A_193_47#_c_989_p N_VGND_c_1794_n 0.0146263f $X=4.975 $Y=0.85 $X2=0
+ $Y2=0
cc_737 N_A_193_47#_c_857_n N_VGND_c_1794_n 0.0147739f $X=6.715 $Y=0.85 $X2=0
+ $Y2=0
cc_738 N_A_193_47#_c_859_n N_VGND_c_1794_n 0.00247098f $X=5.045 $Y=0.87 $X2=0
+ $Y2=0
cc_739 N_A_193_47#_c_860_n N_VGND_c_1794_n 0.00563926f $X=5.045 $Y=0.705 $X2=0
+ $Y2=0
cc_740 N_A_193_47#_c_861_n N_VGND_c_1794_n 0.00134095f $X=6.925 $Y=0.87 $X2=0
+ $Y2=0
cc_741 N_A_1098_183#_c_1070_n N_A_939_413#_c_1160_n 0.00595764f $X=6.395
+ $Y=2.135 $X2=0 $Y2=0
cc_742 N_A_1098_183#_M1006_g N_A_939_413#_M1025_g 0.0139082f $X=5.565 $Y=2.275
+ $X2=0 $Y2=0
cc_743 N_A_1098_183#_c_1081_n N_A_939_413#_M1025_g 0.00378805f $X=6.435 $Y=2.3
+ $X2=0 $Y2=0
cc_744 N_A_1098_183#_c_1070_n N_A_939_413#_M1025_g 0.0122998f $X=6.395 $Y=2.135
+ $X2=0 $Y2=0
cc_745 N_A_1098_183#_M1023_g N_A_939_413#_c_1161_n 0.0109128f $X=5.595 $Y=0.445
+ $X2=0 $Y2=0
cc_746 N_A_1098_183#_c_1067_n N_A_939_413#_c_1161_n 0.00351053f $X=6.27 $Y=0.915
+ $X2=0 $Y2=0
cc_747 N_A_1098_183#_c_1093_n N_A_939_413#_c_1161_n 0.00675936f $X=6.355
+ $Y=0.765 $X2=0 $Y2=0
cc_748 N_A_1098_183#_c_1113_p N_A_939_413#_c_1161_n 0.004701f $X=6.44 $Y=0.45
+ $X2=0 $Y2=0
cc_749 N_A_1098_183#_c_1069_n N_A_939_413#_c_1161_n 0.00333126f $X=6.355
+ $Y=0.915 $X2=0 $Y2=0
cc_750 N_A_1098_183#_c_1071_n N_A_939_413#_c_1161_n 0.00500517f $X=5.595 $Y=0.93
+ $X2=0 $Y2=0
cc_751 N_A_1098_183#_M1006_g N_A_939_413#_c_1162_n 0.00398999f $X=5.565 $Y=2.275
+ $X2=0 $Y2=0
cc_752 N_A_1098_183#_c_1067_n N_A_939_413#_c_1162_n 0.00996228f $X=6.27 $Y=0.915
+ $X2=0 $Y2=0
cc_753 N_A_1098_183#_c_1068_n N_A_939_413#_c_1162_n 2.46578e-19 $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_754 N_A_1098_183#_c_1069_n N_A_939_413#_c_1162_n 0.00234347f $X=6.355
+ $Y=0.915 $X2=0 $Y2=0
cc_755 N_A_1098_183#_c_1070_n N_A_939_413#_c_1162_n 0.00394884f $X=6.395
+ $Y=2.135 $X2=0 $Y2=0
cc_756 N_A_1098_183#_c_1071_n N_A_939_413#_c_1162_n 0.00573363f $X=5.595 $Y=0.93
+ $X2=0 $Y2=0
cc_757 N_A_1098_183#_M1006_g N_A_939_413#_c_1163_n 0.0173592f $X=5.565 $Y=2.275
+ $X2=0 $Y2=0
cc_758 N_A_1098_183#_c_1067_n N_A_939_413#_c_1163_n 0.00400764f $X=6.27 $Y=0.915
+ $X2=0 $Y2=0
cc_759 N_A_1098_183#_c_1071_n N_A_939_413#_c_1163_n 0.00238133f $X=5.595 $Y=0.93
+ $X2=0 $Y2=0
cc_760 N_A_1098_183#_c_1070_n N_A_939_413#_c_1164_n 0.00611615f $X=6.395
+ $Y=2.135 $X2=0 $Y2=0
cc_761 N_A_1098_183#_M1006_g N_A_939_413#_c_1178_n 0.0101048f $X=5.565 $Y=2.275
+ $X2=0 $Y2=0
cc_762 N_A_1098_183#_M1023_g N_A_939_413#_c_1165_n 0.00441151f $X=5.595 $Y=0.445
+ $X2=0 $Y2=0
cc_763 N_A_1098_183#_c_1068_n N_A_939_413#_c_1165_n 0.0243525f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_764 N_A_1098_183#_c_1071_n N_A_939_413#_c_1165_n 0.0095167f $X=5.595 $Y=0.93
+ $X2=0 $Y2=0
cc_765 N_A_1098_183#_M1006_g N_A_939_413#_c_1170_n 0.0153788f $X=5.565 $Y=2.275
+ $X2=0 $Y2=0
cc_766 N_A_1098_183#_c_1070_n N_A_939_413#_c_1170_n 0.00754007f $X=6.395
+ $Y=2.135 $X2=0 $Y2=0
cc_767 N_A_1098_183#_M1006_g N_A_939_413#_c_1166_n 0.0138593f $X=5.565 $Y=2.275
+ $X2=0 $Y2=0
cc_768 N_A_1098_183#_c_1067_n N_A_939_413#_c_1166_n 0.0186614f $X=6.27 $Y=0.915
+ $X2=0 $Y2=0
cc_769 N_A_1098_183#_c_1068_n N_A_939_413#_c_1166_n 0.0112018f $X=5.81 $Y=0.93
+ $X2=0 $Y2=0
cc_770 N_A_1098_183#_c_1070_n N_A_939_413#_c_1166_n 0.0245884f $X=6.395 $Y=2.135
+ $X2=0 $Y2=0
cc_771 N_A_1098_183#_c_1071_n N_A_939_413#_c_1166_n 0.00213749f $X=5.595 $Y=0.93
+ $X2=0 $Y2=0
cc_772 N_A_1098_183#_c_1081_n N_A_1355_413#_c_1380_n 0.0109209f $X=6.435 $Y=2.3
+ $X2=0 $Y2=0
cc_773 N_A_1098_183#_M1006_g N_VPWR_c_1460_n 0.0057281f $X=5.565 $Y=2.275 $X2=0
+ $Y2=0
cc_774 N_A_1098_183#_c_1070_n N_VPWR_c_1460_n 0.0237f $X=6.395 $Y=2.135 $X2=0
+ $Y2=0
cc_775 N_A_1098_183#_M1006_g N_VPWR_c_1466_n 0.00378797f $X=5.565 $Y=2.275 $X2=0
+ $Y2=0
cc_776 N_A_1098_183#_c_1081_n N_VPWR_c_1471_n 0.015079f $X=6.435 $Y=2.3 $X2=0
+ $Y2=0
cc_777 N_A_1098_183#_M1025_d N_VPWR_c_1456_n 0.00285154f $X=6.3 $Y=1.735 $X2=0
+ $Y2=0
cc_778 N_A_1098_183#_M1006_g N_VPWR_c_1456_n 0.00596544f $X=5.565 $Y=2.275 $X2=0
+ $Y2=0
cc_779 N_A_1098_183#_c_1081_n N_VPWR_c_1456_n 0.00439826f $X=6.435 $Y=2.3 $X2=0
+ $Y2=0
cc_780 N_A_1098_183#_c_1067_n N_VGND_M1023_d 0.00306998f $X=6.27 $Y=0.915 $X2=0
+ $Y2=0
cc_781 N_A_1098_183#_M1023_g N_VGND_c_1776_n 0.00585385f $X=5.595 $Y=0.445 $X2=0
+ $Y2=0
cc_782 N_A_1098_183#_M1023_g N_VGND_c_1777_n 0.00603751f $X=5.595 $Y=0.445 $X2=0
+ $Y2=0
cc_783 N_A_1098_183#_c_1093_n N_VGND_c_1777_n 0.00354103f $X=6.355 $Y=0.765
+ $X2=0 $Y2=0
cc_784 N_A_1098_183#_c_1113_p N_VGND_c_1777_n 0.013122f $X=6.44 $Y=0.45 $X2=0
+ $Y2=0
cc_785 N_A_1098_183#_c_1068_n N_VGND_c_1777_n 0.0258565f $X=5.81 $Y=0.93 $X2=0
+ $Y2=0
cc_786 N_A_1098_183#_c_1071_n N_VGND_c_1777_n 0.00122075f $X=5.595 $Y=0.93 $X2=0
+ $Y2=0
cc_787 N_A_1098_183#_c_1113_p N_VGND_c_1786_n 0.00594819f $X=6.44 $Y=0.45 $X2=0
+ $Y2=0
cc_788 N_A_1098_183#_c_1094_n N_VGND_c_1786_n 0.0100275f $X=6.565 $Y=0.45 $X2=0
+ $Y2=0
cc_789 N_A_1098_183#_M1017_d N_VGND_c_1794_n 0.00246577f $X=6.4 $Y=0.235 $X2=0
+ $Y2=0
cc_790 N_A_1098_183#_M1023_g N_VGND_c_1794_n 0.0070154f $X=5.595 $Y=0.445 $X2=0
+ $Y2=0
cc_791 N_A_1098_183#_c_1067_n N_VGND_c_1794_n 0.0042145f $X=6.27 $Y=0.915 $X2=0
+ $Y2=0
cc_792 N_A_1098_183#_c_1113_p N_VGND_c_1794_n 0.00261981f $X=6.44 $Y=0.45 $X2=0
+ $Y2=0
cc_793 N_A_1098_183#_c_1094_n N_VGND_c_1794_n 0.00441842f $X=6.565 $Y=0.45 $X2=0
+ $Y2=0
cc_794 N_A_1098_183#_c_1068_n N_VGND_c_1794_n 0.00269026f $X=5.81 $Y=0.93 $X2=0
+ $Y2=0
cc_795 N_A_939_413#_c_1178_n N_VPWR_M1006_d 0.00236303f $X=5.59 $Y=2.275 $X2=0
+ $Y2=0
cc_796 N_A_939_413#_c_1170_n N_VPWR_M1006_d 0.00412006f $X=5.675 $Y=2.19 $X2=0
+ $Y2=0
cc_797 N_A_939_413#_M1025_g N_VPWR_c_1460_n 0.00314007f $X=6.225 $Y=2.11 $X2=0
+ $Y2=0
cc_798 N_A_939_413#_c_1163_n N_VPWR_c_1460_n 9.53331e-19 $X=6.15 $Y=1.41 $X2=0
+ $Y2=0
cc_799 N_A_939_413#_c_1178_n N_VPWR_c_1460_n 0.0138309f $X=5.59 $Y=2.275 $X2=0
+ $Y2=0
cc_800 N_A_939_413#_c_1170_n N_VPWR_c_1460_n 0.0252383f $X=5.675 $Y=2.19 $X2=0
+ $Y2=0
cc_801 N_A_939_413#_c_1166_n N_VPWR_c_1460_n 0.00741701f $X=5.675 $Y=1.41 $X2=0
+ $Y2=0
cc_802 N_A_939_413#_c_1178_n N_VPWR_c_1466_n 0.0359536f $X=5.59 $Y=2.275 $X2=0
+ $Y2=0
cc_803 N_A_939_413#_M1025_g N_VPWR_c_1471_n 0.00541359f $X=6.225 $Y=2.11 $X2=0
+ $Y2=0
cc_804 N_A_939_413#_M1008_d N_VPWR_c_1456_n 0.00217001f $X=4.695 $Y=2.065 $X2=0
+ $Y2=0
cc_805 N_A_939_413#_M1025_g N_VPWR_c_1456_n 0.00665748f $X=6.225 $Y=2.11 $X2=0
+ $Y2=0
cc_806 N_A_939_413#_c_1178_n N_VPWR_c_1456_n 0.0161666f $X=5.59 $Y=2.275 $X2=0
+ $Y2=0
cc_807 N_A_939_413#_c_1178_n N_A_559_369#_c_1631_n 0.0102204f $X=5.59 $Y=2.275
+ $X2=0 $Y2=0
cc_808 N_A_939_413#_c_1178_n A_1032_413# 0.0045944f $X=5.59 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_809 N_A_939_413#_c_1204_n N_VGND_c_1776_n 0.0255873f $X=5.3 $Y=0.45 $X2=0
+ $Y2=0
cc_810 N_A_939_413#_c_1161_n N_VGND_c_1777_n 0.00816054f $X=6.325 $Y=0.95 $X2=0
+ $Y2=0
cc_811 N_A_939_413#_c_1161_n N_VGND_c_1786_n 0.00407056f $X=6.325 $Y=0.95 $X2=0
+ $Y2=0
cc_812 N_A_939_413#_M1028_d N_VGND_c_1794_n 0.00228264f $X=4.7 $Y=0.235 $X2=0
+ $Y2=0
cc_813 N_A_939_413#_c_1161_n N_VGND_c_1794_n 0.00620172f $X=6.325 $Y=0.95 $X2=0
+ $Y2=0
cc_814 N_A_939_413#_c_1204_n N_VGND_c_1794_n 0.0113257f $X=5.3 $Y=0.45 $X2=0
+ $Y2=0
cc_815 N_A_939_413#_c_1204_n A_1036_47# 0.00455507f $X=5.3 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_816 N_A_939_413#_c_1165_n A_1036_47# 0.00200718f $X=5.385 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_817 N_A_1526_315#_c_1270_n N_A_1355_413#_c_1368_n 0.0193264f $X=9.215
+ $Y=0.995 $X2=0 $Y2=0
cc_818 N_A_1526_315#_c_1272_n N_A_1355_413#_c_1368_n 0.00505396f $X=8.65
+ $Y=0.995 $X2=0 $Y2=0
cc_819 N_A_1526_315#_c_1274_n N_A_1355_413#_c_1368_n 0.00768498f $X=8.55
+ $Y=0.385 $X2=0 $Y2=0
cc_820 N_A_1526_315#_M1010_g N_A_1355_413#_M1002_g 0.0196417f $X=9.215 $Y=1.985
+ $X2=0 $Y2=0
cc_821 N_A_1526_315#_c_1281_n N_A_1355_413#_M1002_g 0.00198604f $X=7.885 $Y=1.74
+ $X2=0 $Y2=0
cc_822 N_A_1526_315#_c_1293_p N_A_1355_413#_M1002_g 0.0104955f $X=8.55 $Y=2.29
+ $X2=0 $Y2=0
cc_823 N_A_1526_315#_c_1282_n N_A_1355_413#_M1002_g 0.00742753f $X=8.65 $Y=1.575
+ $X2=0 $Y2=0
cc_824 N_A_1526_315#_c_1295_p N_A_1355_413#_M1002_g 0.00489897f $X=8.55 $Y=1.68
+ $X2=0 $Y2=0
cc_825 N_A_1526_315#_M1027_g N_A_1355_413#_c_1369_n 0.0149936f $X=7.82 $Y=0.445
+ $X2=0 $Y2=0
cc_826 N_A_1526_315#_c_1280_n N_A_1355_413#_c_1369_n 0.00734699f $X=8.465
+ $Y=1.74 $X2=0 $Y2=0
cc_827 N_A_1526_315#_c_1274_n N_A_1355_413#_c_1369_n 0.00747686f $X=8.55
+ $Y=0.385 $X2=0 $Y2=0
cc_828 N_A_1526_315#_c_1295_p N_A_1355_413#_c_1369_n 0.00407845f $X=8.55 $Y=1.68
+ $X2=0 $Y2=0
cc_829 N_A_1526_315#_c_1300_p N_A_1355_413#_c_1369_n 0.01406f $X=8.65 $Y=1.16
+ $X2=0 $Y2=0
cc_830 N_A_1526_315#_c_1273_n N_A_1355_413#_c_1370_n 0.0155195f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_831 N_A_1526_315#_c_1300_p N_A_1355_413#_c_1370_n 0.00155371f $X=8.65 $Y=1.16
+ $X2=0 $Y2=0
cc_832 N_A_1526_315#_c_1275_n N_A_1355_413#_c_1370_n 0.021601f $X=9.635 $Y=1.16
+ $X2=0 $Y2=0
cc_833 N_A_1526_315#_M1019_g N_A_1355_413#_c_1380_n 0.00194535f $X=7.705
+ $Y=2.275 $X2=0 $Y2=0
cc_834 N_A_1526_315#_M1027_g N_A_1355_413#_c_1383_n 0.00114979f $X=7.82 $Y=0.445
+ $X2=0 $Y2=0
cc_835 N_A_1526_315#_c_1280_n N_A_1355_413#_c_1377_n 0.0262086f $X=8.465 $Y=1.74
+ $X2=0 $Y2=0
cc_836 N_A_1526_315#_c_1281_n N_A_1355_413#_c_1377_n 0.00865902f $X=7.885
+ $Y=1.74 $X2=0 $Y2=0
cc_837 N_A_1526_315#_M1027_g N_A_1355_413#_c_1371_n 0.018366f $X=7.82 $Y=0.445
+ $X2=0 $Y2=0
cc_838 N_A_1526_315#_c_1280_n N_A_1355_413#_c_1371_n 0.0355898f $X=8.465 $Y=1.74
+ $X2=0 $Y2=0
cc_839 N_A_1526_315#_c_1281_n N_A_1355_413#_c_1371_n 0.00739167f $X=7.885
+ $Y=1.74 $X2=0 $Y2=0
cc_840 N_A_1526_315#_c_1274_n N_A_1355_413#_c_1371_n 7.42989e-19 $X=8.55
+ $Y=0.385 $X2=0 $Y2=0
cc_841 N_A_1526_315#_c_1300_p N_A_1355_413#_c_1371_n 0.0278269f $X=8.65 $Y=1.16
+ $X2=0 $Y2=0
cc_842 N_A_1526_315#_M1027_g N_A_1355_413#_c_1372_n 0.00880678f $X=7.82 $Y=0.445
+ $X2=0 $Y2=0
cc_843 N_A_1526_315#_M1027_g N_A_1355_413#_c_1373_n 0.00779225f $X=7.82 $Y=0.445
+ $X2=0 $Y2=0
cc_844 N_A_1526_315#_M1019_g N_VPWR_c_1461_n 0.0115962f $X=7.705 $Y=2.275 $X2=0
+ $Y2=0
cc_845 N_A_1526_315#_c_1280_n N_VPWR_c_1461_n 0.0182102f $X=8.465 $Y=1.74 $X2=0
+ $Y2=0
cc_846 N_A_1526_315#_c_1281_n N_VPWR_c_1461_n 0.0049226f $X=7.885 $Y=1.74 $X2=0
+ $Y2=0
cc_847 N_A_1526_315#_c_1293_p N_VPWR_c_1461_n 0.014785f $X=8.55 $Y=2.29 $X2=0
+ $Y2=0
cc_848 N_A_1526_315#_c_1293_p N_VPWR_c_1462_n 0.0157187f $X=8.55 $Y=2.29 $X2=0
+ $Y2=0
cc_849 N_A_1526_315#_M1010_g N_VPWR_c_1463_n 0.00715342f $X=9.215 $Y=1.985 $X2=0
+ $Y2=0
cc_850 N_A_1526_315#_c_1293_p N_VPWR_c_1463_n 0.0400358f $X=8.55 $Y=2.29 $X2=0
+ $Y2=0
cc_851 N_A_1526_315#_c_1273_n N_VPWR_c_1463_n 0.00982851f $X=9.18 $Y=1.16 $X2=0
+ $Y2=0
cc_852 N_A_1526_315#_c_1295_p N_VPWR_c_1463_n 0.022052f $X=8.55 $Y=1.68 $X2=0
+ $Y2=0
cc_853 N_A_1526_315#_c_1275_n N_VPWR_c_1463_n 7.34886e-19 $X=9.635 $Y=1.16 $X2=0
+ $Y2=0
cc_854 N_A_1526_315#_M1033_g N_VPWR_c_1465_n 0.0101826f $X=9.635 $Y=1.985 $X2=0
+ $Y2=0
cc_855 N_A_1526_315#_M1019_g N_VPWR_c_1471_n 0.00585385f $X=7.705 $Y=2.275 $X2=0
+ $Y2=0
cc_856 N_A_1526_315#_M1010_g N_VPWR_c_1472_n 0.0054411f $X=9.215 $Y=1.985 $X2=0
+ $Y2=0
cc_857 N_A_1526_315#_M1033_g N_VPWR_c_1472_n 0.00522761f $X=9.635 $Y=1.985 $X2=0
+ $Y2=0
cc_858 N_A_1526_315#_M1002_s N_VPWR_c_1456_n 0.00234057f $X=8.425 $Y=1.485 $X2=0
+ $Y2=0
cc_859 N_A_1526_315#_M1019_g N_VPWR_c_1456_n 0.0124099f $X=7.705 $Y=2.275 $X2=0
+ $Y2=0
cc_860 N_A_1526_315#_M1010_g N_VPWR_c_1456_n 0.00972437f $X=9.215 $Y=1.985 $X2=0
+ $Y2=0
cc_861 N_A_1526_315#_M1033_g N_VPWR_c_1456_n 0.00996308f $X=9.635 $Y=1.985 $X2=0
+ $Y2=0
cc_862 N_A_1526_315#_c_1280_n N_VPWR_c_1456_n 0.0145324f $X=8.465 $Y=1.74 $X2=0
+ $Y2=0
cc_863 N_A_1526_315#_c_1281_n N_VPWR_c_1456_n 7.75814e-19 $X=7.885 $Y=1.74 $X2=0
+ $Y2=0
cc_864 N_A_1526_315#_c_1293_p N_VPWR_c_1456_n 0.00997475f $X=8.55 $Y=2.29 $X2=0
+ $Y2=0
cc_865 N_A_1526_315#_M1010_g N_Q_c_1744_n 0.00414943f $X=9.215 $Y=1.985 $X2=0
+ $Y2=0
cc_866 N_A_1526_315#_M1033_g N_Q_c_1744_n 0.00206615f $X=9.635 $Y=1.985 $X2=0
+ $Y2=0
cc_867 N_A_1526_315#_c_1282_n N_Q_c_1744_n 0.00198007f $X=8.65 $Y=1.575 $X2=0
+ $Y2=0
cc_868 N_A_1526_315#_c_1295_p N_Q_c_1744_n 0.00158627f $X=8.55 $Y=1.68 $X2=0
+ $Y2=0
cc_869 N_A_1526_315#_c_1275_n N_Q_c_1744_n 0.00241802f $X=9.635 $Y=1.16 $X2=0
+ $Y2=0
cc_870 N_A_1526_315#_c_1270_n N_Q_c_1742_n 0.00259707f $X=9.215 $Y=0.995 $X2=0
+ $Y2=0
cc_871 N_A_1526_315#_M1010_g N_Q_c_1742_n 0.00275407f $X=9.215 $Y=1.985 $X2=0
+ $Y2=0
cc_872 N_A_1526_315#_c_1271_n N_Q_c_1742_n 0.0047058f $X=9.635 $Y=0.995 $X2=0
+ $Y2=0
cc_873 N_A_1526_315#_M1033_g N_Q_c_1742_n 0.00569148f $X=9.635 $Y=1.985 $X2=0
+ $Y2=0
cc_874 N_A_1526_315#_c_1273_n N_Q_c_1742_n 0.0250466f $X=9.18 $Y=1.16 $X2=0
+ $Y2=0
cc_875 N_A_1526_315#_c_1275_n N_Q_c_1742_n 0.0236868f $X=9.635 $Y=1.16 $X2=0
+ $Y2=0
cc_876 N_A_1526_315#_M1010_g Q 0.00801319f $X=9.215 $Y=1.985 $X2=0 $Y2=0
cc_877 N_A_1526_315#_M1033_g Q 0.00911451f $X=9.635 $Y=1.985 $X2=0 $Y2=0
cc_878 N_A_1526_315#_c_1270_n N_Q_c_1757_n 0.00816502f $X=9.215 $Y=0.995 $X2=0
+ $Y2=0
cc_879 N_A_1526_315#_c_1271_n N_Q_c_1757_n 0.00665089f $X=9.635 $Y=0.995 $X2=0
+ $Y2=0
cc_880 N_A_1526_315#_c_1274_n N_Q_c_1757_n 0.00375716f $X=8.55 $Y=0.385 $X2=0
+ $Y2=0
cc_881 N_A_1526_315#_c_1275_n N_Q_c_1757_n 0.00233371f $X=9.635 $Y=1.16 $X2=0
+ $Y2=0
cc_882 N_A_1526_315#_M1027_g N_VGND_c_1778_n 0.0215676f $X=7.82 $Y=0.445 $X2=0
+ $Y2=0
cc_883 N_A_1526_315#_c_1274_n N_VGND_c_1778_n 0.0187345f $X=8.55 $Y=0.385 $X2=0
+ $Y2=0
cc_884 N_A_1526_315#_c_1274_n N_VGND_c_1779_n 0.0172098f $X=8.55 $Y=0.385 $X2=0
+ $Y2=0
cc_885 N_A_1526_315#_c_1270_n N_VGND_c_1780_n 0.00556109f $X=9.215 $Y=0.995
+ $X2=0 $Y2=0
cc_886 N_A_1526_315#_c_1273_n N_VGND_c_1780_n 0.00956157f $X=9.18 $Y=1.16 $X2=0
+ $Y2=0
cc_887 N_A_1526_315#_c_1274_n N_VGND_c_1780_n 0.0292994f $X=8.55 $Y=0.385 $X2=0
+ $Y2=0
cc_888 N_A_1526_315#_c_1275_n N_VGND_c_1780_n 6.26814e-19 $X=9.635 $Y=1.16 $X2=0
+ $Y2=0
cc_889 N_A_1526_315#_c_1271_n N_VGND_c_1782_n 0.0081377f $X=9.635 $Y=0.995 $X2=0
+ $Y2=0
cc_890 N_A_1526_315#_c_1270_n N_VGND_c_1787_n 0.00543342f $X=9.215 $Y=0.995
+ $X2=0 $Y2=0
cc_891 N_A_1526_315#_c_1271_n N_VGND_c_1787_n 0.00521596f $X=9.635 $Y=0.995
+ $X2=0 $Y2=0
cc_892 N_A_1526_315#_M1015_s N_VGND_c_1794_n 0.00212021f $X=8.425 $Y=0.235 $X2=0
+ $Y2=0
cc_893 N_A_1526_315#_M1027_g N_VGND_c_1794_n 9.61436e-19 $X=7.82 $Y=0.445 $X2=0
+ $Y2=0
cc_894 N_A_1526_315#_c_1270_n N_VGND_c_1794_n 0.00973405f $X=9.215 $Y=0.995
+ $X2=0 $Y2=0
cc_895 N_A_1526_315#_c_1271_n N_VGND_c_1794_n 0.00995869f $X=9.635 $Y=0.995
+ $X2=0 $Y2=0
cc_896 N_A_1526_315#_c_1274_n N_VGND_c_1794_n 0.0127495f $X=8.55 $Y=0.385 $X2=0
+ $Y2=0
cc_897 N_A_1355_413#_M1002_g N_VPWR_c_1461_n 0.0021703f $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_898 N_A_1355_413#_M1002_g N_VPWR_c_1462_n 0.00511679f $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_899 N_A_1355_413#_M1002_g N_VPWR_c_1463_n 0.0059044f $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_900 N_A_1355_413#_c_1380_n N_VPWR_c_1471_n 0.0273845f $X=7.46 $Y=2.25 $X2=0
+ $Y2=0
cc_901 N_A_1355_413#_M1009_d N_VPWR_c_1456_n 0.00219484f $X=6.775 $Y=2.065 $X2=0
+ $Y2=0
cc_902 N_A_1355_413#_M1002_g N_VPWR_c_1456_n 0.0103298f $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_903 N_A_1355_413#_c_1380_n N_VPWR_c_1456_n 0.0276628f $X=7.46 $Y=2.25 $X2=0
+ $Y2=0
cc_904 N_A_1355_413#_c_1380_n A_1439_413# 0.0105858f $X=7.46 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_905 N_A_1355_413#_c_1377_n A_1439_413# 0.00184879f $X=7.545 $Y=2.165
+ $X2=-0.19 $Y2=-0.24
cc_906 N_A_1355_413#_M1002_g N_Q_c_1744_n 5.08641e-19 $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_907 N_A_1355_413#_c_1368_n N_Q_c_1757_n 4.19418e-19 $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_908 N_A_1355_413#_c_1368_n N_VGND_c_1778_n 0.00268732f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_909 N_A_1355_413#_c_1383_n N_VGND_c_1778_n 0.0104892f $X=7.33 $Y=0.45 $X2=0
+ $Y2=0
cc_910 N_A_1355_413#_c_1371_n N_VGND_c_1778_n 0.0154767f $X=8.31 $Y=1.16 $X2=0
+ $Y2=0
cc_911 N_A_1355_413#_c_1373_n N_VGND_c_1778_n 0.00447237f $X=7.48 $Y=0.995 $X2=0
+ $Y2=0
cc_912 N_A_1355_413#_c_1368_n N_VGND_c_1779_n 0.00514019f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_913 N_A_1355_413#_c_1368_n N_VGND_c_1780_n 0.00534404f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_914 N_A_1355_413#_c_1383_n N_VGND_c_1786_n 0.0184388f $X=7.33 $Y=0.45 $X2=0
+ $Y2=0
cc_915 N_A_1355_413#_M1003_d N_VGND_c_1794_n 0.00333348f $X=6.905 $Y=0.235 $X2=0
+ $Y2=0
cc_916 N_A_1355_413#_c_1368_n N_VGND_c_1794_n 0.0103347f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_917 N_A_1355_413#_c_1383_n N_VGND_c_1794_n 0.0182474f $X=7.33 $Y=0.45 $X2=0
+ $Y2=0
cc_918 N_A_1355_413#_c_1383_n A_1484_47# 0.00201232f $X=7.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_919 N_A_1355_413#_c_1373_n A_1484_47# 0.00127737f $X=7.48 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_920 N_VPWR_c_1456_n A_467_369# 0.00274581f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_921 N_VPWR_c_1456_n N_A_559_369#_M1016_d 0.00179277f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1456_n N_A_559_369#_M1008_s 0.00269423f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1458_n N_A_559_369#_c_1632_n 0.00574724f $X=2.045 $Y=2.33 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1459_n N_A_559_369#_c_1632_n 0.0133617f $X=3.84 $Y=2.33 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1470_n N_A_559_369#_c_1632_n 0.0382337f $X=3.755 $Y=2.72 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1456_n N_A_559_369#_c_1632_n 0.0141871f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1459_n N_A_559_369#_c_1656_n 0.00558244f $X=3.84 $Y=2.33 $X2=0
+ $Y2=0
cc_928 N_VPWR_M1005_d N_A_559_369#_c_1628_n 0.00372198f $X=3.68 $Y=1.845 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1459_n N_A_559_369#_c_1628_n 0.0119067f $X=3.84 $Y=2.33 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1466_n N_A_559_369#_c_1628_n 0.00429797f $X=5.93 $Y=2.72 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1470_n N_A_559_369#_c_1628_n 0.00196122f $X=3.755 $Y=2.72 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1456_n N_A_559_369#_c_1628_n 0.00533045f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1459_n N_A_559_369#_c_1631_n 0.0144725f $X=3.84 $Y=2.33 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1466_n N_A_559_369#_c_1631_n 0.0140749f $X=5.93 $Y=2.72 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1456_n N_A_559_369#_c_1631_n 0.00421345f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_936 N_VPWR_c_1456_n A_643_369# 0.00210687f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_937 N_VPWR_c_1456_n A_1032_413# 0.00220641f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_938 N_VPWR_c_1456_n A_1439_413# 0.00377587f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_939 N_VPWR_c_1456_n N_Q_M1010_d 0.00220947f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_940 N_VPWR_c_1463_n N_Q_c_1744_n 0.0546648f $X=8.99 $Y=1.79 $X2=0 $Y2=0
cc_941 N_VPWR_c_1465_n N_Q_c_1742_n 0.0733896f $X=9.86 $Y=1.63 $X2=0 $Y2=0
cc_942 N_VPWR_c_1472_n Q 0.0137796f $X=9.775 $Y=2.72 $X2=0 $Y2=0
cc_943 N_VPWR_c_1456_n Q 0.0122496f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_944 N_VPWR_c_1465_n N_VGND_c_1782_n 0.00769463f $X=9.86 $Y=1.63 $X2=0 $Y2=0
cc_945 N_A_559_369#_c_1632_n A_643_369# 0.00382565f $X=3.415 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_946 N_A_559_369#_c_1656_n A_643_369# 0.00266005f $X=3.5 $Y=2.245 $X2=-0.19
+ $Y2=-0.24
cc_947 N_A_559_369#_c_1629_n A_643_369# 9.25434e-19 $X=3.585 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_948 N_A_559_369#_c_1644_n N_VGND_c_1774_n 0.00106538f $X=3.42 $Y=0.36 $X2=0
+ $Y2=0
cc_949 N_A_559_369#_c_1644_n N_VGND_c_1775_n 0.0135146f $X=3.42 $Y=0.36 $X2=0
+ $Y2=0
cc_950 N_A_559_369#_c_1621_n N_VGND_c_1775_n 0.00565411f $X=3.505 $Y=0.695 $X2=0
+ $Y2=0
cc_951 N_A_559_369#_c_1622_n N_VGND_c_1775_n 0.0142693f $X=4.21 $Y=0.78 $X2=0
+ $Y2=0
cc_952 N_A_559_369#_c_1626_n N_VGND_c_1775_n 0.00958978f $X=4.395 $Y=0.45 $X2=0
+ $Y2=0
cc_953 N_A_559_369#_c_1622_n N_VGND_c_1776_n 0.00402378f $X=4.21 $Y=0.78 $X2=0
+ $Y2=0
cc_954 N_A_559_369#_c_1626_n N_VGND_c_1776_n 0.012161f $X=4.395 $Y=0.45 $X2=0
+ $Y2=0
cc_955 N_A_559_369#_c_1644_n N_VGND_c_1785_n 0.0378786f $X=3.42 $Y=0.36 $X2=0
+ $Y2=0
cc_956 N_A_559_369#_c_1622_n N_VGND_c_1785_n 0.00256455f $X=4.21 $Y=0.78 $X2=0
+ $Y2=0
cc_957 N_A_559_369#_M1022_d N_VGND_c_1794_n 0.00217379f $X=2.82 $Y=0.235 $X2=0
+ $Y2=0
cc_958 N_A_559_369#_M1028_s N_VGND_c_1794_n 0.00195217f $X=4.27 $Y=0.235 $X2=0
+ $Y2=0
cc_959 N_A_559_369#_c_1644_n N_VGND_c_1794_n 0.0126583f $X=3.42 $Y=0.36 $X2=0
+ $Y2=0
cc_960 N_A_559_369#_c_1622_n N_VGND_c_1794_n 0.00517112f $X=4.21 $Y=0.78 $X2=0
+ $Y2=0
cc_961 N_A_559_369#_c_1626_n N_VGND_c_1794_n 0.00544577f $X=4.395 $Y=0.45 $X2=0
+ $Y2=0
cc_962 N_A_559_369#_c_1644_n A_660_47# 0.00210886f $X=3.42 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_963 N_A_559_369#_c_1621_n A_660_47# 0.00222412f $X=3.505 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_964 N_Q_c_1757_n N_VGND_c_1780_n 0.0270681f $X=9.425 $Y=0.395 $X2=0 $Y2=0
cc_965 N_Q_c_1757_n N_VGND_c_1782_n 0.0462989f $X=9.425 $Y=0.395 $X2=0 $Y2=0
cc_966 N_Q_c_1757_n N_VGND_c_1787_n 0.0149988f $X=9.425 $Y=0.395 $X2=0 $Y2=0
cc_967 N_Q_M1011_s N_VGND_c_1794_n 0.00218509f $X=9.29 $Y=0.235 $X2=0 $Y2=0
cc_968 N_Q_c_1757_n N_VGND_c_1794_n 0.0123405f $X=9.425 $Y=0.395 $X2=0 $Y2=0
cc_969 N_VGND_c_1794_n A_486_47# 0.00171756f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_970 N_VGND_c_1794_n A_660_47# 0.00152414f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_971 N_VGND_c_1794_n A_1036_47# 0.00272292f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24
cc_972 N_VGND_c_1794_n A_1484_47# 0.0111093f $X=9.89 $Y=0 $X2=-0.19 $Y2=-0.24

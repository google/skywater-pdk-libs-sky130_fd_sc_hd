* File: sky130_fd_sc_hd__clkdlybuf4s18_2.pex.spice
* Created: Tue Sep  1 19:00:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A 3 5 7 9 13
c30 5 0 2.2234e-19 $X=0.48 $Y=1.305
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.395
+ $Y=1.16 $X2=0.395 $Y2=1.16
r32 9 13 8.57632 $w=2.13e-07 $l=1.6e-07 $layer=LI1_cond $X=0.235 $Y=1.182
+ $X2=0.395 $Y2=1.182
r33 5 12 35.6637 $w=3.29e-07 $l=1.8262e-07 $layer=POLY_cond $X=0.48 $Y=1.305
+ $X2=0.395 $Y2=1.16
r34 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.48 $Y=1.305 $X2=0.48
+ $Y2=1.985
r35 1 12 35.6637 $w=3.29e-07 $l=1.8262e-07 $layer=POLY_cond $X=0.48 $Y=1.015
+ $X2=0.395 $Y2=1.16
r36 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.48 $Y=1.015 $X2=0.48
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_27_47# 1 2 9 13 17 21 23 24 25 26
+ 30 31
c62 30 0 1.74e-19 $X=0.97 $Y=1.16
c63 25 0 1.08211e-19 $X=0.73 $Y=1.545
c64 23 0 1.14128e-19 $X=0.73 $Y=0.82
r65 31 34 35.4445 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.97 $Y=1.16
+ $X2=0.97 $Y2=1.295
r66 31 33 35.4445 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.97 $Y=1.16
+ $X2=0.97 $Y2=1.025
r67 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.16 $X2=0.97 $Y2=1.16
r68 28 30 10.6379 $w=3.23e-07 $l=3e-07 $layer=LI1_cond $X=0.892 $Y=1.46
+ $X2=0.892 $Y2=1.16
r69 27 30 9.04224 $w=3.23e-07 $l=2.55e-07 $layer=LI1_cond $X=0.892 $Y=0.905
+ $X2=0.892 $Y2=1.16
r70 25 28 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=0.73 $Y=1.545
+ $X2=0.892 $Y2=1.46
r71 25 26 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.73 $Y=1.545 $X2=0.43
+ $Y2=1.545
r72 23 27 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=0.73 $Y=0.82
+ $X2=0.892 $Y2=0.905
r73 23 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.73 $Y=0.82
+ $X2=0.415 $Y2=0.82
r74 19 26 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.257 $Y=1.63
+ $X2=0.43 $Y2=1.545
r75 19 21 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=1.63
+ $X2=0.257 $Y2=1.965
r76 15 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.25 $Y=0.735
+ $X2=0.415 $Y2=0.82
r77 15 17 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.25 $Y=0.735 $X2=0.25
+ $Y2=0.435
r78 13 34 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=1.045 $Y=2.075
+ $X2=1.045 $Y2=1.295
r79 9 33 180.75 $w=1.8e-07 $l=4.65e-07 $layer=POLY_cond $X=1.045 $Y=0.56
+ $X2=1.045 $Y2=1.025
r80 2 21 300 $w=1.7e-07 $l=5.4111e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.265 $Y2=1.965
r81 1 17 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.265 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_227_47# 1 2 11 15 19 22 27 28 30
+ 32 35
c63 28 0 1.74e-19 $X=2.04 $Y=1.16
c64 27 0 1.8113e-19 $X=2.04 $Y=1.16
c65 15 0 1.14658e-19 $X=2.025 $Y=2.075
r66 32 34 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=0.435
+ $X2=1.3 $Y2=0.6
r67 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.04
+ $Y=1.16 $X2=2.04 $Y2=1.16
r68 25 35 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=1.165
+ $X2=1.355 $Y2=1.165
r69 25 27 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=1.44 $Y=1.165 $X2=2.04
+ $Y2=1.165
r70 23 35 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.355 $Y=1.255
+ $X2=1.355 $Y2=1.165
r71 23 30 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.355 $Y=1.255
+ $X2=1.355 $Y2=1.8
r72 22 35 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.355 $Y=1.075
+ $X2=1.355 $Y2=1.165
r73 22 34 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.355 $Y=1.075
+ $X2=1.355 $Y2=0.6
r74 19 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=1.965
+ $X2=1.275 $Y2=1.8
r75 13 28 28.1878 $w=1.8e-07 $l=1.55885e-07 $layer=POLY_cond $X=2.025 $Y=1.295
+ $X2=2.07 $Y2=1.16
r76 13 15 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=2.025 $Y=1.295
+ $X2=2.025 $Y2=2.075
r77 9 28 28.1878 $w=1.8e-07 $l=1.55885e-07 $layer=POLY_cond $X=2.025 $Y=1.025
+ $X2=2.07 $Y2=1.16
r78 9 11 180.75 $w=1.8e-07 $l=4.65e-07 $layer=POLY_cond $X=2.025 $Y=1.025
+ $X2=2.025 $Y2=0.56
r79 2 19 300 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.665 $X2=1.275 $Y2=1.965
r80 1 32 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.135
+ $Y=0.235 $X2=1.275 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_334_47# 1 2 9 13 15 19 23 25 28 32
+ 34 35 36 37 39 41 44 45 47
c97 45 0 3.94822e-19 $X=2.675 $Y=1.16
c98 34 0 1.59543e-19 $X=2.375 $Y=0.82
r99 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.16 $X2=2.675 $Y2=1.16
r100 42 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=1.16
+ $X2=2.46 $Y2=1.16
r101 42 44 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.545 $Y=1.16
+ $X2=2.675 $Y2=1.16
r102 40 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.245
+ $X2=2.46 $Y2=1.16
r103 40 41 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.46 $Y=1.245
+ $X2=2.46 $Y2=1.46
r104 39 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.075
+ $X2=2.46 $Y2=1.16
r105 38 39 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.46 $Y=0.905
+ $X2=2.46 $Y2=1.075
r106 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=1.545
+ $X2=2.46 $Y2=1.46
r107 36 37 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.375 $Y=1.545
+ $X2=1.96 $Y2=1.545
r108 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=0.82
+ $X2=2.46 $Y2=0.905
r109 34 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.375 $Y=0.82
+ $X2=1.96 $Y2=0.82
r110 30 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.795 $Y=1.63
+ $X2=1.96 $Y2=1.545
r111 30 32 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.795 $Y=1.63
+ $X2=1.795 $Y2=1.965
r112 26 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.795 $Y=0.735
+ $X2=1.96 $Y2=0.82
r113 26 28 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.795 $Y=0.735
+ $X2=1.795 $Y2=0.435
r114 21 25 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.095 $Y=1.295
+ $X2=3.095 $Y2=1.16
r115 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.095 $Y=1.295
+ $X2=3.095 $Y2=1.985
r116 17 25 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.095 $Y=1.025
+ $X2=3.095 $Y2=1.16
r117 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.095 $Y=1.025
+ $X2=3.095 $Y2=0.445
r118 16 45 2.60871 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=2.74 $Y=1.16
+ $X2=2.625 $Y2=1.16
r119 15 25 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.02 $Y=1.16
+ $X2=3.095 $Y2=1.16
r120 15 16 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=3.02 $Y=1.16
+ $X2=2.74 $Y2=1.16
r121 11 45 32.2453 $w=1.5e-07 $l=1.53704e-07 $layer=POLY_cond $X=2.665 $Y=1.295
+ $X2=2.625 $Y2=1.16
r122 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.665 $Y=1.295
+ $X2=2.665 $Y2=1.985
r123 7 45 32.2453 $w=1.5e-07 $l=1.53704e-07 $layer=POLY_cond $X=2.665 $Y=1.025
+ $X2=2.625 $Y2=1.16
r124 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.665 $Y=1.025
+ $X2=2.665 $Y2=0.445
r125 2 32 300 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_PDIFF $count=2 $X=1.67
+ $Y=1.665 $X2=1.795 $Y2=1.965
r126 1 28 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.235 $X2=1.795 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%VPWR 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
c44 16 0 1.14886e-19 $X=2.35 $Y=1.965
r45 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r48 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r49 39 47 4.27912 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.32 $Y=2.72 $X2=3.5
+ $Y2=2.72
r50 39 41 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.32 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.765 $Y2=2.72
r58 32 34 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.765 $Y2=2.72
r60 27 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r61 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 23 37 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.13 $Y=2.72 $X2=2.07
+ $Y2=2.72
r64 23 24 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=2.13 $Y=2.72
+ $X2=2.337 $Y2=2.72
r65 22 41 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.99 $Y2=2.72
r66 22 24 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.337 $Y2=2.72
r67 18 47 3.04293 $w=2.75e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.457 $Y=2.635
+ $X2=3.5 $Y2=2.72
r68 18 20 28.0777 $w=2.73e-07 $l=6.7e-07 $layer=LI1_cond $X=3.457 $Y=2.635
+ $X2=3.457 $Y2=1.965
r69 14 24 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.337 $Y=2.635
+ $X2=2.337 $Y2=2.72
r70 14 16 18.6057 $w=4.13e-07 $l=6.7e-07 $layer=LI1_cond $X=2.337 $Y=2.635
+ $X2=2.337 $Y2=1.965
r71 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2.72
r72 10 12 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=1.965
r73 3 20 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=3.17
+ $Y=1.485 $X2=3.405 $Y2=1.965
r74 2 16 300 $w=1.7e-07 $l=4.00625e-07 $layer=licon1_PDIFF $count=2 $X=2.115
+ $Y=1.665 $X2=2.35 $Y2=1.965
r75 1 12 300 $w=1.7e-07 $l=5.755e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.765 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%X 1 2 12 13 14 15 16 17 18 30
c42 13 0 1.14658e-19 $X=2.947 $Y=1.525
r43 18 25 6.49077 $w=4.33e-07 $l=2.45e-07 $layer=LI1_cond $X=2.932 $Y=2.21
+ $X2=2.932 $Y2=1.965
r44 17 25 2.51683 $w=4.33e-07 $l=9.5e-08 $layer=LI1_cond $X=2.932 $Y=1.87
+ $X2=2.932 $Y2=1.965
r45 16 34 7.40247 $w=4.43e-07 $l=1.3e-07 $layer=LI1_cond $X=2.927 $Y=0.51
+ $X2=2.927 $Y2=0.64
r46 16 30 1.94232 $w=4.43e-07 $l=7.5e-08 $layer=LI1_cond $X=2.927 $Y=0.51
+ $X2=2.927 $Y2=0.435
r47 14 15 9.98442 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.072 $Y=0.78
+ $X2=3.072 $Y2=0.945
r48 14 34 8.39312 $w=1.83e-07 $l=1.4e-07 $layer=LI1_cond $X=3.057 $Y=0.78
+ $X2=3.057 $Y2=0.64
r49 13 17 9.14007 $w=4.33e-07 $l=3.45e-07 $layer=LI1_cond $X=2.932 $Y=1.525
+ $X2=2.932 $Y2=1.87
r50 12 13 7.22028 $w=4.33e-07 $l=1.05e-07 $layer=LI1_cond $X=2.947 $Y=1.42
+ $X2=2.947 $Y2=1.525
r51 12 15 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.095 $Y=1.42
+ $X2=3.095 $Y2=0.945
r52 2 25 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=2.74
+ $Y=1.485 $X2=2.88 $Y2=1.965
r53 1 30 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=2.74
+ $Y=0.235 $X2=2.88 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%VGND 1 2 3 12 16 18 20 23 24 25 27
+ 39 44 48
c49 39 0 1.59543e-19 $X=3.32 $Y=0
c50 16 0 9.88072e-20 $X=2.34 $Y=0.4
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r54 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 39 47 4.27912 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=3.5
+ $Y2=0
r56 39 41 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=2.99
+ $Y2=0
r57 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r58 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r59 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r60 35 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r61 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r62 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r63 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r64 32 34 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.15
+ $Y2=0
r65 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r66 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.23
+ $Y2=0
r67 25 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r68 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 23 37 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.07
+ $Y2=0
r70 23 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.35
+ $Y2=0
r71 22 41 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.99
+ $Y2=0
r72 22 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.35
+ $Y2=0
r73 18 47 3.04293 $w=2.75e-07 $l=1.04307e-07 $layer=LI1_cond $X=3.457 $Y=0.085
+ $X2=3.5 $Y2=0
r74 18 20 14.6675 $w=2.73e-07 $l=3.5e-07 $layer=LI1_cond $X=3.457 $Y=0.085
+ $X2=3.457 $Y2=0.435
r75 14 24 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0
r76 14 16 9.81134 $w=3.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0.4
r77 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r78 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.4
r79 3 20 182 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.405 $Y2=0.435
r80 2 16 182 $w=1.7e-07 $l=2.96226e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.34 $Y2=0.4
r81 1 12 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.75 $Y2=0.4
.ends


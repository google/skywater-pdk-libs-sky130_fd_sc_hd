* File: sky130_fd_sc_hd__and4bb_1.pex.spice
* Created: Tue Sep  1 18:58:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4BB_1%A_N 3 7 9 12 13
c35 12 0 2.18412e-20 $X=0.59 $Y=1.74
c36 3 0 1.57088e-19 $X=0.61 $Y=0.445
r37 12 15 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.59 $Y=1.74
+ $X2=0.59 $Y2=1.875
r38 12 14 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.59 $Y=1.74
+ $X2=0.59 $Y2=1.605
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.74 $X2=0.59 $Y2=1.74
r40 9 13 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=0.6 $Y=1.87 $X2=0.6
+ $Y2=1.74
r41 7 15 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.61 $Y=2.275 $X2=0.61
+ $Y2=1.875
r42 3 14 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=0.61 $Y=0.445
+ $X2=0.61 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%B_N 3 7 11 12 14
c48 12 0 1.84198e-19 $X=1.06 $Y=1.03
c49 11 0 1.57088e-19 $X=1.06 $Y=1.03
c50 7 0 1.85684e-19 $X=1.04 $Y=2.275
r51 14 22 9.50649 $w=2.08e-07 $l=1.8e-07 $layer=LI1_cond $X=0.71 $Y=0.85
+ $X2=0.71 $Y2=1.03
r52 12 18 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.06 $Y=1.03
+ $X2=1.06 $Y2=1.165
r53 12 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.06 $Y=1.03
+ $X2=1.06 $Y2=0.895
r54 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.03 $X2=1.06 $Y2=1.03
r55 9 22 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.815 $Y=1.03 $X2=0.71
+ $Y2=1.03
r56 9 11 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.815 $Y=1.03
+ $X2=1.06 $Y2=1.03
r57 7 18 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.04 $Y=2.275
+ $X2=1.04 $Y2=1.165
r58 3 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.04 $Y=0.445
+ $X2=1.04 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%A_27_47# 1 2 7 8 11 14 16 17 18 20 22 23 27
+ 33 35 39 41
c92 27 0 3.69882e-19 $X=1.46 $Y=1.66
r93 41 43 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.13 $Y=1.37
+ $X2=1.13 $Y2=1.66
r94 36 39 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=2.3 $X2=0.26
+ $Y2=2.3
r95 30 33 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.46
+ $Y=1.66 $X2=1.46 $Y2=1.66
r97 25 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=1.66
+ $X2=1.13 $Y2=1.66
r98 25 27 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.215 $Y=1.66
+ $X2=1.46 $Y2=1.66
r99 24 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=1.37
+ $X2=0.17 $Y2=1.37
r100 23 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=1.37
+ $X2=1.13 $Y2=1.37
r101 23 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.045 $Y=1.37
+ $X2=0.255 $Y2=1.37
r102 22 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=2.135
+ $X2=0.17 $Y2=2.3
r103 21 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=1.37
r104 21 22 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.17 $Y2=2.135
r105 20 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=1.285
+ $X2=0.17 $Y2=1.37
r106 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r107 19 20 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.285
r108 17 28 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=1.785 $Y=1.66
+ $X2=1.46 $Y2=1.66
r109 17 18 1.70994 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.785 $Y=1.66
+ $X2=1.965 $Y2=1.66
r110 12 18 25.1511 $w=2.55e-07 $l=2.11069e-07 $layer=POLY_cond $X=2.07 $Y=1.825
+ $X2=1.965 $Y2=1.66
r111 12 14 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.07 $Y=1.825
+ $X2=2.07 $Y2=2.275
r112 11 16 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.07 $Y=0.675 $X2=2.07
+ $Y2=0.975
r113 8 18 25.1511 $w=2.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.495
+ $X2=1.965 $Y2=1.66
r114 7 16 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.965 $Y=1.155
+ $X2=1.965 $Y2=0.975
r115 7 8 54.4984 $w=3.6e-07 $l=3.4e-07 $layer=POLY_cond $X=1.965 $Y=1.155
+ $X2=1.965 $Y2=1.495
r116 2 39 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r117 1 33 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%A_223_47# 1 2 9 12 16 19 20 21 22 24 25 27
+ 30 31 33 39
r99 36 37 13.5455 $w=3.98e-07 $l=3.35e-07 $layer=LI1_cond $X=1.365 $Y=0.42
+ $X2=1.365 $Y2=0.755
r100 33 36 2.30489 $w=3.98e-07 $l=8e-08 $layer=LI1_cond $X=1.365 $Y=0.34
+ $X2=1.365 $Y2=0.42
r101 31 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.56 $Y=1.16
+ $X2=2.56 $Y2=1.325
r102 31 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.56 $Y=1.16
+ $X2=2.56 $Y2=0.995
r103 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.16 $X2=2.56 $Y2=1.16
r104 28 30 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=1.16
r105 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.88 $Y=1.405
+ $X2=1.88 $Y2=1.915
r106 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=1.32
+ $X2=1.88 $Y2=1.405
r107 24 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.795 $Y=1.32
+ $X2=1.565 $Y2=1.32
r108 23 33 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.565 $Y=0.34
+ $X2=1.365 $Y2=0.34
r109 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=2.56 $Y2=0.425
r110 22 23 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=1.565 $Y2=0.34
r111 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=2
+ $X2=1.88 $Y2=1.915
r112 20 21 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.795 $Y=2
+ $X2=1.415 $Y2=2
r113 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.48 $Y=1.235
+ $X2=1.565 $Y2=1.32
r114 19 37 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.48 $Y=1.235
+ $X2=1.48 $Y2=0.755
r115 14 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.32 $Y=2.085
+ $X2=1.415 $Y2=2
r116 14 16 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.32 $Y=2.085
+ $X2=1.32 $Y2=2.3
r117 12 40 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.5 $Y=2.275
+ $X2=2.5 $Y2=1.325
r118 9 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.5 $Y=0.675 $X2=2.5
+ $Y2=0.995
r119 2 16 600 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=2.065 $X2=1.31 $Y2=2.3
r120 1 36 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.235 $X2=1.32 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%C 3 6 8 9 10 11 17 19
c45 8 0 1.50285e-19 $X=2.985 $Y=0.51
r46 17 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.16
+ $X2=3.04 $Y2=1.325
r47 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.16
+ $X2=3.04 $Y2=0.995
r48 11 34 12.2899 $w=1.83e-07 $l=2.05e-07 $layer=LI1_cond $X=2.987 $Y=1.53
+ $X2=2.987 $Y2=1.325
r49 10 34 8.74215 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.16
+ $X2=3.01 $Y2=1.325
r50 10 32 8.74215 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.16
+ $X2=3.01 $Y2=0.995
r51 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.16 $X2=3.04 $Y2=1.16
r52 9 32 8.69287 $w=1.83e-07 $l=1.45e-07 $layer=LI1_cond $X=2.987 $Y=0.85
+ $X2=2.987 $Y2=0.995
r53 8 9 20.3833 $w=1.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.987 $Y=0.51
+ $X2=2.987 $Y2=0.85
r54 6 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3 $Y=2.275 $X2=3
+ $Y2=1.325
r55 3 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3 $Y=0.675 $X2=3
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%D 1 3 6 8 9 10 11 17
r45 11 32 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.447 $Y=1.53
+ $X2=3.447 $Y2=1.325
r46 10 32 8.12371 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.477 $Y=1.16
+ $X2=3.477 $Y2=1.325
r47 10 30 8.12371 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.477 $Y=1.16
+ $X2=3.477 $Y2=0.995
r48 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.52
+ $Y=1.16 $X2=3.52 $Y2=1.16
r49 9 30 8.24709 $w=1.93e-07 $l=1.45e-07 $layer=LI1_cond $X=3.447 $Y=0.85
+ $X2=3.447 $Y2=0.995
r50 8 9 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=3.447 $Y=0.51 $X2=3.447
+ $Y2=0.85
r51 4 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.16
r52 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.52 $Y=1.325 $X2=3.52
+ $Y2=2.275
r53 1 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=0.995
+ $X2=3.52 $Y2=1.16
r54 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.52 $Y=0.995 $X2=3.52
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%A_343_93# 1 2 3 12 15 17 22 25 27 31 33 37
+ 38 40 41 43
r91 38 44 50.2341 $w=6.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.177 $Y=1.16
+ $X2=4.177 $Y2=1.325
r92 38 43 50.2341 $w=6.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.177 $Y=1.16
+ $X2=4.177 $Y2=0.995
r93 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4 $Y=1.16
+ $X2=4 $Y2=1.16
r94 35 37 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4 $Y=1.915 $X2=4
+ $Y2=1.16
r95 34 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=2 $X2=3.245
+ $Y2=2
r96 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.915 $Y=2 $X2=4
+ $Y2=1.915
r97 33 34 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.915 $Y=2 $X2=3.33
+ $Y2=2
r98 29 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=2.085
+ $X2=3.245 $Y2=2
r99 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.245 $Y=2.085
+ $X2=3.245 $Y2=2.3
r100 28 40 1.34256 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.375 $Y=2 $X2=2.255
+ $Y2=2
r101 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=2 $X2=3.245
+ $Y2=2
r102 27 28 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.16 $Y=2
+ $X2=2.375 $Y2=2
r103 23 40 5.16603 $w=1.7e-07 $l=1.00995e-07 $layer=LI1_cond $X=2.29 $Y=2.085
+ $X2=2.255 $Y2=2
r104 23 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.29 $Y=2.085
+ $X2=2.29 $Y2=2.3
r105 22 40 5.16603 $w=1.7e-07 $l=1.00995e-07 $layer=LI1_cond $X=2.22 $Y=1.915
+ $X2=2.255 $Y2=2
r106 21 22 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.22 $Y=0.925
+ $X2=2.22 $Y2=1.915
r107 17 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.135 $Y=0.76
+ $X2=2.22 $Y2=0.925
r108 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.135 $Y=0.76
+ $X2=1.86 $Y2=0.76
r109 15 44 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.13 $Y=1.985
+ $X2=4.13 $Y2=1.325
r110 12 43 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.56
+ $X2=4.13 $Y2=0.995
r111 3 31 600 $w=1.7e-07 $l=3.08504e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=2.065 $X2=3.245 $Y2=2.3
r112 2 25 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=2.145
+ $Y=2.065 $X2=2.29 $Y2=2.3
r113 1 19 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.465 $X2=1.86 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%VPWR 1 2 3 4 17 21 25 29 32 33 35 36 37 46
+ 52 53 56 59
c77 53 0 2.18412e-20 $X=4.37 $Y=2.72
r78 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 53 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r81 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r82 50 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=3.92 $Y2=2.72
r83 50 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=4.37 $Y2=2.72
r84 49 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r85 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r86 46 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.92 $Y2=2.72
r87 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.45 $Y2=2.72
r88 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r90 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r91 42 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r92 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=0.82 $Y2=2.72
r94 39 41 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=1.61 $Y2=2.72
r95 37 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 35 44 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.57 $Y=2.72 $X2=2.53
+ $Y2=2.72
r97 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=2.72
+ $X2=2.735 $Y2=2.72
r98 34 48 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.9 $Y=2.72 $X2=3.45
+ $Y2=2.72
r99 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=2.72
+ $X2=2.735 $Y2=2.72
r100 32 41 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.61 $Y2=2.72
r101 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.83 $Y2=2.72
r102 31 44 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.995 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=2.72
+ $X2=1.83 $Y2=2.72
r104 27 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.92 $Y2=2.72
r105 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.92 $Y=2.635
+ $X2=3.92 $Y2=2.34
r106 23 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.635
+ $X2=2.735 $Y2=2.72
r107 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.735 $Y=2.635
+ $X2=2.735 $Y2=2.34
r108 19 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.72
r109 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.83 $Y=2.635
+ $X2=1.83 $Y2=2.34
r110 15 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=2.635
+ $X2=0.82 $Y2=2.72
r111 15 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.82 $Y=2.635
+ $X2=0.82 $Y2=2.34
r112 4 29 600 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_PDIFF $count=1 $X=3.595
+ $Y=2.065 $X2=3.92 $Y2=2.34
r113 3 25 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.065 $X2=2.735 $Y2=2.34
r114 2 21 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=2.065 $X2=1.83 $Y2=2.34
r115 1 17 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.065 $X2=0.82 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%X 1 2 7 8 9 10 11 18
r12 11 29 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=4.385 $Y=2.21
+ $X2=4.385 $Y2=1.96
r13 10 29 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=4.385 $Y=1.87
+ $X2=4.385 $Y2=1.96
r14 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=4.385 $Y=1.53
+ $X2=4.385 $Y2=1.87
r15 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=4.385 $Y=1.19
+ $X2=4.385 $Y2=1.53
r16 7 8 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=4.385 $Y=0.85
+ $X2=4.385 $Y2=1.19
r17 7 18 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=4.385 $Y=0.85
+ $X2=4.385 $Y2=0.42
r18 2 29 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.205
+ $Y=1.485 $X2=4.34 $Y2=1.96
r19 1 18 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.235 $X2=4.34 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_1%VGND 1 2 11 15 17 19 29 30 33 36
c48 15 0 1.50285e-19 $X=3.92 $Y=0.38
r49 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r50 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r52 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r53 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=3.92
+ $Y2=0
r54 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.37
+ $Y2=0
r55 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r56 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r57 23 26 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r58 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r59 22 25 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r60 22 23 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.82
+ $Y2=0
r62 20 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.15
+ $Y2=0
r63 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.92
+ $Y2=0
r64 19 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.45
+ $Y2=0
r65 17 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r66 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=0.085
+ $X2=3.92 $Y2=0
r67 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.92 $Y=0.085
+ $X2=3.92 $Y2=0.38
r68 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=0.085 $X2=0.82
+ $Y2=0
r69 9 11 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0.38
r70 2 15 182 $w=1.7e-07 $l=3.65034e-07 $layer=licon1_NDIFF $count=1 $X=3.595
+ $Y=0.465 $X2=3.92 $Y2=0.38
r71 1 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.685
+ $Y=0.235 $X2=0.82 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__clkinv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=5.45e+11p pd=5.09e+06u as=5.45e+11p ps=5.09e+06u
M1001 VPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.205e+11p ps=2.73e+06u
M1003 Y A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__ha_4.spice
* Created: Thu Aug 27 14:22:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__ha_4.spice.pex"
.subckt sky130_fd_sc_hd__ha_4  VNB VPB A B VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_A_79_21#_M1014_g N_SUM_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A_79_21#_M1020_g N_SUM_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1020_d N_A_79_21#_M1021_g N_SUM_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1031 N_VGND_M1031_d N_A_79_21#_M1031_g N_SUM_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1015 N_A_467_47#_M1015_d N_A_514_199#_M1015_g N_A_79_21#_M1015_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1017 N_A_467_47#_M1017_d N_A_514_199#_M1017_g N_A_79_21#_M1015_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_A_467_47#_M1017_d VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.08775 PD=0.945 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1013_d N_B_M1023_g N_A_467_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.08775 PD=0.945 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1025_d N_B_M1025_g N_A_467_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_A_M1024_g N_A_467_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.18525 PD=0.92 PS=1.87 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75000.2
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1009 A_1325_47# N_A_M1009_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.65 AD=0.0715
+ AS=0.08775 PD=0.87 PS=0.92 NRD=10.152 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_514_199#_M1000_d N_B_M1000_g A_1325_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.0715 PD=0.92 PS=0.87 NRD=0 NRS=10.152 M=1 R=4.33333 SA=75001
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1006 N_A_514_199#_M1000_d N_B_M1006_g A_1167_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75001.4
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1033 A_1167_47# N_A_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.11375 PD=0.92 PS=1 NRD=14.76 NRS=6.456 M=1 R=4.33333 SA=75001.8
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1033_s N_A_514_199#_M1001_g N_COUT_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.11375 AS=0.08775 PD=1 PS=0.92 NRD=6.456 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_514_199#_M1004_g N_COUT_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.8 SB=75001 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1004_d N_A_514_199#_M1010_g N_COUT_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_514_199#_M1012_g N_COUT_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_SUM_M1005_d N_A_79_21#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75008.4 A=0.15 P=2.3 MULT=1
MM1011 N_SUM_M1005_d N_A_79_21#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75008 A=0.15 P=2.3 MULT=1
MM1022 N_SUM_M1022_d N_A_79_21#_M1022_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75007.6 A=0.15 P=2.3 MULT=1
MM1030 N_SUM_M1022_d N_A_79_21#_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.3825 PD=1.27 PS=1.765 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75007.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_79_21#_M1002_d N_A_514_199#_M1002_g N_VPWR_M1030_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.3825 PD=1.27 PS=1.765 NRD=0 NRS=29.5303 M=1 R=6.66667
+ SA=75002.4 SB=75006.3 A=0.15 P=2.3 MULT=1
MM1016 N_A_79_21#_M1002_d N_A_514_199#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.1475 PD=1.27 PS=1.295 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75005.8 A=0.15 P=2.3 MULT=1
MM1026 N_VPWR_M1016_s N_A_M1026_g A_717_297# VPB PHIGHVT L=0.15 W=1 AD=0.1475
+ AS=0.1475 PD=1.295 PS=1.295 NRD=3.9203 NRS=18.2028 M=1 R=6.66667 SA=75003.2
+ SB=75005.4 A=0.15 P=2.3 MULT=1
MM1007 A_717_297# N_B_M1007_g N_A_79_21#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1475 AS=0.135 PD=1.295 PS=1.27 NRD=18.2028 NRS=0 M=1 R=6.66667 SA=75003.7
+ SB=75005 A=0.15 P=2.3 MULT=1
MM1032 A_890_297# N_B_M1032_g N_A_79_21#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2875 AS=0.135 PD=1.575 PS=1.27 NRD=45.7828 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1028 N_VPWR_M1028_d N_A_M1028_g A_890_297# VPB PHIGHVT L=0.15 W=1 AD=0.23
+ AS=0.2875 PD=1.46 PS=1.575 NRD=17.73 NRS=45.7828 M=1 R=6.66667 SA=75004.8
+ SB=75003.8 A=0.15 P=2.3 MULT=1
MM1029 N_A_514_199#_M1029_d N_A_M1029_g N_VPWR_M1028_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.23 PD=1.27 PS=1.46 NRD=0 NRS=17.73 M=1 R=6.66667 SA=75005.4
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_514_199#_M1029_d N_B_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.8
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1018 N_A_514_199#_M1018_d N_B_M1018_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.3
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1034 N_A_514_199#_M1018_d N_A_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.175 PD=1.27 PS=1.35 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75006.7
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1008 N_COUT_M1008_d N_A_514_199#_M1008_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.175 PD=1.27 PS=1.35 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75007.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1019 N_COUT_M1008_d N_A_514_199#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1027 N_COUT_M1027_d N_A_514_199#_M1027_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1035 N_COUT_M1027_d N_A_514_199#_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX36_noxref VNB VPB NWDIODE A=15.3759 P=22.37
c_145 VPB 0 2.91462e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__ha_4.spice.SKY130_FD_SC_HD__HA_4.pxi"
*
.ends
*
*

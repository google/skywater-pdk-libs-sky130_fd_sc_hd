* File: sky130_fd_sc_hd__dfxtp_1.pex.spice
* Created: Tue Sep  1 19:04:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFXTP_1%CLK 1 2 3 5 6 8 11 13
c40 1 0 2.71124e-20 $X=0.305 $Y=1.325
r41 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r42 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r43 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r44 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r45 3 16 88.7086 $w=2.58e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r46 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r47 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r48 1 16 39.2009 $w=2.58e-07 $l=1.75656e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.327 $Y2=1.16
r49 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%A_27_47# 1 2 9 13 17 21 25 27 31 35 39 40 41
+ 44 46 48 51 54 56 57 58 59 60 67 69 74 82 85 89
c239 89 0 1.92554e-19 $X=4.375 $Y=1.41
c240 60 0 3.69553e-20 $X=2.96 $Y=1.87
c241 59 0 8.81722e-20 $X=4.24 $Y=1.87
c242 51 0 1.91737e-19 $X=2.38 $Y=0.87
c243 44 0 1.81794e-19 $X=0.725 $Y=1.795
c244 41 0 3.29888e-20 $X=0.61 $Y=1.88
r245 88 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.41
+ $X2=4.375 $Y2=1.575
r246 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.375
+ $Y=1.41 $X2=4.375 $Y2=1.41
r247 85 88 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=4.375 $Y=1.32
+ $X2=4.375 $Y2=1.41
r248 79 82 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.73 $Y=1.74
+ $X2=2.825 $Y2=1.74
r249 70 89 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=4.385 $Y=1.87
+ $X2=4.385 $Y2=1.41
r250 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.385 $Y=1.87
+ $X2=4.385 $Y2=1.87
r251 67 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.74 $X2=2.825 $Y2=1.74
r252 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.815 $Y=1.87
+ $X2=2.815 $Y2=1.87
r253 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.715 $Y=1.87
+ $X2=0.715 $Y2=1.87
r254 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.96 $Y=1.87
+ $X2=2.815 $Y2=1.87
r255 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.24 $Y=1.87
+ $X2=4.385 $Y2=1.87
r256 59 60 1.58416 $w=1.4e-07 $l=1.28e-06 $layer=MET1_cond $X=4.24 $Y=1.87
+ $X2=2.96 $Y2=1.87
r257 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.86 $Y=1.87
+ $X2=0.715 $Y2=1.87
r258 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.67 $Y=1.87
+ $X2=2.815 $Y2=1.87
r259 57 58 2.24009 $w=1.4e-07 $l=1.81e-06 $layer=MET1_cond $X=2.67 $Y=1.87
+ $X2=0.86 $Y2=1.87
r260 54 67 5.05181 $w=3.63e-07 $l=1.6e-07 $layer=LI1_cond $X=2.655 $Y=1.837
+ $X2=2.815 $Y2=1.837
r261 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.655 $Y=0.955
+ $X2=2.655 $Y2=1.655
r262 51 77 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.38 $Y=0.87
+ $X2=2.38 $Y2=0.735
r263 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=0.87 $X2=2.38 $Y2=0.87
r264 48 53 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.57 $Y=0.845
+ $X2=2.655 $Y2=0.955
r265 48 50 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=2.57 $Y=0.845
+ $X2=2.38 $Y2=0.845
r266 47 74 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r267 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r268 44 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r269 44 46 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r270 43 46 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r271 42 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r272 41 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r273 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r274 39 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r275 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r276 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r277 33 35 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r278 29 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=5.01 $Y=1.245
+ $X2=5.01 $Y2=0.415
r279 28 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.51 $Y=1.32
+ $X2=4.375 $Y2=1.32
r280 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.935 $Y=1.32
+ $X2=5.01 $Y2=1.245
r281 27 28 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.935 $Y=1.32
+ $X2=4.51 $Y2=1.32
r282 25 90 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.38 $Y=2.275
+ $X2=4.38 $Y2=1.575
r283 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.905
+ $X2=2.73 $Y2=1.74
r284 19 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.73 $Y=1.905
+ $X2=2.73 $Y2=2.275
r285 17 77 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.39 $Y=0.415
+ $X2=2.39 $Y2=0.735
r286 11 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r287 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r288 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r289 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r290 2 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r291 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%D 3 7 9 15
r45 12 15 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.565 $Y=1.5
+ $X2=1.83 $Y2=1.5
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.5 $X2=1.565 $Y2=1.5
r47 9 13 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.51 $Y=1.19 $X2=1.51
+ $Y2=1.5
r48 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.665
+ $X2=1.83 $Y2=1.5
r49 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.83 $Y=1.665 $X2=1.83
+ $Y2=2.275
r50 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.335
+ $X2=1.83 $Y2=1.5
r51 1 3 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.83 $Y=1.335 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%A_193_47# 1 2 9 11 15 17 19 22 26 27 30 31
+ 32 33 42 43 45 49 58 62
c179 45 0 1.74123e-19 $X=2.28 $Y=1.29
c180 43 0 2.06462e-20 $X=4.82 $Y=1.53
c181 22 0 1.92554e-19 $X=4.8 $Y=2.275
r182 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.74 $X2=4.885 $Y2=1.74
r183 55 58 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=4.8 $Y=1.74
+ $X2=4.885 $Y2=1.74
r184 48 50 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.28 $Y=1.35
+ $X2=2.28 $Y2=1.485
r185 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.35 $X2=2.28 $Y2=1.35
r186 45 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.28 $Y=1.29 $X2=2.28
+ $Y2=1.35
r187 43 59 7.56291 $w=3.18e-07 $l=2.1e-07 $layer=LI1_cond $X=4.81 $Y=1.53
+ $X2=4.81 $Y2=1.74
r188 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.82 $Y=1.53
+ $X2=4.82 $Y2=1.53
r189 40 49 8.64332 $w=2.38e-07 $l=1.8e-07 $layer=LI1_cond $X=2.28 $Y=1.53
+ $X2=2.28 $Y2=1.35
r190 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.3 $Y=1.53 $X2=2.3
+ $Y2=1.53
r191 36 66 25.7789 $w=1.83e-07 $l=4.3e-07 $layer=LI1_cond $X=1.107 $Y=1.53
+ $X2=1.107 $Y2=1.96
r192 36 62 61.1499 $w=1.83e-07 $l=1.02e-06 $layer=LI1_cond $X=1.107 $Y=1.53
+ $X2=1.107 $Y2=0.51
r193 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.11 $Y=1.53
+ $X2=1.11 $Y2=1.53
r194 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.445 $Y=1.53
+ $X2=2.3 $Y2=1.53
r195 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.675 $Y=1.53
+ $X2=4.82 $Y2=1.53
r196 32 33 2.7599 $w=1.4e-07 $l=2.23e-06 $layer=MET1_cond $X=4.675 $Y=1.53
+ $X2=2.445 $Y2=1.53
r197 31 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.255 $Y=1.53
+ $X2=1.11 $Y2=1.53
r198 30 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.155 $Y=1.53
+ $X2=2.3 $Y2=1.53
r199 30 31 1.11386 $w=1.4e-07 $l=9e-07 $layer=MET1_cond $X=2.155 $Y=1.53
+ $X2=1.255 $Y2=1.53
r200 29 43 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=4.81 $Y=1.035
+ $X2=4.81 $Y2=1.53
r201 27 51 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.59 $Y=0.87
+ $X2=4.48 $Y2=0.87
r202 26 29 5.41706 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=4.737 $Y=0.87
+ $X2=4.737 $Y2=1.035
r203 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.59
+ $Y=0.87 $X2=4.59 $Y2=0.87
r204 20 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.8 $Y=1.875
+ $X2=4.8 $Y2=1.74
r205 20 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.8 $Y=1.875 $X2=4.8
+ $Y2=2.275
r206 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=0.705
+ $X2=4.48 $Y2=0.87
r207 17 19 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.48 $Y=0.705
+ $X2=4.48 $Y2=0.415
r208 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.885 $Y=1.215
+ $X2=2.885 $Y2=0.415
r209 12 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=1.29
+ $X2=2.28 $Y2=1.29
r210 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=1.29
+ $X2=2.885 $Y2=1.215
r211 11 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.81 $Y=1.29
+ $X2=2.445 $Y2=1.29
r212 9 50 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.255 $Y=2.275
+ $X2=2.255 $Y2=1.485
r213 2 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r214 1 62 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%A_634_159# 1 2 9 13 15 18 25 29 31 33 34 39
r90 33 34 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.3
+ $X2=4.075 $Y2=2.135
r91 26 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.035 $Y=0.45
+ $X2=4.19 $Y2=0.45
r92 23 39 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=3.375 $Y=0.93 $X2=3.38
+ $Y2=0.93
r93 23 36 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=3.375 $Y=0.93
+ $X2=3.245 $Y2=0.93
r94 22 25 4.13427 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.375 $Y=0.93
+ $X2=3.49 $Y2=0.93
r95 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.375
+ $Y=0.93 $X2=3.375 $Y2=0.93
r96 19 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.035 $Y=1.065
+ $X2=4.035 $Y2=0.915
r97 19 34 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.035 $Y=1.065
+ $X2=4.035 $Y2=2.135
r98 18 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.035 $Y=0.765
+ $X2=4.035 $Y2=0.915
r99 17 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.535
+ $X2=4.035 $Y2=0.45
r100 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.035 $Y=0.535
+ $X2=4.035 $Y2=0.765
r101 15 31 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=0.915
+ $X2=4.035 $Y2=0.915
r102 15 25 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.95 $Y=0.915
+ $X2=3.49 $Y2=0.915
r103 11 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.38 $Y=0.795
+ $X2=3.38 $Y2=0.93
r104 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.38 $Y=0.795
+ $X2=3.38 $Y2=0.445
r105 7 36 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.245 $Y=1.065
+ $X2=3.245 $Y2=0.93
r106 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=3.245 $Y=1.065
+ $X2=3.245 $Y2=2.275
r107 2 33 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.735 $X2=4.115 $Y2=2.3
r108 1 29 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.05
+ $Y=0.235 $X2=4.19 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%A_466_413# 1 2 8 11 15 16 17 18 19 20 24 29
+ 30 31 33 34
c120 31 0 1.25128e-19 $X=3.08 $Y=1.4
c121 29 0 2.60836e-19 $X=2.995 $Y=1.315
r122 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.41 $X2=3.695 $Y2=1.41
r123 34 36 14.6572 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=3.355 $Y=1.41
+ $X2=3.695 $Y2=1.41
r124 32 34 3.71884 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=1.575
+ $X2=3.355 $Y2=1.41
r125 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.355 $Y=1.575
+ $X2=3.355 $Y2=2.19
r126 30 34 5.59441 $w=2.83e-07 $l=8.9861e-08 $layer=LI1_cond $X=3.27 $Y=1.4
+ $X2=3.355 $Y2=1.41
r127 30 31 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.27 $Y=1.4
+ $X2=3.08 $Y2=1.4
r128 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=1.315
+ $X2=3.08 $Y2=1.4
r129 28 29 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.995 $Y=0.535
+ $X2=2.995 $Y2=1.315
r130 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.91 $Y=0.45
+ $X2=2.995 $Y2=0.535
r131 24 26 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.91 $Y=0.45
+ $X2=2.6 $Y2=0.45
r132 20 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=2.275
+ $X2=3.355 $Y2=2.19
r133 20 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.27 $Y=2.275
+ $X2=2.5 $Y2=2.275
r134 18 37 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.41
+ $X2=3.695 $Y2=1.41
r135 18 19 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.83 $Y=1.41
+ $X2=3.905 $Y2=1.41
r136 16 17 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.94 $Y=0.95
+ $X2=3.94 $Y2=1.1
r137 15 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.975 $Y=0.555
+ $X2=3.975 $Y2=0.95
r138 9 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.905 $Y=1.545
+ $X2=3.905 $Y2=1.41
r139 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.905 $Y=1.545
+ $X2=3.905 $Y2=2.11
r140 8 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.905 $Y=1.275
+ $X2=3.905 $Y2=1.41
r141 8 17 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.905 $Y=1.275
+ $X2=3.905 $Y2=1.1
r142 2 22 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=2.065 $X2=2.5 $Y2=2.275
r143 1 26 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.6 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%A_1059_315# 1 2 9 13 17 19 21 22 25 29 33 36
+ 38 41 42 45 46 47
c90 42 0 2.71678e-19 $X=6.85 $Y=1.16
c91 13 0 2.06462e-20 $X=5.485 $Y=0.445
r92 48 50 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.37 $Y=1.74
+ $X2=5.485 $Y2=1.74
r93 42 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.85 $Y=1.16
+ $X2=6.85 $Y2=1.325
r94 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.16 $X2=6.85 $Y2=1.16
r95 39 47 0.463323 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=6.385 $Y=1.16
+ $X2=6.285 $Y2=1.16
r96 39 41 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.385 $Y=1.16
+ $X2=6.85 $Y2=1.16
r97 38 45 6.82437 $w=2.65e-07 $l=2.21346e-07 $layer=LI1_cond $X=6.28 $Y=1.53
+ $X2=6.205 $Y2=1.717
r98 37 47 7.80489 $w=1.95e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.28 $Y=1.325
+ $X2=6.285 $Y2=1.16
r99 37 38 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=6.28 $Y=1.325
+ $X2=6.28 $Y2=1.53
r100 36 47 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=6.285 $Y=0.995
+ $X2=6.285 $Y2=1.16
r101 36 46 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=6.285 $Y=0.995
+ $X2=6.285 $Y2=0.825
r102 31 46 7.53752 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.22 $Y=0.66
+ $X2=6.22 $Y2=0.825
r103 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.22 $Y=0.66
+ $X2=6.22 $Y2=0.385
r104 27 45 6.82437 $w=2.65e-07 $l=1.88e-07 $layer=LI1_cond $X=6.205 $Y=1.905
+ $X2=6.205 $Y2=1.717
r105 27 29 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=6.205 $Y=1.905
+ $X2=6.205 $Y2=2.34
r106 25 50 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.565 $Y=1.74
+ $X2=5.485 $Y2=1.74
r107 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.565
+ $Y=1.74 $X2=5.565 $Y2=1.74
r108 22 45 0.127723 $w=3.75e-07 $l=1.7e-07 $layer=LI1_cond $X=6.035 $Y=1.717
+ $X2=6.205 $Y2=1.717
r109 22 24 14.444 $w=3.73e-07 $l=4.7e-07 $layer=LI1_cond $X=6.035 $Y=1.717
+ $X2=5.565 $Y2=1.717
r110 19 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.85 $Y=0.995
+ $X2=6.85 $Y2=1.16
r111 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.85 $Y=0.995
+ $X2=6.85 $Y2=0.56
r112 17 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.84 $Y=1.985
+ $X2=6.84 $Y2=1.325
r113 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=1.575
+ $X2=5.485 $Y2=1.74
r114 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=5.485 $Y=1.575
+ $X2=5.485 $Y2=0.445
r115 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.37 $Y=1.905
+ $X2=5.37 $Y2=1.74
r116 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.37 $Y=1.905
+ $X2=5.37 $Y2=2.275
r117 2 45 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.075
+ $Y=1.485 $X2=6.2 $Y2=1.63
r118 2 29 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=6.075
+ $Y=1.485 $X2=6.2 $Y2=2.34
r119 1 33 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=6.095
+ $Y=0.235 $X2=6.22 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%A_891_413# 1 2 9 11 13 14 15 16 20 25 27 30
+ 33
c82 33 0 1.78258e-19 $X=5.225 $Y=1.16
c83 30 0 1.01102e-19 $X=5.93 $Y=1.16
c84 11 0 1.81857e-19 $X=6.43 $Y=0.995
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.93
+ $Y=1.16 $X2=5.93 $Y2=1.16
r86 28 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=1.16
+ $X2=5.225 $Y2=1.16
r87 28 30 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=5.31 $Y=1.16 $X2=5.93
+ $Y2=1.16
r88 26 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=1.325
+ $X2=5.225 $Y2=1.16
r89 26 27 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.225 $Y=1.325
+ $X2=5.225 $Y2=2.165
r90 25 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0.995
+ $X2=5.225 $Y2=1.16
r91 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.225 $Y=0.535
+ $X2=5.225 $Y2=0.995
r92 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=0.45
+ $X2=5.225 $Y2=0.535
r93 20 22 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.14 $Y=0.45
+ $X2=4.705 $Y2=0.45
r94 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=2.25
+ $X2=5.225 $Y2=2.165
r95 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.14 $Y=2.25
+ $X2=4.59 $Y2=2.25
r96 14 31 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=6.345 $Y=1.16
+ $X2=5.93 $Y2=1.16
r97 14 15 5.03009 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=6.345 $Y=1.16
+ $X2=6.425 $Y2=1.16
r98 11 15 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.425 $Y2=1.16
r99 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.995
+ $X2=6.43 $Y2=0.56
r100 7 15 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=6.42 $Y=1.325
+ $X2=6.425 $Y2=1.16
r101 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.42 $Y=1.325
+ $X2=6.42 $Y2=1.985
r102 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=2.065 $X2=4.59 $Y2=2.25
r103 1 22 182 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_NDIFF $count=1 $X=4.555
+ $Y=0.235 $X2=4.705 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 45 47 52 74 75 78 81
c114 75 0 1.81794e-19 $X=7.13 $Y=2.72
c115 1 0 3.29888e-20 $X=0.545 $Y=1.815
r116 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r117 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r119 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r120 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r121 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r122 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r123 66 69 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r124 65 68 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r125 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r126 63 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r127 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 60 63 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 60 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r130 59 62 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r131 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r132 57 81 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.572 $Y2=2.72
r133 57 59 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 56 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 56 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r137 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r138 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 52 81 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.572 $Y2=2.72
r140 52 55 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.15 $Y2=2.72
r141 47 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r142 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r143 45 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r144 45 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 43 71 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=6.21 $Y2=2.72
r146 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=6.63 $Y2=2.72
r147 42 74 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.715 $Y=2.72
+ $X2=7.13 $Y2=2.72
r148 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=2.72
+ $X2=6.63 $Y2=2.72
r149 40 68 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.49 $Y=2.72 $X2=5.29
+ $Y2=2.72
r150 40 41 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=5.49 $Y=2.72
+ $X2=5.647 $Y2=2.72
r151 39 71 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.805 $Y=2.72
+ $X2=6.21 $Y2=2.72
r152 39 41 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=5.805 $Y=2.72
+ $X2=5.647 $Y2=2.72
r153 37 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r154 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.695 $Y2=2.72
r155 36 65 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.91 $Y2=2.72
r156 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.695 $Y2=2.72
r157 32 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.63 $Y=2.635
+ $X2=6.63 $Y2=2.72
r158 32 34 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=6.63 $Y=2.635
+ $X2=6.63 $Y2=1.79
r159 28 41 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.647 $Y=2.635
+ $X2=5.647 $Y2=2.72
r160 28 30 12.2561 $w=3.13e-07 $l=3.35e-07 $layer=LI1_cond $X=5.647 $Y=2.635
+ $X2=5.647 $Y2=2.3
r161 24 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2.72
r162 24 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2
r163 20 81 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.572 $Y=2.635
+ $X2=1.572 $Y2=2.72
r164 20 22 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.572 $Y=2.635
+ $X2=1.572 $Y2=2.34
r165 16 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r166 16 18 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r167 5 34 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=6.495
+ $Y=1.485 $X2=6.63 $Y2=1.79
r168 4 30 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=2.065 $X2=5.585 $Y2=2.3
r169 3 26 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=3.32
+ $Y=2.065 $X2=3.695 $Y2=2
r170 2 22 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.065 $X2=1.62 $Y2=2.34
r171 1 18 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%A_381_47# 1 2 13 15 16 17 18 21
c49 18 0 1.74123e-19 $X=1.972 $Y=2.04
c50 15 0 1.97281e-19 $X=1.932 $Y=0.675
r51 17 18 7.17986 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.972 $Y=1.91
+ $X2=1.972 $Y2=2.04
r52 16 17 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=1.905 $Y=0.805
+ $X2=1.905 $Y2=1.91
r53 15 16 6.65856 $w=2.23e-07 $l=1.3e-07 $layer=LI1_cond $X=1.932 $Y=0.675
+ $X2=1.932 $Y2=0.805
r54 13 18 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2 $Y=2.3 $X2=2
+ $Y2=2.04
r55 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.535
+ $X2=1.96 $Y2=0.45
r56 9 15 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.96 $Y=0.535
+ $X2=1.96 $Y2=0.675
r57 2 13 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.065 $X2=2.04 $Y2=2.3
r58 1 21 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.045 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%Q 1 2 9 14 15 16 19
c31 19 0 1.81857e-19 $X=7.06 $Y=0.395
r32 16 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.06 $Y=0.51
+ $X2=7.06 $Y2=0.395
r33 15 16 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=7.06 $Y=0.74
+ $X2=7.06 $Y2=0.51
r34 13 15 4.62121 $w=3.3e-07 $l=1.82071e-07 $layer=LI1_cond $X=7.19 $Y=0.865
+ $X2=7.06 $Y2=0.74
r35 13 14 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.19 $Y=0.865
+ $X2=7.19 $Y2=1.445
r36 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.05 $Y=1.63 $X2=7.05
+ $Y2=2.31
r37 7 14 4.92547 $w=3.22e-07 $l=1.94422e-07 $layer=LI1_cond $X=7.05 $Y=1.575
+ $X2=7.19 $Y2=1.445
r38 7 9 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=7.05 $Y=1.575 $X2=7.05
+ $Y2=1.63
r39 2 11 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=6.915
+ $Y=1.485 $X2=7.05 $Y2=2.31
r40 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.915
+ $Y=1.485 $X2=7.05 $Y2=1.63
r41 1 19 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=6.925
+ $Y=0.235 $X2=7.06 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__DFXTP_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 42
+ 44 49 54 70 71 74 77 80
c111 71 0 2.71124e-20 $X=7.13 $Y=0
c112 34 0 1.70577e-19 $X=6.64 $Y=0.53
r113 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r114 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r115 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r117 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r118 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r119 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r120 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r121 62 65 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r122 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r123 61 64 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r124 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r125 59 80 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.77 $Y=0 $X2=3.585
+ $Y2=0
r126 59 61 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.77 $Y=0 $X2=3.91
+ $Y2=0
r127 58 81 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r128 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r129 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r130 55 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.58
+ $Y2=0
r131 55 57 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r132 54 80 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.585
+ $Y2=0
r133 54 57 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.4 $Y=0 $X2=2.07
+ $Y2=0
r134 53 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r135 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r136 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r137 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r138 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r139 49 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.58
+ $Y2=0
r140 49 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r141 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r142 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r143 42 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r144 42 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r145 40 67 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.21
+ $Y2=0
r146 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.64
+ $Y2=0
r147 39 70 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.725 $Y=0
+ $X2=7.13 $Y2=0
r148 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.725 $Y=0 $X2=6.64
+ $Y2=0
r149 37 64 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.585 $Y=0 $X2=5.29
+ $Y2=0
r150 37 38 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.585 $Y=0 $X2=5.69
+ $Y2=0
r151 36 67 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.795 $Y=0
+ $X2=6.21 $Y2=0
r152 36 38 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.69
+ $Y2=0
r153 32 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.64 $Y=0.085
+ $X2=6.64 $Y2=0
r154 32 34 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.64 $Y=0.085
+ $X2=6.64 $Y2=0.53
r155 28 38 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.69 $Y=0.085
+ $X2=5.69 $Y2=0
r156 28 30 19.2771 $w=2.08e-07 $l=3.65e-07 $layer=LI1_cond $X=5.69 $Y=0.085
+ $X2=5.69 $Y2=0.45
r157 24 80 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0
r158 24 26 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0.42
r159 20 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r160 20 22 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.38
r161 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r162 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r163 5 34 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.64 $Y2=0.53
r164 4 30 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.235 $X2=5.695 $Y2=0.45
r165 3 26 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.235 $X2=3.595 $Y2=0.42
r166 2 22 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r167 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__dfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=1.2195e+12p ps=1.255e+07u
M1001 a_1283_21# a_1108_47# a_1462_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u
M1002 a_805_47# a_761_289# a_639_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u
M1003 VGND RESET_B a_805_47# VNB nshort w=420000u l=150000u
+  ad=1.0617e+12p pd=9.62e+06u as=0p ps=0u
M1004 a_1462_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Q a_1283_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1006 a_651_413# a_193_47# a_543_47# VPB phighvt w=420000u l=150000u
+  ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u
M1007 VPWR a_1283_21# a_1270_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1008 a_543_47# a_193_47# a_448_47# VNB nshort w=360000u l=150000u
+  ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u
M1009 VPWR a_761_289# a_651_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1270_413# a_27_47# a_1108_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1011 VPWR CLK_N a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1012 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1013 VPWR a_1108_47# a_1283_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1014 a_761_289# a_543_47# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.583e+11p pd=2.37e+06u as=0p ps=0u
M1015 Q a_1283_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1016 a_1283_21# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_639_47# a_27_47# a_543_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1217_47# a_193_47# a_1108_47# VNB nshort w=360000u l=150000u
+  ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u
M1019 a_761_289# a_543_47# VGND VNB nshort w=640000u l=150000u
+  ad=1.998e+11p pd=1.97e+06u as=0p ps=0u
M1020 a_1108_47# a_27_47# a_761_289# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1108_47# a_193_47# a_761_289# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1283_21# a_1217_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1024 a_448_47# D VPWR VPB phighvt w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1025 a_448_47# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_543_47# a_27_47# a_448_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_651_413# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


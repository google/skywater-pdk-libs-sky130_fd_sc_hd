* File: sky130_fd_sc_hd__xnor2_4.pex.spice
* Created: Thu Aug 27 14:49:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XNOR2_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 43 45 48 50 52 55 58 59 60 62 63 68 71 72 84 92
c203 92 0 7.68269e-20 $X=7.375 $Y=1.16
c204 59 0 1.48557e-19 $X=5.56 $Y=1.53
c205 22 0 1.79953e-19 $X=1.805 $Y=0.995
r206 89 90 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.535 $Y=1.16
+ $X2=6.955 $Y2=1.16
r207 82 84 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.675 $Y=1.16
+ $X2=1.805 $Y2=1.16
r208 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r209 80 82 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.675 $Y2=1.16
r210 79 80 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=1.385 $Y2=1.16
r211 77 79 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.965 $Y2=1.16
r212 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.655
+ $Y=1.16 $X2=0.655 $Y2=1.16
r213 74 77 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.545 $Y=1.16
+ $X2=0.655 $Y2=1.16
r214 72 83 29.1136 $w=1.98e-07 $l=5.25e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=1.675 $Y2=1.175
r215 72 78 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=0.655 $Y2=1.175
r216 71 83 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=1.685 $Y=1.175
+ $X2=1.675 $Y2=1.175
r217 69 92 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.26 $Y=1.16
+ $X2=7.375 $Y2=1.16
r218 69 90 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=7.26 $Y=1.16
+ $X2=6.955 $Y2=1.16
r219 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.26
+ $Y=1.16 $X2=7.26 $Y2=1.16
r220 66 89 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=6.24 $Y=1.16
+ $X2=6.535 $Y2=1.16
r221 66 86 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.24 $Y=1.16
+ $X2=6.115 $Y2=1.16
r222 65 68 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=6.24 $Y=1.175
+ $X2=7.26 $Y2=1.175
r223 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.24
+ $Y=1.16 $X2=6.24 $Y2=1.16
r224 63 65 28.2818 $w=1.98e-07 $l=5.1e-07 $layer=LI1_cond $X=5.73 $Y=1.175
+ $X2=6.24 $Y2=1.175
r225 61 63 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.645 $Y=1.275
+ $X2=5.73 $Y2=1.175
r226 61 62 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.645 $Y=1.275
+ $X2=5.645 $Y2=1.445
r227 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.56 $Y=1.53
+ $X2=5.645 $Y2=1.445
r228 59 60 241.717 $w=1.68e-07 $l=3.705e-06 $layer=LI1_cond $X=5.56 $Y=1.53
+ $X2=1.855 $Y2=1.53
r229 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.77 $Y=1.445
+ $X2=1.855 $Y2=1.53
r230 57 71 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.77 $Y=1.275
+ $X2=1.685 $Y2=1.175
r231 57 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.77 $Y=1.275
+ $X2=1.77 $Y2=1.445
r232 53 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.375 $Y=1.325
+ $X2=7.375 $Y2=1.16
r233 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.375 $Y=1.325
+ $X2=7.375 $Y2=1.985
r234 50 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.375 $Y=0.995
+ $X2=7.375 $Y2=1.16
r235 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.375 $Y=0.995
+ $X2=7.375 $Y2=0.56
r236 46 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.955 $Y=1.325
+ $X2=6.955 $Y2=1.16
r237 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.955 $Y=1.325
+ $X2=6.955 $Y2=1.985
r238 43 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.955 $Y=0.995
+ $X2=6.955 $Y2=1.16
r239 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.955 $Y=0.995
+ $X2=6.955 $Y2=0.56
r240 39 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.535 $Y=1.325
+ $X2=6.535 $Y2=1.16
r241 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.535 $Y=1.325
+ $X2=6.535 $Y2=1.985
r242 36 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.535 $Y=0.995
+ $X2=6.535 $Y2=1.16
r243 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.535 $Y=0.995
+ $X2=6.535 $Y2=0.56
r244 32 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=1.325
+ $X2=6.115 $Y2=1.16
r245 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.115 $Y=1.325
+ $X2=6.115 $Y2=1.985
r246 29 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=0.995
+ $X2=6.115 $Y2=1.16
r247 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.115 $Y=0.995
+ $X2=6.115 $Y2=0.56
r248 25 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.325
+ $X2=1.805 $Y2=1.16
r249 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.805 $Y=1.325
+ $X2=1.805 $Y2=1.985
r250 22 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=0.995
+ $X2=1.805 $Y2=1.16
r251 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.805 $Y=0.995
+ $X2=1.805 $Y2=0.56
r252 18 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.16
r253 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.985
r254 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=0.995
+ $X2=1.385 $Y2=1.16
r255 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.385 $Y=0.995
+ $X2=1.385 $Y2=0.56
r256 11 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.325
+ $X2=0.965 $Y2=1.16
r257 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.965 $Y=1.325
+ $X2=0.965 $Y2=1.985
r258 8 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=0.995
+ $X2=0.965 $Y2=1.16
r259 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.965 $Y=0.995
+ $X2=0.965 $Y2=0.56
r260 4 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.325
+ $X2=0.545 $Y2=1.16
r261 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.545 $Y=1.325
+ $X2=0.545 $Y2=1.985
r262 1 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=1.16
r263 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 43 45 48 50 52 55 57 69 79 81
c152 79 0 7.68269e-20 $X=5.225 $Y=1.16
c153 1 0 8.27827e-20 $X=2.225 $Y=0.995
r154 80 81 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.275 $Y=1.16
+ $X2=5.695 $Y2=1.16
r155 78 80 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=5.225 $Y=1.16
+ $X2=5.275 $Y2=1.16
r156 78 79 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.225
+ $Y=1.16 $X2=5.225 $Y2=1.16
r157 76 78 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=4.855 $Y=1.16
+ $X2=5.225 $Y2=1.16
r158 75 79 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=4.545 $Y=1.175
+ $X2=5.225 $Y2=1.175
r159 74 76 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=4.545 $Y=1.16
+ $X2=4.855 $Y2=1.16
r160 74 75 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.545
+ $Y=1.16 $X2=4.545 $Y2=1.16
r161 71 74 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.435 $Y=1.16
+ $X2=4.545 $Y2=1.16
r162 67 69 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.37 $Y=1.16
+ $X2=3.485 $Y2=1.16
r163 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.37
+ $Y=1.16 $X2=3.37 $Y2=1.16
r164 65 67 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=3.065 $Y=1.16
+ $X2=3.37 $Y2=1.16
r165 64 65 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.645 $Y=1.16
+ $X2=3.065 $Y2=1.16
r166 63 68 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=2.35 $Y=1.175
+ $X2=3.37 $Y2=1.175
r167 62 64 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=2.35 $Y=1.16
+ $X2=2.645 $Y2=1.16
r168 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.35
+ $Y=1.16 $X2=2.35 $Y2=1.16
r169 59 62 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.35 $Y2=1.16
r170 57 75 35.2136 $w=1.98e-07 $l=6.35e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=4.545 $Y2=1.175
r171 57 68 29.9455 $w=1.98e-07 $l=5.4e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=3.37 $Y2=1.175
r172 53 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.325
+ $X2=5.695 $Y2=1.16
r173 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.695 $Y=1.325
+ $X2=5.695 $Y2=1.985
r174 50 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=0.995
+ $X2=5.695 $Y2=1.16
r175 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.695 $Y=0.995
+ $X2=5.695 $Y2=0.56
r176 46 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=1.325
+ $X2=5.275 $Y2=1.16
r177 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.275 $Y=1.325
+ $X2=5.275 $Y2=1.985
r178 43 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=0.995
+ $X2=5.275 $Y2=1.16
r179 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.275 $Y=0.995
+ $X2=5.275 $Y2=0.56
r180 39 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.325
+ $X2=4.855 $Y2=1.16
r181 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.855 $Y=1.325
+ $X2=4.855 $Y2=1.985
r182 36 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=0.995
+ $X2=4.855 $Y2=1.16
r183 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.855 $Y=0.995
+ $X2=4.855 $Y2=0.56
r184 32 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=1.325
+ $X2=4.435 $Y2=1.16
r185 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.435 $Y=1.325
+ $X2=4.435 $Y2=1.985
r186 29 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=0.995
+ $X2=4.435 $Y2=1.16
r187 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.435 $Y=0.995
+ $X2=4.435 $Y2=0.56
r188 25 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.325
+ $X2=3.485 $Y2=1.16
r189 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.485 $Y=1.325
+ $X2=3.485 $Y2=1.985
r190 22 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=0.995
+ $X2=3.485 $Y2=1.16
r191 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.485 $Y=0.995
+ $X2=3.485 $Y2=0.56
r192 18 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.325
+ $X2=3.065 $Y2=1.16
r193 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.065 $Y=1.325
+ $X2=3.065 $Y2=1.985
r194 15 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=0.995
+ $X2=3.065 $Y2=1.16
r195 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.065 $Y=0.995
+ $X2=3.065 $Y2=0.56
r196 11 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.325
+ $X2=2.645 $Y2=1.16
r197 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.645 $Y=1.325
+ $X2=2.645 $Y2=1.985
r198 8 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=0.995
+ $X2=2.645 $Y2=1.16
r199 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.645 $Y=0.995
+ $X2=2.645 $Y2=0.56
r200 4 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.325
+ $X2=2.225 $Y2=1.16
r201 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.225 $Y=1.325
+ $X2=2.225 $Y2=1.985
r202 1 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=0.995
+ $X2=2.225 $Y2=1.16
r203 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.225 $Y=0.995
+ $X2=2.225 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%A_38_297# 1 2 3 4 5 6 7 22 24 27 29 31 34 36
+ 38 41 43 45 48 51 54 58 62 64 66 72 76 80 85 86 91 94 96 98 100 102 103 104
+ 105 111 120
c212 111 0 1.48557e-19 $X=6.21 $Y=1.53
c213 62 0 8.27827e-20 $X=1.595 $Y=0.73
r214 117 118 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.755 $Y=1.16
+ $X2=9.175 $Y2=1.16
r215 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=1.53
+ $X2=6.21 $Y2=1.53
r216 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.53
+ $X2=1.15 $Y2=1.53
r217 105 107 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.53
+ $X2=1.15 $Y2=1.53
r218 104 111 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.065 $Y=1.53
+ $X2=6.21 $Y2=1.53
r219 104 105 5.90345 $w=1.4e-07 $l=4.77e-06 $layer=MET1_cond $X=6.065 $Y=1.53
+ $X2=1.295 $Y2=1.53
r220 103 112 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=7.6 $Y=1.53
+ $X2=6.21 $Y2=1.53
r221 92 120 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=9.465 $Y=1.16
+ $X2=9.595 $Y2=1.16
r222 92 118 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=9.465 $Y=1.16
+ $X2=9.175 $Y2=1.16
r223 91 92 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.465
+ $Y=1.16 $X2=9.465 $Y2=1.16
r224 89 117 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=8.445 $Y=1.16
+ $X2=8.755 $Y2=1.16
r225 89 114 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.445 $Y=1.16
+ $X2=8.335 $Y2=1.16
r226 88 91 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=8.445 $Y=1.175
+ $X2=9.465 $Y2=1.175
r227 88 89 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.445
+ $Y=1.16 $X2=8.445 $Y2=1.16
r228 86 88 37.4318 $w=1.98e-07 $l=6.75e-07 $layer=LI1_cond $X=7.77 $Y=1.175
+ $X2=8.445 $Y2=1.175
r229 85 103 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.685 $Y=1.445
+ $X2=7.6 $Y2=1.53
r230 84 86 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.685 $Y=1.275
+ $X2=7.77 $Y2=1.175
r231 84 85 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.685 $Y=1.275
+ $X2=7.685 $Y2=1.445
r232 81 100 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.98 $Y=1.895
+ $X2=2.855 $Y2=1.895
r233 80 102 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=3.57 $Y=1.895
+ $X2=3.695 $Y2=1.895
r234 80 81 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=3.57 $Y=1.895
+ $X2=2.98 $Y2=1.895
r235 77 98 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.14 $Y=1.895
+ $X2=2.015 $Y2=1.895
r236 76 100 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.73 $Y=1.895
+ $X2=2.855 $Y2=1.895
r237 76 77 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=2.73 $Y=1.895
+ $X2=2.14 $Y2=1.895
r238 73 96 1.80668 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.3 $Y=1.895
+ $X2=1.175 $Y2=1.895
r239 72 98 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.89 $Y=1.895
+ $X2=2.015 $Y2=1.895
r240 72 73 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=1.89 $Y=1.895
+ $X2=1.3 $Y2=1.895
r241 67 96 4.63873 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.175 $Y=1.785
+ $X2=1.175 $Y2=1.895
r242 67 69 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=1.785
+ $X2=1.175 $Y2=1.62
r243 66 108 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=1.615
+ $X2=1.175 $Y2=1.53
r244 66 69 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.175 $Y=1.615
+ $X2=1.175 $Y2=1.62
r245 65 94 3.51065 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.46 $Y=1.53
+ $X2=0.272 $Y2=1.53
r246 64 108 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.05 $Y=1.53
+ $X2=1.175 $Y2=1.53
r247 64 65 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.05 $Y=1.53
+ $X2=0.46 $Y2=1.53
r248 60 62 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=0.755 $Y=0.775
+ $X2=1.595 $Y2=0.775
r249 58 60 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=0.32 $Y=0.775
+ $X2=0.755 $Y2=0.775
r250 54 56 20.8976 $w=3.73e-07 $l=6.8e-07 $layer=LI1_cond $X=0.272 $Y=1.62
+ $X2=0.272 $Y2=2.3
r251 52 94 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.272 $Y=1.615
+ $X2=0.272 $Y2=1.53
r252 52 54 0.153659 $w=3.73e-07 $l=5e-09 $layer=LI1_cond $X=0.272 $Y=1.615
+ $X2=0.272 $Y2=1.62
r253 51 94 3.10218 $w=3.05e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.202 $Y=1.445
+ $X2=0.272 $Y2=1.53
r254 50 58 6.83913 $w=2.6e-07 $l=1.79555e-07 $layer=LI1_cond $X=0.202 $Y=0.905
+ $X2=0.32 $Y2=0.775
r255 50 51 26.4817 $w=2.33e-07 $l=5.4e-07 $layer=LI1_cond $X=0.202 $Y=0.905
+ $X2=0.202 $Y2=1.445
r256 46 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.595 $Y=1.325
+ $X2=9.595 $Y2=1.16
r257 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.595 $Y=1.325
+ $X2=9.595 $Y2=1.985
r258 43 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.595 $Y=0.995
+ $X2=9.595 $Y2=1.16
r259 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.595 $Y=0.995
+ $X2=9.595 $Y2=0.56
r260 39 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.175 $Y=1.325
+ $X2=9.175 $Y2=1.16
r261 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.175 $Y=1.325
+ $X2=9.175 $Y2=1.985
r262 36 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.175 $Y=0.995
+ $X2=9.175 $Y2=1.16
r263 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.175 $Y=0.995
+ $X2=9.175 $Y2=0.56
r264 32 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.755 $Y=1.325
+ $X2=8.755 $Y2=1.16
r265 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.755 $Y=1.325
+ $X2=8.755 $Y2=1.985
r266 29 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.755 $Y=0.995
+ $X2=8.755 $Y2=1.16
r267 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.755 $Y=0.995
+ $X2=8.755 $Y2=0.56
r268 25 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.335 $Y=1.325
+ $X2=8.335 $Y2=1.16
r269 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.335 $Y=1.325
+ $X2=8.335 $Y2=1.985
r270 22 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.335 $Y=0.995
+ $X2=8.335 $Y2=1.16
r271 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.335 $Y=0.995
+ $X2=8.335 $Y2=0.56
r272 7 102 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=1.485 $X2=3.695 $Y2=1.96
r273 6 100 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.72
+ $Y=1.485 $X2=2.855 $Y2=1.96
r274 5 98 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.88
+ $Y=1.485 $X2=2.015 $Y2=1.96
r275 4 96 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=1.485 $X2=1.175 $Y2=1.96
r276 4 69 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.485 $X2=1.175 $Y2=1.62
r277 3 56 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.485 $X2=0.335 $Y2=2.3
r278 3 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.485 $X2=0.335 $Y2=1.62
r279 2 62 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.235 $X2=1.595 $Y2=0.73
r280 1 60 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.235 $X2=0.755 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%VPWR 1 2 3 4 5 6 7 8 29 33 37 41 45 49 53 57
+ 60 61 63 64 66 67 69 70 72 73 74 76 97 109 110 113 116 119
r159 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r160 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r161 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r162 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r163 107 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r164 107 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r165 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r166 104 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.67 $Y=2.72
+ $X2=8.545 $Y2=2.72
r167 104 106 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.67 $Y=2.72
+ $X2=8.97 $Y2=2.72
r168 103 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r169 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r170 100 103 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=8.05 $Y2=2.72
r171 99 102 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=8.05 $Y2=2.72
r172 99 100 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r173 97 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.42 $Y=2.72
+ $X2=8.545 $Y2=2.72
r174 97 102 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.42 $Y=2.72
+ $X2=8.05 $Y2=2.72
r175 96 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r176 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r177 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r178 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r179 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r180 89 92 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r181 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r182 87 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r183 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r184 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r185 84 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r186 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r187 81 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.72 $Y=2.72
+ $X2=1.595 $Y2=2.72
r188 81 83 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.72 $Y=2.72
+ $X2=2.07 $Y2=2.72
r189 80 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r190 80 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r191 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r192 77 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.88 $Y=2.72
+ $X2=0.755 $Y2=2.72
r193 77 79 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.88 $Y=2.72
+ $X2=1.15 $Y2=2.72
r194 76 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.595 $Y2=2.72
r195 76 79 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.15 $Y2=2.72
r196 74 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r197 72 106 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.26 $Y=2.72
+ $X2=8.97 $Y2=2.72
r198 72 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.26 $Y=2.72
+ $X2=9.385 $Y2=2.72
r199 71 109 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.51 $Y=2.72
+ $X2=9.89 $Y2=2.72
r200 71 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.51 $Y=2.72
+ $X2=9.385 $Y2=2.72
r201 69 95 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.36 $Y=2.72 $X2=5.29
+ $Y2=2.72
r202 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.36 $Y=2.72
+ $X2=5.485 $Y2=2.72
r203 68 99 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.61 $Y=2.72
+ $X2=5.75 $Y2=2.72
r204 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.61 $Y=2.72
+ $X2=5.485 $Y2=2.72
r205 66 92 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.52 $Y=2.72
+ $X2=4.37 $Y2=2.72
r206 66 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.52 $Y=2.72
+ $X2=4.645 $Y2=2.72
r207 65 95 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.77 $Y=2.72
+ $X2=5.29 $Y2=2.72
r208 65 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.77 $Y=2.72
+ $X2=4.645 $Y2=2.72
r209 63 86 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r210 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.15 $Y=2.72
+ $X2=3.275 $Y2=2.72
r211 62 89 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.4 $Y=2.72 $X2=3.45
+ $Y2=2.72
r212 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.4 $Y=2.72
+ $X2=3.275 $Y2=2.72
r213 60 83 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.07 $Y2=2.72
r214 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.435 $Y2=2.72
r215 59 86 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.56 $Y=2.72
+ $X2=2.99 $Y2=2.72
r216 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.56 $Y=2.72
+ $X2=2.435 $Y2=2.72
r217 55 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.385 $Y=2.635
+ $X2=9.385 $Y2=2.72
r218 55 57 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=9.385 $Y=2.635
+ $X2=9.385 $Y2=2
r219 51 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=2.635
+ $X2=8.545 $Y2=2.72
r220 51 53 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.545 $Y=2.635
+ $X2=8.545 $Y2=2
r221 47 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=2.635
+ $X2=5.485 $Y2=2.72
r222 47 49 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.485 $Y=2.635
+ $X2=5.485 $Y2=2.34
r223 43 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=2.635
+ $X2=4.645 $Y2=2.72
r224 43 45 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.645 $Y=2.635
+ $X2=4.645 $Y2=2.34
r225 39 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=2.635
+ $X2=3.275 $Y2=2.72
r226 39 41 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.275 $Y=2.635
+ $X2=3.275 $Y2=2.34
r227 35 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=2.635
+ $X2=2.435 $Y2=2.72
r228 35 37 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.435 $Y=2.635
+ $X2=2.435 $Y2=2.34
r229 31 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=2.635
+ $X2=1.595 $Y2=2.72
r230 31 33 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.595 $Y=2.635
+ $X2=1.595 $Y2=2.34
r231 27 113 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=2.635
+ $X2=0.755 $Y2=2.72
r232 27 29 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.755 $Y=2.635
+ $X2=0.755 $Y2=2
r233 8 57 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.25
+ $Y=1.485 $X2=9.385 $Y2=2
r234 7 53 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.41
+ $Y=1.485 $X2=8.545 $Y2=2
r235 6 49 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.485 $X2=5.485 $Y2=2.34
r236 5 45 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.485 $X2=4.645 $Y2=2.34
r237 4 41 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.485 $X2=3.275 $Y2=2.34
r238 3 37 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=1.485 $X2=2.435 $Y2=2.34
r239 2 33 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.485 $X2=1.595 $Y2=2.34
r240 1 29 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.62
+ $Y=1.485 $X2=0.755 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%A_820_297# 1 2 3 4 5 18 22 24 25 30 33 35
r61 28 30 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=6.745 $Y=2.34
+ $X2=7.585 $Y2=2.34
r62 26 39 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.99 $Y=2.34
+ $X2=5.885 $Y2=2.34
r63 26 28 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=5.99 $Y=2.34
+ $X2=6.745 $Y2=2.34
r64 25 39 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=2.215
+ $X2=5.885 $Y2=2.34
r65 24 37 3.48996 $w=2.1e-07 $l=1.1e-07 $layer=LI1_cond $X=5.885 $Y=2.005
+ $X2=5.885 $Y2=1.895
r66 24 25 11.0909 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=5.885 $Y=2.005
+ $X2=5.885 $Y2=2.215
r67 23 35 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.19 $Y=1.895
+ $X2=5.065 $Y2=1.895
r68 22 37 3.33133 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=5.78 $Y=1.895
+ $X2=5.885 $Y2=1.895
r69 22 23 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=5.78 $Y=1.895
+ $X2=5.19 $Y2=1.895
r70 19 33 4.18571 $w=2.2e-07 $l=1.58e-07 $layer=LI1_cond $X=4.35 $Y=1.895
+ $X2=4.192 $Y2=1.895
r71 18 35 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.94 $Y=1.895
+ $X2=5.065 $Y2=1.895
r72 18 19 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=4.94 $Y=1.895
+ $X2=4.35 $Y2=1.895
r73 5 30 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.45
+ $Y=1.485 $X2=7.585 $Y2=2.3
r74 4 28 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.61
+ $Y=1.485 $X2=6.745 $Y2=2.3
r75 3 39 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.485 $X2=5.905 $Y2=2.3
r76 3 37 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.485 $X2=5.905 $Y2=1.96
r77 2 35 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.93
+ $Y=1.485 $X2=5.065 $Y2=1.96
r78 1 33 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.1
+ $Y=1.485 $X2=4.225 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%Y 1 2 3 4 5 6 7 22 30 32 34 42 44 47 48 54
+ 57 58
r76 58 63 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=9.857 $Y=1.87
+ $X2=9.857 $Y2=2.3
r77 55 58 6.65495 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=9.857 $Y=1.665
+ $X2=9.857 $Y2=1.87
r78 55 57 4.11246 $w=2.87e-07 $l=1.1e-07 $layer=LI1_cond $X=9.857 $Y=1.665
+ $X2=9.857 $Y2=1.555
r79 51 52 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=8.105 $Y=1.62
+ $X2=8.105 $Y2=1.915
r80 48 51 2.58306 $w=2.88e-07 $l=6.5e-08 $layer=LI1_cond $X=8.105 $Y=1.555
+ $X2=8.105 $Y2=1.62
r81 47 57 4.11246 $w=2.87e-07 $l=1.39929e-07 $layer=LI1_cond $X=9.925 $Y=1.445
+ $X2=9.857 $Y2=1.555
r82 46 47 28.2872 $w=2.18e-07 $l=5.4e-07 $layer=LI1_cond $X=9.925 $Y=0.905
+ $X2=9.925 $Y2=1.445
r83 45 54 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=9.09 $Y=1.555
+ $X2=8.965 $Y2=1.555
r84 44 57 2.32165 $w=2.2e-07 $l=1.77e-07 $layer=LI1_cond $X=9.68 $Y=1.555
+ $X2=9.857 $Y2=1.555
r85 44 45 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=9.68 $Y=1.555
+ $X2=9.09 $Y2=1.555
r86 40 54 0.886536 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.965 $Y=1.665
+ $X2=8.965 $Y2=1.555
r87 40 42 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.965 $Y=1.665
+ $X2=8.965 $Y2=2.3
r88 36 39 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=8.545 $Y=0.775
+ $X2=9.385 $Y2=0.775
r89 34 46 6.87824 $w=2.6e-07 $l=1.76635e-07 $layer=LI1_cond $X=9.815 $Y=0.775
+ $X2=9.925 $Y2=0.905
r90 34 39 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=9.815 $Y=0.775
+ $X2=9.385 $Y2=0.775
r91 33 48 2.35727 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=8.25 $Y=1.555
+ $X2=8.105 $Y2=1.555
r92 32 54 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.84 $Y=1.555
+ $X2=8.965 $Y2=1.555
r93 32 33 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=8.84 $Y=1.555
+ $X2=8.25 $Y2=1.555
r94 28 52 5.16612 $w=2.88e-07 $l=1.3e-07 $layer=LI1_cond $X=8.105 $Y=2.045
+ $X2=8.105 $Y2=1.915
r95 28 30 10.1336 $w=2.88e-07 $l=2.55e-07 $layer=LI1_cond $X=8.105 $Y=2.045
+ $X2=8.105 $Y2=2.3
r96 24 27 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=6.325 $Y=1.915
+ $X2=7.165 $Y2=1.915
r97 22 52 1.37394 $w=2.6e-07 $l=1.45e-07 $layer=LI1_cond $X=7.96 $Y=1.915
+ $X2=8.105 $Y2=1.915
r98 22 27 35.2382 $w=2.58e-07 $l=7.95e-07 $layer=LI1_cond $X=7.96 $Y=1.915
+ $X2=7.165 $Y2=1.915
r99 7 63 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.67
+ $Y=1.485 $X2=9.805 $Y2=2.3
r100 7 57 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.67
+ $Y=1.485 $X2=9.805 $Y2=1.62
r101 6 54 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=8.83
+ $Y=1.485 $X2=8.965 $Y2=1.62
r102 6 42 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.83
+ $Y=1.485 $X2=8.965 $Y2=2.3
r103 5 51 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.98
+ $Y=1.485 $X2=8.125 $Y2=1.62
r104 5 30 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.98
+ $Y=1.485 $X2=8.125 $Y2=2.3
r105 4 27 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=7.03
+ $Y=1.485 $X2=7.165 $Y2=1.96
r106 3 24 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=6.19
+ $Y=1.485 $X2=6.325 $Y2=1.96
r107 2 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=9.25
+ $Y=0.235 $X2=9.385 $Y2=0.73
r108 1 36 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=8.41
+ $Y=0.235 $X2=8.545 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%A_38_47# 1 2 3 4 5 16 22 23 24 28 30 34 40
c68 23 0 1.79953e-19 $X=2.055 $Y=0.725
r69 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.695 $Y=0.725
+ $X2=3.695 $Y2=0.39
r70 31 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0.815
+ $X2=2.855 $Y2=0.815
r71 30 32 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.53 $Y=0.815
+ $X2=3.695 $Y2=0.725
r72 30 31 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.53 $Y=0.815
+ $X2=3.02 $Y2=0.815
r73 26 40 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.855 $Y=0.725
+ $X2=2.855 $Y2=0.815
r74 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.855 $Y=0.725
+ $X2=2.855 $Y2=0.39
r75 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.18 $Y=0.815
+ $X2=2.055 $Y2=0.815
r76 24 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0.815
+ $X2=2.855 $Y2=0.815
r77 24 25 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.69 $Y=0.815
+ $X2=2.18 $Y2=0.815
r78 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.055 $Y=0.725
+ $X2=2.055 $Y2=0.815
r79 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2.055 $Y=0.475
+ $X2=2.055 $Y2=0.365
r80 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.055 $Y=0.475
+ $X2=2.055 $Y2=0.725
r81 18 21 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=0.335 $Y=0.365
+ $X2=1.175 $Y2=0.365
r82 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.93 $Y=0.365
+ $X2=2.055 $Y2=0.365
r83 16 21 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=1.93 $Y=0.365
+ $X2=1.175 $Y2=0.365
r84 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.235 $X2=3.695 $Y2=0.39
r85 4 28 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.72
+ $Y=0.235 $X2=2.855 $Y2=0.39
r86 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.015 $Y2=0.73
r87 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.015 $Y2=0.39
r88 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.235 $X2=1.175 $Y2=0.39
r89 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.235 $X2=0.335 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 46 50
+ 53 54 56 57 59 60 62 63 64 65 66 87 97 98 101 104
r155 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r156 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r157 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r158 95 98 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.89 $Y2=0
r159 95 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r160 94 97 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=8.05 $Y=0 $X2=9.89
+ $Y2=0
r161 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r162 92 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.77 $Y=0
+ $X2=7.635 $Y2=0
r163 92 94 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=8.05
+ $Y2=0
r164 91 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r165 91 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.67 $Y2=0
r166 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r167 88 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=0 $X2=6.745
+ $Y2=0
r168 88 90 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.83 $Y=0 $X2=7.13
+ $Y2=0
r169 87 104 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.5 $Y=0 $X2=7.635
+ $Y2=0
r170 87 90 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.5 $Y=0 $X2=7.13
+ $Y2=0
r171 86 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r172 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r173 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r174 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r175 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r176 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r177 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r178 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r179 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r180 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r181 69 73 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r182 66 74 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=2.07 $Y2=0
r183 66 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r184 64 85 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.82 $Y=0 $X2=5.75
+ $Y2=0
r185 64 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0 $X2=5.905
+ $Y2=0
r186 62 82 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.98 $Y=0 $X2=4.83
+ $Y2=0
r187 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0 $X2=5.065
+ $Y2=0
r188 61 85 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.75
+ $Y2=0
r189 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.065
+ $Y2=0
r190 59 79 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.035 $Y=0
+ $X2=3.91 $Y2=0
r191 59 60 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.035 $Y=0
+ $X2=4.172 $Y2=0
r192 58 82 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.83
+ $Y2=0
r193 58 60 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.172
+ $Y2=0
r194 56 76 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=2.99
+ $Y2=0
r195 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.275
+ $Y2=0
r196 55 79 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.91
+ $Y2=0
r197 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.275
+ $Y2=0
r198 53 73 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.07
+ $Y2=0
r199 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.435
+ $Y2=0
r200 52 76 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.52 $Y=0 $X2=2.99
+ $Y2=0
r201 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0 $X2=2.435
+ $Y2=0
r202 48 104 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.635 $Y=0.085
+ $X2=7.635 $Y2=0
r203 48 50 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.635 $Y=0.085
+ $X2=7.635 $Y2=0.39
r204 44 101 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0.085
+ $X2=6.745 $Y2=0
r205 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.745 $Y=0.085
+ $X2=6.745 $Y2=0.39
r206 43 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=0 $X2=5.905
+ $Y2=0
r207 42 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0 $X2=6.745
+ $Y2=0
r208 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.66 $Y=0 $X2=5.99
+ $Y2=0
r209 38 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0.085
+ $X2=5.905 $Y2=0
r210 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=0.085
+ $X2=5.905 $Y2=0.39
r211 34 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0.085
+ $X2=5.065 $Y2=0
r212 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.065 $Y=0.085
+ $X2=5.065 $Y2=0.39
r213 30 60 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.172 $Y=0.085
+ $X2=4.172 $Y2=0
r214 30 32 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=4.172 $Y=0.085
+ $X2=4.172 $Y2=0.39
r215 26 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=0.085
+ $X2=3.275 $Y2=0
r216 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.275 $Y=0.085
+ $X2=3.275 $Y2=0.39
r217 22 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0
r218 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0.39
r219 7 50 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.45
+ $Y=0.235 $X2=7.585 $Y2=0.39
r220 6 46 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.61
+ $Y=0.235 $X2=6.745 $Y2=0.39
r221 5 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.77
+ $Y=0.235 $X2=5.905 $Y2=0.39
r222 4 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.235 $X2=5.065 $Y2=0.39
r223 3 32 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=4.1
+ $Y=0.235 $X2=4.225 $Y2=0.39
r224 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.14
+ $Y=0.235 $X2=3.275 $Y2=0.39
r225 1 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.235 $X2=2.435 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_4%A_902_47# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 42 44 46 49 54 56 57 58
r118 52 54 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=8.965 $Y=0.39
+ $X2=9.805 $Y2=0.39
r119 50 60 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.21 $Y=0.39
+ $X2=8.085 $Y2=0.39
r120 50 52 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.21 $Y=0.39
+ $X2=8.965 $Y2=0.39
r121 47 49 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.085 $Y=0.735
+ $X2=8.085 $Y2=0.73
r122 46 60 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.085 $Y=0.475
+ $X2=8.085 $Y2=0.39
r123 46 49 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.085 $Y=0.475
+ $X2=8.085 $Y2=0.73
r124 45 58 8.43672 $w=1.75e-07 $l=2.17486e-07 $layer=LI1_cond $X=7.43 $Y=0.82
+ $X2=7.215 $Y2=0.815
r125 44 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.96 $Y=0.82
+ $X2=8.085 $Y2=0.735
r126 44 45 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.96 $Y=0.82
+ $X2=7.43 $Y2=0.82
r127 40 58 0.806278 $w=3.3e-07 $l=1.1225e-07 $layer=LI1_cond $X=7.165 $Y=0.725
+ $X2=7.215 $Y2=0.815
r128 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.165 $Y=0.725
+ $X2=7.165 $Y2=0.39
r129 39 57 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.49 $Y=0.815
+ $X2=6.325 $Y2=0.815
r130 38 58 8.43672 $w=1.75e-07 $l=2.15e-07 $layer=LI1_cond $X=7 $Y=0.815
+ $X2=7.215 $Y2=0.815
r131 38 39 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7 $Y=0.815 $X2=6.49
+ $Y2=0.815
r132 34 57 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.325 $Y=0.725
+ $X2=6.325 $Y2=0.815
r133 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.325 $Y=0.725
+ $X2=6.325 $Y2=0.39
r134 33 56 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.65 $Y=0.815
+ $X2=5.485 $Y2=0.815
r135 32 57 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.16 $Y=0.815
+ $X2=6.325 $Y2=0.815
r136 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.16 $Y=0.815
+ $X2=5.65 $Y2=0.815
r137 28 56 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.485 $Y=0.725
+ $X2=5.485 $Y2=0.815
r138 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.485 $Y=0.725
+ $X2=5.485 $Y2=0.39
r139 26 56 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=0.815
+ $X2=5.485 $Y2=0.815
r140 26 27 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.32 $Y=0.815
+ $X2=4.81 $Y2=0.815
r141 22 27 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.645 $Y=0.725
+ $X2=4.81 $Y2=0.815
r142 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.645 $Y=0.725
+ $X2=4.645 $Y2=0.39
r143 7 54 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.67
+ $Y=0.235 $X2=9.805 $Y2=0.39
r144 6 52 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.83
+ $Y=0.235 $X2=8.965 $Y2=0.39
r145 5 60 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=8
+ $Y=0.235 $X2=8.125 $Y2=0.39
r146 5 49 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=8
+ $Y=0.235 $X2=8.125 $Y2=0.73
r147 4 42 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.03
+ $Y=0.235 $X2=7.165 $Y2=0.39
r148 3 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.19
+ $Y=0.235 $X2=6.325 $Y2=0.39
r149 2 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.35
+ $Y=0.235 $X2=5.485 $Y2=0.39
r150 1 24 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.51
+ $Y=0.235 $X2=4.645 $Y2=0.39
.ends


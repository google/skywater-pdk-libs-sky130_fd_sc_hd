* File: sky130_fd_sc_hd__a2bb2oi_1.spice
* Created: Thu Aug 27 14:03:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2bb2oi_1.spice.pex"
.subckt sky130_fd_sc_hd__a2bb2oi_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1008 N_A_109_47#_M1008_d N_A1_N_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_N_M1006_g N_A_109_47#_M1008_d VNB NSHORT L=0.15
+ W=0.65 AD=0.28275 AS=0.08775 PD=1.52 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_A_109_47#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.28275 PD=0.92 PS=1.52 NRD=0 NRS=47.076 M=1 R=4.33333
+ SA=75001.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1001 A_481_47# N_B2_M1001_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75002 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g A_481_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75002.5 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1007 A_109_297# N_A1_N_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.105
+ AS=0.26 PD=1.21 PS=2.52 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75000.5
+ A=0.15 P=2.3 MULT=1
MM1005 N_A_109_47#_M1005_d N_A2_N_M1005_g A_109_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_397_297#_M1003_d N_A_109_47#_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.34 PD=1.27 PS=2.68 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75000.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_B2_M1000_g N_A_397_297#_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_A_397_297#_M1009_d N_B1_M1009_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a2bb2oi_1.spice.SKY130_FD_SC_HD__A2BB2OI_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__einvn_8.spice
* Created: Thu Aug 27 14:20:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__einvn_8.pex.spice"
.subckt sky130_fd_sc_hd__einvn_8  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1030 N_VGND_M1030_d N_TE_B_M1030_g N_A_27_47#_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_215_47#_M1008_d N_A_27_47#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75006.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_215_47#_M1009_d N_A_27_47#_M1009_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75006.1 A=0.0975 P=1.6 MULT=1
MM1012 N_A_215_47#_M1009_d N_A_27_47#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75005.7 A=0.0975 P=1.6 MULT=1
MM1014 N_A_215_47#_M1014_d N_A_27_47#_M1014_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1015 N_A_215_47#_M1014_d N_A_27_47#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1017 N_A_215_47#_M1017_d N_A_27_47#_M1017_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1018 N_A_215_47#_M1017_d N_A_27_47#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75004 A=0.0975 P=1.6 MULT=1
MM1021 N_A_215_47#_M1021_d N_A_27_47#_M1021_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.105625 AS=0.08775 PD=0.975 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_215_47#_M1021_d N_A_M1002_g N_Z_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.08775 PD=0.975 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75003.6 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1003 N_A_215_47#_M1003_d N_A_M1003_g N_Z_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1004 N_A_215_47#_M1003_d N_A_M1004_g N_Z_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1011 N_A_215_47#_M1011_d N_A_M1011_g N_Z_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1027 N_A_215_47#_M1011_d N_A_M1027_g N_Z_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1031 N_A_215_47#_M1031_d N_A_M1031_g N_Z_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1032 N_A_215_47#_M1031_d N_A_M1032_g N_Z_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1033 N_A_215_47#_M1033_d N_A_M1033_g N_Z_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1023 N_VPWR_M1023_d N_TE_B_M1023_g N_A_27_47#_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165206 AS=0.26 PD=1.36598 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1023_d N_TE_B_M1000_g N_A_204_309#_M1000_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.155294 AS=0.1269 PD=1.28402 PS=1.21 NRD=10.4607 NRS=0 M=1
+ R=6.26667 SA=75000.7 SB=75003.1 A=0.141 P=2.18 MULT=1
MM1005 N_VPWR_M1005_d N_TE_B_M1005_g N_A_204_309#_M1000_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75001.1 SB=75002.7 A=0.141 P=2.18 MULT=1
MM1006 N_VPWR_M1005_d N_TE_B_M1006_g N_A_204_309#_M1006_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75001.5 SB=75002.3 A=0.141 P=2.18 MULT=1
MM1010 N_VPWR_M1010_d N_TE_B_M1010_g N_A_204_309#_M1006_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75001.9 SB=75001.9 A=0.141 P=2.18 MULT=1
MM1013 N_VPWR_M1010_d N_TE_B_M1013_g N_A_204_309#_M1013_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75002.3 SB=75001.4 A=0.141 P=2.18 MULT=1
MM1016 N_VPWR_M1016_d N_TE_B_M1016_g N_A_204_309#_M1013_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75002.8 SB=75001 A=0.141 P=2.18 MULT=1
MM1024 N_VPWR_M1016_d N_TE_B_M1024_g N_A_204_309#_M1024_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667
+ SA=75003.2 SB=75000.6 A=0.141 P=2.18 MULT=1
MM1028 N_VPWR_M1028_d N_TE_B_M1028_g N_A_204_309#_M1024_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.2444 AS=0.1269 PD=2.4 PS=1.21 NRD=0 NRS=0 M=1 R=6.26667 SA=75003.6
+ SB=75000.2 A=0.141 P=2.18 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g N_A_204_309#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1007 N_Z_M1001_d N_A_M1007_g N_A_204_309#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1019 N_Z_M1019_d N_A_M1019_g N_A_204_309#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1020 N_Z_M1019_d N_A_M1020_g N_A_204_309#_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1022 N_Z_M1022_d N_A_M1022_g N_A_204_309#_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1025 N_Z_M1022_d N_A_M1025_g N_A_204_309#_M1025_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1026 N_Z_M1026_d N_A_M1026_g N_A_204_309#_M1025_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1029 N_Z_M1026_d N_A_M1029_g N_A_204_309#_M1029_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX34_noxref VNB VPB NWDIODE A=13.8993 P=20.53
*
.include "sky130_fd_sc_hd__einvn_8.pxi.spice"
*
.ends
*
*

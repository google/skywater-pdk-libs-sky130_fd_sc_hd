* File: sky130_fd_sc_hd__clkinvlp_4.pex.spice
* Created: Thu Aug 27 14:13:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKINVLP_4%A 3 7 11 15 19 23 27 31 33 34 48
c69 33 0 1.46135e-19 $X=0.23 $Y=0.85
r70 47 48 85.682 $w=3.3e-07 $l=4.9e-07 $layer=POLY_cond $X=1.625 $Y=1.16
+ $X2=2.115 $Y2=1.16
r71 46 47 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.585 $Y=1.16
+ $X2=1.625 $Y2=1.16
r72 45 46 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.265 $Y=1.16
+ $X2=1.585 $Y2=1.16
r73 44 45 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.055 $Y=1.16
+ $X2=1.265 $Y2=1.16
r74 43 44 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.835 $Y=1.16
+ $X2=1.055 $Y2=1.16
r75 42 43 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.525 $Y=1.16
+ $X2=0.835 $Y2=1.16
r76 41 42 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.16
+ $X2=0.525 $Y2=1.16
r77 38 41 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.315 $Y=1.16
+ $X2=0.475 $Y2=1.16
r78 34 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=1.16 $X2=0.315 $Y2=1.16
r79 33 34 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.255 $Y=0.85
+ $X2=0.255 $Y2=1.16
r80 29 48 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.325
+ $X2=2.115 $Y2=1.16
r81 29 31 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.115 $Y=1.325
+ $X2=2.115 $Y2=1.985
r82 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=0.995
+ $X2=1.625 $Y2=1.16
r83 25 27 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.625 $Y=0.995
+ $X2=1.625 $Y2=0.51
r84 21 46 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.325
+ $X2=1.585 $Y2=1.16
r85 21 23 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.585 $Y=1.325
+ $X2=1.585 $Y2=1.985
r86 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=0.995
+ $X2=1.265 $Y2=1.16
r87 17 19 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.265 $Y=0.995
+ $X2=1.265 $Y2=0.51
r88 13 44 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.325
+ $X2=1.055 $Y2=1.16
r89 13 15 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.055 $Y=1.325
+ $X2=1.055 $Y2=1.985
r90 9 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=0.995
+ $X2=0.835 $Y2=1.16
r91 9 11 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.835 $Y=0.995
+ $X2=0.835 $Y2=0.51
r92 5 42 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.16
r93 5 7 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.985
r94 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r95 1 3 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINVLP_4%VPWR 1 2 3 10 12 18 22 24 29 30 31 37 46
r40 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 40 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r42 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 37 45 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.487 $Y2=2.72
r44 37 39 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 36 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 33 42 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r48 33 35 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 31 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 31 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 29 35 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.155 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=2.72
+ $X2=1.32 $Y2=2.72
r53 28 39 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.485 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=2.72
+ $X2=1.32 $Y2=2.72
r55 24 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.38 $Y=1.63 $X2=2.38
+ $Y2=2.34
r56 22 45 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.487 $Y2=2.72
r57 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.38 $Y2=2.34
r58 18 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.32 $Y=1.63 $X2=1.32
+ $Y2=2.34
r59 16 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=2.635
+ $X2=1.32 $Y2=2.72
r60 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.32 $Y=2.635
+ $X2=1.32 $Y2=2.34
r61 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r62 10 42 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r63 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r64 3 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.485 $X2=2.38 $Y2=2.34
r65 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.485 $X2=2.38 $Y2=1.63
r66 2 21 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.485 $X2=1.32 $Y2=2.34
r67 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.485 $X2=1.32 $Y2=1.63
r68 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r69 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINVLP_4%Y 1 2 3 10 14 18 19 20 21 22 23 51
r40 49 51 7.45698 $w=4.23e-07 $l=2.75e-07 $layer=LI1_cond $X=0.775 $Y=0.467
+ $X2=1.05 $Y2=0.467
r41 30 49 1.7104 $w=3.6e-07 $l=2.13e-07 $layer=LI1_cond $X=0.775 $Y=0.68
+ $X2=0.775 $Y2=0.467
r42 23 44 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.775 $Y=2.21
+ $X2=0.775 $Y2=2.34
r43 22 23 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.775 $Y=1.87
+ $X2=0.775 $Y2=2.21
r44 22 38 7.68295 $w=3.58e-07 $l=2.4e-07 $layer=LI1_cond $X=0.775 $Y=1.87
+ $X2=0.775 $Y2=1.63
r45 21 38 3.20123 $w=3.58e-07 $l=1e-07 $layer=LI1_cond $X=0.775 $Y=1.53
+ $X2=0.775 $Y2=1.63
r46 21 34 7.52289 $w=3.58e-07 $l=2.35e-07 $layer=LI1_cond $X=0.775 $Y=1.53
+ $X2=0.775 $Y2=1.295
r47 20 31 4.17112 $w=3.6e-07 $l=1.4e-07 $layer=LI1_cond $X=0.775 $Y=1.155
+ $X2=0.775 $Y2=1.015
r48 20 34 4.17112 $w=3.6e-07 $l=1.4e-07 $layer=LI1_cond $X=0.775 $Y=1.155
+ $X2=0.775 $Y2=1.295
r49 19 31 5.28203 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=0.85
+ $X2=0.775 $Y2=1.015
r50 19 30 5.44209 $w=3.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.775 $Y=0.85
+ $X2=0.775 $Y2=0.68
r51 18 49 2.30489 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.467
+ $X2=0.775 $Y2=0.467
r52 14 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.85 $Y=1.63 $X2=1.85
+ $Y2=2.34
r53 12 14 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.85 $Y=1.295
+ $X2=1.85 $Y2=1.63
r54 11 20 2.26131 $w=2.8e-07 $l=1.8e-07 $layer=LI1_cond $X=0.955 $Y=1.155
+ $X2=0.775 $Y2=1.155
r55 10 12 6.87623 $w=2.8e-07 $l=2.24332e-07 $layer=LI1_cond $X=1.685 $Y=1.155
+ $X2=1.85 $Y2=1.295
r56 10 11 30.0458 $w=2.78e-07 $l=7.3e-07 $layer=LI1_cond $X=1.685 $Y=1.155
+ $X2=0.955 $Y2=1.155
r57 3 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.485 $X2=1.85 $Y2=2.34
r58 3 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.485 $X2=1.85 $Y2=1.63
r59 2 44 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.485 $X2=0.79 $Y2=2.34
r60 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.485 $X2=0.79 $Y2=1.63
r61 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINVLP_4%VGND 1 2 7 9 13 16 17 18 28 29
c31 7 0 1.46135e-19 $X=0.26 $Y=0.085
r32 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r33 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r34 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r35 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r36 22 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r37 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r38 20 32 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r39 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r40 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r41 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r42 16 25 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.61
+ $Y2=0
r43 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.84
+ $Y2=0
r44 15 28 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.53
+ $Y2=0
r45 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.84
+ $Y2=0
r46 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r47 11 13 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.51
r48 7 32 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r49 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.43
r50 2 13 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=1.84 $Y2=0.51
r51 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends


* File: sky130_fd_sc_hd__nor4_1.spice.SKY130_FD_SC_HD__NOR4_1.pxi
* Created: Thu Aug 27 14:32:41 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4_1%D N_D_c_45_n N_D_M1007_g N_D_M1005_g D D N_D_c_47_n
+ PM_SKY130_FD_SC_HD__NOR4_1%D
x_PM_SKY130_FD_SC_HD__NOR4_1%C N_C_M1004_g N_C_M1003_g N_C_c_75_n N_C_c_76_n C
+ N_C_c_77_n N_C_c_81_n PM_SKY130_FD_SC_HD__NOR4_1%C
x_PM_SKY130_FD_SC_HD__NOR4_1%B N_B_c_121_n N_B_M1002_g N_B_M1000_g N_B_c_122_n
+ N_B_c_123_n B PM_SKY130_FD_SC_HD__NOR4_1%B
x_PM_SKY130_FD_SC_HD__NOR4_1%A N_A_c_162_n N_A_M1001_g N_A_M1006_g A N_A_c_164_n
+ PM_SKY130_FD_SC_HD__NOR4_1%A
x_PM_SKY130_FD_SC_HD__NOR4_1%Y N_Y_M1007_d N_Y_M1002_d N_Y_M1005_s N_Y_c_194_n
+ N_Y_c_190_n N_Y_c_211_n N_Y_c_192_n N_Y_c_221_n Y PM_SKY130_FD_SC_HD__NOR4_1%Y
x_PM_SKY130_FD_SC_HD__NOR4_1%VPWR N_VPWR_M1006_d N_VPWR_c_246_n N_VPWR_c_247_n
+ VPWR N_VPWR_c_248_n N_VPWR_c_245_n PM_SKY130_FD_SC_HD__NOR4_1%VPWR
x_PM_SKY130_FD_SC_HD__NOR4_1%VGND N_VGND_M1007_s N_VGND_M1003_d N_VGND_M1001_d
+ N_VGND_c_272_n N_VGND_c_273_n N_VGND_c_274_n N_VGND_c_275_n N_VGND_c_276_n
+ VGND N_VGND_c_277_n N_VGND_c_278_n N_VGND_c_279_n N_VGND_c_280_n
+ PM_SKY130_FD_SC_HD__NOR4_1%VGND
cc_1 VNB N_D_c_45_n 0.0196026f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB D 0.0213668f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_D_c_47_n 0.0365032f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_C_c_75_n 0.00306446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_C_c_76_n 0.0209081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_C_c_77_n 0.0170942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_121_n 0.016263f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_B_c_122_n 0.019478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_c_123_n 0.0047678f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_10 VNB B 8.26803e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_c_162_n 0.0185152f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_12 VNB A 0.0253118f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_13 VNB N_A_c_164_n 0.0369005f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_14 VNB N_Y_c_190_n 0.00293422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_245_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_272_n 0.00988671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_273_n 0.0184315f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_18 VNB N_VGND_c_274_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_19 VNB N_VGND_c_275_n 0.0102656f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=0.85
cc_20 VNB N_VGND_c_276_n 0.0125842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_277_n 0.0177782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_278_n 0.0121123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_279_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_280_n 0.141132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_D_M1005_g 0.0252354f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_26 VPB D 0.00299612f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_27 VPB N_D_c_47_n 0.00976713f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_28 VPB N_C_M1004_g 0.0192016f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_29 VPB N_C_c_75_n 0.0012565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_C_c_76_n 0.00478764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_C_c_81_n 0.00373943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_B_M1000_g 0.0192797f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB N_B_c_122_n 0.00560678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB B 0.00120416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_M1006_g 0.0221377f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB A 0.0148428f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_37 VPB N_A_c_164_n 0.0112741f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_38 VPB N_Y_c_190_n 0.00105672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_192_n 0.00742573f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=0.85
cc_40 VPB Y 0.0310196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_246_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_42 VPB N_VPWR_c_247_n 0.030224f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_43 VPB N_VPWR_c_248_n 0.0568135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_245_n 0.0429403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 N_D_M1005_g N_C_M1004_g 0.0594214f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_46 N_D_c_47_n N_C_c_75_n 3.91349e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_47 N_D_c_47_n N_C_c_76_n 0.0161574f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_48 N_D_c_45_n N_C_c_77_n 0.0209519f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_49 N_D_c_45_n N_Y_c_194_n 0.00924059f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_50 D N_Y_c_194_n 0.00646135f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_51 N_D_c_45_n N_Y_c_190_n 0.00344066f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_52 N_D_M1005_g N_Y_c_190_n 0.00822876f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_53 D N_Y_c_190_n 0.0354406f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_54 N_D_c_47_n N_Y_c_190_n 0.00776423f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_55 N_D_M1005_g N_Y_c_192_n 0.0138543f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_56 D N_Y_c_192_n 0.0190584f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_D_c_47_n N_Y_c_192_n 0.00291752f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_58 N_D_M1005_g Y 0.015112f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_59 N_D_M1005_g N_VPWR_c_248_n 0.00541964f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_60 N_D_M1005_g N_VPWR_c_245_n 0.0106574f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_61 D N_VGND_M1007_s 0.00402345f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_62 N_D_c_45_n N_VGND_c_273_n 0.00450677f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_63 D N_VGND_c_273_n 0.021476f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_64 N_D_c_47_n N_VGND_c_273_n 0.00125865f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_65 N_D_c_45_n N_VGND_c_274_n 0.00163214f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_66 N_D_c_45_n N_VGND_c_277_n 0.00542994f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_67 N_D_c_45_n N_VGND_c_280_n 0.0105094f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_68 D N_VGND_c_280_n 0.00102136f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_69 N_C_c_77_n N_B_c_121_n 0.0250335f $X=0.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_70 N_C_M1004_g N_B_M1000_g 0.0321711f $X=0.88 $Y=1.985 $X2=0 $Y2=0
cc_71 N_C_c_75_n N_B_M1000_g 6.94586e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_72 N_C_c_81_n N_B_M1000_g 0.00133462f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_73 N_C_c_75_n N_B_c_122_n 0.00277064f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_74 N_C_c_76_n N_B_c_122_n 0.0208957f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_75 N_C_c_81_n N_B_c_122_n 2.47458e-19 $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_76 N_C_c_75_n N_B_c_123_n 0.0140108f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C_c_76_n N_B_c_123_n 5.71225e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_78 N_C_c_81_n N_B_c_123_n 0.00301186f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_79 N_C_M1004_g B 4.19685e-19 $X=0.88 $Y=1.985 $X2=0 $Y2=0
cc_80 N_C_c_75_n B 0.00699672f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_81 N_C_c_81_n B 0.0100784f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_82 N_C_c_75_n N_Y_c_194_n 8.46486e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_83 N_C_c_76_n N_Y_c_194_n 0.00236955f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_84 N_C_M1004_g N_Y_c_190_n 9.90588e-19 $X=0.88 $Y=1.985 $X2=0 $Y2=0
cc_85 N_C_c_75_n N_Y_c_190_n 0.0306798f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_86 N_C_c_76_n N_Y_c_190_n 0.00205802f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_87 N_C_c_77_n N_Y_c_190_n 0.00336265f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_88 N_C_c_81_n N_Y_c_190_n 0.0060866f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_89 N_C_c_75_n N_Y_c_211_n 0.0135231f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_90 N_C_c_77_n N_Y_c_211_n 0.0107092f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_91 N_C_c_81_n N_Y_c_211_n 0.00461545f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_92 N_C_M1004_g N_Y_c_192_n 0.00127917f $X=0.88 $Y=1.985 $X2=0 $Y2=0
cc_93 N_C_c_81_n N_Y_c_192_n 0.0121833f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_94 N_C_M1004_g Y 0.00239003f $X=0.88 $Y=1.985 $X2=0 $Y2=0
cc_95 N_C_c_81_n Y 0.0219504f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_96 N_C_c_81_n A_191_297# 0.0273559f $X=1.157 $Y=1.615 $X2=-0.19 $Y2=-0.24
cc_97 N_C_M1004_g N_VPWR_c_248_n 0.00585385f $X=0.88 $Y=1.985 $X2=0 $Y2=0
cc_98 N_C_c_81_n N_VPWR_c_248_n 0.0160407f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_99 N_C_M1004_g N_VPWR_c_245_n 0.0110983f $X=0.88 $Y=1.985 $X2=0 $Y2=0
cc_100 N_C_c_81_n N_VPWR_c_245_n 0.0097455f $X=1.157 $Y=1.615 $X2=0 $Y2=0
cc_101 N_C_c_77_n N_VGND_c_274_n 0.00902243f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_102 N_C_c_77_n N_VGND_c_277_n 0.00355956f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_103 N_C_c_77_n N_VGND_c_280_n 0.00442282f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_104 N_B_c_121_n N_A_c_162_n 0.0233891f $X=1.41 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_105 N_B_M1000_g N_A_M1006_g 0.0557039f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B_c_122_n A 5.58023e-19 $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B_c_123_n A 0.00980363f $X=1.575 $Y=1.245 $X2=0 $Y2=0
cc_108 B A 0.0189062f $X=1.525 $Y=1.785 $X2=0 $Y2=0
cc_109 N_B_c_122_n N_A_c_164_n 0.0212338f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B_c_123_n N_A_c_164_n 0.00153916f $X=1.575 $Y=1.245 $X2=0 $Y2=0
cc_111 B N_A_c_164_n 0.0129772f $X=1.525 $Y=1.785 $X2=0 $Y2=0
cc_112 N_B_c_121_n N_Y_c_211_n 0.0103436f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_122_n N_Y_c_211_n 0.00122295f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B_c_123_n N_Y_c_211_n 0.0119758f $X=1.575 $Y=1.245 $X2=0 $Y2=0
cc_115 N_B_c_123_n N_Y_c_221_n 0.00939151f $X=1.575 $Y=1.245 $X2=0 $Y2=0
cc_116 B A_297_297# 0.0127489f $X=1.525 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_117 N_B_M1000_g N_VPWR_c_248_n 0.00541964f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_118 B N_VPWR_c_248_n 0.013407f $X=1.525 $Y=1.785 $X2=0 $Y2=0
cc_119 N_B_M1000_g N_VPWR_c_245_n 0.0100523f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_120 B N_VPWR_c_245_n 0.00896636f $X=1.525 $Y=1.785 $X2=0 $Y2=0
cc_121 N_B_c_121_n N_VGND_c_274_n 0.00774927f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_121_n N_VGND_c_276_n 8.33085e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_121_n N_VGND_c_278_n 0.00341689f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_121_n N_VGND_c_280_n 0.00405445f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_125 A N_VPWR_M1006_d 0.00404422f $X=1.985 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_126 N_A_M1006_g N_VPWR_c_247_n 0.00450677f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_127 A N_VPWR_c_247_n 0.022894f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_128 N_A_c_164_n N_VPWR_c_247_n 9.13389e-19 $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_M1006_g N_VPWR_c_248_n 0.00585385f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_M1006_g N_VPWR_c_245_n 0.0115954f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_131 A N_VGND_M1001_d 0.00389911f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_132 N_A_c_162_n N_VGND_c_274_n 8.33085e-19 $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_162_n N_VGND_c_276_n 0.00988319f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_134 A N_VGND_c_276_n 0.0206507f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_135 N_A_c_164_n N_VGND_c_276_n 8.93814e-19 $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_162_n N_VGND_c_278_n 0.0046653f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_162_n N_VGND_c_280_n 0.00799591f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_138 A N_VGND_c_280_n 0.00151946f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_139 N_Y_c_190_n A_109_297# 2.95377e-19 $X=0.59 $Y=1.495 $X2=-0.19 $Y2=-0.24
cc_140 N_Y_c_192_n A_109_297# 0.00452621f $X=0.59 $Y=1.58 $X2=-0.19 $Y2=-0.24
cc_141 Y N_VPWR_c_248_n 0.0195303f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_142 N_Y_M1005_s N_VPWR_c_245_n 0.00209863f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_143 Y N_VPWR_c_245_n 0.012527f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_144 N_Y_c_211_n N_VGND_M1003_d 0.00455769f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_145 N_Y_c_211_n N_VGND_c_274_n 0.0160859f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_146 N_Y_c_194_n N_VGND_c_277_n 0.0108093f $X=0.59 $Y=0.825 $X2=0 $Y2=0
cc_147 N_Y_c_211_n N_VGND_c_277_n 0.00240209f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_148 N_Y_c_211_n N_VGND_c_278_n 0.00232396f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_149 N_Y_c_221_n N_VGND_c_278_n 0.00600088f $X=1.62 $Y=0.55 $X2=0 $Y2=0
cc_150 N_Y_M1007_d N_VGND_c_280_n 0.00348005f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_151 N_Y_M1002_d N_VGND_c_280_n 0.00423098f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_152 N_Y_c_194_n N_VGND_c_280_n 0.0118726f $X=0.59 $Y=0.825 $X2=0 $Y2=0
cc_153 N_Y_c_211_n N_VGND_c_280_n 0.00982733f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_154 N_Y_c_221_n N_VGND_c_280_n 0.00592513f $X=1.62 $Y=0.55 $X2=0 $Y2=0
cc_155 A_109_297# N_VPWR_c_245_n 0.0111139f $X=0.545 $Y=1.485 $X2=0.682 $Y2=0.55
cc_156 A_191_297# N_VPWR_c_245_n 0.00739666f $X=0.955 $Y=1.485 $X2=0 $Y2=0
cc_157 A_297_297# N_VPWR_c_245_n 0.00429012f $X=1.485 $Y=1.485 $X2=0 $Y2=0

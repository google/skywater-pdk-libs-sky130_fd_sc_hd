* File: sky130_fd_sc_hd__nand3_4.spice.SKY130_FD_SC_HD__NAND3_4.pxi
* Created: Thu Aug 27 14:29:39 2020
* 
x_PM_SKY130_FD_SC_HD__NAND3_4%C N_C_M1008_g N_C_M1002_g N_C_M1010_g N_C_M1003_g
+ N_C_M1013_g N_C_M1014_g N_C_c_106_n N_C_M1023_g N_C_M1020_g C C C C
+ PM_SKY130_FD_SC_HD__NAND3_4%C
x_PM_SKY130_FD_SC_HD__NAND3_4%B N_B_M1011_g N_B_M1000_g N_B_M1015_g N_B_M1004_g
+ N_B_M1018_g N_B_M1017_g N_B_M1019_g N_B_M1021_g B B B B N_B_c_200_n
+ PM_SKY130_FD_SC_HD__NAND3_4%B
x_PM_SKY130_FD_SC_HD__NAND3_4%A N_A_M1006_g N_A_M1001_g N_A_M1009_g N_A_M1005_g
+ N_A_M1012_g N_A_M1007_g N_A_M1016_g N_A_M1022_g A A A A N_A_c_286_n
+ N_A_c_287_n PM_SKY130_FD_SC_HD__NAND3_4%A
x_PM_SKY130_FD_SC_HD__NAND3_4%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1020_s
+ N_VPWR_M1004_s N_VPWR_M1021_s N_VPWR_M1001_s N_VPWR_M1005_s N_VPWR_M1022_s
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n
+ N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n
+ N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n
+ N_VPWR_c_367_n N_VPWR_c_368_n VPWR N_VPWR_c_369_n N_VPWR_c_370_n
+ N_VPWR_c_351_n N_VPWR_c_372_n N_VPWR_c_373_n PM_SKY130_FD_SC_HD__NAND3_4%VPWR
x_PM_SKY130_FD_SC_HD__NAND3_4%Y N_Y_M1006_d N_Y_M1012_d N_Y_M1002_d N_Y_M1014_d
+ N_Y_M1000_d N_Y_M1017_d N_Y_M1001_d N_Y_M1007_d N_Y_c_447_n N_Y_c_464_n
+ N_Y_c_448_n N_Y_c_471_n N_Y_c_449_n N_Y_c_476_n N_Y_c_450_n N_Y_c_491_n
+ N_Y_c_451_n N_Y_c_507_n N_Y_c_452_n N_Y_c_514_n N_Y_c_453_n N_Y_c_454_n
+ N_Y_c_455_n N_Y_c_456_n N_Y_c_457_n Y Y Y N_Y_c_446_n
+ PM_SKY130_FD_SC_HD__NAND3_4%Y
x_PM_SKY130_FD_SC_HD__NAND3_4%A_27_47# N_A_27_47#_M1008_d N_A_27_47#_M1010_d
+ N_A_27_47#_M1023_d N_A_27_47#_M1015_s N_A_27_47#_M1019_s N_A_27_47#_c_578_n
+ N_A_27_47#_c_579_n N_A_27_47#_c_580_n N_A_27_47#_c_597_n N_A_27_47#_c_581_n
+ N_A_27_47#_c_582_n N_A_27_47#_c_583_n N_A_27_47#_c_584_n N_A_27_47#_c_585_n
+ N_A_27_47#_c_586_n N_A_27_47#_c_587_n PM_SKY130_FD_SC_HD__NAND3_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND3_4%VGND N_VGND_M1008_s N_VGND_M1013_s N_VGND_c_663_n
+ N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n N_VGND_c_668_n
+ VGND N_VGND_c_669_n N_VGND_c_670_n PM_SKY130_FD_SC_HD__NAND3_4%VGND
x_PM_SKY130_FD_SC_HD__NAND3_4%A_445_47# N_A_445_47#_M1011_d N_A_445_47#_M1018_d
+ N_A_445_47#_M1006_s N_A_445_47#_M1009_s N_A_445_47#_M1016_s
+ N_A_445_47#_c_735_n PM_SKY130_FD_SC_HD__NAND3_4%A_445_47#
cc_1 VNB N_C_M1008_g 0.0230765f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_C_M1010_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_C_M1003_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_4 VNB N_C_M1013_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_5 VNB N_C_M1014_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_6 VNB N_C_c_106_n 0.0849196f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.025
cc_7 VNB N_C_M1023_g 0.0175697f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_8 VNB N_C_M1020_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_9 VNB C 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_10 VNB N_B_M1011_g 0.0175697f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_11 VNB N_B_M1000_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_12 VNB N_B_M1015_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_13 VNB N_B_M1004_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_14 VNB N_B_M1018_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_15 VNB N_B_M1017_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_16 VNB N_B_M1019_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_17 VNB N_B_M1021_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_18 VNB B 0.0057433f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_19 VNB N_B_c_200_n 0.0626315f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_20 VNB N_A_M1006_g 0.023925f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_A_M1001_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_22 VNB N_A_M1009_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_23 VNB N_A_M1005_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_24 VNB N_A_M1012_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_25 VNB N_A_M1007_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_26 VNB N_A_M1016_g 0.021463f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_27 VNB N_A_M1022_g 5.40111e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_28 VNB A 0.0040376f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_29 VNB N_A_c_286_n 0.032981f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_30 VNB N_A_c_287_n 0.0615271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_351_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB Y 0.0383338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_446_n 0.015438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_578_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_35 VNB N_A_27_47#_c_579_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_c_580_n 0.00922665f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.295
cc_37 VNB N_A_27_47#_c_581_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_582_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_39 VNB N_A_27_47#_c_583_n 0.00359609f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_40 VNB N_A_27_47#_c_584_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_27_47#_c_585_n 0.00219816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_586_n 0.00792198f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_43 VNB N_A_27_47#_c_587_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_44 VNB N_VGND_c_663_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_45 VNB N_VGND_c_664_n 0.00415222f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_46 VNB N_VGND_c_665_n 0.0171909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_666_n 0.00323658f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_48 VNB N_VGND_c_667_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_49 VNB N_VGND_c_668_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_669_n 0.115396f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_51 VNB N_VGND_c_670_n 0.320571f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_52 VNB N_A_445_47#_c_735_n 0.0196325f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_53 VPB N_C_M1002_g 0.0263683f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_54 VPB N_C_M1003_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_55 VPB N_C_M1014_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_56 VPB N_C_c_106_n 0.00805825f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.025
cc_57 VPB N_C_M1020_g 0.0194869f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_58 VPB N_B_M1000_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_59 VPB N_B_M1004_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_60 VPB N_B_M1017_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_61 VPB N_B_M1021_g 0.026721f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_62 VPB N_A_M1001_g 0.026721f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_63 VPB N_A_M1005_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_64 VPB N_A_M1007_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_65 VPB N_A_M1022_g 0.0238675f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_66 VPB N_VPWR_c_352_n 0.00994749f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.025
cc_67 VPB N_VPWR_c_353_n 0.0459243f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_68 VPB N_VPWR_c_354_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_69 VPB N_VPWR_c_355_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_356_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_71 VPB N_VPWR_c_357_n 0.0153464f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_72 VPB N_VPWR_c_358_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_73 VPB N_VPWR_c_359_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_360_n 0.0296314f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_75 VPB N_VPWR_c_361_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.175
cc_76 VPB N_VPWR_c_362_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_363_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_364_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_365_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_366_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_367_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_368_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_369_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_370_n 0.016145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_351_n 0.057553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_372_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_373_n 0.00506799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_Y_c_447_n 0.00223815f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.025
cc_89 VPB N_Y_c_448_n 0.00219943f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.295
cc_90 VPB N_Y_c_449_n 0.0035864f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_91 VPB N_Y_c_450_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_92 VPB N_Y_c_451_n 0.014171f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_93 VPB N_Y_c_452_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Y_c_453_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_Y_c_454_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_Y_c_455_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_Y_c_456_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_457_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB Y 0.00788001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB Y 0.0322602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 N_C_M1023_g N_B_M1011_g 0.024325f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_102 N_C_M1020_g N_B_M1000_g 0.024325f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_103 N_C_c_106_n B 0.00184043f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_104 C B 0.0118174f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_105 N_C_c_106_n N_B_c_200_n 0.024325f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_106 N_C_M1002_g N_VPWR_c_353_n 0.0041053f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_C_c_106_n N_VPWR_c_353_n 0.00550986f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_108 C N_VPWR_c_353_n 0.0190809f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_109 N_C_M1003_g N_VPWR_c_354_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_110 N_C_M1014_g N_VPWR_c_354_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_111 N_C_M1020_g N_VPWR_c_355_n 0.00146448f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_112 N_C_M1002_g N_VPWR_c_361_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_113 N_C_M1003_g N_VPWR_c_361_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_114 N_C_M1014_g N_VPWR_c_363_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_115 N_C_M1020_g N_VPWR_c_363_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_116 N_C_M1002_g N_VPWR_c_351_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_117 N_C_M1003_g N_VPWR_c_351_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_118 N_C_M1014_g N_VPWR_c_351_n 0.00950154f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_119 N_C_M1020_g N_VPWR_c_351_n 0.00952874f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_120 N_C_M1002_g N_Y_c_447_n 0.00331821f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_121 N_C_M1003_g N_Y_c_447_n 0.00149073f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_122 N_C_c_106_n N_Y_c_447_n 0.00206439f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_123 C N_Y_c_447_n 0.026643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_124 N_C_M1002_g N_Y_c_464_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_125 N_C_M1003_g N_Y_c_464_n 0.00975139f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C_M1014_g N_Y_c_464_n 6.1949e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_127 N_C_M1003_g N_Y_c_448_n 0.0120357f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_128 N_C_M1014_g N_Y_c_448_n 0.0120357f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_129 N_C_c_106_n N_Y_c_448_n 0.0019951f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_130 C N_Y_c_448_n 0.0366837f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_131 N_C_M1003_g N_Y_c_471_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_132 N_C_M1014_g N_Y_c_471_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C_M1020_g N_Y_c_471_n 0.00975139f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_134 N_C_M1020_g N_Y_c_449_n 0.0132678f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_135 C N_Y_c_449_n 0.00101487f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_136 N_C_M1020_g N_Y_c_476_n 6.1949e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_137 N_C_M1014_g N_Y_c_453_n 0.00149073f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_138 N_C_c_106_n N_Y_c_453_n 0.00206439f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_139 N_C_M1020_g N_Y_c_453_n 0.00149073f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_140 C N_Y_c_453_n 0.026643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_141 N_C_M1008_g N_A_27_47#_c_578_n 0.00641402f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_142 N_C_M1010_g N_A_27_47#_c_578_n 5.25091e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_143 N_C_M1008_g N_A_27_47#_c_579_n 0.00850187f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_144 N_C_M1010_g N_A_27_47#_c_579_n 0.00850187f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_145 N_C_c_106_n N_A_27_47#_c_579_n 0.00205431f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_146 C N_A_27_47#_c_579_n 0.0359512f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_147 N_C_M1008_g N_A_27_47#_c_580_n 0.00126954f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_148 N_C_c_106_n N_A_27_47#_c_580_n 0.00693855f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_149 C N_A_27_47#_c_580_n 0.0254514f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_150 N_C_M1008_g N_A_27_47#_c_597_n 5.25176e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_151 N_C_M1010_g N_A_27_47#_c_597_n 0.00641402f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_152 N_C_M1013_g N_A_27_47#_c_597_n 0.0065125f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_153 N_C_M1023_g N_A_27_47#_c_597_n 7.07818e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_154 N_C_M1010_g N_A_27_47#_c_581_n 0.00110555f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_155 N_C_M1013_g N_A_27_47#_c_581_n 0.00110555f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_156 N_C_c_106_n N_A_27_47#_c_581_n 0.00213429f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_157 C N_A_27_47#_c_581_n 0.0265408f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_158 N_C_M1013_g N_A_27_47#_c_582_n 0.00850187f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_159 N_C_c_106_n N_A_27_47#_c_582_n 0.00205431f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_160 N_C_M1023_g N_A_27_47#_c_582_n 0.00939924f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_161 C N_A_27_47#_c_582_n 0.0308372f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_162 N_C_M1013_g N_A_27_47#_c_583_n 2.32235e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_163 N_C_M1023_g N_A_27_47#_c_583_n 0.00351435f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_164 N_C_M1008_g N_VGND_c_663_n 0.00268723f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_165 N_C_M1010_g N_VGND_c_663_n 0.00146448f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_166 N_C_M1013_g N_VGND_c_664_n 0.00146448f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_167 N_C_M1023_g N_VGND_c_664_n 0.00268723f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_168 N_C_M1008_g N_VGND_c_665_n 0.00424416f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_169 N_C_M1010_g N_VGND_c_667_n 0.00424416f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_170 N_C_M1013_g N_VGND_c_667_n 0.00424416f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_171 N_C_M1023_g N_VGND_c_669_n 0.00436969f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_172 N_C_M1008_g N_VGND_c_670_n 0.00669028f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_173 N_C_M1010_g N_VGND_c_670_n 0.00573607f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_174 N_C_M1013_g N_VGND_c_670_n 0.00573607f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_175 N_C_M1023_g N_VGND_c_670_n 0.0059446f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_176 N_C_M1023_g N_A_445_47#_c_735_n 6.89492e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_177 B A 0.0121822f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_178 N_B_c_200_n A 8.71733e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_179 B N_A_c_286_n 8.07044e-19 $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_180 N_B_c_200_n N_A_c_286_n 0.00741568f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B_M1000_g N_VPWR_c_355_n 0.00146448f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B_M1004_g N_VPWR_c_356_n 0.00146448f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B_M1017_g N_VPWR_c_356_n 0.00146448f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B_M1021_g N_VPWR_c_357_n 0.0033532f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B_M1000_g N_VPWR_c_365_n 0.00541359f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B_M1004_g N_VPWR_c_365_n 0.00541359f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B_M1017_g N_VPWR_c_369_n 0.00541359f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B_M1021_g N_VPWR_c_369_n 0.00541359f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B_M1000_g N_VPWR_c_351_n 0.00952874f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B_M1004_g N_VPWR_c_351_n 0.00950154f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_191 N_B_M1017_g N_VPWR_c_351_n 0.00950154f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B_M1021_g N_VPWR_c_351_n 0.0108276f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B_M1000_g N_Y_c_471_n 6.1949e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B_M1000_g N_Y_c_449_n 0.0119784f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_195 B N_Y_c_449_n 0.0149743f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_196 N_B_M1000_g N_Y_c_476_n 0.00975139f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B_M1004_g N_Y_c_476_n 0.00975139f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B_M1017_g N_Y_c_476_n 6.1949e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B_M1004_g N_Y_c_450_n 0.0120357f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B_M1017_g N_Y_c_450_n 0.0120357f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_201 B N_Y_c_450_n 0.0366837f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_202 N_B_c_200_n N_Y_c_450_n 0.0019951f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B_M1004_g N_Y_c_491_n 6.1949e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_204 N_B_M1017_g N_Y_c_491_n 0.00975139f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B_M1021_g N_Y_c_491_n 0.0145598f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B_M1021_g N_Y_c_451_n 0.0147646f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_207 B N_Y_c_451_n 0.0126419f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_208 N_B_M1000_g N_Y_c_454_n 0.00149073f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B_M1004_g N_Y_c_454_n 0.00149073f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_210 B N_Y_c_454_n 0.026643f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_211 N_B_c_200_n N_Y_c_454_n 0.00206439f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B_M1017_g N_Y_c_455_n 0.00149073f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B_M1021_g N_Y_c_455_n 0.00149073f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_214 B N_Y_c_455_n 0.026643f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_215 N_B_c_200_n N_Y_c_455_n 0.00206439f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B_M1011_g N_A_27_47#_c_583_n 0.0031423f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_217 N_B_M1015_g N_A_27_47#_c_583_n 2.32132e-19 $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_218 B N_A_27_47#_c_583_n 0.111538f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_219 N_B_M1011_g N_A_27_47#_c_584_n 0.00823396f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_220 N_B_M1015_g N_A_27_47#_c_584_n 0.00743915f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_221 N_B_c_200_n N_A_27_47#_c_584_n 0.00205431f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B_M1011_g N_A_27_47#_c_585_n 2.32132e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_223 N_B_M1015_g N_A_27_47#_c_585_n 0.00286631f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_224 N_B_M1018_g N_A_27_47#_c_585_n 0.00286631f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_225 N_B_M1019_g N_A_27_47#_c_585_n 2.32132e-19 $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_226 N_B_c_200_n N_A_27_47#_c_585_n 0.00207461f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B_M1018_g N_A_27_47#_c_586_n 2.32132e-19 $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_228 N_B_M1019_g N_A_27_47#_c_586_n 0.00302029f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_229 N_B_M1018_g N_A_27_47#_c_587_n 0.00743915f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_230 N_B_M1019_g N_A_27_47#_c_587_n 0.00743915f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_231 N_B_c_200_n N_A_27_47#_c_587_n 0.00205431f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B_M1011_g N_VGND_c_669_n 0.00420703f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_233 N_B_M1015_g N_VGND_c_669_n 0.00357877f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_234 N_B_M1018_g N_VGND_c_669_n 0.00357877f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_235 N_B_M1019_g N_VGND_c_669_n 0.00357877f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_236 N_B_M1011_g N_VGND_c_670_n 0.00590125f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B_M1015_g N_VGND_c_670_n 0.00522516f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B_M1018_g N_VGND_c_670_n 0.00522516f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B_M1019_g N_VGND_c_670_n 0.00660224f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B_M1011_g N_A_445_47#_c_735_n 0.00501478f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_241 N_B_M1015_g N_A_445_47#_c_735_n 0.00956495f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B_M1018_g N_A_445_47#_c_735_n 0.00956495f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_243 N_B_M1019_g N_A_445_47#_c_735_n 0.012419f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_244 N_A_M1001_g N_VPWR_c_357_n 0.0033532f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_M1005_g N_VPWR_c_358_n 0.00146448f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A_M1007_g N_VPWR_c_358_n 0.00146448f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_M1007_g N_VPWR_c_359_n 0.00541359f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_M1022_g N_VPWR_c_359_n 0.00541359f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_M1022_g N_VPWR_c_360_n 0.00322031f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_M1001_g N_VPWR_c_367_n 0.00541359f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A_M1005_g N_VPWR_c_367_n 0.00541359f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_M1001_g N_VPWR_c_351_n 0.0108276f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_M1005_g N_VPWR_c_351_n 0.00950154f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A_M1007_g N_VPWR_c_351_n 0.00950154f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A_M1022_g N_VPWR_c_351_n 0.0108276f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A_M1001_g N_Y_c_451_n 0.0147646f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_257 A N_Y_c_451_n 0.0400987f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_258 N_A_c_286_n N_Y_c_451_n 0.00729564f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_M1001_g N_Y_c_507_n 0.0145598f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_M1005_g N_Y_c_507_n 0.00975139f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A_M1007_g N_Y_c_507_n 6.1949e-19 $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A_M1005_g N_Y_c_452_n 0.0120357f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_M1007_g N_Y_c_452_n 0.0120357f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_264 A N_Y_c_452_n 0.0366837f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_265 N_A_c_287_n N_Y_c_452_n 0.0019951f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_M1005_g N_Y_c_514_n 6.1949e-19 $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A_M1007_g N_Y_c_514_n 0.00975139f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A_M1022_g N_Y_c_514_n 0.0145598f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A_M1001_g N_Y_c_456_n 0.00149073f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_M1005_g N_Y_c_456_n 0.00149073f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_271 A N_Y_c_456_n 0.026643f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_272 N_A_c_287_n N_Y_c_456_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_M1007_g N_Y_c_457_n 0.00149073f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A_M1022_g N_Y_c_457_n 0.00149073f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_275 A N_Y_c_457_n 0.026643f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_276 N_A_c_287_n N_Y_c_457_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_M1006_g Y 0.00636949f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A_M1009_g Y 0.0107009f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A_M1012_g Y 0.0107009f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_280 N_A_M1016_g Y 0.0289239f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_281 A Y 0.0924613f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_282 N_A_c_287_n Y 0.00622382f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A_M1022_g Y 0.0160095f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A_M1006_g N_A_27_47#_c_586_n 0.0042433f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A_M1006_g N_VGND_c_669_n 0.00357877f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_M1009_g N_VGND_c_669_n 0.00357877f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_M1012_g N_VGND_c_669_n 0.00357877f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A_M1016_g N_VGND_c_669_n 0.00357877f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A_M1006_g N_VGND_c_670_n 0.00655123f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_M1009_g N_VGND_c_670_n 0.00522516f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A_M1012_g N_VGND_c_670_n 0.00522516f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A_M1016_g N_VGND_c_670_n 0.00655123f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_M1006_g N_A_445_47#_c_735_n 0.0108017f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A_M1009_g N_A_445_47#_c_735_n 0.00918728f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_295 N_A_M1012_g N_A_445_47#_c_735_n 0.00918728f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_296 N_A_M1016_g N_A_445_47#_c_735_n 0.00918728f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_297 A N_A_445_47#_c_735_n 0.0144225f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_298 N_A_c_286_n N_A_445_47#_c_735_n 0.00531811f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_299 N_VPWR_c_351_n N_Y_M1002_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_300 N_VPWR_c_351_n N_Y_M1014_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_c_351_n N_Y_M1000_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_302 N_VPWR_c_351_n N_Y_M1017_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_303 N_VPWR_c_351_n N_Y_M1001_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_304 N_VPWR_c_351_n N_Y_M1007_d 0.00215201f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_305 N_VPWR_c_353_n N_Y_c_447_n 0.0108343f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_306 N_VPWR_c_361_n N_Y_c_464_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_307 N_VPWR_c_351_n N_Y_c_464_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_308 N_VPWR_M1003_s N_Y_c_448_n 0.00167154f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_309 N_VPWR_c_354_n N_Y_c_448_n 0.0129161f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_310 N_VPWR_c_363_n N_Y_c_471_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_311 N_VPWR_c_351_n N_Y_c_471_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_312 N_VPWR_M1020_s N_Y_c_449_n 0.00167154f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_313 N_VPWR_c_355_n N_Y_c_449_n 0.0129161f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_314 N_VPWR_c_365_n N_Y_c_476_n 0.0189039f $X=2.695 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_c_351_n N_Y_c_476_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_316 N_VPWR_M1004_s N_Y_c_450_n 0.00167154f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_317 N_VPWR_c_356_n N_Y_c_450_n 0.0129161f $X=2.78 $Y=2 $X2=0 $Y2=0
cc_318 N_VPWR_c_369_n N_Y_c_491_n 0.0189039f $X=3.535 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_c_351_n N_Y_c_491_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_M1021_s N_Y_c_451_n 0.00296777f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_321 N_VPWR_M1001_s N_Y_c_451_n 0.00296777f $X=4.015 $Y=1.485 $X2=0 $Y2=0
cc_322 N_VPWR_c_357_n N_Y_c_451_n 0.0568271f $X=3.62 $Y=2 $X2=0 $Y2=0
cc_323 N_VPWR_c_367_n N_Y_c_507_n 0.0189039f $X=4.895 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_c_351_n N_Y_c_507_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_325 N_VPWR_M1005_s N_Y_c_452_n 0.00167154f $X=4.845 $Y=1.485 $X2=0 $Y2=0
cc_326 N_VPWR_c_358_n N_Y_c_452_n 0.0129161f $X=4.98 $Y=2 $X2=0 $Y2=0
cc_327 N_VPWR_c_359_n N_Y_c_514_n 0.0189039f $X=5.735 $Y=2.72 $X2=0 $Y2=0
cc_328 N_VPWR_c_351_n N_Y_c_514_n 0.0122217f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_329 N_VPWR_M1022_s Y 0.00317399f $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_330 N_VPWR_c_360_n Y 0.0214182f $X=5.82 $Y=2 $X2=0 $Y2=0
cc_331 N_VPWR_c_353_n N_A_27_47#_c_580_n 7.91944e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_332 N_Y_c_449_n N_A_27_47#_c_582_n 0.00939305f $X=2.195 $Y=1.555 $X2=0 $Y2=0
cc_333 N_Y_c_451_n N_A_27_47#_c_586_n 0.00869712f $X=4.395 $Y=1.555 $X2=0 $Y2=0
cc_334 Y N_A_27_47#_c_586_n 0.0082021f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_335 Y N_VGND_c_669_n 0.00224394f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_336 N_Y_c_446_n N_VGND_c_669_n 0.00448298f $X=6.24 $Y=0.905 $X2=0 $Y2=0
cc_337 N_Y_M1006_d N_VGND_c_670_n 0.00216833f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_338 N_Y_M1012_d N_VGND_c_670_n 0.00216833f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_339 Y N_VGND_c_670_n 0.00659949f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_340 N_Y_c_446_n N_VGND_c_670_n 0.00681927f $X=6.24 $Y=0.905 $X2=0 $Y2=0
cc_341 Y N_A_445_47#_M1009_s 0.00162409f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_342 Y N_A_445_47#_M1016_s 0.00335828f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_343 N_Y_M1006_d N_A_445_47#_c_735_n 0.0030596f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_344 N_Y_M1012_d N_A_445_47#_c_735_n 0.0030596f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_345 Y N_A_445_47#_c_735_n 0.0853982f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_579_n N_VGND_M1008_s 0.00162006f $X=0.935 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_347 N_A_27_47#_c_582_n N_VGND_M1013_s 0.00162006f $X=1.775 $Y=0.78 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_579_n N_VGND_c_663_n 0.0122414f $X=0.935 $Y=0.82 $X2=0 $Y2=0
cc_349 N_A_27_47#_c_582_n N_VGND_c_664_n 0.0122414f $X=1.775 $Y=0.78 $X2=0 $Y2=0
cc_350 N_A_27_47#_c_578_n N_VGND_c_665_n 0.0213324f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_351 N_A_27_47#_c_579_n N_VGND_c_665_n 0.00193763f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_579_n N_VGND_c_667_n 0.00193763f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_597_n N_VGND_c_667_n 0.0188551f $X=1.1 $Y=0.4 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_582_n N_VGND_c_667_n 0.00193763f $X=1.775 $Y=0.78 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_582_n N_VGND_c_669_n 0.00193763f $X=1.775 $Y=0.78 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_583_n N_VGND_c_669_n 0.00468912f $X=2.105 $Y=0.78 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_584_n N_VGND_c_669_n 0.00117399f $X=2.615 $Y=0.78 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_M1008_d N_VGND_c_670_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_M1010_d N_VGND_c_670_n 0.00215201f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_M1023_d N_VGND_c_670_n 0.00323135f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_M1015_s N_VGND_c_670_n 0.00216833f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_M1019_s N_VGND_c_670_n 0.00210147f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_578_n N_VGND_c_670_n 0.0126042f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_364 N_A_27_47#_c_579_n N_VGND_c_670_n 0.00825759f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_597_n N_VGND_c_670_n 0.0122069f $X=1.1 $Y=0.4 $X2=0 $Y2=0
cc_366 N_A_27_47#_c_582_n N_VGND_c_670_n 0.00825759f $X=1.775 $Y=0.78 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_583_n N_VGND_c_670_n 0.00902546f $X=2.105 $Y=0.78 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_584_n N_VGND_c_670_n 0.00282588f $X=2.615 $Y=0.78 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_584_n N_A_445_47#_M1011_d 0.00191689f $X=2.615 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_370 N_A_27_47#_c_587_n N_A_445_47#_M1018_d 0.00191689f $X=3.455 $Y=0.78 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_M1015_s N_A_445_47#_c_735_n 0.0030596f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_M1019_s N_A_445_47#_c_735_n 0.00511748f $X=3.485 $Y=0.235
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_584_n N_A_445_47#_c_735_n 0.0149721f $X=2.615 $Y=0.78 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_585_n N_A_445_47#_c_735_n 0.0153745f $X=2.945 $Y=0.78 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_586_n N_A_445_47#_c_735_n 0.0198093f $X=3.62 $Y=0.74 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_587_n N_A_445_47#_c_735_n 0.0191683f $X=3.455 $Y=0.78 $X2=0
+ $Y2=0
cc_377 N_VGND_c_670_n N_A_445_47#_M1011_d 0.00215227f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_378 N_VGND_c_670_n N_A_445_47#_M1018_d 0.00215227f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_670_n N_A_445_47#_M1006_s 0.00209344f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_670_n N_A_445_47#_M1009_s 0.00215227f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_c_670_n N_A_445_47#_M1016_s 0.00217543f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_669_n N_A_445_47#_c_735_n 0.219048f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_c_670_n N_A_445_47#_c_735_n 0.137165f $X=6.21 $Y=0 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nand4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 0.725000 3.640000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.780000 1.655000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.735000 1.720000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 1.075000 1.320000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.909000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.120000 1.495000 2.670000 1.665000 ;
        RECT 1.120000 1.665000 1.450000 2.465000 ;
        RECT 2.140000 1.665000 2.470000 2.465000 ;
        RECT 2.420000 0.255000 2.930000 0.825000 ;
        RECT 2.420000 0.825000 2.670000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.140000 0.085000 ;
        RECT 0.595000  0.085000 0.900000 0.545000 ;
        RECT 3.100000  0.085000 3.450000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.140000 2.805000 ;
        RECT 0.595000 1.835000 0.925000 2.635000 ;
        RECT 1.640000 1.835000 1.970000 2.635000 ;
        RECT 2.680000 2.175000 3.450000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.485000 0.425000 0.715000 ;
      RECT 0.085000 0.715000 1.270000 0.905000 ;
      RECT 0.085000 0.905000 0.260000 2.065000 ;
      RECT 0.085000 2.065000 0.425000 2.465000 ;
      RECT 1.080000 0.365000 2.250000 0.555000 ;
      RECT 1.080000 0.555000 1.270000 0.715000 ;
      RECT 1.970000 0.555000 2.250000 1.325000 ;
      RECT 2.840000 0.995000 3.090000 1.835000 ;
      RECT 2.840000 1.835000 4.055000 2.005000 ;
      RECT 3.620000 0.255000 4.055000 0.545000 ;
      RECT 3.635000 2.005000 4.055000 2.465000 ;
      RECT 3.810000 0.545000 4.055000 1.835000 ;
  END
END sky130_fd_sc_hd__nand4bb_1
END LIBRARY

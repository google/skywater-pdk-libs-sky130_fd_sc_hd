* File: sky130_fd_sc_hd__a41o_1.spice.SKY130_FD_SC_HD__A41O_1.pxi
* Created: Thu Aug 27 14:06:01 2020
* 
x_PM_SKY130_FD_SC_HD__A41O_1%A_79_21# N_A_79_21#_M1004_d N_A_79_21#_M1001_s
+ N_A_79_21#_M1011_g N_A_79_21#_M1007_g N_A_79_21#_c_65_n N_A_79_21#_c_66_n
+ N_A_79_21#_c_67_n N_A_79_21#_c_94_p N_A_79_21#_c_72_n N_A_79_21#_c_101_p
+ N_A_79_21#_c_73_n N_A_79_21#_c_76_p N_A_79_21#_c_68_n
+ PM_SKY130_FD_SC_HD__A41O_1%A_79_21#
x_PM_SKY130_FD_SC_HD__A41O_1%B1 N_B1_c_131_n N_B1_M1004_g N_B1_M1001_g B1 B1
+ N_B1_c_133_n PM_SKY130_FD_SC_HD__A41O_1%B1
x_PM_SKY130_FD_SC_HD__A41O_1%A1 N_A1_c_165_n N_A1_M1002_g N_A1_M1010_g A1
+ N_A1_c_167_n PM_SKY130_FD_SC_HD__A41O_1%A1
x_PM_SKY130_FD_SC_HD__A41O_1%A2 N_A2_M1005_g N_A2_M1008_g N_A2_c_199_n
+ N_A2_c_200_n A2 A2 N_A2_c_201_n N_A2_c_213_n PM_SKY130_FD_SC_HD__A41O_1%A2
x_PM_SKY130_FD_SC_HD__A41O_1%A3 N_A3_M1006_g N_A3_M1003_g A3 A3 A3 A3
+ N_A3_c_241_n N_A3_c_242_n A3 PM_SKY130_FD_SC_HD__A41O_1%A3
x_PM_SKY130_FD_SC_HD__A41O_1%A4 N_A4_c_277_n N_A4_M1009_g N_A4_M1000_g A4 A4
+ N_A4_c_279_n PM_SKY130_FD_SC_HD__A41O_1%A4
x_PM_SKY130_FD_SC_HD__A41O_1%X N_X_M1011_s N_X_M1007_s X X X X X X N_X_c_304_n X
+ X PM_SKY130_FD_SC_HD__A41O_1%X
x_PM_SKY130_FD_SC_HD__A41O_1%VPWR N_VPWR_M1007_d N_VPWR_M1010_d N_VPWR_M1003_d
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n VPWR N_VPWR_c_323_n
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_319_n N_VPWR_c_328_n
+ N_VPWR_c_329_n N_VPWR_c_330_n PM_SKY130_FD_SC_HD__A41O_1%VPWR
x_PM_SKY130_FD_SC_HD__A41O_1%A_297_297# N_A_297_297#_M1001_d
+ N_A_297_297#_M1008_d N_A_297_297#_M1000_d N_A_297_297#_c_386_n
+ N_A_297_297#_c_394_n N_A_297_297#_c_389_n N_A_297_297#_c_392_n
+ N_A_297_297#_c_399_n PM_SKY130_FD_SC_HD__A41O_1%A_297_297#
x_PM_SKY130_FD_SC_HD__A41O_1%VGND N_VGND_M1011_d N_VGND_M1009_d N_VGND_c_420_n
+ N_VGND_c_421_n N_VGND_c_422_n VGND N_VGND_c_423_n N_VGND_c_424_n
+ N_VGND_c_425_n N_VGND_c_426_n PM_SKY130_FD_SC_HD__A41O_1%VGND
cc_1 VNB N_A_79_21#_c_65_n 9.98293e-19 $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_2 VNB N_A_79_21#_c_66_n 0.0297635f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_3 VNB N_A_79_21#_c_67_n 0.0111928f $X=-0.19 $Y=-0.24 $X2=1.115 $Y2=0.82
cc_4 VNB N_A_79_21#_c_68_n 0.0204737f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=0.995
cc_5 VNB N_B1_c_131_n 0.0201268f $X=-0.19 $Y=-0.24 $X2=1.19 $Y2=0.235
cc_6 VNB B1 0.00209895f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_7 VNB N_B1_c_133_n 0.0323034f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_8 VNB N_A1_c_165_n 0.0186918f $X=-0.19 $Y=-0.24 $X2=1.19 $Y2=0.235
cc_9 VNB A1 0.00972855f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A1_c_167_n 0.0205835f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_11 VNB N_A2_c_199_n 9.449e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_12 VNB N_A2_c_200_n 0.0225369f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_13 VNB N_A2_c_201_n 0.0163858f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_14 VNB A3 0.00188705f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB A3 0.00425273f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_16 VNB N_A3_c_241_n 0.0205482f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_17 VNB N_A3_c_242_n 0.0174945f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.82
cc_18 VNB A3 7.68134e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A4_c_277_n 0.0218222f $X=-0.19 $Y=-0.24 $X2=1.19 $Y2=0.235
cc_20 VNB A4 0.00243804f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_A4_c_279_n 0.0440674f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.825
cc_22 VNB X 0.0338278f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_23 VNB N_X_c_304_n 0.0105828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_319_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_420_n 0.00559666f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_26 VNB N_VGND_c_421_n 0.0102094f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_27 VNB N_VGND_c_422_n 0.0262961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_423_n 0.0178772f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_29 VNB N_VGND_c_424_n 0.0608045f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.91
cc_30 VNB N_VGND_c_425_n 0.00632006f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.16
cc_31 VNB N_VGND_c_426_n 0.199093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_79_21#_M1007_g 0.0263894f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_33 VPB N_A_79_21#_c_65_n 0.00153334f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_34 VPB N_A_79_21#_c_66_n 0.0070917f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_35 VPB N_A_79_21#_c_72_n 0.0121808f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.91
cc_36 VPB N_A_79_21#_c_73_n 0.00523849f $X=-0.19 $Y=1.305 $X2=1.2 $Y2=2
cc_37 VPB N_B1_M1001_g 0.022117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB B1 0.00488162f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_39 VPB N_B1_c_133_n 0.0101114f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_40 VPB N_A1_M1010_g 0.0182177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB A1 0.00124009f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_42 VPB N_A1_c_167_n 0.0046065f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_43 VPB N_A2_M1008_g 0.0197833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A2_c_199_n 0.00172012f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_45 VPB N_A2_c_200_n 0.00463657f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_46 VPB N_A3_M1003_g 0.0195405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A3_c_241_n 0.00453751f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_48 VPB A3 0.00115543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A4_M1000_g 0.0227754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB A4 0.012924f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_51 VPB N_A4_c_279_n 0.0107861f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.825
cc_52 VPB X 0.0350296f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_53 VPB X 0.0105794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_320_n 0.00862158f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_55 VPB N_VPWR_c_321_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_56 VPB N_VPWR_c_322_n 0.0051673f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.82
cc_57 VPB N_VPWR_c_323_n 0.0178428f $X=-0.19 $Y=1.305 $X2=1.2 $Y2=2
cc_58 VPB N_VPWR_c_324_n 0.0280808f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=0.385
cc_59 VPB N_VPWR_c_325_n 0.018193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_326_n 0.0183302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_319_n 0.0479428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_328_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_329_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_330_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_65_n N_B1_c_131_n 0.00161465f $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_79_21#_c_67_n N_B1_c_131_n 0.00949491f $X=1.115 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_67 N_A_79_21#_c_76_p N_B1_c_131_n 0.00887628f $X=1.365 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_68 N_A_79_21#_c_68_n N_B1_c_131_n 0.0167276f $X=0.565 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_69 N_A_79_21#_c_65_n N_B1_M1001_g 0.00426467f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_72_n N_B1_M1001_g 0.00320272f $X=1.035 $Y=1.91 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_73_n N_B1_M1001_g 0.00476434f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_72 N_A_79_21#_M1001_s B1 0.00380279f $X=1.075 $Y=1.485 $X2=0 $Y2=0
cc_73 N_A_79_21#_M1007_g B1 0.00159773f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_65_n B1 0.0274523f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_66_n B1 0.00181932f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_67_n B1 0.0271342f $X=1.115 $Y=0.82 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_72_n B1 0.0220166f $X=1.035 $Y=1.91 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_65_n N_B1_c_133_n 7.94331e-19 $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_66_n N_B1_c_133_n 0.0139293f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_67_n N_B1_c_133_n 0.0107163f $X=1.115 $Y=0.82 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_72_n N_B1_c_133_n 0.00110259f $X=1.035 $Y=1.91 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_67_n N_A1_c_165_n 0.00425738f $X=1.115 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_79_21#_c_76_p N_A1_c_165_n 0.00712121f $X=1.365 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_79_21#_c_65_n X 0.054279f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_94_p X 0.00792678f $X=0.685 $Y=0.82 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_68_n X 0.0146741f $X=0.565 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_68_n N_X_c_304_n 0.00439012f $X=0.565 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_79_21#_M1007_g X 0.00455601f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_73_n X 3.01625e-19 $X=1.2 $Y=2 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_65_n N_VPWR_M1007_d 0.00524561f $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_79_21#_c_72_n N_VPWR_M1007_d 0.0054329f $X=1.035 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_79_21#_c_101_p N_VPWR_M1007_d 9.06359e-19 $X=0.685 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_79_21#_M1007_g N_VPWR_c_320_n 0.0044954f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_72_n N_VPWR_c_320_n 0.0119307f $X=1.035 $Y=1.91 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_101_p N_VPWR_c_320_n 0.00678689f $X=0.685 $Y=1.91 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_73_n N_VPWR_c_320_n 0.0188543f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_97 N_A_79_21#_M1007_g N_VPWR_c_323_n 0.00513419f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_101_p N_VPWR_c_323_n 8.16647e-19 $X=0.685 $Y=1.91 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_72_n N_VPWR_c_324_n 0.00288053f $X=1.035 $Y=1.91 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_73_n N_VPWR_c_324_n 0.0166218f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_101 N_A_79_21#_M1001_s N_VPWR_c_319_n 0.00211564f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_M1007_g N_VPWR_c_319_n 0.0108728f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_72_n N_VPWR_c_319_n 0.00567086f $X=1.035 $Y=1.91 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_101_p N_VPWR_c_319_n 0.00244861f $X=0.685 $Y=1.91 $X2=0
+ $Y2=0
cc_105 N_A_79_21#_c_73_n N_VPWR_c_319_n 0.0121298f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_67_n N_VGND_M1011_d 0.00418635f $X=1.115 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_79_21#_c_94_p N_VGND_M1011_d 8.97268e-19 $X=0.685 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_79_21#_c_66_n N_VGND_c_420_n 4.85811e-19 $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_67_n N_VGND_c_420_n 0.0187205f $X=1.115 $Y=0.82 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_94_p N_VGND_c_420_n 0.00719606f $X=0.685 $Y=0.82 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_76_p N_VGND_c_420_n 0.0192053f $X=1.365 $Y=0.385 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_68_n N_VGND_c_420_n 0.0054486f $X=0.565 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_94_p N_VGND_c_423_n 8.04923e-19 $X=0.685 $Y=0.82 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_68_n N_VGND_c_423_n 0.00513885f $X=0.565 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_A_79_21#_c_67_n N_VGND_c_424_n 0.00222393f $X=1.115 $Y=0.82 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_76_p N_VGND_c_424_n 0.0205472f $X=1.365 $Y=0.385 $X2=0 $Y2=0
cc_117 N_A_79_21#_M1004_d N_VGND_c_426_n 0.010584f $X=1.19 $Y=0.235 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_67_n N_VGND_c_426_n 0.00553482f $X=1.115 $Y=0.82 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_94_p N_VGND_c_426_n 0.00246127f $X=0.685 $Y=0.82 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_76_p N_VGND_c_426_n 0.0150402f $X=1.365 $Y=0.385 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_68_n N_VGND_c_426_n 0.0100991f $X=0.565 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B1_c_131_n N_A1_c_165_n 0.010303f $X=1.115 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_123 N_B1_M1001_g N_A1_M1010_g 0.0266823f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_124 B1 A1 0.0295499f $X=1.09 $Y=1.105 $X2=0 $Y2=0
cc_125 N_B1_c_133_n A1 0.00608409f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B1_c_133_n N_A1_c_167_n 0.0208073f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B1_M1001_g N_VPWR_c_320_n 0.00283988f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_128 N_B1_M1001_g N_VPWR_c_324_n 0.00542953f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_129 N_B1_M1001_g N_VPWR_c_319_n 0.0109803f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_130 N_B1_c_131_n N_VGND_c_420_n 0.00696921f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_c_131_n N_VGND_c_424_n 0.00404518f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_c_131_n N_VGND_c_426_n 0.00674866f $X=1.115 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A1_M1010_g N_A2_M1008_g 0.0456295f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_134 A1 N_A2_M1008_g 0.00160758f $X=1.55 $Y=1.445 $X2=0 $Y2=0
cc_135 N_A1_c_165_n N_A2_c_199_n 0.00224964f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_136 A1 N_A2_c_199_n 0.0150642f $X=1.55 $Y=1.445 $X2=0 $Y2=0
cc_137 N_A1_c_167_n N_A2_c_199_n 0.00106653f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_138 A1 N_A2_c_200_n 0.00106544f $X=1.55 $Y=1.445 $X2=0 $Y2=0
cc_139 N_A1_c_167_n N_A2_c_200_n 0.0198587f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A1_c_165_n N_A2_c_201_n 0.0423649f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A1_c_165_n N_A2_c_213_n 0.0120277f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_142 A1 N_A2_c_213_n 0.00698426f $X=1.55 $Y=1.445 $X2=0 $Y2=0
cc_143 N_A1_c_167_n N_A2_c_213_n 8.38682e-19 $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A1_M1010_g N_VPWR_c_321_n 0.00302074f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1010_g N_VPWR_c_324_n 0.00441875f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1010_g N_VPWR_c_319_n 0.00591459f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_147 A1 N_A_297_297#_M1001_d 0.00195309f $X=1.55 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_148 N_A1_M1010_g N_A_297_297#_c_386_n 0.010913f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_149 A1 N_A_297_297#_c_386_n 0.00823625f $X=1.55 $Y=1.445 $X2=0 $Y2=0
cc_150 N_A1_c_167_n N_A_297_297#_c_386_n 7.75645e-19 $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_151 A1 N_A_297_297#_c_389_n 0.0136607f $X=1.55 $Y=1.445 $X2=0 $Y2=0
cc_152 N_A1_c_165_n N_VGND_c_424_n 0.00389067f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_165_n N_VGND_c_426_n 0.00605686f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A2_M1008_g N_A3_M1003_g 0.0229064f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A2_c_199_n A3 0.0151147f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A2_c_199_n A3 0.0172698f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_200_n A3 0.00102703f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A2_c_199_n N_A3_c_241_n 0.0011547f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_c_200_n N_A3_c_241_n 0.0196859f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A2_c_199_n N_A3_c_242_n 0.00337011f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A2_c_201_n N_A3_c_242_n 0.0320378f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_M1008_g A3 0.00163369f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_M1008_g N_VPWR_c_321_n 0.00302074f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A2_M1008_g N_VPWR_c_325_n 0.00441875f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A2_M1008_g N_VPWR_c_319_n 0.00605519f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A2_M1008_g N_A_297_297#_c_386_n 0.0127439f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A2_c_199_n N_A_297_297#_c_386_n 0.00419677f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A2_c_199_n N_A_297_297#_c_392_n 0.002579f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A2_c_200_n N_A_297_297#_c_392_n 4.339e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A2_c_201_n N_VGND_c_424_n 0.00389067f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A2_c_213_n N_VGND_c_424_n 0.0257279f $X=2.225 $Y=0.507 $X2=0 $Y2=0
cc_172 N_A2_c_201_n N_VGND_c_426_n 0.00561644f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A2_c_213_n N_VGND_c_426_n 0.0304095f $X=2.225 $Y=0.507 $X2=0 $Y2=0
cc_174 N_A2_c_213_n A_381_47# 0.00789698f $X=2.225 $Y=0.507 $X2=-0.19 $Y2=-0.24
cc_175 N_A2_c_199_n A_465_47# 0.00379633f $X=2.31 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_176 A2 A_465_47# 0.00980836f $X=2.47 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_177 A3 N_A4_c_277_n 0.00339611f $X=2.9 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_178 N_A3_c_242_n N_A4_c_277_n 0.0281211f $X=2.79 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_179 N_A3_M1003_g N_A4_M1000_g 0.0349354f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_180 A3 N_A4_M1000_g 0.00339611f $X=2.985 $Y=1.19 $X2=0 $Y2=0
cc_181 A3 A4 0.0312766f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A3_c_241_n A4 2.49049e-19 $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_183 A3 N_A4_c_279_n 0.00339611f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A3_c_241_n N_A4_c_279_n 0.0207732f $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_185 A3 N_VPWR_M1003_d 0.00296711f $X=2.985 $Y=1.19 $X2=0 $Y2=0
cc_186 N_A3_M1003_g N_VPWR_c_322_n 0.00294145f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A3_M1003_g N_VPWR_c_325_n 0.00441875f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A3_M1003_g N_VPWR_c_319_n 0.00627106f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A3_M1003_g N_A_297_297#_c_394_n 0.0120453f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A3_c_241_n N_A_297_297#_c_394_n 3.67145e-19 $X=2.79 $Y=1.16 $X2=0 $Y2=0
cc_191 A3 N_A_297_297#_c_394_n 0.0250575f $X=2.985 $Y=1.19 $X2=0 $Y2=0
cc_192 N_A3_c_242_n N_VGND_c_422_n 0.00183532f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_193 A3 N_VGND_c_424_n 0.00734712f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_194 N_A3_c_242_n N_VGND_c_424_n 0.00585385f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_195 A3 N_VGND_c_426_n 0.00722417f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_196 N_A3_c_242_n N_VGND_c_426_n 0.0111601f $X=2.79 $Y=0.995 $X2=0 $Y2=0
cc_197 A3 A_561_47# 0.0124505f $X=2.9 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_198 N_A4_M1000_g N_VPWR_c_322_n 0.00294145f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A4_M1000_g N_VPWR_c_326_n 0.00441875f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A4_M1000_g N_VPWR_c_319_n 0.00705747f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_201 A4 N_A_297_297#_M1000_d 0.00487515f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A4_M1000_g N_A_297_297#_c_394_n 0.015073f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_203 A4 N_A_297_297#_c_399_n 0.0145976f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_204 N_A4_c_279_n N_A_297_297#_c_399_n 6.87511e-19 $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A4_c_277_n N_VGND_c_422_n 0.0149367f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_206 A4 N_VGND_c_422_n 0.0195285f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_207 N_A4_c_279_n N_VGND_c_422_n 0.00216025f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A4_c_277_n N_VGND_c_424_n 0.0046653f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A4_c_277_n N_VGND_c_426_n 0.00814192f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_210 X N_VPWR_c_323_n 0.0172332f $X=0.235 $Y=2.21 $X2=0 $Y2=0
cc_211 N_X_M1007_s N_VPWR_c_319_n 0.00211564f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_212 X N_VPWR_c_319_n 0.0124665f $X=0.235 $Y=2.21 $X2=0 $Y2=0
cc_213 N_X_c_304_n N_VGND_c_423_n 0.0168043f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_214 N_X_M1011_s N_VGND_c_426_n 0.00212021f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_215 N_X_c_304_n N_VGND_c_426_n 0.0124421f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_216 N_VPWR_c_319_n N_A_297_297#_M1001_d 0.00414531f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_217 N_VPWR_c_319_n N_A_297_297#_M1008_d 0.003474f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_c_319_n N_A_297_297#_M1000_d 0.00377405f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_219 N_VPWR_M1010_d N_A_297_297#_c_386_n 0.00761236f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_321_n N_A_297_297#_c_386_n 0.0102407f $X=2.04 $Y=2.34 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_324_n N_A_297_297#_c_386_n 0.0023033f $X=1.915 $Y=2.72 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_325_n N_A_297_297#_c_386_n 0.0023033f $X=2.845 $Y=2.72 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_319_n N_A_297_297#_c_386_n 0.010153f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_M1003_d N_A_297_297#_c_394_n 0.00467301f $X=2.805 $Y=1.485 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_322_n N_A_297_297#_c_394_n 0.0141794f $X=2.97 $Y=2.34 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_325_n N_A_297_297#_c_394_n 0.00328576f $X=2.845 $Y=2.72 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_326_n N_A_297_297#_c_394_n 0.00251892f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_319_n N_A_297_297#_c_394_n 0.0132513f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_324_n N_A_297_297#_c_389_n 0.0113839f $X=1.915 $Y=2.72 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_319_n N_A_297_297#_c_389_n 0.00646745f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_325_n N_A_297_297#_c_392_n 0.0115924f $X=2.845 $Y=2.72 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_319_n N_A_297_297#_c_392_n 0.00646745f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_326_n N_A_297_297#_c_399_n 0.0115924f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_319_n N_A_297_297#_c_399_n 0.00646745f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_235 N_VGND_c_426_n A_381_47# 0.00240861f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_236 N_VGND_c_426_n A_465_47# 0.00311298f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_237 N_VGND_c_426_n A_561_47# 0.00720093f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a2bb2o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 0.995000 1.675000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 0.995000 2.135000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.730000 0.765000 3.990000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.355000 3.530000 1.655000 ;
        RECT 3.270000 0.765000 3.530000 1.355000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.780000 0.810000 ;
        RECT 0.525000 0.810000 0.695000 1.525000 ;
        RECT 0.525000 1.525000 0.780000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.140000 0.085000 ;
        RECT 0.185000  0.085000 0.355000 0.930000 ;
        RECT 0.950000  0.085000 1.380000 0.530000 ;
        RECT 1.955000  0.085000 2.690000 0.485000 ;
        RECT 3.605000  0.085000 4.005000 0.595000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.140000 2.805000 ;
        RECT 0.185000 1.445000 0.355000 2.635000 ;
        RECT 0.950000 2.235000 1.280000 2.635000 ;
        RECT 3.375000 2.175000 3.625000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.865000 0.995000 1.120000 1.325000 ;
      RECT 0.950000 1.325000 1.120000 1.805000 ;
      RECT 0.950000 1.805000 1.710000 1.975000 ;
      RECT 1.540000 1.975000 1.710000 2.200000 ;
      RECT 1.540000 2.200000 2.670000 2.370000 ;
      RECT 1.615000 0.255000 1.785000 0.655000 ;
      RECT 1.615000 0.655000 2.510000 0.825000 ;
      RECT 1.975000 1.545000 2.510000 1.715000 ;
      RECT 1.975000 1.715000 2.145000 1.905000 ;
      RECT 2.340000 0.825000 2.510000 1.545000 ;
      RECT 2.440000 1.895000 2.850000 2.065000 ;
      RECT 2.440000 2.065000 2.670000 2.200000 ;
      RECT 2.500000 2.370000 2.670000 2.465000 ;
      RECT 2.680000 0.700000 3.030000 0.870000 ;
      RECT 2.680000 0.870000 2.850000 1.895000 ;
      RECT 2.860000 0.255000 3.030000 0.700000 ;
      RECT 2.875000 2.255000 3.205000 2.425000 ;
      RECT 3.035000 1.835000 3.965000 2.005000 ;
      RECT 3.035000 2.005000 3.205000 2.255000 ;
      RECT 3.795000 2.005000 3.965000 2.465000 ;
  END
END sky130_fd_sc_hd__a2bb2o_2

* File: sky130_fd_sc_hd__and3b_1.pex.spice
* Created: Thu Aug 27 14:07:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND3B_1%A_N 2 5 8 10 11 12 13 18 20
c25 11 0 1.17844e-19 $X=0.23 $Y=1.19
r26 18 20 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.327 $Y=1.16
+ $X2=0.327 $Y2=0.995
r27 12 13 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.255 $Y=1.53
+ $X2=0.255 $Y2=1.87
r28 11 12 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r29 11 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r30 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.695
r31 5 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
r32 2 10 53.1843 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.327 $Y=1.478
+ $X2=0.327 $Y2=1.695
r33 1 18 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=0.327 $Y=1.212
+ $X2=0.327 $Y2=1.16
r34 1 2 34.0085 $w=4.35e-07 $l=2.66e-07 $layer=POLY_cond $X=0.327 $Y=1.212
+ $X2=0.327 $Y2=1.478
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_1%A_109_93# 1 2 9 13 15 17 21 30
c43 30 0 1.17844e-19 $X=1.405 $Y=1.16
c44 21 0 2.08126e-19 $X=1.195 $Y=1.16
r45 29 30 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.38 $Y=1.16
+ $X2=1.405 $Y2=1.16
r46 25 26 15.7687 $w=2.94e-07 $l=3.8e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=0.68 $Y2=1.12
r47 22 29 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.195 $Y=1.16
+ $X2=1.38 $Y2=1.16
r48 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.16 $X2=1.195 $Y2=1.16
r49 19 26 1.68758 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.12
+ $X2=0.68 $Y2=1.12
r50 19 21 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=0.845 $Y=1.12
+ $X2=1.195 $Y2=1.12
r51 15 26 7.33909 $w=2.94e-07 $l=1.25e-07 $layer=LI1_cond $X=0.68 $Y=1.245
+ $X2=0.68 $Y2=1.12
r52 15 17 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=0.68 $Y=1.245
+ $X2=0.68 $Y2=2.26
r53 11 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=0.995
+ $X2=1.405 $Y2=1.16
r54 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.405 $Y=0.995
+ $X2=1.405 $Y2=0.475
r55 7 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.325
+ $X2=1.38 $Y2=1.16
r56 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.38 $Y=1.325 $X2=1.38
+ $Y2=1.765
r57 2 17 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.26
r58 1 25 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.68 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_1%B 3 8 10 11 14
c38 8 0 3.59332e-20 $X=1.8 $Y=1.765
c39 3 0 1.72192e-19 $X=1.765 $Y=0.475
r40 14 16 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.867 $Y=2.3
+ $X2=1.867 $Y2=2.135
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.875
+ $Y=2.3 $X2=1.875 $Y2=2.3
r42 11 15 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=2.07 $Y=2.295
+ $X2=1.875 $Y2=2.295
r43 9 10 68.3433 $w=1.85e-07 $l=1.85e-07 $layer=POLY_cond $X=1.782 $Y=1.015
+ $X2=1.782 $Y2=1.2
r44 8 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.8 $Y=1.765 $X2=1.8
+ $Y2=2.135
r45 8 10 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.8 $Y=1.765 $X2=1.8
+ $Y2=1.2
r46 3 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.765 $Y=0.475
+ $X2=1.765 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_1%C 3 7 9 10 14
r47 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=1.325
r48 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.16
+ $X2=2.23 $Y2=0.995
r49 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.16 $X2=2.23 $Y2=1.16
r50 10 15 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=2.19 $Y=0.85
+ $X2=2.19 $Y2=1.16
r51 10 22 6.54281 $w=4.08e-07 $l=1.25e-07 $layer=LI1_cond $X=2.19 $Y=0.85
+ $X2=2.19 $Y2=0.725
r52 9 22 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=2.085 $Y=0.51
+ $X2=2.085 $Y2=0.725
r53 7 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.275 $Y=1.695
+ $X2=2.275 $Y2=1.325
r54 3 16 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.17 $Y=0.475
+ $X2=2.17 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_1%A_209_311# 1 2 3 12 15 19 21 25 26 28 29 30
+ 33 34 40
r86 36 38 16.5476 $w=2.75e-07 $l=3.73e-07 $layer=LI1_cond $X=1.687 $Y=1.595
+ $X2=2.06 $Y2=1.595
r87 34 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.71 $Y2=1.325
r88 34 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.71 $Y2=0.995
r89 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.16 $X2=2.71 $Y2=1.16
r90 31 33 13.2781 $w=2.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.68 $Y=1.425
+ $X2=2.68 $Y2=1.16
r91 30 38 5.87701 $w=4.65e-07 $l=1.7528e-07 $layer=LI1_cond $X=2.207 $Y=1.657
+ $X2=2.06 $Y2=1.595
r92 29 31 5.48862 $w=4.99e-07 $l=2.83732e-07 $layer=LI1_cond $X=2.565 $Y=1.657
+ $X2=2.68 $Y2=1.425
r93 29 30 9.20852 $w=4.63e-07 $l=3.58e-07 $layer=LI1_cond $X=2.565 $Y=1.657
+ $X2=2.207 $Y2=1.657
r94 28 36 1.19494 $w=2.55e-07 $l=1.7e-07 $layer=LI1_cond $X=1.687 $Y=1.425
+ $X2=1.687 $Y2=1.595
r95 27 28 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=1.687 $Y=0.57
+ $X2=1.687 $Y2=1.425
r96 25 36 7.40164 $w=2.75e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.56 $Y=1.51
+ $X2=1.687 $Y2=1.595
r97 25 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.56 $Y=1.51
+ $X2=1.255 $Y2=1.51
r98 21 27 6.81977 $w=2.65e-07 $l=1.85957e-07 $layer=LI1_cond $X=1.56 $Y=0.437
+ $X2=1.687 $Y2=0.57
r99 21 23 15.8733 $w=2.63e-07 $l=3.65e-07 $layer=LI1_cond $X=1.56 $Y=0.437
+ $X2=1.195 $Y2=0.437
r100 17 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.13 $Y=1.595
+ $X2=1.255 $Y2=1.51
r101 17 19 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.13 $Y=1.595
+ $X2=1.13 $Y2=1.76
r102 15 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.75 $Y=1.985
+ $X2=2.75 $Y2=1.325
r103 12 40 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.56
+ $X2=2.75 $Y2=0.995
r104 3 38 600 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_PDIFF $count=1 $X=1.875
+ $Y=1.555 $X2=2.06 $Y2=1.725
r105 2 19 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.555 $X2=1.17 $Y2=1.76
r106 1 23 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.265 $X2=1.195 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_1%VPWR 1 2 3 10 12 18 23 25 27 32 39 40 46 51
r53 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 40 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 37 51 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=2.65 $Y=2.72
+ $X2=2.542 $Y2=2.72
r57 37 39 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.65 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 36 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 36 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 33 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.62 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 32 51 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.542 $Y2=2.72
r63 32 35 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.07 $Y2=2.72
r64 31 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 28 43 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r67 28 30 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 27 33 8.47627 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=1.312 $Y=2.72
+ $X2=1.62 $Y2=2.72
r69 27 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 27 46 17.5371 $w=6.13e-07 $l=5.9e-07 $layer=LI1_cond $X=1.312 $Y=2.72
+ $X2=1.312 $Y2=2.13
r71 27 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 25 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 20 23 3.96938 $w=1.88e-07 $l=6.8e-08 $layer=LI1_cond $X=1.522 $Y=1.86
+ $X2=1.59 $Y2=1.86
r75 16 51 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.542 $Y=2.635
+ $X2=2.542 $Y2=2.72
r76 16 18 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=2.542 $Y=2.635
+ $X2=2.542 $Y2=2.34
r77 14 20 0.589566 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=1.522 $Y=1.955
+ $X2=1.522 $Y2=1.86
r78 14 46 9.95338 $w=1.93e-07 $l=1.75e-07 $layer=LI1_cond $X=1.522 $Y=1.955
+ $X2=1.522 $Y2=2.13
r79 10 43 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r80 10 12 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.29
r81 3 18 600 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.485 $X2=2.54 $Y2=2.34
r82 2 23 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=1.455
+ $Y=1.555 $X2=1.59 $Y2=1.85
r83 1 12 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_1%X 1 2 9 10 12 13 14 22
r18 14 22 11.734 $w=2.73e-07 $l=2.8e-07 $layer=LI1_cond $X=2.997 $Y=2.21
+ $X2=2.997 $Y2=1.93
r19 11 13 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=3.005 $Y=0.605
+ $X2=3.005 $Y2=0.51
r20 11 12 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.005 $Y=0.605
+ $X2=3.005 $Y2=0.735
r21 10 12 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.05 $Y=1.765
+ $X2=3.05 $Y2=0.735
r22 9 22 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=2.997 $Y=1.902
+ $X2=2.997 $Y2=1.93
r23 9 10 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.997 $Y=1.902
+ $X2=2.997 $Y2=1.765
r24 2 22 300 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_PDIFF $count=2 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.93
r25 1 13 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__AND3B_1%VGND 1 2 7 9 13 15 17 27 28 34
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r39 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r40 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r41 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.54
+ $Y2=0
r42 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.99
+ $Y2=0
r43 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r44 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r45 21 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r46 20 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r47 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 18 31 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r49 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r50 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.54
+ $Y2=0
r51 17 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.07
+ $Y2=0
r52 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r53 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r54 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0
r55 11 13 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0.46
r56 7 31 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r57 7 9 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.73
r58 2 13 182 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.265 $X2=2.54 $Y2=0.46
r59 1 9 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.73
.ends


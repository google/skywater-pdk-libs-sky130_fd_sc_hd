* File: sky130_fd_sc_hd__dfrbp_1.spice.SKY130_FD_SC_HD__DFRBP_1.pxi
* Created: Thu Aug 27 14:14:19 2020
* 
x_PM_SKY130_FD_SC_HD__DFRBP_1%CLK N_CLK_c_217_n N_CLK_c_221_n N_CLK_c_218_n
+ N_CLK_M1027_g N_CLK_c_222_n N_CLK_M1014_g N_CLK_c_223_n CLK CLK
+ PM_SKY130_FD_SC_HD__DFRBP_1%CLK
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_27_47# N_A_27_47#_M1027_s N_A_27_47#_M1014_s
+ N_A_27_47#_M1015_g N_A_27_47#_M1000_g N_A_27_47#_M1009_g N_A_27_47#_c_259_n
+ N_A_27_47#_c_260_n N_A_27_47#_c_261_n N_A_27_47#_M1007_g N_A_27_47#_c_262_n
+ N_A_27_47#_M1025_g N_A_27_47#_M1021_g N_A_27_47#_c_264_n N_A_27_47#_c_265_n
+ N_A_27_47#_c_266_n N_A_27_47#_c_283_n N_A_27_47#_c_284_n N_A_27_47#_c_267_n
+ N_A_27_47#_c_268_n N_A_27_47#_c_269_n N_A_27_47#_c_270_n N_A_27_47#_c_271_n
+ N_A_27_47#_c_272_n N_A_27_47#_c_273_n N_A_27_47#_c_274_n N_A_27_47#_c_275_n
+ N_A_27_47#_c_276_n PM_SKY130_FD_SC_HD__DFRBP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DFRBP_1%D N_D_M1029_g N_D_M1028_g N_D_c_494_n N_D_c_498_n
+ D N_D_c_495_n PM_SKY130_FD_SC_HD__DFRBP_1%D
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_193_47# N_A_193_47#_M1015_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1030_g N_A_193_47#_M1020_g N_A_193_47#_c_547_n
+ N_A_193_47#_M1023_g N_A_193_47#_M1012_g N_A_193_47#_c_548_n
+ N_A_193_47#_c_549_n N_A_193_47#_c_550_n N_A_193_47#_c_558_n
+ N_A_193_47#_c_559_n N_A_193_47#_c_551_n N_A_193_47#_c_552_n
+ N_A_193_47#_c_560_n N_A_193_47#_c_561_n N_A_193_47#_c_562_n
+ N_A_193_47#_c_563_n N_A_193_47#_c_564_n N_A_193_47#_c_565_n
+ N_A_193_47#_c_566_n N_A_193_47#_c_567_n N_A_193_47#_c_568_n
+ N_A_193_47#_c_553_n PM_SKY130_FD_SC_HD__DFRBP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_761_289# N_A_761_289#_M1022_d
+ N_A_761_289#_M1017_d N_A_761_289#_M1010_g N_A_761_289#_M1003_g
+ N_A_761_289#_c_762_n N_A_761_289#_c_763_n N_A_761_289#_c_784_n
+ N_A_761_289#_c_759_n N_A_761_289#_c_786_n N_A_761_289#_c_771_n
+ N_A_761_289#_c_791_n N_A_761_289#_c_773_n N_A_761_289#_c_809_p
+ N_A_761_289#_c_774_n N_A_761_289#_c_775_n
+ PM_SKY130_FD_SC_HD__DFRBP_1%A_761_289#
x_PM_SKY130_FD_SC_HD__DFRBP_1%RESET_B N_RESET_B_M1004_g N_RESET_B_M1031_g
+ N_RESET_B_M1005_g N_RESET_B_M1018_g RESET_B RESET_B N_RESET_B_c_871_n
+ N_RESET_B_c_872_n N_RESET_B_c_873_n N_RESET_B_c_874_n N_RESET_B_c_875_n
+ N_RESET_B_c_876_n N_RESET_B_c_877_n N_RESET_B_c_878_n N_RESET_B_c_879_n
+ N_RESET_B_c_880_n PM_SKY130_FD_SC_HD__DFRBP_1%RESET_B
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_543_47# N_A_543_47#_M1009_d N_A_543_47#_M1030_d
+ N_A_543_47#_M1022_g N_A_543_47#_c_1028_n N_A_543_47#_c_1029_n
+ N_A_543_47#_M1017_g N_A_543_47#_c_1037_n N_A_543_47#_c_1058_n
+ N_A_543_47#_c_1030_n N_A_543_47#_c_1023_n N_A_543_47#_c_1024_n
+ N_A_543_47#_c_1025_n N_A_543_47#_c_1026_n N_A_543_47#_c_1027_n
+ PM_SKY130_FD_SC_HD__DFRBP_1%A_543_47#
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_1283_21# N_A_1283_21#_M1001_d
+ N_A_1283_21#_M1018_d N_A_1283_21#_M1026_g N_A_1283_21#_M1008_g
+ N_A_1283_21#_M1011_g N_A_1283_21#_c_1150_n N_A_1283_21#_M1019_g
+ N_A_1283_21#_c_1151_n N_A_1283_21#_c_1152_n N_A_1283_21#_c_1153_n
+ N_A_1283_21#_c_1154_n N_A_1283_21#_M1006_g N_A_1283_21#_M1024_g
+ N_A_1283_21#_c_1155_n N_A_1283_21#_c_1170_n N_A_1283_21#_c_1171_n
+ N_A_1283_21#_c_1156_n N_A_1283_21#_c_1157_n N_A_1283_21#_c_1200_n
+ N_A_1283_21#_c_1205_n N_A_1283_21#_c_1284_p N_A_1283_21#_c_1172_n
+ N_A_1283_21#_c_1173_n N_A_1283_21#_c_1158_n N_A_1283_21#_c_1159_n
+ N_A_1283_21#_c_1174_n N_A_1283_21#_c_1160_n N_A_1283_21#_c_1161_n
+ N_A_1283_21#_c_1162_n PM_SKY130_FD_SC_HD__DFRBP_1%A_1283_21#
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_1108_47# N_A_1108_47#_M1023_d
+ N_A_1108_47#_M1025_d N_A_1108_47#_M1016_g N_A_1108_47#_M1001_g
+ N_A_1108_47#_c_1346_n N_A_1108_47#_c_1349_n N_A_1108_47#_c_1339_n
+ N_A_1108_47#_c_1342_n N_A_1108_47#_c_1343_n N_A_1108_47#_c_1344_n
+ N_A_1108_47#_c_1345_n PM_SKY130_FD_SC_HD__DFRBP_1%A_1108_47#
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_1847_47# N_A_1847_47#_M1006_s
+ N_A_1847_47#_M1024_s N_A_1847_47#_M1002_g N_A_1847_47#_M1013_g
+ N_A_1847_47#_c_1444_n N_A_1847_47#_c_1449_n N_A_1847_47#_c_1445_n
+ N_A_1847_47#_c_1446_n N_A_1847_47#_c_1463_n N_A_1847_47#_c_1447_n
+ PM_SKY130_FD_SC_HD__DFRBP_1%A_1847_47#
x_PM_SKY130_FD_SC_HD__DFRBP_1%VPWR N_VPWR_M1014_d N_VPWR_M1028_s N_VPWR_M1010_d
+ N_VPWR_M1017_s N_VPWR_M1008_d N_VPWR_M1016_d N_VPWR_M1024_d N_VPWR_c_1493_n
+ N_VPWR_c_1494_n N_VPWR_c_1495_n N_VPWR_c_1496_n N_VPWR_c_1497_n
+ N_VPWR_c_1498_n N_VPWR_c_1499_n N_VPWR_c_1500_n N_VPWR_c_1501_n
+ N_VPWR_c_1502_n N_VPWR_c_1503_n N_VPWR_c_1504_n VPWR N_VPWR_c_1505_n
+ N_VPWR_c_1506_n N_VPWR_c_1507_n N_VPWR_c_1508_n N_VPWR_c_1492_n
+ N_VPWR_c_1510_n N_VPWR_c_1511_n N_VPWR_c_1512_n N_VPWR_c_1513_n
+ N_VPWR_c_1514_n PM_SKY130_FD_SC_HD__DFRBP_1%VPWR
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_448_47# N_A_448_47#_M1029_d N_A_448_47#_M1028_d
+ N_A_448_47#_c_1648_n N_A_448_47#_c_1665_n N_A_448_47#_c_1656_n
+ PM_SKY130_FD_SC_HD__DFRBP_1%A_448_47#
x_PM_SKY130_FD_SC_HD__DFRBP_1%A_651_413# N_A_651_413#_M1007_d
+ N_A_651_413#_M1031_d N_A_651_413#_c_1682_n N_A_651_413#_c_1683_n
+ N_A_651_413#_c_1684_n N_A_651_413#_c_1685_n
+ PM_SKY130_FD_SC_HD__DFRBP_1%A_651_413#
x_PM_SKY130_FD_SC_HD__DFRBP_1%Q N_Q_M1019_d N_Q_M1011_d N_Q_c_1721_n
+ N_Q_c_1722_n Q N_Q_c_1720_n Q PM_SKY130_FD_SC_HD__DFRBP_1%Q
x_PM_SKY130_FD_SC_HD__DFRBP_1%Q_N N_Q_N_M1002_d N_Q_N_M1013_d N_Q_N_c_1748_n
+ N_Q_N_c_1751_n N_Q_N_c_1752_n N_Q_N_c_1749_n Q_N Q_N
+ PM_SKY130_FD_SC_HD__DFRBP_1%Q_N
x_PM_SKY130_FD_SC_HD__DFRBP_1%VGND N_VGND_M1027_d N_VGND_M1029_s N_VGND_M1004_d
+ N_VGND_M1026_d N_VGND_M1019_s N_VGND_M1006_d N_VGND_c_1764_n N_VGND_c_1765_n
+ N_VGND_c_1766_n N_VGND_c_1767_n N_VGND_c_1768_n N_VGND_c_1769_n
+ N_VGND_c_1770_n N_VGND_c_1771_n N_VGND_c_1772_n N_VGND_c_1773_n
+ N_VGND_c_1774_n N_VGND_c_1775_n N_VGND_c_1776_n N_VGND_c_1777_n
+ N_VGND_c_1778_n VGND N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n
+ N_VGND_c_1782_n N_VGND_c_1783_n PM_SKY130_FD_SC_HD__DFRBP_1%VGND
cc_1 VNB N_CLK_c_217_n 0.0577303f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.325
cc_2 VNB N_CLK_c_218_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0158337f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_27_47#_M1015_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_5 VNB N_A_27_47#_M1009_g 0.0209769f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_6 VNB N_A_27_47#_c_259_n 0.00890826f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_7 VNB N_A_27_47#_c_260_n 0.0150251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_261_n 0.00188961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_262_n 0.0380394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1021_g 0.0280213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_264_n 0.0111414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_265_n 7.34103e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_266_n 0.00783792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_267_n 0.0271377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_268_n 0.00215116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_269_n 0.0264033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_270_n 6.62431e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_271_n 0.0023967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_272_n 0.00191399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_273_n 0.0231886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_274_n 0.0236925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_275_n 0.00799011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_276_n 0.00574157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_D_M1029_g 0.0533319f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_25 VNB N_D_c_494_n 0.0139927f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_26 VNB N_D_c_495_n 0.0188284f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_27 VNB N_A_193_47#_M1020_g 0.0237069f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_28 VNB N_A_193_47#_c_547_n 0.0181872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_c_548_n 0.00292129f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_30 VNB N_A_193_47#_c_549_n 0.00474375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_193_47#_c_550_n 0.0376939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_193_47#_c_551_n 0.00318417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_552_n 0.027804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_c_553_n 0.0131434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_761_289#_M1003_g 0.0470937f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_36 VNB N_A_761_289#_c_759_n 0.00648449f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_37 VNB N_RESET_B_M1031_g 0.00906477f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_38 VNB N_RESET_B_M1005_g 0.0270317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_M1018_g 9.0366e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_40 VNB RESET_B 0.00278754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_RESET_B_c_871_n 0.00606631f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.16
cc_42 VNB N_RESET_B_c_872_n 0.010211f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_43 VNB N_RESET_B_c_873_n 0.0158918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_RESET_B_c_874_n 6.54108e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_875_n 0.0012119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_c_876_n 0.0033021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_877_n 0.0257225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_878_n 0.0174472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_879_n 0.0250293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_880_n 0.00240216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_543_47#_M1022_g 0.0193117f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_52 VNB N_A_543_47#_c_1023_n 0.0116433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_543_47#_c_1024_n 0.00578907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_543_47#_c_1025_n 0.00317656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_543_47#_c_1026_n 0.00141599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_543_47#_c_1027_n 0.0285537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1283_21#_M1026_g 0.02143f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_58 VNB N_A_1283_21#_M1008_g 0.00982494f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_59 VNB N_A_1283_21#_c_1150_n 0.0236735f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_60 VNB N_A_1283_21#_c_1151_n 0.0442415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1283_21#_c_1152_n 0.0157199f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_62 VNB N_A_1283_21#_c_1153_n 0.0304581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1283_21#_c_1154_n 0.017939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1283_21#_c_1155_n 0.0258772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1283_21#_c_1156_n 0.00209314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1283_21#_c_1157_n 6.41492e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1283_21#_c_1158_n 0.00280904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1283_21#_c_1159_n 0.0062084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1283_21#_c_1160_n 0.0073052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1283_21#_c_1161_n 0.0161291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1283_21#_c_1162_n 0.0464685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1108_47#_M1001_g 0.0448001f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_73 VNB N_A_1108_47#_c_1339_n 0.00617495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1847_47#_c_1444_n 0.00662965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1847_47#_c_1445_n 0.00575059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1847_47#_c_1446_n 0.0256191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1847_47#_c_1447_n 0.0202221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VPWR_c_1492_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_448_47#_c_1648_n 0.0051081f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_80 VNB N_Q_c_1720_n 0.00683788f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_81 VNB N_Q_N_c_1748_n 0.0154962f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_82 VNB N_Q_N_c_1749_n 0.00479254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB Q_N 0.0240401f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_84 VNB N_VGND_c_1764_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1765_n 0.0192467f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_86 VNB N_VGND_c_1766_n 0.00858778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1767_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1768_n 0.00480551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1769_n 0.00468725f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1770_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1771_n 0.0711727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1772_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1773_n 0.0475682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1774_n 0.00362291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1775_n 0.0357945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1776_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1777_n 0.0349491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1778_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1779_n 0.0147253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1780_n 0.0204935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1781_n 0.513854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1782_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1783_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VPB N_CLK_c_217_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.325
cc_105 VPB N_CLK_c_221_n 0.0162394f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_106 VPB N_CLK_c_222_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_107 VPB N_CLK_c_223_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_108 VPB CLK 0.0152002f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_109 VPB N_A_27_47#_M1000_g 0.0393762f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_110 VPB N_A_27_47#_c_260_n 0.0162228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_261_n 0.00553413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_27_47#_M1007_g 0.0491475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_27_47#_c_262_n 0.0112552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_27_47#_M1025_g 0.0463897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_27_47#_c_283_n 0.00118305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_27_47#_c_284_n 0.0297336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_268_n 4.26143e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_27_47#_c_271_n 0.00320885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_272_n 3.60888e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_273_n 0.012023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_275_n 0.00283708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_276_n 9.66093e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_D_M1028_g 0.0392567f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_124 VPB N_D_c_494_n 0.0355299f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_125 VPB N_D_c_498_n 0.0197975f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB D 0.0281043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_D_c_495_n 0.00129394f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_128 VPB N_A_193_47#_M1030_g 0.0211021f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_129 VPB N_A_193_47#_M1012_g 0.0185283f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_130 VPB N_A_193_47#_c_548_n 0.00403367f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_131 VPB N_A_193_47#_c_549_n 0.00387694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_193_47#_c_558_n 0.00222651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_193_47#_c_559_n 0.00160169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_193_47#_c_560_n 0.012684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_193_47#_c_561_n 0.00221097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_193_47#_c_562_n 0.0160841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_193_47#_c_563_n 0.00178929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_193_47#_c_564_n 0.005939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_193_47#_c_565_n 0.00225318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_193_47#_c_566_n 0.0267174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_193_47#_c_567_n 0.0305358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_193_47#_c_568_n 0.00788798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_193_47#_c_553_n 0.0113511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_761_289#_M1010_g 0.0280169f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_145 VPB N_A_761_289#_M1003_g 0.00821552f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_146 VPB N_A_761_289#_c_762_n 0.0139674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_761_289#_c_763_n 0.0282266f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_148 VPB N_A_761_289#_c_759_n 0.00172612f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_149 VPB N_RESET_B_M1031_g 0.0573733f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_150 VPB N_RESET_B_M1018_g 0.0509764f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_151 VPB N_RESET_B_c_880_n 0.00388678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_543_47#_c_1028_n 0.0276965f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_153 VPB N_A_543_47#_c_1029_n 0.0174138f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_154 VPB N_A_543_47#_c_1030_n 0.00704944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_543_47#_c_1024_n 0.00782024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_543_47#_c_1025_n 0.00346469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_543_47#_c_1026_n 0.00113493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_543_47#_c_1027_n 0.0226938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_1283_21#_M1008_g 0.0502048f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_160 VPB N_A_1283_21#_M1011_g 0.0249724f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.16
cc_161 VPB N_A_1283_21#_c_1151_n 0.0242502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_1283_21#_c_1152_n 0.00237174f $X=-0.19 $Y=1.305 $X2=0.265
+ $Y2=1.53
cc_163 VPB N_A_1283_21#_c_1153_n 5.42563e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_1283_21#_M1024_g 0.0252926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_1283_21#_c_1155_n 0.0111379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_1283_21#_c_1170_n 0.0126997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_1283_21#_c_1171_n 0.0137966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1283_21#_c_1172_n 0.00465963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_1283_21#_c_1173_n 0.00304108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1283_21#_c_1174_n 0.00891481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_1283_21#_c_1161_n 0.00907377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1108_47#_M1016_g 0.0253068f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_173 VPB N_A_1108_47#_M1001_g 0.0114779f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_174 VPB N_A_1108_47#_c_1342_n 0.0110964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1108_47#_c_1343_n 0.00205899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1108_47#_c_1344_n 0.0229549f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1108_47#_c_1345_n 0.0286887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1847_47#_M1013_g 0.0232251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1847_47#_c_1449_n 0.0107428f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.16
cc_180 VPB N_A_1847_47#_c_1445_n 0.0055902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_1847_47#_c_1446_n 0.00618542f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1493_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1494_n 0.00927346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1495_n 0.00273179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1496_n 0.00650484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1497_n 0.0022316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1498_n 0.00472845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1499_n 0.0475825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1500_n 0.00507461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1501_n 0.0394977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1502_n 0.0035344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1503_n 0.034562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1504_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1505_n 0.0146985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1506_n 0.0265368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1507_n 0.0170787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1508_n 0.0210182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1492_n 0.0712388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1510_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1511_n 0.00477715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1512_n 0.00572697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1513_n 0.0122509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1514_n 0.0135196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_448_47#_c_1648_n 0.00778159f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_205 VPB N_A_651_413#_c_1682_n 4.85478e-19 $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_206 VPB N_A_651_413#_c_1683_n 0.00848337f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.665
cc_207 VPB N_A_651_413#_c_1684_n 0.00246665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_651_413#_c_1685_n 7.0682e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_Q_c_1721_n 0.0127741f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_210 VPB N_Q_c_1722_n 0.00466507f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_211 VPB N_Q_c_1720_n 0.00208449f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_212 VPB N_Q_N_c_1751_n 0.00604747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_Q_N_c_1752_n 0.028786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB Q_N 0.00716904f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_215 N_CLK_c_217_n N_A_27_47#_M1015_g 0.00510767f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_216 N_CLK_c_218_n N_A_27_47#_M1015_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_217 CLK N_A_27_47#_M1015_g 3.09846e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_218 N_CLK_c_221_n N_A_27_47#_M1000_g 0.00531917f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_219 N_CLK_c_223_n N_A_27_47#_M1000_g 0.0275602f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_220 CLK N_A_27_47#_M1000_g 5.73308e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_221 N_CLK_c_217_n N_A_27_47#_c_265_n 0.00787672f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_222 N_CLK_c_218_n N_A_27_47#_c_265_n 0.00695273f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_223 CLK N_A_27_47#_c_265_n 0.00736322f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_224 N_CLK_c_217_n N_A_27_47#_c_266_n 0.0070116f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_225 CLK N_A_27_47#_c_266_n 0.0220292f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_226 N_CLK_c_222_n N_A_27_47#_c_283_n 0.0128403f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_227 N_CLK_c_223_n N_A_27_47#_c_283_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_228 CLK N_A_27_47#_c_283_n 0.00728212f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_229 N_CLK_c_217_n N_A_27_47#_c_284_n 4.93713e-19 $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_230 N_CLK_c_222_n N_A_27_47#_c_284_n 2.20356e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_231 N_CLK_c_223_n N_A_27_47#_c_284_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_232 CLK N_A_27_47#_c_284_n 0.0231715f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_233 CLK N_A_27_47#_c_268_n 0.00784263f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_234 N_CLK_c_217_n N_A_27_47#_c_271_n 0.00475399f $X=0.305 $Y=1.325 $X2=0
+ $Y2=0
cc_235 N_CLK_c_221_n N_A_27_47#_c_271_n 7.09762e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_236 N_CLK_c_223_n N_A_27_47#_c_271_n 0.00454961f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_237 CLK N_A_27_47#_c_271_n 0.048988f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_238 N_CLK_c_217_n N_A_27_47#_c_273_n 0.0179788f $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_239 CLK N_A_27_47#_c_273_n 0.00143822f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_240 N_CLK_c_222_n N_VPWR_c_1493_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_241 N_CLK_c_222_n N_VPWR_c_1505_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_222_n N_VPWR_c_1492_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_243 N_CLK_c_218_n N_VGND_c_1764_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_244 N_CLK_c_217_n N_VGND_c_1779_n 4.74473e-19 $X=0.305 $Y=1.325 $X2=0 $Y2=0
cc_245 N_CLK_c_218_n N_VGND_c_1779_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_246 N_CLK_c_218_n N_VGND_c_1781_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_247 N_A_27_47#_M1009_g N_D_M1029_g 0.0124137f $X=2.64 $Y=0.415 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_259_n N_D_M1029_g 0.00561622f $X=2.642 $Y=1.245 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_267_n N_D_M1029_g 0.00237886f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_270_n N_D_M1029_g 0.00141197f $X=2.675 $Y=1.19 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_274_n N_D_M1029_g 0.0194268f $X=2.585 $Y=0.93 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_275_n N_D_M1029_g 0.00359265f $X=2.585 $Y=0.93 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_267_n N_D_c_494_n 0.00328759f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_273_n N_D_c_494_n 0.00307512f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_261_n N_D_c_498_n 0.00561622f $X=2.72 $Y=1.32 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_267_n N_D_c_498_n 0.00121575f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_267_n D 0.00176122f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_267_n N_D_c_495_n 0.0454089f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_259 N_A_27_47#_M1007_g N_A_193_47#_M1030_g 0.0202456f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1009_g N_A_193_47#_M1020_g 0.0132876f $X=2.64 $Y=0.415 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_M1021_g N_A_193_47#_c_547_n 0.0127456f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_M1025_g N_A_193_47#_M1012_g 0.0170357f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_260_n N_A_193_47#_c_548_n 0.0110546f $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1007_g N_A_193_47#_c_548_n 0.00405215f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_269_n N_A_193_47#_c_548_n 0.0110887f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_270_n N_A_193_47#_c_548_n 5.58797e-19 $X=2.675 $Y=1.19 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_274_n N_A_193_47#_c_548_n 0.00150746f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_275_n N_A_193_47#_c_548_n 0.0290824f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_262_n N_A_193_47#_c_549_n 0.00866804f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_270 N_A_27_47#_M1021_g N_A_193_47#_c_549_n 3.88889e-19 $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_269_n N_A_193_47#_c_549_n 0.0145489f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_272_n N_A_193_47#_c_549_n 5.12182e-19 $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_276_n N_A_193_47#_c_549_n 0.045569f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1021_g N_A_193_47#_c_550_n 0.021218f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_269_n N_A_193_47#_c_550_n 0.00188252f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_276_n N_A_193_47#_c_550_n 0.00185788f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_262_n N_A_193_47#_c_558_n 0.00133124f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_278 N_A_27_47#_M1025_g N_A_193_47#_c_558_n 0.0109104f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_269_n N_A_193_47#_c_558_n 0.00491458f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_276_n N_A_193_47#_c_558_n 0.00841432f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_260_n N_A_193_47#_c_551_n 0.00114671f $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_269_n N_A_193_47#_c_551_n 0.00894827f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_274_n N_A_193_47#_c_551_n 7.0175e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_275_n N_A_193_47#_c_551_n 0.0184123f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_260_n N_A_193_47#_c_552_n 0.0226065f $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_269_n N_A_193_47#_c_552_n 0.00261571f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_274_n N_A_193_47#_c_552_n 0.0175107f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_275_n N_A_193_47#_c_552_n 8.36786e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_267_n N_A_193_47#_c_560_n 0.0494564f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_269_n N_A_193_47#_c_560_n 0.00684111f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_270_n N_A_193_47#_c_560_n 0.0133153f $X=2.675 $Y=1.19 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_275_n N_A_193_47#_c_560_n 0.00548636f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1000_g N_A_193_47#_c_561_n 0.00307706f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_283_n N_A_193_47#_c_561_n 0.00527405f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_284_n N_A_193_47#_c_561_n 3.65662e-19 $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_267_n N_A_193_47#_c_561_n 0.0136396f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_271_n N_A_193_47#_c_561_n 0.00104863f $X=0.695 $Y=1.19 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1007_g N_A_193_47#_c_562_n 0.00283709f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1025_g N_A_193_47#_c_562_n 0.00608452f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_300 N_A_27_47#_c_269_n N_A_193_47#_c_562_n 0.121215f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_260_n N_A_193_47#_c_563_n 3.78985e-19 $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1007_g N_A_193_47#_c_563_n 0.00277626f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_269_n N_A_193_47#_c_563_n 0.0129897f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_260_n N_A_193_47#_c_564_n 8.09221e-19 $X=3.105 $Y=1.32 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_261_n N_A_193_47#_c_564_n 0.00542966f $X=2.72 $Y=1.32 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1007_g N_A_193_47#_c_564_n 0.00325095f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_269_n N_A_193_47#_c_564_n 0.00524922f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_270_n N_A_193_47#_c_564_n 2.72172e-19 $X=2.675 $Y=1.19 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_275_n N_A_193_47#_c_564_n 0.00817823f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1025_g N_A_193_47#_c_565_n 0.00147605f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_311 N_A_27_47#_c_272_n N_A_193_47#_c_565_n 0.0139913f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_276_n N_A_193_47#_c_565_n 7.23087e-19 $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_261_n N_A_193_47#_c_566_n 0.0187505f $X=2.72 $Y=1.32 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_M1007_g N_A_193_47#_c_566_n 0.0138904f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_274_n N_A_193_47#_c_566_n 6.13774e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_275_n N_A_193_47#_c_566_n 0.00142642f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_262_n N_A_193_47#_c_567_n 0.00311561f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_318 N_A_27_47#_M1025_g N_A_193_47#_c_567_n 0.0207208f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_272_n N_A_193_47#_c_567_n 0.00104369f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_276_n N_A_193_47#_c_567_n 4.78088e-19 $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_262_n N_A_193_47#_c_568_n 0.00367588f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_M1025_g N_A_193_47#_c_568_n 0.00525218f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_323 N_A_27_47#_c_272_n N_A_193_47#_c_568_n 0.00244943f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_276_n N_A_193_47#_c_568_n 0.0147695f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1015_g N_A_193_47#_c_553_n 0.0227708f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_265_n N_A_193_47#_c_553_n 0.01251f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_283_n N_A_193_47#_c_553_n 0.00874344f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_267_n N_A_193_47#_c_553_n 0.0193882f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_268_n N_A_193_47#_c_553_n 0.0021977f $X=0.84 $Y=1.19 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_271_n N_A_193_47#_c_553_n 0.0685829f $X=0.695 $Y=1.19 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_260_n N_A_761_289#_M1003_g 0.00256582f $X=3.105 $Y=1.32
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_269_n N_A_761_289#_M1003_g 0.0022411f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_M1007_g N_A_761_289#_c_762_n 6.41799e-19 $X=3.18 $Y=2.275
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_269_n N_A_761_289#_c_762_n 0.00791634f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_M1007_g N_A_761_289#_c_763_n 0.01719f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_269_n N_A_761_289#_c_759_n 0.0128787f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_M1025_g N_A_761_289#_c_771_n 0.00242771f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_269_n N_A_761_289#_c_771_n 0.00205194f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_M1025_g N_A_761_289#_c_773_n 0.00383854f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_269_n N_A_761_289#_c_774_n 7.74909e-19 $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_M1025_g N_A_761_289#_c_775_n 2.31682e-19 $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_c_269_n N_RESET_B_M1031_g 0.00162058f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_269_n N_RESET_B_c_871_n 0.0589913f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_269_n N_RESET_B_c_872_n 0.00492178f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_262_n N_RESET_B_c_873_n 5.35574e-19 $X=5.845 $Y=1.395 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_269_n N_RESET_B_c_873_n 0.12382f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_272_n N_RESET_B_c_873_n 0.0255775f $X=6.11 $Y=1.19 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_276_n N_RESET_B_c_873_n 0.0184793f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_269_n N_RESET_B_c_877_n 0.00221649f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_M1025_g N_A_543_47#_c_1028_n 0.0268099f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_269_n N_A_543_47#_c_1028_n 0.00359773f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_M1007_g N_A_543_47#_c_1037_n 0.0169036f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_260_n N_A_543_47#_c_1030_n 0.00114222f $X=3.105 $Y=1.32
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_M1007_g N_A_543_47#_c_1030_n 0.0167379f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_269_n N_A_543_47#_c_1030_n 4.47512e-19 $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_269_n N_A_543_47#_c_1023_n 0.0135671f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_269_n N_A_543_47#_c_1024_n 0.0379321f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_260_n N_A_543_47#_c_1025_n 0.00382694f $X=3.105 $Y=1.32
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_269_n N_A_543_47#_c_1025_n 0.0134122f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_269_n N_A_543_47#_c_1026_n 0.0100049f $X=5.965 $Y=1.19 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_269_n N_A_543_47#_c_1027_n 0.00476255f $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_M1021_g N_A_1283_21#_M1026_g 0.0308149f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_276_n N_A_1283_21#_M1026_g 6.8514e-19 $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_262_n N_A_1283_21#_M1008_g 0.00175162f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_M1025_g N_A_1283_21#_M1008_g 0.00178563f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_366 N_A_27_47#_c_262_n N_A_1283_21#_c_1162_n 0.0089256f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_c_262_n N_A_1108_47#_c_1346_n 8.21465e-19 $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_M1021_g N_A_1108_47#_c_1346_n 0.0109079f $X=6.01 $Y=0.415
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_276_n N_A_1108_47#_c_1346_n 0.0215171f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_M1025_g N_A_1108_47#_c_1349_n 0.00464335f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_262_n N_A_1108_47#_c_1339_n 0.00235645f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_M1021_g N_A_1108_47#_c_1339_n 0.00182809f $X=6.01 $Y=0.415
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_272_n N_A_1108_47#_c_1339_n 0.00772758f $X=6.11 $Y=1.19
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_276_n N_A_1108_47#_c_1339_n 0.0429822f $X=6.07 $Y=1.11 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_262_n N_A_1108_47#_c_1342_n 0.00164867f $X=5.845 $Y=1.395
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_M1025_g N_A_1108_47#_c_1342_n 0.00219772f $X=5.845 $Y=2.275
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_276_n N_A_1108_47#_c_1342_n 8.53289e-19 $X=6.07 $Y=1.11
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_c_283_n N_VPWR_M1014_d 0.00167655f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_379 N_A_27_47#_M1000_g N_VPWR_c_1493_n 0.00939211f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_283_n N_VPWR_c_1493_n 0.0175536f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_381 N_A_27_47#_c_284_n N_VPWR_c_1493_n 0.0127425f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_382 N_A_27_47#_M1025_g N_VPWR_c_1496_n 0.00111281f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_M1007_g N_VPWR_c_1499_n 0.00357863f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_M1025_g N_VPWR_c_1501_n 0.0055505f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_283_n N_VPWR_c_1505_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_386 N_A_27_47#_c_284_n N_VPWR_c_1505_n 0.0181185f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_387 N_A_27_47#_M1000_g N_VPWR_c_1506_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_M1000_g N_VPWR_c_1492_n 0.00859122f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1007_g N_VPWR_c_1492_n 0.00600164f $X=3.18 $Y=2.275 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_M1025_g N_VPWR_c_1492_n 0.00644128f $X=5.845 $Y=2.275 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_283_n N_VPWR_c_1492_n 0.00507261f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_284_n N_VPWR_c_1492_n 0.00973967f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_M1009_g N_A_448_47#_c_1648_n 0.00138047f $X=2.64 $Y=0.415
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_259_n N_A_448_47#_c_1648_n 3.20092e-19 $X=2.642 $Y=1.245
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_267_n N_A_448_47#_c_1648_n 0.0205223f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_270_n N_A_448_47#_c_1648_n 0.00258354f $X=2.675 $Y=1.19
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_274_n N_A_448_47#_c_1648_n 3.50691e-19 $X=2.585 $Y=0.93
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_275_n N_A_448_47#_c_1648_n 0.0463537f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_270_n N_A_448_47#_c_1656_n 6.44071e-19 $X=2.675 $Y=1.19
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_274_n N_A_448_47#_c_1656_n 4.7648e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_275_n N_A_448_47#_c_1656_n 0.0060732f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_M1007_g N_A_651_413#_c_1682_n 8.91651e-19 $X=3.18 $Y=2.275
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_269_n N_A_651_413#_c_1683_n 2.79618e-19 $X=5.965 $Y=1.19
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_M1007_g N_A_651_413#_c_1684_n 4.86622e-19 $X=3.18 $Y=2.275
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_265_n N_VGND_M1027_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_406 N_A_27_47#_M1015_g N_VGND_c_1764_n 0.0111875f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_265_n N_VGND_c_1764_n 0.0166634f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_408 N_A_27_47#_c_268_n N_VGND_c_1764_n 9.27814e-19 $X=0.84 $Y=1.19 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_273_n N_VGND_c_1764_n 5.7379e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_M1015_g N_VGND_c_1765_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_M1015_g N_VGND_c_1766_n 0.00430756f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_M1009_g N_VGND_c_1771_n 0.00585385f $X=2.64 $Y=0.415 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_274_n N_VGND_c_1771_n 2.72564e-19 $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_M1021_g N_VGND_c_1773_n 0.00357877f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_264_n N_VGND_c_1779_n 0.0108577f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_416 N_A_27_47#_c_265_n N_VGND_c_1779_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_M1027_s N_VGND_c_1781_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_M1015_g N_VGND_c_1781_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_M1009_g N_VGND_c_1781_n 0.00642996f $X=2.64 $Y=0.415 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_M1021_g N_VGND_c_1781_n 0.00565064f $X=6.01 $Y=0.415 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_264_n N_VGND_c_1781_n 0.00916732f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_265_n N_VGND_c_1781_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_275_n N_VGND_c_1781_n 0.00714893f $X=2.585 $Y=0.93 $X2=0
+ $Y2=0
cc_424 N_D_M1028_g N_A_193_47#_M1030_g 0.014327f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_425 N_D_c_498_n N_A_193_47#_c_548_n 0.00459927f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_426 N_D_M1028_g N_A_193_47#_c_560_n 0.00135182f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_427 N_D_c_494_n N_A_193_47#_c_560_n 0.00295589f $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_428 D N_A_193_47#_c_560_n 0.0339847f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_429 D N_A_193_47#_c_561_n 0.00279509f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_430 N_D_c_498_n N_A_193_47#_c_564_n 0.00143055f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_431 N_D_c_498_n N_A_193_47#_c_566_n 0.0151527f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_432 N_D_c_494_n N_A_193_47#_c_553_n 8.20589e-19 $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_433 D N_A_193_47#_c_553_n 0.0745399f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_434 N_D_c_495_n N_A_193_47#_c_553_n 0.0518322f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_435 N_D_M1028_g N_VPWR_c_1494_n 0.0044954f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_436 N_D_c_494_n N_VPWR_c_1494_n 0.00536585f $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_437 D N_VPWR_c_1494_n 0.0228549f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_438 N_D_M1028_g N_VPWR_c_1499_n 0.00420613f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_439 D N_VPWR_c_1506_n 0.0211539f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_440 N_D_M1028_g N_VPWR_c_1492_n 0.00685455f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_441 D N_VPWR_c_1492_n 0.00588351f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_442 N_D_M1029_g N_A_448_47#_c_1648_n 0.0279651f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_443 N_D_M1028_g N_A_448_47#_c_1648_n 0.0259313f $X=2.225 $Y=2.275 $X2=0 $Y2=0
cc_444 N_D_c_494_n N_A_448_47#_c_1648_n 0.00781441f $X=2.09 $Y=1.465 $X2=0 $Y2=0
cc_445 N_D_c_498_n N_A_448_47#_c_1648_n 0.0131062f $X=2.09 $Y=1.3 $X2=0 $Y2=0
cc_446 D N_A_448_47#_c_1648_n 0.0365307f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_447 N_D_c_495_n N_A_448_47#_c_1648_n 0.0623934f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_448 N_D_M1029_g N_A_448_47#_c_1665_n 0.00588428f $X=2.165 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_D_M1029_g N_A_448_47#_c_1656_n 0.00163056f $X=2.165 $Y=0.445 $X2=0
+ $Y2=0
cc_450 N_D_c_495_n N_VGND_M1029_s 0.00431154f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_451 N_D_c_495_n N_VGND_c_1765_n 0.00272126f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_452 N_D_M1029_g N_VGND_c_1766_n 0.00675175f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_453 N_D_c_495_n N_VGND_c_1766_n 0.0275242f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_454 N_D_M1029_g N_VGND_c_1771_n 0.00367956f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_455 N_D_M1029_g N_VGND_c_1781_n 0.00677951f $X=2.165 $Y=0.445 $X2=0 $Y2=0
cc_456 N_D_c_495_n N_VGND_c_1781_n 0.005702f $X=1.79 $Y=1.465 $X2=0 $Y2=0
cc_457 N_A_193_47#_c_558_n N_A_761_289#_M1017_d 2.38738e-19 $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_458 N_A_193_47#_c_559_n N_A_761_289#_M1017_d 0.00203554f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_459 N_A_193_47#_c_562_n N_A_761_289#_M1017_d 0.00257222f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_460 N_A_193_47#_c_562_n N_A_761_289#_M1010_g 0.0023317f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_461 N_A_193_47#_M1020_g N_A_761_289#_M1003_g 0.00811432f $X=3.12 $Y=0.415
+ $X2=0 $Y2=0
cc_462 N_A_193_47#_c_552_n N_A_761_289#_M1003_g 0.00345535f $X=3.095 $Y=0.9
+ $X2=0 $Y2=0
cc_463 N_A_193_47#_c_562_n N_A_761_289#_c_762_n 0.0223886f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_464 N_A_193_47#_c_562_n N_A_761_289#_c_763_n 0.00270169f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_465 N_A_193_47#_c_547_n N_A_761_289#_c_784_n 0.00348356f $X=5.465 $Y=0.705
+ $X2=0 $Y2=0
cc_466 N_A_193_47#_c_559_n N_A_761_289#_c_759_n 0.00219387f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_467 N_A_193_47#_c_562_n N_A_761_289#_c_786_n 0.00749812f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_468 N_A_193_47#_c_559_n N_A_761_289#_c_771_n 0.0134011f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_469 N_A_193_47#_c_562_n N_A_761_289#_c_771_n 0.0181068f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_470 N_A_193_47#_c_565_n N_A_761_289#_c_771_n 0.00186336f $X=6.11 $Y=1.87
+ $X2=0 $Y2=0
cc_471 N_A_193_47#_c_568_n N_A_761_289#_c_771_n 0.00477525f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_472 N_A_193_47#_c_562_n N_A_761_289#_c_791_n 0.00696518f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_473 N_A_193_47#_c_549_n N_A_761_289#_c_774_n 0.0522946f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_474 N_A_193_47#_c_550_n N_A_761_289#_c_774_n 0.00348356f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_475 N_A_193_47#_c_559_n N_A_761_289#_c_775_n 0.0105163f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_476 N_A_193_47#_c_562_n N_RESET_B_M1031_g 0.00286324f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_477 N_A_193_47#_c_549_n N_RESET_B_c_873_n 0.0127742f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_478 N_A_193_47#_c_550_n N_RESET_B_c_873_n 0.00393129f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_479 N_A_193_47#_c_547_n N_A_543_47#_M1022_g 0.0103966f $X=5.465 $Y=0.705
+ $X2=0 $Y2=0
cc_480 N_A_193_47#_c_549_n N_A_543_47#_c_1028_n 7.67033e-19 $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_481 N_A_193_47#_c_550_n N_A_543_47#_c_1028_n 0.00138652f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_482 N_A_193_47#_c_559_n N_A_543_47#_c_1028_n 0.0016569f $X=5.675 $Y=1.58
+ $X2=0 $Y2=0
cc_483 N_A_193_47#_c_562_n N_A_543_47#_c_1029_n 0.0027309f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_484 N_A_193_47#_M1030_g N_A_543_47#_c_1037_n 0.00421429f $X=2.685 $Y=2.275
+ $X2=0 $Y2=0
cc_485 N_A_193_47#_c_560_n N_A_543_47#_c_1037_n 4.97575e-19 $X=2.845 $Y=1.87
+ $X2=0 $Y2=0
cc_486 N_A_193_47#_c_562_n N_A_543_47#_c_1037_n 0.00304089f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_487 N_A_193_47#_c_563_n N_A_543_47#_c_1037_n 0.0046344f $X=3.135 $Y=1.87
+ $X2=0 $Y2=0
cc_488 N_A_193_47#_c_564_n N_A_543_47#_c_1037_n 0.0208127f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_489 N_A_193_47#_c_566_n N_A_543_47#_c_1037_n 4.68077e-19 $X=2.695 $Y=1.74
+ $X2=0 $Y2=0
cc_490 N_A_193_47#_M1020_g N_A_543_47#_c_1058_n 0.00973778f $X=3.12 $Y=0.415
+ $X2=0 $Y2=0
cc_491 N_A_193_47#_c_551_n N_A_543_47#_c_1058_n 0.0121475f $X=3.095 $Y=0.9 $X2=0
+ $Y2=0
cc_492 N_A_193_47#_c_552_n N_A_543_47#_c_1058_n 0.00324607f $X=3.095 $Y=0.9
+ $X2=0 $Y2=0
cc_493 N_A_193_47#_M1030_g N_A_543_47#_c_1030_n 8.68564e-19 $X=2.685 $Y=2.275
+ $X2=0 $Y2=0
cc_494 N_A_193_47#_c_548_n N_A_543_47#_c_1030_n 0.0155497f $X=2.99 $Y=1.575
+ $X2=0 $Y2=0
cc_495 N_A_193_47#_c_562_n N_A_543_47#_c_1030_n 0.0157004f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_496 N_A_193_47#_c_563_n N_A_543_47#_c_1030_n 0.00273426f $X=3.135 $Y=1.87
+ $X2=0 $Y2=0
cc_497 N_A_193_47#_c_564_n N_A_543_47#_c_1030_n 0.0280664f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_498 N_A_193_47#_c_566_n N_A_543_47#_c_1030_n 2.1939e-19 $X=2.695 $Y=1.74
+ $X2=0 $Y2=0
cc_499 N_A_193_47#_M1020_g N_A_543_47#_c_1023_n 0.00647277f $X=3.12 $Y=0.415
+ $X2=0 $Y2=0
cc_500 N_A_193_47#_c_548_n N_A_543_47#_c_1023_n 0.00810958f $X=2.99 $Y=1.575
+ $X2=0 $Y2=0
cc_501 N_A_193_47#_c_551_n N_A_543_47#_c_1023_n 0.0159961f $X=3.095 $Y=0.9 $X2=0
+ $Y2=0
cc_502 N_A_193_47#_c_552_n N_A_543_47#_c_1023_n 0.00150777f $X=3.095 $Y=0.9
+ $X2=0 $Y2=0
cc_503 N_A_193_47#_c_548_n N_A_543_47#_c_1025_n 0.0123239f $X=2.99 $Y=1.575
+ $X2=0 $Y2=0
cc_504 N_A_193_47#_c_551_n N_A_543_47#_c_1025_n 7.96251e-19 $X=3.095 $Y=0.9
+ $X2=0 $Y2=0
cc_505 N_A_193_47#_c_562_n N_A_543_47#_c_1025_n 0.00748451f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_506 N_A_193_47#_c_550_n N_A_543_47#_c_1027_n 0.0103966f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_507 N_A_193_47#_M1012_g N_A_1283_21#_M1008_g 0.0335217f $X=6.275 $Y=2.275
+ $X2=0 $Y2=0
cc_508 N_A_193_47#_c_567_n N_A_1283_21#_M1008_g 0.0198765f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_509 N_A_193_47#_c_568_n N_A_1283_21#_M1008_g 0.00149229f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_510 N_A_193_47#_c_549_n N_A_1108_47#_c_1346_n 0.0060004f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_511 N_A_193_47#_c_550_n N_A_1108_47#_c_1346_n 0.00264523f $X=5.59 $Y=0.87
+ $X2=0 $Y2=0
cc_512 N_A_193_47#_M1012_g N_A_1108_47#_c_1349_n 0.0120896f $X=6.275 $Y=2.275
+ $X2=0 $Y2=0
cc_513 N_A_193_47#_c_558_n N_A_1108_47#_c_1349_n 7.08603e-19 $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_514 N_A_193_47#_c_562_n N_A_1108_47#_c_1349_n 9.42387e-19 $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_515 N_A_193_47#_c_565_n N_A_1108_47#_c_1349_n 0.00337735f $X=6.11 $Y=1.87
+ $X2=0 $Y2=0
cc_516 N_A_193_47#_c_567_n N_A_1108_47#_c_1349_n 3.21714e-19 $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_517 N_A_193_47#_c_568_n N_A_1108_47#_c_1349_n 0.02818f $X=6.265 $Y=1.74 $X2=0
+ $Y2=0
cc_518 N_A_193_47#_c_567_n N_A_1108_47#_c_1342_n 0.00200126f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_519 N_A_193_47#_c_568_n N_A_1108_47#_c_1342_n 0.0205187f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_520 N_A_193_47#_M1012_g N_A_1108_47#_c_1343_n 0.00233339f $X=6.275 $Y=2.275
+ $X2=0 $Y2=0
cc_521 N_A_193_47#_c_565_n N_A_1108_47#_c_1343_n 0.00209221f $X=6.11 $Y=1.87
+ $X2=0 $Y2=0
cc_522 N_A_193_47#_c_567_n N_A_1108_47#_c_1343_n 4.36865e-19 $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_523 N_A_193_47#_c_568_n N_A_1108_47#_c_1343_n 0.0162391f $X=6.265 $Y=1.74
+ $X2=0 $Y2=0
cc_524 N_A_193_47#_c_562_n N_VPWR_M1017_s 0.00127798f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_525 N_A_193_47#_c_553_n N_VPWR_c_1493_n 0.012721f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_526 N_A_193_47#_c_560_n N_VPWR_c_1494_n 0.00656454f $X=2.845 $Y=1.87 $X2=0
+ $Y2=0
cc_527 N_A_193_47#_c_553_n N_VPWR_c_1494_n 4.4131e-19 $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_528 N_A_193_47#_c_562_n N_VPWR_c_1495_n 0.00139202f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_c_562_n N_VPWR_c_1496_n 0.00326091f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_530 N_A_193_47#_M1030_g N_VPWR_c_1499_n 0.00427876f $X=2.685 $Y=2.275 $X2=0
+ $Y2=0
cc_531 N_A_193_47#_c_564_n N_VPWR_c_1499_n 0.00166184f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_532 N_A_193_47#_M1012_g N_VPWR_c_1501_n 0.00357877f $X=6.275 $Y=2.275 $X2=0
+ $Y2=0
cc_533 N_A_193_47#_c_553_n N_VPWR_c_1506_n 0.0120448f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_534 N_A_193_47#_M1030_g N_VPWR_c_1492_n 0.0059104f $X=2.685 $Y=2.275 $X2=0
+ $Y2=0
cc_535 N_A_193_47#_M1012_g N_VPWR_c_1492_n 0.00526867f $X=6.275 $Y=2.275 $X2=0
+ $Y2=0
cc_536 N_A_193_47#_c_560_n N_VPWR_c_1492_n 0.0759296f $X=2.845 $Y=1.87 $X2=0
+ $Y2=0
cc_537 N_A_193_47#_c_561_n N_VPWR_c_1492_n 0.0154052f $X=1.245 $Y=1.87 $X2=0
+ $Y2=0
cc_538 N_A_193_47#_c_562_n N_VPWR_c_1492_n 0.131729f $X=5.965 $Y=1.87 $X2=0
+ $Y2=0
cc_539 N_A_193_47#_c_563_n N_VPWR_c_1492_n 0.0159609f $X=3.135 $Y=1.87 $X2=0
+ $Y2=0
cc_540 N_A_193_47#_c_564_n N_VPWR_c_1492_n 0.00140124f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_541 N_A_193_47#_c_565_n N_VPWR_c_1492_n 0.0158397f $X=6.11 $Y=1.87 $X2=0
+ $Y2=0
cc_542 N_A_193_47#_c_566_n N_VPWR_c_1492_n 4.39969e-19 $X=2.695 $Y=1.74 $X2=0
+ $Y2=0
cc_543 N_A_193_47#_c_553_n N_VPWR_c_1492_n 0.0029375f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_544 N_A_193_47#_M1030_g N_A_448_47#_c_1648_n 0.00392609f $X=2.685 $Y=2.275
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_c_560_n N_A_448_47#_c_1648_n 0.0288873f $X=2.845 $Y=1.87
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_c_563_n N_A_448_47#_c_1648_n 0.00100139f $X=3.135 $Y=1.87
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_c_564_n N_A_448_47#_c_1648_n 0.0185011f $X=2.99 $Y=1.87 $X2=0
+ $Y2=0
cc_548 N_A_193_47#_c_566_n N_A_448_47#_c_1648_n 9.81315e-19 $X=2.695 $Y=1.74
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_562_n N_A_651_413#_c_1683_n 0.0297495f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_550 N_A_193_47#_c_562_n N_A_651_413#_c_1684_n 0.00857493f $X=5.965 $Y=1.87
+ $X2=0 $Y2=0
cc_551 N_A_193_47#_c_553_n N_VGND_c_1765_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_552 N_A_193_47#_c_553_n N_VGND_c_1766_n 0.00457032f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_553 N_A_193_47#_M1020_g N_VGND_c_1771_n 0.00368123f $X=3.12 $Y=0.415 $X2=0
+ $Y2=0
cc_554 N_A_193_47#_c_547_n N_VGND_c_1773_n 0.0051118f $X=5.465 $Y=0.705 $X2=0
+ $Y2=0
cc_555 N_A_193_47#_c_549_n N_VGND_c_1773_n 0.00183172f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_556 N_A_193_47#_c_550_n N_VGND_c_1773_n 2.13253e-19 $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_557 N_A_193_47#_M1015_d N_VGND_c_1781_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_558 N_A_193_47#_M1020_g N_VGND_c_1781_n 0.00618454f $X=3.12 $Y=0.415 $X2=0
+ $Y2=0
cc_559 N_A_193_47#_c_547_n N_VGND_c_1781_n 0.00654107f $X=5.465 $Y=0.705 $X2=0
+ $Y2=0
cc_560 N_A_193_47#_c_549_n N_VGND_c_1781_n 0.00150843f $X=5.59 $Y=0.87 $X2=0
+ $Y2=0
cc_561 N_A_193_47#_c_553_n N_VGND_c_1781_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_562 N_A_761_289#_M1010_g N_RESET_B_M1031_g 0.0224927f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_563 N_A_761_289#_M1003_g N_RESET_B_M1031_g 0.0177106f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_564 N_A_761_289#_c_762_n N_RESET_B_M1031_g 0.0115545f $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_565 N_A_761_289#_c_763_n N_RESET_B_M1031_g 0.0220442f $X=3.94 $Y=1.61 $X2=0
+ $Y2=0
cc_566 N_A_761_289#_c_759_n N_RESET_B_M1031_g 4.12396e-19 $X=5.19 $Y=1.525 $X2=0
+ $Y2=0
cc_567 N_A_761_289#_c_786_n N_RESET_B_M1031_g 0.00253836f $X=5.19 $Y=1.835 $X2=0
+ $Y2=0
cc_568 N_A_761_289#_c_791_n N_RESET_B_M1031_g 9.1253e-19 $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_569 N_A_761_289#_M1003_g N_RESET_B_c_871_n 0.00269192f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_570 N_A_761_289#_M1003_g N_RESET_B_c_872_n 0.0139529f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_571 N_A_761_289#_c_759_n N_RESET_B_c_872_n 0.0051548f $X=5.19 $Y=1.525 $X2=0
+ $Y2=0
cc_572 N_A_761_289#_c_774_n N_RESET_B_c_872_n 0.00197464f $X=5.145 $Y=0.835
+ $X2=0 $Y2=0
cc_573 N_A_761_289#_M1022_d N_RESET_B_c_873_n 3.28012e-19 $X=5.045 $Y=0.235
+ $X2=0 $Y2=0
cc_574 N_A_761_289#_c_762_n N_RESET_B_c_873_n 2.43406e-19 $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_575 N_A_761_289#_c_759_n N_RESET_B_c_873_n 0.00696464f $X=5.19 $Y=1.525 $X2=0
+ $Y2=0
cc_576 N_A_761_289#_c_809_p N_RESET_B_c_873_n 0.00227253f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_577 N_A_761_289#_c_774_n N_RESET_B_c_873_n 0.0121464f $X=5.145 $Y=0.835 $X2=0
+ $Y2=0
cc_578 N_A_761_289#_M1003_g N_RESET_B_c_878_n 0.0635296f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_579 N_A_761_289#_c_809_p N_RESET_B_c_878_n 9.82944e-19 $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_580 N_A_761_289#_c_784_n N_A_543_47#_M1022_g 0.0061779f $X=5.145 $Y=0.705
+ $X2=0 $Y2=0
cc_581 N_A_761_289#_c_759_n N_A_543_47#_M1022_g 0.0120311f $X=5.19 $Y=1.525
+ $X2=0 $Y2=0
cc_582 N_A_761_289#_c_809_p N_A_543_47#_M1022_g 0.00225962f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_583 N_A_761_289#_c_774_n N_A_543_47#_M1022_g 0.00423512f $X=5.145 $Y=0.835
+ $X2=0 $Y2=0
cc_584 N_A_761_289#_c_762_n N_A_543_47#_c_1028_n 0.00207011f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_585 N_A_761_289#_c_759_n N_A_543_47#_c_1028_n 0.00860889f $X=5.19 $Y=1.525
+ $X2=0 $Y2=0
cc_586 N_A_761_289#_c_774_n N_A_543_47#_c_1028_n 8.88512e-19 $X=5.145 $Y=0.835
+ $X2=0 $Y2=0
cc_587 N_A_761_289#_c_775_n N_A_543_47#_c_1028_n 0.00482334f $X=5.19 $Y=1.61
+ $X2=0 $Y2=0
cc_588 N_A_761_289#_c_786_n N_A_543_47#_c_1029_n 0.00308571f $X=5.19 $Y=1.835
+ $X2=0 $Y2=0
cc_589 N_A_761_289#_c_771_n N_A_543_47#_c_1029_n 0.0106757f $X=5.495 $Y=1.92
+ $X2=0 $Y2=0
cc_590 N_A_761_289#_c_791_n N_A_543_47#_c_1029_n 0.00298755f $X=5.275 $Y=1.92
+ $X2=0 $Y2=0
cc_591 N_A_761_289#_c_773_n N_A_543_47#_c_1029_n 0.00453769f $X=5.58 $Y=2.3
+ $X2=0 $Y2=0
cc_592 N_A_761_289#_c_775_n N_A_543_47#_c_1029_n 0.00385118f $X=5.19 $Y=1.61
+ $X2=0 $Y2=0
cc_593 N_A_761_289#_M1010_g N_A_543_47#_c_1037_n 0.00124715f $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_594 N_A_761_289#_M1003_g N_A_543_47#_c_1058_n 0.00466363f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_595 N_A_761_289#_M1010_g N_A_543_47#_c_1030_n 4.99336e-19 $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_596 N_A_761_289#_M1003_g N_A_543_47#_c_1030_n 0.00150033f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_597 N_A_761_289#_c_762_n N_A_543_47#_c_1030_n 0.00842454f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_598 N_A_761_289#_c_763_n N_A_543_47#_c_1030_n 0.0048158f $X=3.94 $Y=1.61
+ $X2=0 $Y2=0
cc_599 N_A_761_289#_M1003_g N_A_543_47#_c_1023_n 0.0114869f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_600 N_A_761_289#_M1003_g N_A_543_47#_c_1024_n 0.0109334f $X=3.95 $Y=0.445
+ $X2=0 $Y2=0
cc_601 N_A_761_289#_c_762_n N_A_543_47#_c_1024_n 0.063308f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_602 N_A_761_289#_c_763_n N_A_543_47#_c_1024_n 0.00338177f $X=3.94 $Y=1.61
+ $X2=0 $Y2=0
cc_603 N_A_761_289#_c_762_n N_A_543_47#_c_1026_n 0.0116159f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_604 N_A_761_289#_c_759_n N_A_543_47#_c_1026_n 0.0244986f $X=5.19 $Y=1.525
+ $X2=0 $Y2=0
cc_605 N_A_761_289#_c_762_n N_A_543_47#_c_1027_n 0.00751143f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_606 N_A_761_289#_c_773_n N_A_1108_47#_c_1349_n 0.0206716f $X=5.58 $Y=2.3
+ $X2=0 $Y2=0
cc_607 N_A_761_289#_c_762_n N_VPWR_M1017_s 0.00130684f $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_608 N_A_761_289#_c_786_n N_VPWR_M1017_s 0.00241466f $X=5.19 $Y=1.835 $X2=0
+ $Y2=0
cc_609 N_A_761_289#_c_791_n N_VPWR_M1017_s 0.00353974f $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_610 N_A_761_289#_M1010_g N_VPWR_c_1495_n 0.0044935f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_611 N_A_761_289#_c_762_n N_VPWR_c_1496_n 0.00261535f $X=5.105 $Y=1.61 $X2=0
+ $Y2=0
cc_612 N_A_761_289#_c_771_n N_VPWR_c_1496_n 0.003184f $X=5.495 $Y=1.92 $X2=0
+ $Y2=0
cc_613 N_A_761_289#_c_791_n N_VPWR_c_1496_n 0.008938f $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_614 N_A_761_289#_c_773_n N_VPWR_c_1496_n 0.0216047f $X=5.58 $Y=2.3 $X2=0
+ $Y2=0
cc_615 N_A_761_289#_M1010_g N_VPWR_c_1499_n 0.00432313f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_616 N_A_761_289#_c_771_n N_VPWR_c_1501_n 0.00199878f $X=5.495 $Y=1.92 $X2=0
+ $Y2=0
cc_617 N_A_761_289#_c_773_n N_VPWR_c_1501_n 0.0117479f $X=5.58 $Y=2.3 $X2=0
+ $Y2=0
cc_618 N_A_761_289#_M1017_d N_VPWR_c_1492_n 0.00326756f $X=5.425 $Y=1.645 $X2=0
+ $Y2=0
cc_619 N_A_761_289#_M1010_g N_VPWR_c_1492_n 0.00628822f $X=3.88 $Y=2.275 $X2=0
+ $Y2=0
cc_620 N_A_761_289#_c_771_n N_VPWR_c_1492_n 0.00181326f $X=5.495 $Y=1.92 $X2=0
+ $Y2=0
cc_621 N_A_761_289#_c_791_n N_VPWR_c_1492_n 4.80263e-19 $X=5.275 $Y=1.92 $X2=0
+ $Y2=0
cc_622 N_A_761_289#_c_773_n N_VPWR_c_1492_n 0.00306902f $X=5.58 $Y=2.3 $X2=0
+ $Y2=0
cc_623 N_A_761_289#_M1010_g N_A_651_413#_c_1682_n 7.77269e-19 $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_624 N_A_761_289#_M1010_g N_A_651_413#_c_1683_n 0.0117327f $X=3.88 $Y=2.275
+ $X2=0 $Y2=0
cc_625 N_A_761_289#_c_762_n N_A_651_413#_c_1683_n 0.0556558f $X=5.105 $Y=1.61
+ $X2=0 $Y2=0
cc_626 N_A_761_289#_c_763_n N_A_651_413#_c_1683_n 0.00332707f $X=3.94 $Y=1.61
+ $X2=0 $Y2=0
cc_627 N_A_761_289#_c_791_n N_A_651_413#_c_1683_n 0.00487217f $X=5.275 $Y=1.92
+ $X2=0 $Y2=0
cc_628 N_A_761_289#_c_809_p N_VGND_c_1767_n 0.0177195f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_629 N_A_761_289#_M1003_g N_VGND_c_1771_n 0.00585385f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_630 N_A_761_289#_c_809_p N_VGND_c_1773_n 0.0185505f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_631 N_A_761_289#_M1022_d N_VGND_c_1781_n 0.00246666f $X=5.045 $Y=0.235 $X2=0
+ $Y2=0
cc_632 N_A_761_289#_M1003_g N_VGND_c_1781_n 0.00633204f $X=3.95 $Y=0.445 $X2=0
+ $Y2=0
cc_633 N_A_761_289#_c_809_p N_VGND_c_1781_n 0.00609105f $X=5.2 $Y=0.36 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_872_n N_A_543_47#_M1022_g 0.00182794f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_873_n N_A_543_47#_M1022_g 0.00503251f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_874_n N_A_543_47#_M1022_g 4.85534e-19 $X=4.395 $Y=0.85 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_877_n N_A_543_47#_M1022_g 0.0070799f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_878_n N_A_543_47#_M1022_g 0.0129551f $X=4.37 $Y=0.765 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_871_n N_A_543_47#_c_1023_n 0.00858647f $X=4.28 $Y=0.85 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_872_n N_A_543_47#_c_1023_n 0.0146357f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_641 N_RESET_B_M1031_g N_A_543_47#_c_1024_n 0.00939437f $X=4.365 $Y=2.275
+ $X2=0 $Y2=0
cc_642 N_RESET_B_c_871_n N_A_543_47#_c_1024_n 0.00116894f $X=4.28 $Y=0.85 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_872_n N_A_543_47#_c_1024_n 0.0505984f $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_873_n N_A_543_47#_c_1024_n 0.00103298f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_645 N_RESET_B_c_877_n N_A_543_47#_c_1024_n 0.00314155f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_646 N_RESET_B_M1031_g N_A_543_47#_c_1026_n 8.07088e-19 $X=4.365 $Y=2.275
+ $X2=0 $Y2=0
cc_647 N_RESET_B_c_872_n N_A_543_47#_c_1026_n 7.26099e-19 $X=4.25 $Y=0.85 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_873_n N_A_543_47#_c_1026_n 0.00420388f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_877_n N_A_543_47#_c_1026_n 5.16993e-19 $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_650 N_RESET_B_M1031_g N_A_543_47#_c_1027_n 0.0181811f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_873_n N_A_543_47#_c_1027_n 8.21109e-19 $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_877_n N_A_543_47#_c_1027_n 0.00600523f $X=4.37 $Y=0.93 $X2=0
+ $Y2=0
cc_653 N_RESET_B_M1005_g N_A_1283_21#_M1026_g 0.0101625f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_654 N_RESET_B_c_873_n N_A_1283_21#_M1026_g 8.78915e-19 $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_655 N_RESET_B_M1018_g N_A_1283_21#_M1008_g 0.0333609f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_876_n N_A_1283_21#_M1008_g 0.00197455f $X=7.19 $Y=1.165 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_879_n N_A_1283_21#_M1008_g 0.00410139f $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_880_n N_A_1283_21#_M1008_g 0.00166565f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_880_n N_A_1283_21#_c_1155_n 2.17163e-19 $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_660 N_RESET_B_M1005_g N_A_1283_21#_c_1156_n 3.49601e-19 $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_661 RESET_B N_A_1283_21#_c_1156_n 0.00296317f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_662 N_RESET_B_c_873_n N_A_1283_21#_c_1156_n 0.0109517f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_663 N_RESET_B_c_875_n N_A_1283_21#_c_1156_n 0.00740908f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_664 N_RESET_B_c_879_n N_A_1283_21#_c_1156_n 4.00963e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_880_n N_A_1283_21#_c_1156_n 0.006652f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_666 N_RESET_B_M1005_g N_A_1283_21#_c_1157_n 0.00733777f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_667 RESET_B N_A_1283_21#_c_1157_n 0.0043842f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_668 N_RESET_B_c_875_n N_A_1283_21#_c_1157_n 4.41459e-19 $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_669 N_RESET_B_M1005_g N_A_1283_21#_c_1200_n 0.00588467f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_670 RESET_B N_A_1283_21#_c_1200_n 0.0122946f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_671 N_RESET_B_c_875_n N_A_1283_21#_c_1200_n 0.00297971f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_672 N_RESET_B_c_879_n N_A_1283_21#_c_1200_n 9.38055e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_673 N_RESET_B_c_880_n N_A_1283_21#_c_1200_n 0.00166967f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_674 N_RESET_B_M1005_g N_A_1283_21#_c_1205_n 0.00390919f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_675 N_RESET_B_M1018_g N_A_1283_21#_c_1173_n 0.00230253f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_676 RESET_B N_A_1283_21#_c_1159_n 0.0127158f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_677 N_RESET_B_c_875_n N_A_1283_21#_c_1159_n 6.44878e-19 $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_678 N_RESET_B_c_880_n N_A_1283_21#_c_1174_n 0.0036174f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_679 N_RESET_B_M1005_g N_A_1283_21#_c_1160_n 0.00557763f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_680 RESET_B N_A_1283_21#_c_1160_n 0.0119774f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_681 N_RESET_B_c_873_n N_A_1283_21#_c_1160_n 0.0122086f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_682 N_RESET_B_c_875_n N_A_1283_21#_c_1160_n 0.00988863f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_683 N_RESET_B_c_879_n N_A_1283_21#_c_1160_n 4.8034e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_684 N_RESET_B_c_880_n N_A_1283_21#_c_1160_n 0.00872348f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_685 RESET_B N_A_1283_21#_c_1161_n 0.015514f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_686 N_RESET_B_c_875_n N_A_1283_21#_c_1161_n 0.00108995f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_687 N_RESET_B_c_876_n N_A_1283_21#_c_1161_n 0.00125428f $X=7.19 $Y=1.165
+ $X2=0 $Y2=0
cc_688 N_RESET_B_c_880_n N_A_1283_21#_c_1161_n 0.0232032f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_689 N_RESET_B_M1005_g N_A_1283_21#_c_1162_n 0.00837678f $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_873_n N_A_1283_21#_c_1162_n 0.00336334f $X=7.045 $Y=0.85
+ $X2=0 $Y2=0
cc_691 N_RESET_B_c_875_n N_A_1283_21#_c_1162_n 0.00369633f $X=7.19 $Y=0.965
+ $X2=0 $Y2=0
cc_692 N_RESET_B_c_879_n N_A_1283_21#_c_1162_n 0.0123335f $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_693 N_RESET_B_c_880_n N_A_1283_21#_c_1162_n 5.46251e-19 $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_694 N_RESET_B_M1018_g N_A_1108_47#_M1016_g 0.0209789f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_695 N_RESET_B_M1005_g N_A_1108_47#_M1001_g 0.0345821f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_696 N_RESET_B_M1018_g N_A_1108_47#_M1001_g 0.00874253f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_697 RESET_B N_A_1108_47#_M1001_g 0.00842841f $X=7.405 $Y=0.765 $X2=0 $Y2=0
cc_698 N_RESET_B_c_879_n N_A_1108_47#_M1001_g 0.0210473f $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_699 N_RESET_B_c_880_n N_A_1108_47#_M1001_g 0.00864073f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_700 N_RESET_B_c_873_n N_A_1108_47#_c_1346_n 0.012043f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_701 N_RESET_B_M1005_g N_A_1108_47#_c_1339_n 3.06785e-19 $X=7.235 $Y=0.445
+ $X2=0 $Y2=0
cc_702 N_RESET_B_c_873_n N_A_1108_47#_c_1339_n 0.0190486f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_703 N_RESET_B_c_876_n N_A_1108_47#_c_1339_n 0.00350005f $X=7.19 $Y=1.165
+ $X2=0 $Y2=0
cc_704 N_RESET_B_c_880_n N_A_1108_47#_c_1339_n 0.00372747f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_705 N_RESET_B_M1018_g N_A_1108_47#_c_1342_n 0.00109897f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_873_n N_A_1108_47#_c_1342_n 0.00621195f $X=7.045 $Y=0.85
+ $X2=0 $Y2=0
cc_707 N_RESET_B_c_880_n N_A_1108_47#_c_1342_n 0.00451828f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_708 N_RESET_B_M1018_g N_A_1108_47#_c_1343_n 0.00180441f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_709 N_RESET_B_M1018_g N_A_1108_47#_c_1344_n 0.0144262f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_710 N_RESET_B_c_876_n N_A_1108_47#_c_1344_n 0.00392251f $X=7.19 $Y=1.165
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_879_n N_A_1108_47#_c_1344_n 6.25544e-19 $X=7.27 $Y=1.12 $X2=0
+ $Y2=0
cc_712 N_RESET_B_c_880_n N_A_1108_47#_c_1344_n 0.0397801f $X=7.525 $Y=1.22 $X2=0
+ $Y2=0
cc_713 N_RESET_B_M1018_g N_A_1108_47#_c_1345_n 0.0217285f $X=7.235 $Y=2.275
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_880_n N_A_1108_47#_c_1345_n 0.00253996f $X=7.525 $Y=1.22
+ $X2=0 $Y2=0
cc_715 N_RESET_B_M1031_g N_VPWR_c_1495_n 0.00862424f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_716 N_RESET_B_M1031_g N_VPWR_c_1496_n 0.00315462f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_717 N_RESET_B_M1018_g N_VPWR_c_1497_n 0.00837484f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_718 N_RESET_B_M1031_g N_VPWR_c_1507_n 0.00345093f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_719 N_RESET_B_M1031_g N_VPWR_c_1492_n 0.00519819f $X=4.365 $Y=2.275 $X2=0
+ $Y2=0
cc_720 N_RESET_B_M1018_g N_VPWR_c_1492_n 0.00799591f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_721 N_RESET_B_M1018_g N_VPWR_c_1513_n 0.0046653f $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_722 N_RESET_B_M1018_g N_VPWR_c_1514_n 7.28498e-19 $X=7.235 $Y=2.275 $X2=0
+ $Y2=0
cc_723 N_RESET_B_M1031_g N_A_651_413#_c_1683_n 0.0122302f $X=4.365 $Y=2.275
+ $X2=0 $Y2=0
cc_724 N_RESET_B_M1031_g N_A_651_413#_c_1685_n 0.00113125f $X=4.365 $Y=2.275
+ $X2=0 $Y2=0
cc_725 N_RESET_B_c_873_n N_VGND_M1004_d 0.0025426f $X=7.045 $Y=0.85 $X2=0 $Y2=0
cc_726 N_RESET_B_c_872_n N_VGND_c_1767_n 0.0066953f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_727 N_RESET_B_c_873_n N_VGND_c_1767_n 0.00423599f $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_728 N_RESET_B_c_877_n N_VGND_c_1767_n 6.55014e-19 $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_729 N_RESET_B_c_878_n N_VGND_c_1767_n 0.0117447f $X=4.37 $Y=0.765 $X2=0 $Y2=0
cc_730 N_RESET_B_M1005_g N_VGND_c_1768_n 0.00402543f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_731 N_RESET_B_c_873_n N_VGND_c_1768_n 8.29415e-19 $X=7.045 $Y=0.85 $X2=0
+ $Y2=0
cc_732 N_RESET_B_c_877_n N_VGND_c_1771_n 0.00162298f $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_733 N_RESET_B_c_878_n N_VGND_c_1771_n 0.00585385f $X=4.37 $Y=0.765 $X2=0
+ $Y2=0
cc_734 N_RESET_B_M1005_g N_VGND_c_1775_n 0.0036601f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_735 N_RESET_B_M1005_g N_VGND_c_1781_n 0.00599573f $X=7.235 $Y=0.445 $X2=0
+ $Y2=0
cc_736 N_RESET_B_c_871_n N_VGND_c_1781_n 0.0362506f $X=4.28 $Y=0.85 $X2=0 $Y2=0
cc_737 N_RESET_B_c_872_n N_VGND_c_1781_n 0.00772058f $X=4.25 $Y=0.85 $X2=0 $Y2=0
cc_738 N_RESET_B_c_873_n N_VGND_c_1781_n 0.139055f $X=7.045 $Y=0.85 $X2=0 $Y2=0
cc_739 N_RESET_B_c_875_n N_VGND_c_1781_n 0.0148902f $X=7.19 $Y=0.965 $X2=0 $Y2=0
cc_740 N_RESET_B_c_877_n N_VGND_c_1781_n 0.00136687f $X=4.37 $Y=0.93 $X2=0 $Y2=0
cc_741 N_RESET_B_c_878_n N_VGND_c_1781_n 0.00606683f $X=4.37 $Y=0.765 $X2=0
+ $Y2=0
cc_742 RESET_B A_1462_47# 0.00176151f $X=7.405 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_743 N_A_543_47#_c_1029_n N_VPWR_c_1496_n 0.0111275f $X=5.35 $Y=1.57 $X2=0
+ $Y2=0
cc_744 N_A_543_47#_c_1027_n N_VPWR_c_1496_n 0.00129214f $X=4.85 $Y=1.17 $X2=0
+ $Y2=0
cc_745 N_A_543_47#_c_1037_n N_VPWR_c_1499_n 0.0397779f $X=3.245 $Y=2.3 $X2=0
+ $Y2=0
cc_746 N_A_543_47#_c_1029_n N_VPWR_c_1501_n 0.00290206f $X=5.35 $Y=1.57 $X2=0
+ $Y2=0
cc_747 N_A_543_47#_M1030_d N_VPWR_c_1492_n 0.00221211f $X=2.76 $Y=2.065 $X2=0
+ $Y2=0
cc_748 N_A_543_47#_c_1029_n N_VPWR_c_1492_n 0.00346038f $X=5.35 $Y=1.57 $X2=0
+ $Y2=0
cc_749 N_A_543_47#_c_1037_n N_VPWR_c_1492_n 0.0114478f $X=3.245 $Y=2.3 $X2=0
+ $Y2=0
cc_750 N_A_543_47#_c_1037_n N_A_448_47#_c_1648_n 0.0221744f $X=3.245 $Y=2.3
+ $X2=0 $Y2=0
cc_751 N_A_543_47#_c_1037_n N_A_651_413#_M1007_d 0.00470561f $X=3.245 $Y=2.3
+ $X2=-0.19 $Y2=-0.24
cc_752 N_A_543_47#_c_1030_n N_A_651_413#_M1007_d 6.28858e-19 $X=3.33 $Y=2.135
+ $X2=-0.19 $Y2=-0.24
cc_753 N_A_543_47#_c_1037_n N_A_651_413#_c_1682_n 0.019526f $X=3.245 $Y=2.3
+ $X2=0 $Y2=0
cc_754 N_A_543_47#_c_1030_n N_A_651_413#_c_1682_n 0.00726918f $X=3.33 $Y=2.135
+ $X2=0 $Y2=0
cc_755 N_A_543_47#_c_1029_n N_A_651_413#_c_1683_n 0.00137742f $X=5.35 $Y=1.57
+ $X2=0 $Y2=0
cc_756 N_A_543_47#_c_1024_n N_A_651_413#_c_1683_n 4.0432e-19 $X=4.765 $Y=1.27
+ $X2=0 $Y2=0
cc_757 N_A_543_47#_c_1030_n N_A_651_413#_c_1684_n 0.0132883f $X=3.33 $Y=2.135
+ $X2=0 $Y2=0
cc_758 N_A_543_47#_c_1025_n N_A_651_413#_c_1684_n 0.0035943f $X=3.6 $Y=1.27
+ $X2=0 $Y2=0
cc_759 N_A_543_47#_c_1029_n N_A_651_413#_c_1685_n 0.00269162f $X=5.35 $Y=1.57
+ $X2=0 $Y2=0
cc_760 N_A_543_47#_M1022_g N_VGND_c_1767_n 0.00677972f $X=4.97 $Y=0.555 $X2=0
+ $Y2=0
cc_761 N_A_543_47#_c_1024_n N_VGND_c_1767_n 0.00223331f $X=4.765 $Y=1.27 $X2=0
+ $Y2=0
cc_762 N_A_543_47#_c_1026_n N_VGND_c_1767_n 6.77929e-19 $X=4.85 $Y=1.17 $X2=0
+ $Y2=0
cc_763 N_A_543_47#_c_1027_n N_VGND_c_1767_n 0.001314f $X=4.85 $Y=1.17 $X2=0
+ $Y2=0
cc_764 N_A_543_47#_c_1058_n N_VGND_c_1771_n 0.0387784f $X=3.43 $Y=0.39 $X2=0
+ $Y2=0
cc_765 N_A_543_47#_M1022_g N_VGND_c_1773_n 0.00542163f $X=4.97 $Y=0.555 $X2=0
+ $Y2=0
cc_766 N_A_543_47#_M1009_d N_VGND_c_1781_n 0.00309942f $X=2.715 $Y=0.235 $X2=0
+ $Y2=0
cc_767 N_A_543_47#_M1022_g N_VGND_c_1781_n 0.00686855f $X=4.97 $Y=0.555 $X2=0
+ $Y2=0
cc_768 N_A_543_47#_c_1058_n N_VGND_c_1781_n 0.0303432f $X=3.43 $Y=0.39 $X2=0
+ $Y2=0
cc_769 N_A_543_47#_c_1058_n A_639_47# 0.0148617f $X=3.43 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_770 N_A_543_47#_c_1023_n A_639_47# 0.00606072f $X=3.515 $Y=1.185 $X2=-0.19
+ $Y2=-0.24
cc_771 N_A_1283_21#_M1011_g N_A_1108_47#_M1016_g 0.00535021f $X=8.475 $Y=1.985
+ $X2=0 $Y2=0
cc_772 N_A_1283_21#_c_1172_n N_A_1108_47#_M1016_g 0.0120138f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_773 N_A_1283_21#_c_1174_n N_A_1108_47#_M1016_g 0.00192548f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_774 N_A_1283_21#_M1011_g N_A_1108_47#_M1001_g 0.00177448f $X=8.475 $Y=1.985
+ $X2=0 $Y2=0
cc_775 N_A_1283_21#_c_1155_n N_A_1108_47#_M1001_g 0.013342f $X=8.4 $Y=1.16 $X2=0
+ $Y2=0
cc_776 N_A_1283_21#_c_1157_n N_A_1108_47#_M1001_g 6.19895e-19 $X=7.15 $Y=0.695
+ $X2=0 $Y2=0
cc_777 N_A_1283_21#_c_1200_n N_A_1108_47#_M1001_g 0.0116638f $X=7.815 $Y=0.38
+ $X2=0 $Y2=0
cc_778 N_A_1283_21#_c_1159_n N_A_1108_47#_M1001_g 0.0037075f $X=7.975 $Y=0.82
+ $X2=0 $Y2=0
cc_779 N_A_1283_21#_c_1174_n N_A_1108_47#_M1001_g 0.00279337f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_780 N_A_1283_21#_c_1161_n N_A_1108_47#_M1001_g 0.0066004f $X=8.075 $Y=1.072
+ $X2=0 $Y2=0
cc_781 N_A_1283_21#_M1026_g N_A_1108_47#_c_1346_n 0.00955366f $X=6.49 $Y=0.445
+ $X2=0 $Y2=0
cc_782 N_A_1283_21#_c_1157_n N_A_1108_47#_c_1346_n 3.21819e-19 $X=7.15 $Y=0.695
+ $X2=0 $Y2=0
cc_783 N_A_1283_21#_M1008_g N_A_1108_47#_c_1349_n 0.0102686f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_784 N_A_1283_21#_M1026_g N_A_1108_47#_c_1339_n 0.00739655f $X=6.49 $Y=0.445
+ $X2=0 $Y2=0
cc_785 N_A_1283_21#_c_1156_n N_A_1108_47#_c_1339_n 0.0190293f $X=6.79 $Y=0.98
+ $X2=0 $Y2=0
cc_786 N_A_1283_21#_c_1157_n N_A_1108_47#_c_1339_n 0.00468097f $X=7.15 $Y=0.695
+ $X2=0 $Y2=0
cc_787 N_A_1283_21#_c_1160_n N_A_1108_47#_c_1339_n 0.0122822f $X=7.15 $Y=0.78
+ $X2=0 $Y2=0
cc_788 N_A_1283_21#_c_1162_n N_A_1108_47#_c_1339_n 0.0104269f $X=6.695 $Y=0.98
+ $X2=0 $Y2=0
cc_789 N_A_1283_21#_M1008_g N_A_1108_47#_c_1342_n 0.0164997f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_790 N_A_1283_21#_c_1156_n N_A_1108_47#_c_1342_n 0.00480564f $X=6.79 $Y=0.98
+ $X2=0 $Y2=0
cc_791 N_A_1283_21#_c_1162_n N_A_1108_47#_c_1342_n 0.00270124f $X=6.695 $Y=0.98
+ $X2=0 $Y2=0
cc_792 N_A_1283_21#_M1008_g N_A_1108_47#_c_1343_n 0.0114588f $X=6.695 $Y=2.275
+ $X2=0 $Y2=0
cc_793 N_A_1283_21#_c_1173_n N_A_1108_47#_c_1343_n 0.00493675f $X=7.53 $Y=2
+ $X2=0 $Y2=0
cc_794 N_A_1283_21#_c_1156_n N_A_1108_47#_c_1344_n 0.00570594f $X=6.79 $Y=0.98
+ $X2=0 $Y2=0
cc_795 N_A_1283_21#_c_1172_n N_A_1108_47#_c_1344_n 0.0202553f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_796 N_A_1283_21#_c_1173_n N_A_1108_47#_c_1344_n 0.0138731f $X=7.53 $Y=2 $X2=0
+ $Y2=0
cc_797 N_A_1283_21#_c_1174_n N_A_1108_47#_c_1344_n 0.0141871f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_798 N_A_1283_21#_c_1161_n N_A_1108_47#_c_1344_n 2.98117e-19 $X=8.075 $Y=1.072
+ $X2=0 $Y2=0
cc_799 N_A_1283_21#_c_1162_n N_A_1108_47#_c_1344_n 8.76062e-19 $X=6.695 $Y=0.98
+ $X2=0 $Y2=0
cc_800 N_A_1283_21#_M1011_g N_A_1108_47#_c_1345_n 0.00394467f $X=8.475 $Y=1.985
+ $X2=0 $Y2=0
cc_801 N_A_1283_21#_c_1172_n N_A_1108_47#_c_1345_n 0.00285904f $X=7.99 $Y=2
+ $X2=0 $Y2=0
cc_802 N_A_1283_21#_c_1173_n N_A_1108_47#_c_1345_n 2.53623e-19 $X=7.53 $Y=2
+ $X2=0 $Y2=0
cc_803 N_A_1283_21#_c_1174_n N_A_1108_47#_c_1345_n 0.00447201f $X=8.075 $Y=1.915
+ $X2=0 $Y2=0
cc_804 N_A_1283_21#_c_1170_n N_A_1847_47#_M1013_g 0.00475126f $X=9.542 $Y=1.515
+ $X2=0 $Y2=0
cc_805 N_A_1283_21#_c_1171_n N_A_1847_47#_M1013_g 0.0187208f $X=9.542 $Y=1.665
+ $X2=0 $Y2=0
cc_806 N_A_1283_21#_c_1150_n N_A_1847_47#_c_1444_n 0.00121302f $X=8.63 $Y=0.995
+ $X2=0 $Y2=0
cc_807 N_A_1283_21#_c_1153_n N_A_1847_47#_c_1444_n 0.00985065f $X=9.515 $Y=1.325
+ $X2=0 $Y2=0
cc_808 N_A_1283_21#_c_1154_n N_A_1847_47#_c_1444_n 0.00263294f $X=9.57 $Y=0.73
+ $X2=0 $Y2=0
cc_809 N_A_1283_21#_M1024_g N_A_1847_47#_c_1449_n 0.0130372f $X=9.57 $Y=2.165
+ $X2=0 $Y2=0
cc_810 N_A_1283_21#_c_1170_n N_A_1847_47#_c_1449_n 0.0080198f $X=9.542 $Y=1.515
+ $X2=0 $Y2=0
cc_811 N_A_1283_21#_c_1171_n N_A_1847_47#_c_1449_n 0.00686175f $X=9.542 $Y=1.665
+ $X2=0 $Y2=0
cc_812 N_A_1283_21#_c_1153_n N_A_1847_47#_c_1445_n 0.0133342f $X=9.515 $Y=1.325
+ $X2=0 $Y2=0
cc_813 N_A_1283_21#_c_1171_n N_A_1847_47#_c_1445_n 0.00159098f $X=9.542 $Y=1.665
+ $X2=0 $Y2=0
cc_814 N_A_1283_21#_c_1153_n N_A_1847_47#_c_1446_n 0.0177772f $X=9.515 $Y=1.325
+ $X2=0 $Y2=0
cc_815 N_A_1283_21#_c_1151_n N_A_1847_47#_c_1463_n 0.0200944f $X=9.44 $Y=1.16
+ $X2=0 $Y2=0
cc_816 N_A_1283_21#_c_1153_n N_A_1847_47#_c_1463_n 0.00652717f $X=9.515 $Y=1.325
+ $X2=0 $Y2=0
cc_817 N_A_1283_21#_c_1153_n N_A_1847_47#_c_1447_n 0.00324727f $X=9.515 $Y=1.325
+ $X2=0 $Y2=0
cc_818 N_A_1283_21#_c_1154_n N_A_1847_47#_c_1447_n 0.0191731f $X=9.57 $Y=0.73
+ $X2=0 $Y2=0
cc_819 N_A_1283_21#_c_1172_n N_VPWR_M1016_d 0.00650738f $X=7.99 $Y=2 $X2=0 $Y2=0
cc_820 N_A_1283_21#_c_1174_n N_VPWR_M1016_d 0.00570121f $X=8.075 $Y=1.915 $X2=0
+ $Y2=0
cc_821 N_A_1283_21#_M1008_g N_VPWR_c_1497_n 0.00383525f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_822 N_A_1283_21#_c_1171_n N_VPWR_c_1498_n 0.0107735f $X=9.542 $Y=1.665 $X2=0
+ $Y2=0
cc_823 N_A_1283_21#_M1008_g N_VPWR_c_1501_n 0.00357668f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_824 N_A_1283_21#_M1011_g N_VPWR_c_1503_n 0.0046653f $X=8.475 $Y=1.985 $X2=0
+ $Y2=0
cc_825 N_A_1283_21#_M1024_g N_VPWR_c_1503_n 0.00542953f $X=9.57 $Y=2.165 $X2=0
+ $Y2=0
cc_826 N_A_1283_21#_M1018_d N_VPWR_c_1492_n 0.00416801f $X=7.31 $Y=2.065 $X2=0
+ $Y2=0
cc_827 N_A_1283_21#_M1008_g N_VPWR_c_1492_n 0.00559732f $X=6.695 $Y=2.275 $X2=0
+ $Y2=0
cc_828 N_A_1283_21#_M1011_g N_VPWR_c_1492_n 0.00916934f $X=8.475 $Y=1.985 $X2=0
+ $Y2=0
cc_829 N_A_1283_21#_M1024_g N_VPWR_c_1492_n 0.0112147f $X=9.57 $Y=2.165 $X2=0
+ $Y2=0
cc_830 N_A_1283_21#_c_1284_p N_VPWR_c_1492_n 0.00608739f $X=7.445 $Y=2.21 $X2=0
+ $Y2=0
cc_831 N_A_1283_21#_c_1172_n N_VPWR_c_1492_n 0.00652875f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_832 N_A_1283_21#_c_1284_p N_VPWR_c_1513_n 0.00701792f $X=7.445 $Y=2.21 $X2=0
+ $Y2=0
cc_833 N_A_1283_21#_c_1172_n N_VPWR_c_1513_n 0.00260015f $X=7.99 $Y=2 $X2=0
+ $Y2=0
cc_834 N_A_1283_21#_M1011_g N_VPWR_c_1514_n 0.0106278f $X=8.475 $Y=1.985 $X2=0
+ $Y2=0
cc_835 N_A_1283_21#_c_1172_n N_VPWR_c_1514_n 0.0309612f $X=7.99 $Y=2 $X2=0 $Y2=0
cc_836 N_A_1283_21#_M1024_g N_Q_c_1721_n 0.00167298f $X=9.57 $Y=2.165 $X2=0
+ $Y2=0
cc_837 N_A_1283_21#_M1011_g N_Q_c_1722_n 8.05623e-19 $X=8.475 $Y=1.985 $X2=0
+ $Y2=0
cc_838 N_A_1283_21#_c_1152_n N_Q_c_1722_n 0.00176856f $X=8.705 $Y=1.16 $X2=0
+ $Y2=0
cc_839 N_A_1283_21#_c_1171_n N_Q_c_1722_n 7.40758e-19 $X=9.542 $Y=1.665 $X2=0
+ $Y2=0
cc_840 N_A_1283_21#_c_1174_n N_Q_c_1722_n 0.00893991f $X=8.075 $Y=1.915 $X2=0
+ $Y2=0
cc_841 N_A_1283_21#_M1011_g N_Q_c_1720_n 0.00323657f $X=8.475 $Y=1.985 $X2=0
+ $Y2=0
cc_842 N_A_1283_21#_c_1150_n N_Q_c_1720_n 0.012358f $X=8.63 $Y=0.995 $X2=0 $Y2=0
cc_843 N_A_1283_21#_c_1151_n N_Q_c_1720_n 0.0266971f $X=9.44 $Y=1.16 $X2=0 $Y2=0
cc_844 N_A_1283_21#_c_1152_n N_Q_c_1720_n 0.0072045f $X=8.705 $Y=1.16 $X2=0
+ $Y2=0
cc_845 N_A_1283_21#_c_1153_n N_Q_c_1720_n 0.00115744f $X=9.515 $Y=1.325 $X2=0
+ $Y2=0
cc_846 N_A_1283_21#_c_1154_n N_Q_c_1720_n 0.00209756f $X=9.57 $Y=0.73 $X2=0
+ $Y2=0
cc_847 N_A_1283_21#_c_1170_n N_Q_c_1720_n 7.40758e-19 $X=9.542 $Y=1.515 $X2=0
+ $Y2=0
cc_848 N_A_1283_21#_c_1159_n N_Q_c_1720_n 0.00163683f $X=7.975 $Y=0.82 $X2=0
+ $Y2=0
cc_849 N_A_1283_21#_c_1174_n N_Q_c_1720_n 0.00471114f $X=8.075 $Y=1.915 $X2=0
+ $Y2=0
cc_850 N_A_1283_21#_c_1161_n N_Q_c_1720_n 0.0256177f $X=8.075 $Y=1.072 $X2=0
+ $Y2=0
cc_851 N_A_1283_21#_c_1157_n N_VGND_M1026_d 0.00259202f $X=7.15 $Y=0.695 $X2=0
+ $Y2=0
cc_852 N_A_1283_21#_c_1205_n N_VGND_M1026_d 0.0020638f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_853 N_A_1283_21#_M1026_g N_VGND_c_1768_n 0.00552213f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_854 N_A_1283_21#_c_1157_n N_VGND_c_1768_n 0.0043583f $X=7.15 $Y=0.695 $X2=0
+ $Y2=0
cc_855 N_A_1283_21#_c_1205_n N_VGND_c_1768_n 0.0139352f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_856 N_A_1283_21#_c_1160_n N_VGND_c_1768_n 0.0135486f $X=7.15 $Y=0.78 $X2=0
+ $Y2=0
cc_857 N_A_1283_21#_c_1162_n N_VGND_c_1768_n 0.00108751f $X=6.695 $Y=0.98 $X2=0
+ $Y2=0
cc_858 N_A_1283_21#_c_1150_n N_VGND_c_1769_n 0.00716592f $X=8.63 $Y=0.995 $X2=0
+ $Y2=0
cc_859 N_A_1283_21#_c_1152_n N_VGND_c_1769_n 0.00300999f $X=8.705 $Y=1.16 $X2=0
+ $Y2=0
cc_860 N_A_1283_21#_c_1155_n N_VGND_c_1769_n 7.50078e-19 $X=8.4 $Y=1.16 $X2=0
+ $Y2=0
cc_861 N_A_1283_21#_c_1158_n N_VGND_c_1769_n 0.0125643f $X=7.975 $Y=0.465 $X2=0
+ $Y2=0
cc_862 N_A_1283_21#_c_1159_n N_VGND_c_1769_n 0.021059f $X=7.975 $Y=0.82 $X2=0
+ $Y2=0
cc_863 N_A_1283_21#_c_1161_n N_VGND_c_1769_n 0.0065826f $X=8.075 $Y=1.072 $X2=0
+ $Y2=0
cc_864 N_A_1283_21#_c_1154_n N_VGND_c_1770_n 0.00779477f $X=9.57 $Y=0.73 $X2=0
+ $Y2=0
cc_865 N_A_1283_21#_M1026_g N_VGND_c_1773_n 0.00403211f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_866 N_A_1283_21#_c_1200_n N_VGND_c_1775_n 0.0253037f $X=7.815 $Y=0.38 $X2=0
+ $Y2=0
cc_867 N_A_1283_21#_c_1205_n N_VGND_c_1775_n 0.00758764f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_868 N_A_1283_21#_c_1158_n N_VGND_c_1775_n 0.0178412f $X=7.975 $Y=0.465 $X2=0
+ $Y2=0
cc_869 N_A_1283_21#_c_1160_n N_VGND_c_1775_n 0.00275249f $X=7.15 $Y=0.78 $X2=0
+ $Y2=0
cc_870 N_A_1283_21#_c_1150_n N_VGND_c_1777_n 0.00542163f $X=8.63 $Y=0.995 $X2=0
+ $Y2=0
cc_871 N_A_1283_21#_c_1153_n N_VGND_c_1777_n 0.00105583f $X=9.515 $Y=1.325 $X2=0
+ $Y2=0
cc_872 N_A_1283_21#_c_1154_n N_VGND_c_1777_n 0.00585385f $X=9.57 $Y=0.73 $X2=0
+ $Y2=0
cc_873 N_A_1283_21#_M1001_d N_VGND_c_1781_n 0.00212393f $X=7.765 $Y=0.235 $X2=0
+ $Y2=0
cc_874 N_A_1283_21#_M1026_g N_VGND_c_1781_n 0.00628912f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_875 N_A_1283_21#_c_1150_n N_VGND_c_1781_n 0.0122813f $X=8.63 $Y=0.995 $X2=0
+ $Y2=0
cc_876 N_A_1283_21#_c_1153_n N_VGND_c_1781_n 0.00138273f $X=9.515 $Y=1.325 $X2=0
+ $Y2=0
cc_877 N_A_1283_21#_c_1154_n N_VGND_c_1781_n 0.0123744f $X=9.57 $Y=0.73 $X2=0
+ $Y2=0
cc_878 N_A_1283_21#_c_1200_n N_VGND_c_1781_n 0.012114f $X=7.815 $Y=0.38 $X2=0
+ $Y2=0
cc_879 N_A_1283_21#_c_1205_n N_VGND_c_1781_n 0.00279545f $X=7.235 $Y=0.38 $X2=0
+ $Y2=0
cc_880 N_A_1283_21#_c_1158_n N_VGND_c_1781_n 0.0120802f $X=7.975 $Y=0.465 $X2=0
+ $Y2=0
cc_881 N_A_1283_21#_c_1160_n N_VGND_c_1781_n 0.00245528f $X=7.15 $Y=0.78 $X2=0
+ $Y2=0
cc_882 N_A_1283_21#_c_1162_n N_VGND_c_1781_n 8.11688e-19 $X=6.695 $Y=0.98 $X2=0
+ $Y2=0
cc_883 N_A_1283_21#_c_1200_n A_1462_47# 0.00399694f $X=7.815 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_884 N_A_1108_47#_M1016_g N_VPWR_c_1497_n 7.44815e-19 $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_885 N_A_1108_47#_c_1349_n N_VPWR_c_1497_n 0.0234228f $X=6.6 $Y=2.295 $X2=0
+ $Y2=0
cc_886 N_A_1108_47#_c_1344_n N_VPWR_c_1497_n 0.00898242f $X=7.655 $Y=1.66 $X2=0
+ $Y2=0
cc_887 N_A_1108_47#_c_1349_n N_VPWR_c_1501_n 0.0505746f $X=6.6 $Y=2.295 $X2=0
+ $Y2=0
cc_888 N_A_1108_47#_M1025_d N_VPWR_c_1492_n 0.00178215f $X=5.92 $Y=2.065 $X2=0
+ $Y2=0
cc_889 N_A_1108_47#_M1016_g N_VPWR_c_1492_n 0.00428496f $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_890 N_A_1108_47#_c_1349_n N_VPWR_c_1492_n 0.0242715f $X=6.6 $Y=2.295 $X2=0
+ $Y2=0
cc_891 N_A_1108_47#_M1016_g N_VPWR_c_1513_n 0.00367706f $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_892 N_A_1108_47#_M1016_g N_VPWR_c_1514_n 0.00793125f $X=7.655 $Y=2.275 $X2=0
+ $Y2=0
cc_893 N_A_1108_47#_c_1349_n A_1270_413# 0.00433468f $X=6.6 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_894 N_A_1108_47#_c_1346_n N_VGND_c_1768_n 0.0213874f $X=6.365 $Y=0.395 $X2=0
+ $Y2=0
cc_895 N_A_1108_47#_M1001_g N_VGND_c_1769_n 0.00271669f $X=7.69 $Y=0.445 $X2=0
+ $Y2=0
cc_896 N_A_1108_47#_c_1346_n N_VGND_c_1773_n 0.0567494f $X=6.365 $Y=0.395 $X2=0
+ $Y2=0
cc_897 N_A_1108_47#_M1001_g N_VGND_c_1775_n 0.00366111f $X=7.69 $Y=0.445 $X2=0
+ $Y2=0
cc_898 N_A_1108_47#_M1023_d N_VGND_c_1781_n 0.00272411f $X=5.54 $Y=0.235 $X2=0
+ $Y2=0
cc_899 N_A_1108_47#_M1001_g N_VGND_c_1781_n 0.00675738f $X=7.69 $Y=0.445 $X2=0
+ $Y2=0
cc_900 N_A_1108_47#_c_1346_n N_VGND_c_1781_n 0.0161501f $X=6.365 $Y=0.395 $X2=0
+ $Y2=0
cc_901 N_A_1108_47#_c_1346_n A_1217_47# 0.00484766f $X=6.365 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_902 N_A_1847_47#_M1013_g N_VPWR_c_1498_n 0.00278284f $X=10.055 $Y=1.985 $X2=0
+ $Y2=0
cc_903 N_A_1847_47#_c_1449_n N_VPWR_c_1498_n 0.0534728f $X=9.36 $Y=2 $X2=0 $Y2=0
cc_904 N_A_1847_47#_c_1445_n N_VPWR_c_1498_n 0.0139084f $X=9.97 $Y=1.16 $X2=0
+ $Y2=0
cc_905 N_A_1847_47#_c_1446_n N_VPWR_c_1498_n 0.00217151f $X=9.97 $Y=1.16 $X2=0
+ $Y2=0
cc_906 N_A_1847_47#_c_1449_n N_VPWR_c_1503_n 0.016757f $X=9.36 $Y=2 $X2=0 $Y2=0
cc_907 N_A_1847_47#_M1013_g N_VPWR_c_1508_n 0.00585385f $X=10.055 $Y=1.985 $X2=0
+ $Y2=0
cc_908 N_A_1847_47#_M1024_s N_VPWR_c_1492_n 0.00211564f $X=9.235 $Y=1.845 $X2=0
+ $Y2=0
cc_909 N_A_1847_47#_M1013_g N_VPWR_c_1492_n 0.0118334f $X=10.055 $Y=1.985 $X2=0
+ $Y2=0
cc_910 N_A_1847_47#_c_1449_n N_VPWR_c_1492_n 0.0121755f $X=9.36 $Y=2 $X2=0 $Y2=0
cc_911 N_A_1847_47#_c_1444_n N_Q_c_1720_n 0.0489841f $X=9.36 $Y=0.51 $X2=0 $Y2=0
cc_912 N_A_1847_47#_c_1449_n N_Q_c_1720_n 0.0857608f $X=9.36 $Y=2 $X2=0 $Y2=0
cc_913 N_A_1847_47#_c_1463_n N_Q_c_1720_n 0.024084f $X=9.36 $Y=1.16 $X2=0 $Y2=0
cc_914 N_A_1847_47#_M1013_g N_Q_N_c_1751_n 0.00384193f $X=10.055 $Y=1.985 $X2=0
+ $Y2=0
cc_915 N_A_1847_47#_c_1449_n N_Q_N_c_1751_n 0.00120542f $X=9.36 $Y=2 $X2=0 $Y2=0
cc_916 N_A_1847_47#_c_1445_n Q_N 0.0266145f $X=9.97 $Y=1.16 $X2=0 $Y2=0
cc_917 N_A_1847_47#_c_1447_n Q_N 0.0195346f $X=9.982 $Y=0.995 $X2=0 $Y2=0
cc_918 N_A_1847_47#_c_1444_n N_VGND_c_1770_n 0.0083492f $X=9.36 $Y=0.51 $X2=0
+ $Y2=0
cc_919 N_A_1847_47#_c_1445_n N_VGND_c_1770_n 0.00878358f $X=9.97 $Y=1.16 $X2=0
+ $Y2=0
cc_920 N_A_1847_47#_c_1446_n N_VGND_c_1770_n 0.00198753f $X=9.97 $Y=1.16 $X2=0
+ $Y2=0
cc_921 N_A_1847_47#_c_1447_n N_VGND_c_1770_n 0.00305279f $X=9.982 $Y=0.995 $X2=0
+ $Y2=0
cc_922 N_A_1847_47#_c_1444_n N_VGND_c_1777_n 0.0109259f $X=9.36 $Y=0.51 $X2=0
+ $Y2=0
cc_923 N_A_1847_47#_c_1447_n N_VGND_c_1780_n 0.00585385f $X=9.982 $Y=0.995 $X2=0
+ $Y2=0
cc_924 N_A_1847_47#_M1006_s N_VGND_c_1781_n 0.00272276f $X=9.235 $Y=0.235 $X2=0
+ $Y2=0
cc_925 N_A_1847_47#_c_1444_n N_VGND_c_1781_n 0.00910216f $X=9.36 $Y=0.51 $X2=0
+ $Y2=0
cc_926 N_A_1847_47#_c_1447_n N_VGND_c_1781_n 0.0119159f $X=9.982 $Y=0.995 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1492_n N_A_448_47#_M1028_d 0.00255917f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1494_n N_A_448_47#_c_1648_n 0.00413503f $X=2.015 $Y=2.34 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1499_n N_A_448_47#_c_1648_n 0.0177638f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1492_n N_A_448_47#_c_1648_n 0.00643929f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1492_n N_A_651_413#_M1007_d 0.00515242f $X=10.35 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_932 N_VPWR_c_1492_n N_A_651_413#_M1031_d 0.00220707f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1499_n N_A_651_413#_c_1682_n 0.0071865f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1492_n N_A_651_413#_c_1682_n 0.00287341f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1495_n N_A_651_413#_c_1683_n 0.0205079f $X=4.155 $Y=2.29 $X2=0
+ $Y2=0
cc_936 N_VPWR_c_1499_n N_A_651_413#_c_1683_n 0.00357601f $X=3.99 $Y=2.72 $X2=0
+ $Y2=0
cc_937 N_VPWR_c_1507_n N_A_651_413#_c_1683_n 0.00256078f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1492_n N_A_651_413#_c_1683_n 0.00495172f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_939 N_VPWR_c_1496_n N_A_651_413#_c_1685_n 0.0106232f $X=5.14 $Y=2.34 $X2=0
+ $Y2=0
cc_940 N_VPWR_c_1507_n N_A_651_413#_c_1685_n 0.0071865f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1492_n N_A_651_413#_c_1685_n 0.00287341f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_942 N_VPWR_c_1492_n A_1270_413# 0.00216831f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_943 N_VPWR_c_1492_n N_Q_M1011_d 0.00399293f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_944 N_VPWR_c_1503_n N_Q_c_1721_n 0.0283694f $X=9.76 $Y=2.72 $X2=0 $Y2=0
cc_945 N_VPWR_c_1492_n N_Q_c_1721_n 0.0155202f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_946 N_VPWR_c_1492_n N_Q_N_M1013_d 0.00401809f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_947 N_VPWR_c_1508_n N_Q_N_c_1752_n 0.00923202f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_948 N_VPWR_c_1492_n N_Q_N_c_1752_n 0.00900352f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_949 N_A_448_47#_c_1665_n N_VGND_c_1771_n 0.00763796f $X=2.215 $Y=0.39 $X2=0
+ $Y2=0
cc_950 N_A_448_47#_c_1656_n N_VGND_c_1771_n 0.0137117f $X=2.375 $Y=0.39 $X2=0
+ $Y2=0
cc_951 N_A_448_47#_M1029_d N_VGND_c_1781_n 0.00276506f $X=2.24 $Y=0.235 $X2=0
+ $Y2=0
cc_952 N_A_448_47#_c_1665_n N_VGND_c_1781_n 0.00579413f $X=2.215 $Y=0.39 $X2=0
+ $Y2=0
cc_953 N_A_448_47#_c_1656_n N_VGND_c_1781_n 0.0115463f $X=2.375 $Y=0.39 $X2=0
+ $Y2=0
cc_954 N_Q_c_1720_n N_VGND_c_1777_n 0.0186592f $X=8.84 $Y=0.4 $X2=0 $Y2=0
cc_955 N_Q_M1019_d N_VGND_c_1781_n 0.00210124f $X=8.705 $Y=0.235 $X2=0 $Y2=0
cc_956 N_Q_c_1720_n N_VGND_c_1781_n 0.0123045f $X=8.84 $Y=0.4 $X2=0 $Y2=0
cc_957 N_Q_N_c_1748_n N_VGND_c_1780_n 0.0165374f $X=10.307 $Y=0.668 $X2=0 $Y2=0
cc_958 N_Q_N_M1002_d N_VGND_c_1781_n 0.00387432f $X=10.13 $Y=0.235 $X2=0 $Y2=0
cc_959 N_Q_N_c_1748_n N_VGND_c_1781_n 0.00968619f $X=10.307 $Y=0.668 $X2=0 $Y2=0
cc_960 N_VGND_c_1781_n A_639_47# 0.0110359f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_961 N_VGND_c_1781_n A_805_47# 0.00196925f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_962 N_VGND_c_1781_n A_1217_47# 0.00217995f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24
cc_963 N_VGND_c_1781_n A_1462_47# 0.00196947f $X=10.35 $Y=0 $X2=-0.19 $Y2=-0.24

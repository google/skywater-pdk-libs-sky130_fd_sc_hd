* File: sky130_fd_sc_hd__o2111a_1.pxi.spice
* Created: Tue Sep  1 19:19:51 2020
* 
x_PM_SKY130_FD_SC_HD__O2111A_1%A_79_21# N_A_79_21#_M1004_s N_A_79_21#_M1008_d
+ N_A_79_21#_M1006_d N_A_79_21#_M1011_g N_A_79_21#_M1010_g N_A_79_21#_c_70_n
+ N_A_79_21#_c_74_p N_A_79_21#_c_101_p N_A_79_21#_c_65_n N_A_79_21#_c_86_p
+ N_A_79_21#_c_87_p N_A_79_21#_c_66_n N_A_79_21#_c_67_n N_A_79_21#_c_81_p
+ N_A_79_21#_c_91_p N_A_79_21#_c_68_n PM_SKY130_FD_SC_HD__O2111A_1%A_79_21#
x_PM_SKY130_FD_SC_HD__O2111A_1%D1 N_D1_M1008_g N_D1_M1004_g D1 D1 D1
+ N_D1_c_136_n N_D1_c_137_n PM_SKY130_FD_SC_HD__O2111A_1%D1
x_PM_SKY130_FD_SC_HD__O2111A_1%C1 N_C1_M1005_g N_C1_M1002_g C1 C1 C1
+ N_C1_c_176_n PM_SKY130_FD_SC_HD__O2111A_1%C1
x_PM_SKY130_FD_SC_HD__O2111A_1%B1 N_B1_M1001_g N_B1_M1006_g B1 B1 B1
+ N_B1_c_213_n N_B1_c_214_n PM_SKY130_FD_SC_HD__O2111A_1%B1
x_PM_SKY130_FD_SC_HD__O2111A_1%A2 N_A2_M1007_g N_A2_M1000_g N_A2_c_253_n
+ N_A2_c_254_n A2 A2 A2 A2 N_A2_c_255_n PM_SKY130_FD_SC_HD__O2111A_1%A2
x_PM_SKY130_FD_SC_HD__O2111A_1%A1 N_A1_M1009_g N_A1_M1003_g A1 A1 N_A1_c_296_n
+ PM_SKY130_FD_SC_HD__O2111A_1%A1
x_PM_SKY130_FD_SC_HD__O2111A_1%X N_X_M1011_s N_X_M1010_s X X X X X X N_X_c_320_n
+ PM_SKY130_FD_SC_HD__O2111A_1%X
x_PM_SKY130_FD_SC_HD__O2111A_1%VPWR N_VPWR_M1010_d N_VPWR_M1002_d N_VPWR_M1003_d
+ N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n VPWR
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_331_n
+ PM_SKY130_FD_SC_HD__O2111A_1%VPWR
x_PM_SKY130_FD_SC_HD__O2111A_1%VGND N_VGND_M1011_d N_VGND_M1007_d N_VGND_c_390_n
+ N_VGND_c_391_n VGND N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n
+ N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n PM_SKY130_FD_SC_HD__O2111A_1%VGND
x_PM_SKY130_FD_SC_HD__O2111A_1%A_512_47# N_A_512_47#_M1001_d N_A_512_47#_M1009_d
+ N_A_512_47#_c_454_n N_A_512_47#_c_449_n N_A_512_47#_c_451_n
+ N_A_512_47#_c_450_n PM_SKY130_FD_SC_HD__O2111A_1%A_512_47#
cc_1 VNB N_A_79_21#_c_65_n 0.00554217f $X=-0.19 $Y=-0.24 $X2=1.2 $Y2=0.38
cc_2 VNB N_A_79_21#_c_66_n 0.0308748f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.16
cc_3 VNB N_A_79_21#_c_67_n 0.017721f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.115
cc_4 VNB N_A_79_21#_c_68_n 0.021625f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=0.995
cc_5 VNB N_D1_M1008_g 5.04987e-19 $X=-0.19 $Y=-0.24 $X2=2.805 $Y2=1.485
cc_6 VNB N_D1_M1004_g 0.0228397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB D1 0.00282647f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_D1_c_136_n 0.0292438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_D1_c_137_n 0.00412398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_C1_M1005_g 0.0190817f $X=-0.19 $Y=-0.24 $X2=2.805 $Y2=1.485
cc_11 VNB N_C1_M1002_g 5.59567e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB C1 0.00106266f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_C1_c_176_n 0.0298367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B1_M1001_g 0.0207464f $X=-0.19 $Y=-0.24 $X2=2.805 $Y2=1.485
cc_15 VNB N_B1_M1006_g 5.58651e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB B1 0.00143634f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B1_c_213_n 9.92772e-19 $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=1.58
cc_18 VNB N_B1_c_214_n 0.0373697f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.58
cc_19 VNB N_A2_M1007_g 0.0208339f $X=-0.19 $Y=-0.24 $X2=2.805 $Y2=1.485
cc_20 VNB N_A2_M1000_g 3.99901e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_253_n 0.00185733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_c_254_n 0.0255515f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_23 VNB N_A2_c_255_n 0.00288823f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.665
cc_24 VNB N_A1_M1009_g 0.0235892f $X=-0.19 $Y=-0.24 $X2=2.805 $Y2=1.485
cc_25 VNB N_A1_c_296_n 0.0407468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_320_n 0.045668f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=1.58
cc_27 VNB N_VPWR_c_331_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_390_n 0.00626006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_391_n 0.00258113f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_30 VNB N_VGND_c_392_n 0.0156941f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.325
cc_31 VNB N_VGND_c_393_n 0.0666005f $X=-0.19 $Y=-0.24 $X2=1.195 $Y2=0.38
cc_32 VNB N_VGND_c_394_n 0.0145038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_395_n 0.221966f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.115
cc_34 VNB N_VGND_c_396_n 0.00481106f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=1.115
cc_35 VNB N_VGND_c_397_n 0.0043067f $X=-0.19 $Y=-0.24 $X2=3.055 $Y2=1.58
cc_36 VNB N_A_512_47#_c_449_n 0.00818757f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_37 VNB N_A_512_47#_c_450_n 0.0174597f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_38 VPB N_A_79_21#_M1010_g 0.0245297f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB N_A_79_21#_c_70_n 0.00313924f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.495
cc_40 VPB N_A_79_21#_c_66_n 0.00730438f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.16
cc_41 VPB N_A_79_21#_c_67_n 0.00240564f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.115
cc_42 VPB N_D1_M1008_g 0.0251125f $X=-0.19 $Y=1.305 $X2=2.805 $Y2=1.485
cc_43 VPB N_D1_c_137_n 0.00335563f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_C1_M1002_g 0.0248137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB C1 0.00156017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_B1_M1006_g 0.0242351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_B1_c_213_n 0.00211829f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=1.58
cc_48 VPB N_A2_M1000_g 0.0199597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A2_c_253_n 0.00315506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB A2 9.15875e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_51 VPB N_A1_M1003_g 0.0230274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB A1 0.0136918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A1_c_296_n 0.00840754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_X_c_320_n 0.0466291f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=1.58
cc_55 VPB N_VPWR_c_332_n 0.0165811f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_56 VPB N_VPWR_c_333_n 0.00186974f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_57 VPB N_VPWR_c_334_n 0.0100134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_335_n 0.029168f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=1.495
cc_59 VPB N_VPWR_c_336_n 0.0153973f $X=-0.19 $Y=1.305 $X2=1.195 $Y2=0.38
cc_60 VPB N_VPWR_c_337_n 0.0248029f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.96
cc_61 VPB N_VPWR_c_338_n 0.0159475f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.115
cc_62 VPB N_VPWR_c_339_n 0.0113081f $X=-0.19 $Y=1.305 $X2=3.095 $Y2=1.66
cc_63 VPB N_VPWR_c_331_n 0.0436605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_70_n N_D1_M1008_g 0.00432957f $X=0.78 $Y=1.495 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_74_p N_D1_M1008_g 0.0169667f $X=1.505 $Y=1.58 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_66_n N_D1_M1008_g 4.58994e-19 $X=0.61 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_66_n N_D1_M1004_g 3.71634e-19 $X=0.61 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_67_n N_D1_M1004_g 0.00214201f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_67_n D1 0.00651521f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_66_n N_D1_c_136_n 0.00488976f $X=0.61 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_67_n N_D1_c_136_n 0.00414319f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_81_p N_D1_c_136_n 6.22126e-19 $X=1.67 $Y=1.58 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_74_p N_D1_c_137_n 0.0140703f $X=1.505 $Y=1.58 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_66_n N_D1_c_137_n 3.37508e-19 $X=0.61 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_67_n N_D1_c_137_n 0.0191063f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_81_p N_D1_c_137_n 0.019854f $X=1.67 $Y=1.58 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_86_p N_C1_M1002_g 0.0108806f $X=1.67 $Y=1.96 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_87_p N_C1_M1002_g 0.0172542f $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_87_p C1 0.0193718f $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_87_p N_C1_c_176_n 8.50787e-19 $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_87_p N_B1_M1006_g 0.0163853f $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_91_p N_B1_M1006_g 0.00920472f $X=3.095 $Y=1.66 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_87_p N_B1_c_213_n 0.0189658f $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_87_p N_B1_c_214_n 0.00267499f $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_91_p N_A2_c_253_n 0.0107317f $X=3.095 $Y=1.66 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_91_p N_A2_c_254_n 9.31119e-19 $X=3.095 $Y=1.66 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_70_n N_X_c_320_n 0.00782965f $X=0.78 $Y=1.495 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_67_n N_X_c_320_n 0.0352101f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_68_n N_X_c_320_n 0.0263298f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_70_n N_VPWR_M1010_d 2.31461e-19 $X=0.78 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_79_21#_c_74_p N_VPWR_M1010_d 0.0136956f $X=1.505 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_79_21#_c_101_p N_VPWR_M1010_d 0.00531074f $X=0.865 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_79_21#_c_87_p N_VPWR_M1002_d 0.0183245f $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_86_p N_VPWR_c_332_n 0.0226819f $X=1.67 $Y=1.96 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_86_p N_VPWR_c_333_n 0.0484077f $X=1.67 $Y=1.96 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_87_p N_VPWR_c_333_n 0.05002f $X=2.93 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_91_p N_VPWR_c_333_n 0.0506514f $X=3.095 $Y=1.66 $X2=0 $Y2=0
cc_98 N_A_79_21#_M1010_g N_VPWR_c_336_n 0.00507333f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_91_p N_VPWR_c_337_n 0.0172305f $X=3.095 $Y=1.66 $X2=0 $Y2=0
cc_100 N_A_79_21#_M1010_g N_VPWR_c_338_n 0.0139844f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_74_p N_VPWR_c_338_n 0.0333167f $X=1.505 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_101_p N_VPWR_c_338_n 0.0152373f $X=0.865 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_66_n N_VPWR_c_338_n 9.39525e-19 $X=0.61 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_67_n N_VPWR_c_338_n 0.00475199f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_105 N_A_79_21#_M1008_d N_VPWR_c_331_n 0.00722019f $X=1.46 $Y=1.485 $X2=0
+ $Y2=0
cc_106 N_A_79_21#_M1006_d N_VPWR_c_331_n 0.00954674f $X=2.805 $Y=1.485 $X2=0
+ $Y2=0
cc_107 N_A_79_21#_M1010_g N_VPWR_c_331_n 0.00946032f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_79_21#_c_86_p N_VPWR_c_331_n 0.0126319f $X=1.67 $Y=1.96 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_91_p N_VPWR_c_331_n 0.00955092f $X=3.095 $Y=1.66 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_67_n N_VGND_M1011_d 0.00339065f $X=0.78 $Y=1.115 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_79_21#_c_65_n N_VGND_c_390_n 0.0247334f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_66_n N_VGND_c_390_n 0.00100453f $X=0.61 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_67_n N_VGND_c_390_n 0.01813f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_68_n N_VGND_c_390_n 0.00939154f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_68_n N_VGND_c_392_n 0.00544582f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_65_n N_VGND_c_393_n 0.0223377f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_67_n N_VGND_c_393_n 0.0027257f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_118 N_A_79_21#_M1004_s N_VGND_c_395_n 0.00298283f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_119 N_A_79_21#_c_65_n N_VGND_c_395_n 0.0130015f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_67_n N_VGND_c_395_n 0.00543589f $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_68_n N_VGND_c_395_n 0.0100745f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_87_p N_A_512_47#_c_451_n 0.00181877f $X=2.93 $Y=1.58 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_c_91_p N_A_512_47#_c_451_n 0.00405147f $X=3.095 $Y=1.66 $X2=0
+ $Y2=0
cc_124 N_D1_M1004_g N_C1_M1005_g 0.0255411f $X=1.455 $Y=0.56 $X2=0 $Y2=0
cc_125 D1 N_C1_M1005_g 0.00438327f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_126 N_D1_M1008_g N_C1_M1002_g 0.0293793f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_127 N_D1_c_137_n N_C1_M1002_g 2.31097e-19 $X=1.64 $Y=1.2 $X2=0 $Y2=0
cc_128 D1 C1 0.0486467f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_129 N_D1_c_136_n C1 2.42476e-19 $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_130 N_D1_c_137_n C1 0.01916f $X=1.64 $Y=1.2 $X2=0 $Y2=0
cc_131 D1 N_C1_c_176_n 3.47908e-19 $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_132 N_D1_c_136_n N_C1_c_176_n 0.0121114f $X=1.43 $Y=1.16 $X2=0 $Y2=0
cc_133 N_D1_c_137_n N_C1_c_176_n 0.00164714f $X=1.64 $Y=1.2 $X2=0 $Y2=0
cc_134 N_D1_M1008_g N_VPWR_c_332_n 0.00487821f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_135 N_D1_M1008_g N_VPWR_c_333_n 0.00108643f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_136 N_D1_M1008_g N_VPWR_c_338_n 0.0136305f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_137 N_D1_M1008_g N_VPWR_c_331_n 0.00866926f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_138 N_D1_M1004_g N_VGND_c_390_n 0.00258869f $X=1.455 $Y=0.56 $X2=0 $Y2=0
cc_139 N_D1_M1004_g N_VGND_c_393_n 0.00585385f $X=1.455 $Y=0.56 $X2=0 $Y2=0
cc_140 D1 N_VGND_c_393_n 0.00688149f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_141 N_D1_M1004_g N_VGND_c_395_n 0.0123142f $X=1.455 $Y=0.56 $X2=0 $Y2=0
cc_142 D1 N_VGND_c_395_n 0.00742772f $X=1.535 $Y=0.425 $X2=0 $Y2=0
cc_143 D1 A_306_47# 0.0101938f $X=1.535 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_144 N_C1_M1005_g N_B1_M1001_g 0.0290299f $X=1.97 $Y=0.56 $X2=0 $Y2=0
cc_145 C1 N_B1_M1001_g 0.0044714f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_146 N_C1_M1002_g N_B1_M1006_g 0.0120241f $X=1.97 $Y=1.985 $X2=0 $Y2=0
cc_147 N_C1_M1005_g B1 6.31774e-19 $X=1.97 $Y=0.56 $X2=0 $Y2=0
cc_148 C1 B1 0.0517409f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_149 N_C1_c_176_n N_B1_c_213_n 9.02556e-19 $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_150 C1 N_B1_c_214_n 0.00100889f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_151 N_C1_c_176_n N_B1_c_214_n 0.0163132f $X=2.03 $Y=1.16 $X2=0 $Y2=0
cc_152 N_C1_M1002_g N_VPWR_c_332_n 0.00486043f $X=1.97 $Y=1.985 $X2=0 $Y2=0
cc_153 N_C1_M1002_g N_VPWR_c_333_n 0.0132613f $X=1.97 $Y=1.985 $X2=0 $Y2=0
cc_154 N_C1_M1002_g N_VPWR_c_338_n 0.00107663f $X=1.97 $Y=1.985 $X2=0 $Y2=0
cc_155 N_C1_M1002_g N_VPWR_c_331_n 0.00866921f $X=1.97 $Y=1.985 $X2=0 $Y2=0
cc_156 N_C1_M1005_g N_VGND_c_393_n 0.00425863f $X=1.97 $Y=0.56 $X2=0 $Y2=0
cc_157 C1 N_VGND_c_393_n 0.00881455f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_158 N_C1_M1005_g N_VGND_c_395_n 0.00700304f $X=1.97 $Y=0.56 $X2=0 $Y2=0
cc_159 C1 N_VGND_c_395_n 0.00898535f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_160 C1 A_409_47# 0.00615909f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_161 N_B1_M1001_g N_A2_M1007_g 0.00857689f $X=2.485 $Y=0.56 $X2=0 $Y2=0
cc_162 B1 N_A2_M1007_g 0.00203551f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_163 N_B1_c_213_n N_A2_M1007_g 5.32297e-19 $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B1_M1006_g N_A2_M1000_g 0.022019f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B1_M1006_g N_A2_c_253_n 2.49602e-19 $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_166 N_B1_c_213_n N_A2_c_253_n 0.0108187f $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_167 N_B1_c_214_n N_A2_c_253_n 8.90622e-19 $X=2.73 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B1_c_213_n N_A2_c_254_n 5.29616e-19 $X=2.62 $Y=1.16 $X2=0 $Y2=0
cc_169 N_B1_c_214_n N_A2_c_254_n 0.0145849f $X=2.73 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_M1006_g A2 0.00105217f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B1_M1006_g N_VPWR_c_333_n 0.0198569f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_172 N_B1_M1006_g N_VPWR_c_337_n 0.00173838f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B1_M1006_g N_VPWR_c_331_n 0.00387135f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B1_M1001_g N_VGND_c_393_n 0.00432565f $X=2.485 $Y=0.56 $X2=0 $Y2=0
cc_175 B1 N_VGND_c_393_n 0.00788921f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_176 N_B1_M1001_g N_VGND_c_395_n 0.00761145f $X=2.485 $Y=0.56 $X2=0 $Y2=0
cc_177 B1 N_VGND_c_395_n 0.0081173f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_178 B1 N_A_512_47#_M1001_d 0.00577491f $X=2.445 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_179 N_B1_M1001_g N_A_512_47#_c_454_n 0.00395001f $X=2.485 $Y=0.56 $X2=0 $Y2=0
cc_180 B1 N_A_512_47#_c_454_n 0.0234191f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_181 N_B1_M1001_g N_A_512_47#_c_451_n 6.15707e-19 $X=2.485 $Y=0.56 $X2=0 $Y2=0
cc_182 B1 N_A_512_47#_c_451_n 0.0135863f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_183 N_A2_M1007_g N_A1_M1009_g 0.0284142f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A2_M1000_g N_A1_M1003_g 0.0479841f $X=3.305 $Y=1.985 $X2=0 $Y2=0
cc_185 A2 N_A1_M1003_g 0.00399262f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_186 N_A2_c_254_n A1 4.61796e-19 $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_187 A2 A1 0.0185915f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_188 N_A2_c_255_n A1 0.0204697f $X=3.442 $Y=1.325 $X2=0 $Y2=0
cc_189 N_A2_c_254_n N_A1_c_296_n 0.0479841f $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A2_c_255_n N_A1_c_296_n 0.00190503f $X=3.442 $Y=1.325 $X2=0 $Y2=0
cc_191 N_A2_M1000_g N_VPWR_c_333_n 0.00122602f $X=3.305 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A2_M1000_g N_VPWR_c_335_n 0.00176946f $X=3.305 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A2_M1000_g N_VPWR_c_337_n 0.00543342f $X=3.305 $Y=1.985 $X2=0 $Y2=0
cc_194 A2 N_VPWR_c_337_n 0.00818262f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_195 N_A2_M1000_g N_VPWR_c_331_n 0.00989397f $X=3.305 $Y=1.985 $X2=0 $Y2=0
cc_196 A2 N_VPWR_c_331_n 0.00672871f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_197 A2 A_676_297# 0.00104458f $X=3.365 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_198 N_A2_M1007_g N_VGND_c_391_n 0.00306721f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A2_M1007_g N_VGND_c_393_n 0.00435108f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A2_M1007_g N_VGND_c_395_n 0.00641885f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A2_M1007_g N_A_512_47#_c_449_n 0.0101766f $X=3.245 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A2_c_253_n N_A_512_47#_c_449_n 0.010401f $X=3.35 $Y=1.2 $X2=0 $Y2=0
cc_203 N_A2_c_254_n N_A_512_47#_c_449_n 0.00148964f $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A2_c_255_n N_A_512_47#_c_449_n 0.0125972f $X=3.442 $Y=1.325 $X2=0 $Y2=0
cc_205 N_A2_c_253_n N_A_512_47#_c_451_n 0.00595765f $X=3.35 $Y=1.2 $X2=0 $Y2=0
cc_206 N_A2_c_254_n N_A_512_47#_c_451_n 0.00239859f $X=3.215 $Y=1.16 $X2=0 $Y2=0
cc_207 A1 N_VPWR_M1003_d 0.0031427f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_208 N_A1_M1003_g N_VPWR_c_335_n 0.0122285f $X=3.665 $Y=1.985 $X2=0 $Y2=0
cc_209 A1 N_VPWR_c_335_n 0.0214721f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_210 N_A1_c_296_n N_VPWR_c_335_n 0.00102056f $X=3.87 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A1_M1003_g N_VPWR_c_337_n 0.00544582f $X=3.665 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A1_M1003_g N_VPWR_c_331_n 0.00906165f $X=3.665 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A1_M1009_g N_VGND_c_391_n 0.0088385f $X=3.665 $Y=0.56 $X2=0 $Y2=0
cc_214 N_A1_M1009_g N_VGND_c_394_n 0.00347311f $X=3.665 $Y=0.56 $X2=0 $Y2=0
cc_215 N_A1_M1009_g N_VGND_c_395_n 0.0050404f $X=3.665 $Y=0.56 $X2=0 $Y2=0
cc_216 N_A1_M1009_g N_A_512_47#_c_449_n 0.0167007f $X=3.665 $Y=0.56 $X2=0 $Y2=0
cc_217 A1 N_A_512_47#_c_449_n 0.0222797f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_218 N_A1_c_296_n N_A_512_47#_c_449_n 0.00585725f $X=3.87 $Y=1.16 $X2=0 $Y2=0
cc_219 N_X_c_320_n N_VPWR_c_336_n 0.0176389f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_220 N_X_M1010_s N_VPWR_c_331_n 0.00348182f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_221 N_X_c_320_n N_VPWR_c_331_n 0.00993603f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_222 N_X_c_320_n N_VGND_c_392_n 0.0176389f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_223 N_X_M1011_s N_VGND_c_395_n 0.00348182f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_224 N_X_c_320_n N_VGND_c_395_n 0.00993603f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_225 N_VPWR_c_331_n A_676_297# 0.00364937f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_226 N_VGND_c_395_n A_306_47# 0.00851809f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_227 N_VGND_c_395_n A_409_47# 0.0105275f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_228 N_VGND_c_395_n N_A_512_47#_M1001_d 0.0113694f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_229 N_VGND_c_395_n N_A_512_47#_M1009_d 0.00235517f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_393_n N_A_512_47#_c_454_n 0.018535f $X=3.33 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_c_395_n N_A_512_47#_c_454_n 0.0110646f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_M1007_d N_A_512_47#_c_449_n 0.00335756f $X=3.32 $Y=0.235 $X2=0
+ $Y2=0
cc_233 N_VGND_c_391_n N_A_512_47#_c_449_n 0.0142193f $X=3.455 $Y=0.37 $X2=0
+ $Y2=0
cc_234 N_VGND_c_393_n N_A_512_47#_c_449_n 0.00224628f $X=3.33 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_394_n N_A_512_47#_c_449_n 0.00207753f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_c_395_n N_A_512_47#_c_449_n 0.00879055f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_394_n N_A_512_47#_c_450_n 0.0182296f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_395_n N_A_512_47#_c_450_n 0.0101041f $X=3.91 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__sdfbbp_1.pex.spice
* Created: Tue Sep  1 19:29:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%CLK 4 5 7 8 10 13 17 19 20 24 26
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r47 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r49 15 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_27_47# 1 2 9 13 15 17 20 26 28 29 32 36
+ 40 41 42 45 47 51 52 55 56 57 58 59 68 73 80 81 85 86 87
c264 85 0 2.05666e-19 $X=8.445 $Y=1.74
c265 52 0 9.71454e-20 $X=4.71 $Y=0.87
c266 45 0 1.78014e-19 $X=0.72 $Y=1.795
c267 26 0 3.84972e-20 $X=8.505 $Y=2.275
r268 85 88 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.74
+ $X2=8.445 $Y2=1.905
r269 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.74
+ $X2=8.445 $Y2=1.575
r270 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.445
+ $Y=1.74 $X2=8.445 $Y2=1.74
r271 80 83 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.04 $Y=1.74
+ $X2=5.04 $Y2=1.875
r272 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=1.74 $X2=5.04 $Y2=1.74
r273 68 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=1.87
+ $X2=8.51 $Y2=1.87
r274 66 81 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=1.765
+ $X2=5.04 $Y2=1.765
r275 66 93 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=4.83 $Y=1.765
+ $X2=4.735 $Y2=1.765
r276 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.87
+ $X2=4.83 $Y2=1.87
r277 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.87
+ $X2=0.69 $Y2=1.87
r278 59 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=1.87
+ $X2=4.83 $Y2=1.87
r279 58 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.365 $Y=1.87
+ $X2=8.51 $Y2=1.87
r280 58 59 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=8.365 $Y=1.87
+ $X2=4.975 $Y2=1.87
r281 57 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.87
+ $X2=0.69 $Y2=1.87
r282 56 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=4.83 $Y2=1.87
r283 56 57 4.76484 $w=1.4e-07 $l=3.85e-06 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=0.835 $Y2=1.87
r284 52 75 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=4.71 $Y=0.87
+ $X2=4.58 $Y2=0.87
r285 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.71
+ $Y=0.87 $X2=4.71 $Y2=0.87
r286 49 93 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.735 $Y=1.575
+ $X2=4.735 $Y2=1.765
r287 49 51 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=4.735 $Y=1.575
+ $X2=4.735 $Y2=0.87
r288 48 73 31.1043 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=0.75 $Y=1.235
+ $X2=0.89 $Y2=1.235
r289 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.235 $X2=0.75 $Y2=1.235
r290 45 62 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.795
+ $X2=0.72 $Y2=1.88
r291 45 47 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.72 $Y=1.795
+ $X2=0.72 $Y2=1.235
r292 44 47 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.72 $Y=0.805
+ $X2=0.72 $Y2=1.235
r293 43 55 3.4683 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.257 $Y2=1.88
r294 42 62 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.72 $Y2=1.88
r295 42 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.345 $Y2=1.88
r296 40 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.72 $Y2=0.805
r297 40 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.345 $Y2=0.72
r298 34 41 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.345 $Y2=0.72
r299 34 36 7.92208 $w=1.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.257 $Y2=0.51
r300 30 32 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.035 $Y=1.245
+ $X2=9.035 $Y2=0.415
r301 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.96 $Y=1.32
+ $X2=9.035 $Y2=1.245
r302 28 29 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=8.96 $Y=1.32
+ $X2=8.58 $Y2=1.32
r303 26 88 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.505 $Y=2.275
+ $X2=8.505 $Y2=1.905
r304 22 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.505 $Y=1.395
+ $X2=8.58 $Y2=1.32
r305 22 87 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.505 $Y=1.395
+ $X2=8.505 $Y2=1.575
r306 20 83 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.01 $Y=2.275
+ $X2=5.01 $Y2=1.875
r307 15 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.58 $Y=0.705
+ $X2=4.58 $Y2=0.87
r308 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.58 $Y=0.705
+ $X2=4.58 $Y2=0.415
r309 11 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r310 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r311 7 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r312 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r313 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r314 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%SCD 3 7 9 10 17
c37 9 0 5.96503e-20 $X=1.61 $Y=1.19
c38 7 0 1.53494e-19 $X=1.83 $Y=2.135
c39 3 0 7.69389e-20 $X=1.83 $Y=0.445
r40 14 17 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.635 $Y=1.49
+ $X2=1.83 $Y2=1.49
r41 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.49 $X2=1.635 $Y2=1.49
r42 9 10 12.3476 $w=2.78e-07 $l=3e-07 $layer=LI1_cond $X=1.58 $Y=1.19 $X2=1.58
+ $Y2=1.49
r43 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.655
+ $X2=1.83 $Y2=1.49
r44 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.83 $Y=1.655 $X2=1.83
+ $Y2=2.135
r45 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.49
r46 1 3 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.83 $Y=1.325 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_423_315# 1 2 7 9 10 11 14 17 21 23 25 26
+ 30 31 33 34 40 46
c104 34 0 4.64297e-20 $X=2.905 $Y=1.66
c105 25 0 2.25267e-19 $X=3.475 $Y=0.71
c106 11 0 5.96503e-20 $X=2.265 $Y=1.65
c107 10 0 1.65209e-19 $X=2.695 $Y=1.65
r108 37 39 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=1.74
+ $X2=2.905 $Y2=1.905
r109 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.74 $X2=2.845 $Y2=1.74
r110 34 37 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=2.905 $Y=1.66
+ $X2=2.905 $Y2=1.74
r111 33 40 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.56 $Y=1.575
+ $X2=3.56 $Y2=1.095
r112 31 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=0.93
+ $X2=3.685 $Y2=0.765
r113 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=0.93 $X2=3.685 $Y2=0.93
r114 28 40 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=3.622 $Y=0.948
+ $X2=3.622 $Y2=1.095
r115 28 30 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=3.622 $Y=0.948
+ $X2=3.622 $Y2=0.93
r116 27 30 5.27389 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=3.622 $Y=0.795
+ $X2=3.622 $Y2=0.93
r117 25 27 19.9305 $w=8.7e-08 $l=1.84673e-07 $layer=LI1_cond $X=3.475 $Y=0.71
+ $X2=3.622 $Y2=0.795
r118 25 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.475 $Y=0.71
+ $X2=3.125 $Y2=0.71
r119 24 34 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.065 $Y=1.66
+ $X2=2.905 $Y2=1.66
r120 23 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.475 $Y=1.66
+ $X2=3.56 $Y2=1.575
r121 23 24 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.475 $Y=1.66
+ $X2=3.065 $Y2=1.66
r122 19 26 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.025 $Y=0.625
+ $X2=3.125 $Y2=0.71
r123 19 21 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=3.025 $Y=0.625
+ $X2=3.025 $Y2=0.47
r124 17 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.98 $Y=2.3
+ $X2=2.98 $Y2=1.905
r125 14 46 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.745 $Y=0.445
+ $X2=3.745 $Y2=0.765
r126 10 38 18.9432 $w=2.85e-07 $l=9e-08 $layer=POLY_cond $X=2.837 $Y=1.65
+ $X2=2.837 $Y2=1.74
r127 10 11 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.695 $Y=1.65
+ $X2=2.265 $Y2=1.65
r128 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.19 $Y=1.725
+ $X2=2.265 $Y2=1.65
r129 7 9 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.19 $Y=1.725
+ $X2=2.19 $Y2=2.135
r130 2 17 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=2.065 $X2=2.98 $Y2=2.3
r131 1 21 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%SCE 1 3 4 6 8 10 11 13 14 16 18 19 20 26 29
+ 30 31 35
c98 35 0 7.23866e-20 $X=2.25 $Y=0.81
c99 26 0 1.18777e-19 $X=2.25 $Y=0.93
c100 19 0 4.83365e-20 $X=3.257 $Y=0.81
c101 4 0 4.64297e-20 $X=3.175 $Y=0.81
r102 30 31 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.07 $Y=1.19
+ $X2=2.07 $Y2=1.53
r103 27 35 21.6629 $w=2.67e-07 $l=1.2e-07 $layer=POLY_cond $X=2.25 $Y=0.93
+ $X2=2.25 $Y2=0.81
r104 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=0.93 $X2=2.25 $Y2=0.93
r105 22 30 9.16716 $w=2.18e-07 $l=1.75e-07 $layer=LI1_cond $X=2.07 $Y=1.015
+ $X2=2.07 $Y2=1.19
r106 22 29 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=2.07 $Y=0.845
+ $X2=2.07 $Y2=0.51
r107 22 26 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.07 $Y=0.93
+ $X2=2.25 $Y2=0.93
r108 16 18 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.685 $Y=1.985
+ $X2=3.685 $Y2=2.275
r109 15 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=1.91
+ $X2=3.265 $Y2=1.91
r110 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.61 $Y=1.91
+ $X2=3.685 $Y2=1.985
r111 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.61 $Y=1.91
+ $X2=3.34 $Y2=1.91
r112 11 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.985
+ $X2=3.265 $Y2=1.91
r113 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.265 $Y=1.985
+ $X2=3.265 $Y2=2.275
r114 10 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.835
+ $X2=3.265 $Y2=1.91
r115 9 19 20.4101 $w=1.5e-07 $l=7.88987e-08 $layer=POLY_cond $X=3.265 $Y=0.885
+ $X2=3.257 $Y2=0.81
r116 9 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.265 $Y=0.885
+ $X2=3.265 $Y2=1.835
r117 6 19 20.4101 $w=1.5e-07 $l=7.84219e-08 $layer=POLY_cond $X=3.25 $Y=0.735
+ $X2=3.257 $Y2=0.81
r118 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.25 $Y=0.735
+ $X2=3.25 $Y2=0.445
r119 5 35 16.2448 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.385 $Y=0.81
+ $X2=2.25 $Y2=0.81
r120 4 19 5.30422 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=3.175 $Y=0.81
+ $X2=3.257 $Y2=0.81
r121 4 5 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.175 $Y=0.81
+ $X2=2.385 $Y2=0.81
r122 1 35 22.72 $w=2.67e-07 $l=8.87412e-08 $layer=POLY_cond $X=2.22 $Y=0.735
+ $X2=2.25 $Y2=0.81
r123 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.22 $Y=0.735
+ $X2=2.22 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%D 3 7 9 10 17
c42 3 0 1.09936e-19 $X=4.105 $Y=0.445
r43 14 17 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.94 $Y=1.49
+ $X2=4.105 $Y2=1.49
r44 9 10 39.9273 $w=1.98e-07 $l=7.2e-07 $layer=LI1_cond $X=3.925 $Y=1.49
+ $X2=3.925 $Y2=2.21
r45 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.49 $X2=3.94 $Y2=1.49
r46 5 17 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=1.49
r47 5 7 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=2.275
r48 1 17 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.105 $Y=1.355
+ $X2=4.105 $Y2=1.49
r49 1 3 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.105 $Y=1.355
+ $X2=4.105 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_193_47# 1 2 9 11 12 15 18 19 21 24 28 29
+ 31 33 34 36 37 39 40 41 48 52 56 57 68
c231 39 0 9.71454e-20 $X=5.327 $Y=1.12
c232 31 0 1.22107e-19 $X=8.937 $Y=1.305
c233 29 0 1.7288e-19 $X=8.615 $Y=0.87
c234 9 0 4.43992e-20 $X=4.59 $Y=2.275
r235 56 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.93
+ $X2=5.19 $Y2=1.095
r236 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.93
+ $X2=5.19 $Y2=0.765
r237 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.19
+ $Y=0.93 $X2=5.19 $Y2=0.93
r238 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=1.19
+ $X2=8.51 $Y2=1.19
r239 48 50 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=5.29 $Y=0.85
+ $X2=5.29 $Y2=0.965
r240 48 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0.85
+ $X2=5.29 $Y2=0.85
r241 44 72 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.96
r242 44 68 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.51
r243 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0.85
+ $X2=1.15 $Y2=0.85
r244 40 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=8.51 $Y2=1.19
r245 40 41 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=5.435 $Y2=1.19
r246 39 41 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=5.327 $Y=1.12
+ $X2=5.435 $Y2=1.19
r247 39 50 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=5.327 $Y=1.12
+ $X2=5.327 $Y2=0.965
r248 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=0.85
+ $X2=1.15 $Y2=0.85
r249 36 48 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=0.85
+ $X2=5.29 $Y2=0.85
r250 36 37 4.76484 $w=1.4e-07 $l=3.85e-06 $layer=MET1_cond $X=5.145 $Y=0.85
+ $X2=1.295 $Y2=0.85
r251 34 66 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.955 $Y=1.74
+ $X2=8.955 $Y2=1.875
r252 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.955
+ $Y=1.74 $X2=8.955 $Y2=1.74
r253 31 53 26.3101 $w=1.78e-07 $l=4.27e-07 $layer=LI1_cond $X=8.937 $Y=1.215
+ $X2=8.51 $Y2=1.215
r254 31 33 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=8.937 $Y=1.305
+ $X2=8.937 $Y2=1.74
r255 29 60 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=8.615 $Y=0.87
+ $X2=8.495 $Y2=0.87
r256 28 53 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=8.562 $Y=0.87
+ $X2=8.562 $Y2=1.125
r257 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.615
+ $Y=0.87 $X2=8.615 $Y2=0.87
r258 24 66 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=8.925 $Y=2.275
+ $X2=8.925 $Y2=1.875
r259 19 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.495 $Y=0.705
+ $X2=8.495 $Y2=0.87
r260 19 21 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.495 $Y=0.705
+ $X2=8.495 $Y2=0.415
r261 18 59 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.13 $Y=1.245
+ $X2=5.13 $Y2=1.095
r262 15 58 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.13 $Y=0.415
+ $X2=5.13 $Y2=0.765
r263 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.055 $Y=1.32
+ $X2=5.13 $Y2=1.245
r264 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=5.055 $Y=1.32
+ $X2=4.665 $Y2=1.32
r265 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.59 $Y=1.395
+ $X2=4.665 $Y2=1.32
r266 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=4.59 $Y=1.395
+ $X2=4.59 $Y2=2.275
r267 2 72 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r268 1 68 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_1107_21# 1 2 9 13 17 19 21 22 26 28 30 31
+ 32 35 36 41 45 49
c146 45 0 9.73505e-20 $X=7.96 $Y=0.98
r147 49 56 9.60507 $w=2.76e-07 $l=5.5e-08 $layer=POLY_cond $X=7.96 $Y=1.15
+ $X2=8.015 $Y2=1.15
r148 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.96
+ $Y=1.15 $X2=7.96 $Y2=1.15
r149 45 48 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.96 $Y=0.98
+ $X2=7.96 $Y2=1.15
r150 43 44 14.2969 $w=2.56e-07 $l=3e-07 $layer=LI1_cond $X=6.865 $Y=0.68
+ $X2=6.865 $Y2=0.98
r151 36 53 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.74
+ $X2=5.695 $Y2=1.905
r152 36 52 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.74
+ $X2=5.695 $Y2=1.575
r153 35 38 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.76 $Y=1.74
+ $X2=5.76 $Y2=1.91
r154 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.72
+ $Y=1.74 $X2=5.72 $Y2=1.74
r155 33 44 3.13337 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.03 $Y=0.98
+ $X2=6.865 $Y2=0.98
r156 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=0.98
+ $X2=7.96 $Y2=0.98
r157 32 33 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=7.795 $Y=0.98
+ $X2=7.03 $Y2=0.98
r158 30 44 5.42994 $w=2.56e-07 $l=1.00995e-07 $layer=LI1_cond $X=6.9 $Y=1.065
+ $X2=6.865 $Y2=0.98
r159 30 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.9 $Y=1.065
+ $X2=6.9 $Y2=1.785
r160 29 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.91
+ $X2=6.47 $Y2=1.91
r161 28 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.815 $Y=1.91
+ $X2=6.9 $Y2=1.785
r162 28 29 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=6.815 $Y=1.91
+ $X2=6.555 $Y2=1.91
r163 24 41 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.47 $Y=2.035
+ $X2=6.47 $Y2=1.91
r164 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.47 $Y=2.035
+ $X2=6.47 $Y2=2.21
r165 23 38 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=1.91
+ $X2=5.76 $Y2=1.91
r166 22 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=1.91
+ $X2=6.47 $Y2=1.91
r167 22 23 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=6.385 $Y=1.91
+ $X2=5.885 $Y2=1.91
r168 19 56 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.015 $Y=0.985
+ $X2=8.015 $Y2=1.15
r169 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.015 $Y=0.985
+ $X2=8.015 $Y2=0.555
r170 15 49 30.5616 $w=2.76e-07 $l=2.43926e-07 $layer=POLY_cond $X=7.785 $Y=1.315
+ $X2=7.96 $Y2=1.15
r171 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=7.785 $Y=1.315
+ $X2=7.785 $Y2=2.065
r172 13 53 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.61 $Y=2.275
+ $X2=5.61 $Y2=1.905
r173 9 52 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=5.61 $Y=0.445
+ $X2=5.61 $Y2=1.575
r174 2 41 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.065 $X2=6.47 $Y2=1.87
r175 2 26 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.065 $X2=6.47 $Y2=2.21
r176 1 43 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=6.73
+ $Y=0.235 $X2=6.865 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%SET_B 1 3 7 11 15 17 19 20 26 27 33
c129 33 0 1.51196e-19 $X=9.93 $Y=0.98
c130 19 0 1.30137e-19 $X=9.745 $Y=0.85
c131 15 0 1.0852e-19 $X=10.055 $Y=2.275
r132 33 36 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.962 $Y=0.98
+ $X2=9.962 $Y2=1.145
r133 33 35 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.962 $Y=0.98
+ $X2=9.962 $Y2=0.815
r134 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.93
+ $Y=0.98 $X2=9.93 $Y2=0.98
r135 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0.85
+ $X2=9.89 $Y2=0.85
r136 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.355 $Y=0.85
+ $X2=6.21 $Y2=0.85
r137 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.745 $Y=0.85
+ $X2=9.89 $Y2=0.85
r138 19 20 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=9.745 $Y=0.85
+ $X2=6.355 $Y2=0.85
r139 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.05
+ $Y=0.98 $X2=6.05 $Y2=0.98
r140 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0.85
+ $X2=6.21 $Y2=0.85
r141 15 36 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=10.055 $Y=2.275
+ $X2=10.055 $Y2=1.145
r142 11 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.055 $Y=0.445
+ $X2=10.055 $Y2=0.815
r143 5 30 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=6.18 $Y=0.815
+ $X2=6.085 $Y2=0.98
r144 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.18 $Y=0.815
+ $X2=6.18 $Y2=0.445
r145 1 30 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=6.14 $Y=1.145
+ $X2=6.085 $Y2=0.98
r146 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.14 $Y=1.145
+ $X2=6.14 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_931_47# 1 2 9 13 15 19 24 26 27 32 35
c105 35 0 1.30137e-19 $X=6.56 $Y=1.32
c106 32 0 4.43992e-20 $X=5.715 $Y=1.3
r107 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=1.32
+ $X2=6.59 $Y2=1.485
r108 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=1.32
+ $X2=6.59 $Y2=1.155
r109 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.56
+ $Y=1.32 $X2=6.56 $Y2=1.32
r110 31 32 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=5.63 $Y=1.3
+ $X2=5.715 $Y2=1.3
r111 29 31 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=5.38 $Y=1.3
+ $X2=5.63 $Y2=1.3
r112 27 34 8.9562 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=1.32
+ $X2=6.56 $Y2=1.32
r113 27 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.395 $Y=1.32
+ $X2=5.715 $Y2=1.32
r114 26 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.63 $Y=1.195
+ $X2=5.63 $Y2=1.3
r115 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.63 $Y=0.465
+ $X2=5.63 $Y2=1.195
r116 23 29 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.38 $Y=1.405
+ $X2=5.38 $Y2=1.3
r117 23 24 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.38 $Y=1.405
+ $X2=5.38 $Y2=2.25
r118 19 25 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.545 $Y=0.365
+ $X2=5.63 $Y2=0.465
r119 19 21 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=5.545 $Y=0.365
+ $X2=4.865 $Y2=0.365
r120 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.295 $Y=2.335
+ $X2=5.38 $Y2=2.25
r121 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.295 $Y=2.335
+ $X2=4.8 $Y2=2.335
r122 13 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.68 $Y=2.065
+ $X2=6.68 $Y2=1.485
r123 9 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.655 $Y=0.555
+ $X2=6.655 $Y2=1.155
r124 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=2.065 $X2=4.8 $Y2=2.335
r125 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.235 $X2=4.865 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_1400_21# 1 2 7 9 10 12 16 20 22 23 24 26
+ 30 33 41 42 45 48 53 56
c158 53 0 6.74557e-20 $X=10.95 $Y=1.32
c159 41 0 2.58372e-20 $X=11.125 $Y=1.53
c160 26 0 1.52865e-19 $X=11.68 $Y=1.66
c161 7 0 9.73505e-20 $X=7.075 $Y=0.95
r162 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.165
+ $Y=1.32 $X2=11.165 $Y2=1.32
r163 53 55 33.5372 $w=3.09e-07 $l=2.15e-07 $layer=POLY_cond $X=10.95 $Y=1.32
+ $X2=11.165 $Y2=1.32
r164 52 53 8.57929 $w=3.09e-07 $l=5.5e-08 $layer=POLY_cond $X=10.895 $Y=1.32
+ $X2=10.95 $Y2=1.32
r165 49 56 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=11.217 $Y=1.53
+ $X2=11.217 $Y2=1.32
r166 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=1.53
+ $X2=11.27 $Y2=1.53
r167 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=1.53
+ $X2=8.05 $Y2=1.53
r168 42 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.195 $Y=1.53
+ $X2=8.05 $Y2=1.53
r169 41 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.125 $Y=1.53
+ $X2=11.27 $Y2=1.53
r170 41 42 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.125 $Y=1.53
+ $X2=8.195 $Y2=1.53
r171 40 49 1.88582 $w=2.73e-07 $l=4.5e-08 $layer=LI1_cond $X=11.217 $Y=1.575
+ $X2=11.217 $Y2=1.53
r172 39 56 16.5533 $w=2.73e-07 $l=3.95e-07 $layer=LI1_cond $X=11.217 $Y=0.925
+ $X2=11.217 $Y2=1.32
r173 37 45 27.1304 $w=2.38e-07 $l=5.65e-07 $layer=LI1_cond $X=7.485 $Y=1.535
+ $X2=8.05 $Y2=1.535
r174 36 37 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=7.32 $Y=1.535
+ $X2=7.485 $Y2=1.535
r175 33 36 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.32 $Y=1.32
+ $X2=7.32 $Y2=1.535
r176 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.32
+ $Y=1.32 $X2=7.32 $Y2=1.32
r177 28 30 18.0227 $w=1.98e-07 $l=3.25e-07 $layer=LI1_cond $X=11.665 $Y=0.755
+ $X2=11.665 $Y2=0.43
r178 24 40 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=11.355 $Y=1.66
+ $X2=11.217 $Y2=1.575
r179 24 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.355 $Y=1.66
+ $X2=11.68 $Y2=1.66
r180 23 39 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=11.355 $Y=0.84
+ $X2=11.217 $Y2=0.925
r181 22 28 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.665 $Y2=0.755
r182 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.355 $Y2=0.84
r183 18 53 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.95 $Y=1.155
+ $X2=10.95 $Y2=1.32
r184 18 20 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=10.95 $Y=1.155
+ $X2=10.95 $Y2=0.555
r185 14 52 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.895 $Y=1.485
+ $X2=10.895 $Y2=1.32
r186 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.895 $Y=1.485
+ $X2=10.895 $Y2=2.065
r187 10 34 38.5938 $w=3.29e-07 $l=2.19499e-07 $layer=POLY_cond $X=7.1 $Y=1.485
+ $X2=7.227 $Y2=1.32
r188 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.1 $Y=1.485
+ $X2=7.1 $Y2=2.065
r189 7 34 68.6272 $w=3.29e-07 $l=4.39477e-07 $layer=POLY_cond $X=7.075 $Y=0.95
+ $X2=7.227 $Y2=1.32
r190 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.075 $Y=0.95
+ $X2=7.075 $Y2=0.555
r191 2 26 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=11.555
+ $Y=1.505 $X2=11.68 $Y2=1.66
r192 1 30 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=11.555
+ $Y=0.235 $X2=11.68 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_1887_21# 1 2 9 13 15 17 20 22 23 25 27 28
+ 30 31 33 36 38 41 45 46 48 49 52 54 57 58 61 62 64 67 71
c182 46 0 1.29033e-19 $X=9.635 $Y=1.74
c183 20 0 1.52865e-19 $X=12.375 $Y=1.985
c184 9 0 8.93206e-20 $X=9.51 $Y=0.445
r185 72 79 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=12.34 $Y=1.16
+ $X2=12.375 $Y2=1.16
r186 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.34
+ $Y=1.16 $X2=12.34 $Y2=1.16
r187 68 71 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=12.245 $Y=1.16
+ $X2=12.34 $Y2=1.16
r188 60 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=1.325
+ $X2=12.245 $Y2=1.16
r189 60 61 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.245 $Y=1.325
+ $X2=12.245 $Y2=1.915
r190 59 67 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=10.905 $Y=2
+ $X2=10.817 $Y2=2
r191 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.16 $Y=2
+ $X2=12.245 $Y2=1.915
r192 58 59 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=12.16 $Y=2
+ $X2=10.905 $Y2=2
r193 57 67 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.817 $Y=1.915
+ $X2=10.817 $Y2=2
r194 56 64 0.574824 $w=1.75e-07 $l=1.17346e-07 $layer=LI1_cond $X=10.817
+ $Y=0.815 $X2=10.74 $Y2=0.73
r195 56 57 69.7143 $w=1.73e-07 $l=1.1e-06 $layer=LI1_cond $X=10.817 $Y=0.815
+ $X2=10.817 $Y2=1.915
r196 55 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.41 $Y=2
+ $X2=10.325 $Y2=2
r197 54 67 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=10.73 $Y=2
+ $X2=10.817 $Y2=2
r198 54 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.73 $Y=2 $X2=10.41
+ $Y2=2
r199 50 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.325 $Y=2.085
+ $X2=10.325 $Y2=2
r200 50 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.325 $Y=2.085
+ $X2=10.325 $Y2=2.21
r201 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.24 $Y=2
+ $X2=10.325 $Y2=2
r202 48 49 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=10.24 $Y=2 $X2=9.8
+ $Y2=2
r203 46 76 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.602 $Y=1.74
+ $X2=9.602 $Y2=1.905
r204 46 75 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=9.602 $Y=1.74
+ $X2=9.602 $Y2=1.575
r205 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.635
+ $Y=1.74 $X2=9.635 $Y2=1.74
r206 43 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.675 $Y=1.915
+ $X2=9.8 $Y2=2
r207 43 45 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=9.675 $Y=1.915
+ $X2=9.675 $Y2=1.74
r208 39 41 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=13.19 $Y=1.61
+ $X2=13.315 $Y2=1.61
r209 34 36 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=13.19 $Y=0.805
+ $X2=13.315 $Y2=0.805
r210 31 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.315 $Y=1.685
+ $X2=13.315 $Y2=1.61
r211 31 33 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=13.315 $Y=1.685
+ $X2=13.315 $Y2=2.085
r212 28 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.315 $Y=0.73
+ $X2=13.315 $Y2=0.805
r213 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.315 $Y=0.73
+ $X2=13.315 $Y2=0.445
r214 27 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.19 $Y=1.535
+ $X2=13.19 $Y2=1.61
r215 26 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.19 $Y=1.295
+ $X2=13.19 $Y2=1.16
r216 26 27 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=13.19 $Y=1.295
+ $X2=13.19 $Y2=1.535
r217 25 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.19 $Y=1.025
+ $X2=13.19 $Y2=1.16
r218 24 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.19 $Y=0.88
+ $X2=13.19 $Y2=0.805
r219 24 25 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=13.19 $Y=0.88
+ $X2=13.19 $Y2=1.025
r220 23 79 19.5642 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=12.475 $Y=1.16
+ $X2=12.375 $Y2=1.16
r221 22 38 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=13.115 $Y=1.16
+ $X2=13.19 $Y2=1.16
r222 22 23 142.191 $w=2.7e-07 $l=6.4e-07 $layer=POLY_cond $X=13.115 $Y=1.16
+ $X2=12.475 $Y2=1.16
r223 18 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.375 $Y=1.325
+ $X2=12.375 $Y2=1.16
r224 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.375 $Y=1.325
+ $X2=12.375 $Y2=1.985
r225 15 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.375 $Y=0.995
+ $X2=12.375 $Y2=1.16
r226 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.375 $Y=0.995
+ $X2=12.375 $Y2=0.56
r227 13 76 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.515 $Y=2.275
+ $X2=9.515 $Y2=1.905
r228 9 75 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=9.51 $Y=0.445
+ $X2=9.51 $Y2=1.575
r229 2 52 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=2.065 $X2=10.325 $Y2=2.21
r230 1 64 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=10.605
+ $Y=0.235 $X2=10.74 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_1714_47# 1 2 9 13 15 19 24 26 27 29 31 32
c98 32 0 2.58372e-20 $X=10.475 $Y=1.24
c99 31 0 1.75976e-19 $X=10.475 $Y=1.24
c100 26 0 3.84972e-20 $X=9.295 $Y=2.25
r101 32 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.475 $Y=1.24
+ $X2=10.475 $Y2=1.405
r102 32 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.475 $Y=1.24
+ $X2=10.475 $Y2=1.075
r103 31 34 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=10.45 $Y=1.24
+ $X2=10.45 $Y2=1.32
r104 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.475
+ $Y=1.24 $X2=10.475 $Y2=1.24
r105 28 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.38 $Y=1.32
+ $X2=9.295 $Y2=1.32
r106 27 34 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=10.34 $Y=1.32
+ $X2=10.45 $Y2=1.32
r107 27 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.34 $Y=1.32
+ $X2=9.38 $Y2=1.32
r108 25 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=1.405
+ $X2=9.295 $Y2=1.32
r109 25 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=9.295 $Y=1.405
+ $X2=9.295 $Y2=2.25
r110 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=1.235
+ $X2=9.295 $Y2=1.32
r111 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=9.295 $Y=0.465
+ $X2=9.295 $Y2=1.235
r112 19 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.21 $Y=0.365
+ $X2=9.295 $Y2=0.465
r113 19 21 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=9.21 $Y=0.365
+ $X2=8.78 $Y2=0.365
r114 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.21 $Y=2.335
+ $X2=9.295 $Y2=2.25
r115 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.21 $Y=2.335
+ $X2=8.715 $Y2=2.335
r116 13 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.535 $Y=2.065
+ $X2=10.535 $Y2=1.405
r117 9 37 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=10.53 $Y=0.555
+ $X2=10.53 $Y2=1.075
r118 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=8.58
+ $Y=2.065 $X2=8.715 $Y2=2.335
r119 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.57
+ $Y=0.235 $X2=8.78 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%RESET_B 3 7 9 15
r36 12 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=11.7 $Y=1.18
+ $X2=11.89 $Y2=1.18
r37 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.7
+ $Y=1.18 $X2=11.7 $Y2=1.18
r38 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.89 $Y=1.345
+ $X2=11.89 $Y2=1.18
r39 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.89 $Y=1.345
+ $X2=11.89 $Y2=1.825
r40 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.89 $Y=1.015
+ $X2=11.89 $Y2=1.18
r41 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=11.89 $Y=1.015
+ $X2=11.89 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_2596_47# 1 2 9 12 16 20 24 25 27 29
c52 27 0 1.39343e-19 $X=13.117 $Y=1.16
r53 25 30 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.725 $Y=1.16
+ $X2=13.725 $Y2=1.325
r54 25 29 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.725 $Y=1.16
+ $X2=13.725 $Y2=0.995
r55 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.71
+ $Y=1.16 $X2=13.71 $Y2=1.16
r56 22 27 1.17559 $w=3.3e-07 $l=1.58e-07 $layer=LI1_cond $X=13.275 $Y=1.16
+ $X2=13.117 $Y2=1.16
r57 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=13.275 $Y=1.16
+ $X2=13.71 $Y2=1.16
r58 18 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=13.117 $Y=1.325
+ $X2=13.117 $Y2=1.16
r59 18 20 21.4025 $w=3.13e-07 $l=5.85e-07 $layer=LI1_cond $X=13.117 $Y=1.325
+ $X2=13.117 $Y2=1.91
r60 14 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=13.117 $Y=0.995
+ $X2=13.117 $Y2=1.16
r61 14 16 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=13.117 $Y=0.995
+ $X2=13.117 $Y2=0.51
r62 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.79 $Y=1.985
+ $X2=13.79 $Y2=1.325
r63 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.79 $Y=0.56
+ $X2=13.79 $Y2=0.995
r64 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.98
+ $Y=1.765 $X2=13.105 $Y2=1.91
r65 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=12.98
+ $Y=0.235 $X2=13.105 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 53
+ 54 55 59 60 62 64 70 75 83 95 106 110 117 118 121 124 127 130 133 144 146
c211 118 0 3.07047e-19 $X=14.03 $Y=2.72
r212 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r213 142 144 9.28831 $w=5.48e-07 $l=1.4e-07 $layer=LI1_cond $X=12.19 $Y=2.53
+ $X2=12.33 $Y2=2.53
r214 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r215 140 142 0.543672 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=12.165 $Y=2.53
+ $X2=12.19 $Y2=2.53
r216 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r217 133 136 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=9.81 $Y=2.34
+ $X2=9.81 $Y2=2.72
r218 130 131 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r219 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r220 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r221 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r222 118 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=13.57 $Y2=2.72
r223 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r224 115 146 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=13.745 $Y=2.72
+ $X2=13.597 $Y2=2.72
r225 115 117 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.745 $Y=2.72
+ $X2=14.03 $Y2=2.72
r226 114 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r227 114 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=12.19 $Y2=2.72
r228 113 144 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=13.11 $Y=2.72
+ $X2=12.33 $Y2=2.72
r229 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r230 110 146 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=13.45 $Y=2.72
+ $X2=13.597 $Y2=2.72
r231 110 113 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.45 $Y=2.72
+ $X2=13.11 $Y2=2.72
r232 109 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r233 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r234 106 140 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=12.055 $Y=2.53
+ $X2=12.165 $Y2=2.53
r235 106 108 17.0713 $w=5.48e-07 $l=7.85e-07 $layer=LI1_cond $X=12.055 $Y=2.53
+ $X2=11.27 $Y2=2.53
r236 105 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r237 105 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=9.89 $Y2=2.72
r238 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r239 102 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10 $Y=2.72
+ $X2=9.81 $Y2=2.72
r240 102 104 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=10 $Y=2.72
+ $X2=10.81 $Y2=2.72
r241 101 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r242 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r243 98 101 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r244 97 100 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r245 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r246 95 136 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.81 $Y2=2.72
r247 95 100 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.43 $Y2=2.72
r248 94 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r249 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r250 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r251 91 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r252 90 93 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r253 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r254 88 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=5.895 $Y2=2.72
r255 88 90 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.085 $Y=2.72
+ $X2=6.21 $Y2=2.72
r256 87 131 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.75 $Y2=2.72
r257 87 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r258 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r259 84 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=2.72
+ $X2=3.475 $Y2=2.72
r260 84 86 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.64 $Y=2.72
+ $X2=3.91 $Y2=2.72
r261 83 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=5.895 $Y2=2.72
r262 83 86 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=5.705 $Y=2.72
+ $X2=3.91 $Y2=2.72
r263 82 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r264 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r265 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r266 79 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r267 78 81 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r268 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r269 76 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r270 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r271 75 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=2.72
+ $X2=3.475 $Y2=2.72
r272 75 81 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.31 $Y=2.72
+ $X2=2.99 $Y2=2.72
r273 74 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r274 74 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r275 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r276 71 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r277 71 73 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r278 70 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r279 70 73 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r280 64 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r281 62 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r282 60 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r283 60 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r284 59 104 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=10.94 $Y=2.72
+ $X2=10.81 $Y2=2.72
r285 58 59 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=11.105 $Y=2.53
+ $X2=10.94 $Y2=2.53
r286 55 108 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=11.215 $Y=2.53
+ $X2=11.27 $Y2=2.53
r287 55 58 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=11.215 $Y=2.53
+ $X2=11.105 $Y2=2.53
r288 53 93 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.13 $Y2=2.72
r289 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=2.72
+ $X2=7.34 $Y2=2.72
r290 52 97 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=7.59 $Y2=2.72
r291 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=2.72
+ $X2=7.34 $Y2=2.72
r292 48 146 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=13.597 $Y=2.635
+ $X2=13.597 $Y2=2.72
r293 48 50 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=13.597 $Y=2.635
+ $X2=13.597 $Y2=1.94
r294 44 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.34 $Y=2.635
+ $X2=7.34 $Y2=2.72
r295 44 46 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.34 $Y=2.635
+ $X2=7.34 $Y2=2
r296 40 130 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.895 $Y=2.635
+ $X2=5.895 $Y2=2.72
r297 40 42 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=5.895 $Y=2.635
+ $X2=5.895 $Y2=2.29
r298 36 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=2.635
+ $X2=3.475 $Y2=2.72
r299 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.475 $Y=2.635
+ $X2=3.475 $Y2=2.3
r300 32 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r301 32 34 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=1.97
r302 28 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r303 28 30 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r304 9 50 300 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=2 $X=13.39
+ $Y=1.765 $X2=13.58 $Y2=1.94
r305 8 140 600 $w=1.7e-07 $l=9.29637e-07 $layer=licon1_PDIFF $count=1 $X=11.965
+ $Y=1.505 $X2=12.165 $Y2=2.34
r306 7 58 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=10.97
+ $Y=1.645 $X2=11.105 $Y2=2.34
r307 6 133 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=9.59
+ $Y=2.065 $X2=9.785 $Y2=2.34
r308 5 46 300 $w=1.7e-07 $l=4.29651e-07 $layer=licon1_PDIFF $count=2 $X=7.175
+ $Y=1.645 $X2=7.34 $Y2=2
r309 4 42 600 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=2.065 $X2=5.87 $Y2=2.29
r310 3 38 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=2.065 $X2=3.475 $Y2=2.3
r311 2 34 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.815 $X2=1.62 $Y2=1.97
r312 1 30 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_453_363# 1 2 3 4 18 20 21 25 27 30 31 34
+ 37 43
c114 31 0 1.15331e-19 $X=3.135 $Y=1.19
c115 27 0 4.64318e-20 $X=2.755 $Y=1.22
c116 21 0 1.53494e-19 $X=2.4 $Y=1.875
c117 18 0 7.69389e-20 $X=2.67 $Y=1.075
r118 38 47 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=4.342 $Y=1.19
+ $X2=4.342 $Y2=2.3
r119 38 43 36.8782 $w=2.23e-07 $l=7.2e-07 $layer=LI1_cond $X=4.342 $Y=1.19
+ $X2=4.342 $Y2=0.47
r120 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=1.19
+ $X2=4.37 $Y2=1.19
r121 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.19
+ $X2=2.99 $Y2=1.19
r122 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.19
+ $X2=2.99 $Y2=1.19
r123 30 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.19
+ $X2=4.37 $Y2=1.19
r124 30 31 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=4.225 $Y=1.19
+ $X2=3.135 $Y2=1.19
r125 28 29 11.4982 $w=2.26e-07 $l=2.13e-07 $layer=LI1_cond $X=2.457 $Y=1.22
+ $X2=2.67 $Y2=1.22
r126 27 34 9.33876 $w=2.88e-07 $l=2.35e-07 $layer=LI1_cond $X=2.755 $Y=1.22
+ $X2=2.99 $Y2=1.22
r127 27 29 4.20283 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=1.22
+ $X2=2.67 $Y2=1.22
r128 23 25 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=2.435 $Y=0.43
+ $X2=2.67 $Y2=0.43
r129 20 21 4.36643 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=1.96 $X2=2.4
+ $Y2=1.875
r130 18 29 2.4068 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.67 $Y=1.075
+ $X2=2.67 $Y2=1.22
r131 17 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0.595
+ $X2=2.67 $Y2=0.43
r132 17 18 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.67 $Y=0.595
+ $X2=2.67 $Y2=1.075
r133 15 28 1.0459 $w=2.15e-07 $l=1.45e-07 $layer=LI1_cond $X=2.457 $Y=1.365
+ $X2=2.457 $Y2=1.22
r134 15 21 27.337 $w=2.13e-07 $l=5.1e-07 $layer=LI1_cond $X=2.457 $Y=1.365
+ $X2=2.457 $Y2=1.875
r135 4 47 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=2.065 $X2=4.315 $Y2=2.3
r136 3 20 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.815 $X2=2.4 $Y2=1.96
r137 2 43 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.235 $X2=4.315 $Y2=0.47
r138 1 23 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.235 $X2=2.435 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%Q_N 1 2 9 10 11 12 13 18 21
r31 18 21 2.69684 $w=2.85e-07 $l=6.3e-08 $layer=LI1_cond $X=12.642 $Y=0.573
+ $X2=12.642 $Y2=0.51
r32 12 13 15.9725 $w=2.83e-07 $l=3.95e-07 $layer=LI1_cond $X=12.642 $Y=1.815
+ $X2=12.642 $Y2=2.21
r33 11 30 6.85431 $w=2.83e-07 $l=1.31e-07 $layer=LI1_cond $X=12.642 $Y=0.584
+ $X2=12.642 $Y2=0.715
r34 11 18 0.444803 $w=2.83e-07 $l=1.1e-08 $layer=LI1_cond $X=12.642 $Y=0.584
+ $X2=12.642 $Y2=0.573
r35 11 21 0.470877 $w=2.85e-07 $l=1.1e-08 $layer=LI1_cond $X=12.642 $Y=0.499
+ $X2=12.642 $Y2=0.51
r36 10 30 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=12.695 $Y=1.63
+ $X2=12.695 $Y2=0.715
r37 9 12 1.73877 $w=2.83e-07 $l=4.3e-08 $layer=LI1_cond $X=12.642 $Y=1.772
+ $X2=12.642 $Y2=1.815
r38 9 10 7.29911 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=12.642 $Y=1.772
+ $X2=12.642 $Y2=1.63
r39 2 12 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=12.45
+ $Y=1.485 $X2=12.585 $Y2=1.815
r40 1 21 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=12.45
+ $Y=0.235 $X2=12.585 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%Q 1 2 10 11 12 13 14 15
r16 14 15 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=14.045 $Y=1.82
+ $X2=14.045 $Y2=2.21
r17 11 14 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=14.045 $Y=1.735
+ $X2=14.045 $Y2=1.82
r18 11 12 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=14.045 $Y=1.735
+ $X2=14.045 $Y2=1.605
r19 10 12 41.1948 $w=2.08e-07 $l=7.8e-07 $layer=LI1_cond $X=14.07 $Y=0.825
+ $X2=14.07 $Y2=1.605
r20 9 13 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=14.045 $Y=0.695
+ $X2=14.045 $Y2=0.51
r21 9 10 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=14.045 $Y=0.695
+ $X2=14.045 $Y2=0.825
r22 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=13.865
+ $Y=1.485 $X2=14 $Y2=1.82
r23 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=13.865
+ $Y=0.235 $X2=14 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 61 62 64 65 66 68 70 76 81 105 112 119 120 123 126 129 132 135
c208 120 0 2.71124e-20 $X=14.03 $Y=0
c209 81 0 1.20723e-19 $X=3.37 $Y=0
c210 47 0 1.51196e-19 $X=9.735 $Y=0.36
r211 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r212 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r213 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r214 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r215 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r216 120 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=13.57 $Y2=0
r217 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r218 117 135 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.745 $Y=0
+ $X2=13.6 $Y2=0
r219 117 119 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.745 $Y=0
+ $X2=14.03 $Y2=0
r220 116 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=13.57 $Y2=0
r221 116 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=12.19 $Y2=0
r222 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r223 113 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.33 $Y=0
+ $X2=12.165 $Y2=0
r224 113 115 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=12.33 $Y=0
+ $X2=13.11 $Y2=0
r225 112 135 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.6 $Y2=0
r226 112 115 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.11 $Y2=0
r227 111 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r228 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r229 108 111 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r230 107 110 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r231 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r232 105 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12 $Y=0
+ $X2=12.165 $Y2=0
r233 105 110 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12 $Y=0 $X2=11.73
+ $Y2=0
r234 104 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r235 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r236 101 104 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.43 $Y2=0
r237 100 103 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=9.43 $Y2=0
r238 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r239 98 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r240 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r241 95 98 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r242 94 97 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=7.59
+ $Y2=0
r243 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r244 92 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r245 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r246 89 92 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r247 89 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=3.45 $Y2=0
r248 88 91 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.75
+ $Y2=0
r249 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r250 86 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.535
+ $Y2=0
r251 86 88 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.91
+ $Y2=0
r252 85 130 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r253 85 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r254 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r255 82 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=1.58 $Y2=0
r256 82 84 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r257 81 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.37 $Y=0
+ $X2=3.535 $Y2=0
r258 81 84 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=3.37 $Y=0 $X2=2.07
+ $Y2=0
r259 80 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r260 80 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r261 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r262 77 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r263 77 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r264 76 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.58 $Y2=0
r265 76 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r266 70 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r267 68 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r268 66 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r269 66 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r270 64 103 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=9.56 $Y=0 $X2=9.43
+ $Y2=0
r271 64 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.56 $Y=0 $X2=9.69
+ $Y2=0
r272 63 107 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=9.82 $Y=0 $X2=9.89
+ $Y2=0
r273 63 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.82 $Y=0 $X2=9.69
+ $Y2=0
r274 61 97 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.59
+ $Y2=0
r275 61 62 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.807
+ $Y2=0
r276 60 100 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.975 $Y=0
+ $X2=8.05 $Y2=0
r277 60 62 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.975 $Y=0
+ $X2=7.807 $Y2=0
r278 58 91 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.885 $Y=0
+ $X2=5.75 $Y2=0
r279 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=0 $X2=5.97
+ $Y2=0
r280 57 94 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.055 $Y=0
+ $X2=6.21 $Y2=0
r281 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=0 $X2=5.97
+ $Y2=0
r282 53 135 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=13.6 $Y=0.085
+ $X2=13.6 $Y2=0
r283 53 55 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=13.6 $Y=0.085
+ $X2=13.6 $Y2=0.38
r284 49 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.165 $Y=0.085
+ $X2=12.165 $Y2=0
r285 49 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=12.165 $Y=0.085
+ $X2=12.165 $Y2=0.38
r286 45 65 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=0.085
+ $X2=9.69 $Y2=0
r287 45 47 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=9.69 $Y=0.085
+ $X2=9.69 $Y2=0.36
r288 41 62 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.807 $Y=0.085
+ $X2=7.807 $Y2=0
r289 41 43 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=7.807 $Y=0.085
+ $X2=7.807 $Y2=0.38
r290 37 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0
r291 37 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0.36
r292 33 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0
r293 33 35 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0.36
r294 29 126 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r295 29 31 17.7476 $w=2.48e-07 $l=3.85e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.47
r296 25 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r297 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r298 8 55 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=13.39
+ $Y=0.235 $X2=13.58 $Y2=0.38
r299 7 51 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=11.965
+ $Y=0.235 $X2=12.165 $Y2=0.38
r300 6 47 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=9.585
+ $Y=0.235 $X2=9.735 $Y2=0.36
r301 5 43 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.68
+ $Y=0.235 $X2=7.805 $Y2=0.38
r302 4 39 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.97 $Y2=0.36
r303 3 35 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.535 $Y2=0.36
r304 2 31 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.47
r305 1 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_1251_47# 1 2 7 11 16
r25 14 16 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.39 $Y=0.36
+ $X2=6.555 $Y2=0.36
r26 9 11 7.10956 $w=1.93e-07 $l=1.25e-07 $layer=LI1_cond $X=7.297 $Y=0.425
+ $X2=7.297 $Y2=0.55
r27 7 9 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=7.2 $Y=0.34
+ $X2=7.297 $Y2=0.425
r28 7 16 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=7.2 $Y=0.34
+ $X2=6.555 $Y2=0.34
r29 2 11 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=7.15
+ $Y=0.235 $X2=7.285 $Y2=0.55
r30 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.235 $X2=6.39 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFBBP_1%A_2026_47# 1 2 7 12
r20 10 12 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=10.265 $Y=0.36
+ $X2=10.43 $Y2=0.36
r21 7 12 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=11.075 $Y=0.34
+ $X2=10.43 $Y2=0.34
r22 2 7 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=11.025
+ $Y=0.235 $X2=11.16 $Y2=0.42
r23 1 10 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=10.13
+ $Y=0.235 $X2=10.265 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__clkdlybuf4s25_1.spice
* Created: Thu Aug 27 14:11:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkdlybuf4s25_1.pex.spice"
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_27_47#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0964037 AS=0.1134 PD=0.836075 PS=1.38 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1005 N_A_244_47#_M1005_d N_A_27_47#_M1005_g N_VGND_M1001_d VNB NSHORT L=0.25
+ W=0.65 AD=0.17225 AS=0.149196 PD=1.83 PS=1.29393 NRD=0 NRS=15.684 M=1 R=2.6
+ SA=125001 SB=125000 A=0.1625 P=1.8 MULT=1
MM1002 N_VGND_M1002_d N_A_244_47#_M1002_g N_A_355_47#_M1002_s VNB NSHORT L=0.25
+ W=0.65 AD=0.225495 AS=0.17225 PD=1.53084 PS=1.83 NRD=46.152 NRS=0 M=1 R=2.6
+ SA=125000 SB=125001 A=0.1625 P=1.8 MULT=1
MM1006 N_X_M1006_d N_A_355_47#_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.2079 AS=0.145705 PD=1.83 PS=0.989159 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.1 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.211703 AS=0.27 PD=1.55495 PS=2.54 NRD=12.7853 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_A_244_47#_M1007_d N_A_27_47#_M1007_g N_VPWR_M1004_d VPB PHIGHVT L=0.25
+ W=0.82 AD=0.2173 AS=0.173597 PD=2.17 PS=1.27505 NRD=0 NRS=16.8041 M=1 R=3.28
+ SA=125001 SB=125000 A=0.205 P=2.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_244_47#_M1000_g N_A_355_47#_M1000_s VPB PHIGHVT L=0.25
+ W=0.82 AD=0.24564 AS=0.2173 PD=1.45077 PS=2.17 NRD=60.0456 NRS=0 M=1 R=3.28
+ SA=125000 SB=125001 A=0.205 P=2.14 MULT=1
MM1003 N_X_M1003_d N_A_355_47#_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.495 AS=0.29956 PD=2.99 PS=1.76923 NRD=0 NRS=15.7403 M=1 R=6.66667
+ SA=75000.9 SB=75000.4 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_34 VNB 0 5.32225e-20 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__clkdlybuf4s25_1.pxi.spice"
*
.ends
*
*

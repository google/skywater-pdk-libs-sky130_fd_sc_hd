* File: sky130_fd_sc_hd__dfstp_4.pxi.spice
* Created: Thu Aug 27 14:15:29 2020
* 
x_PM_SKY130_FD_SC_HD__DFSTP_4%CLK N_CLK_c_248_n N_CLK_c_243_n N_CLK_M1036_g
+ N_CLK_c_249_n N_CLK_M1019_g N_CLK_c_244_n N_CLK_c_250_n CLK CLK N_CLK_c_246_n
+ N_CLK_c_247_n PM_SKY130_FD_SC_HD__DFSTP_4%CLK
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_27_47# N_A_27_47#_M1036_s N_A_27_47#_M1019_s
+ N_A_27_47#_M1022_g N_A_27_47#_M1000_g N_A_27_47#_c_288_n N_A_27_47#_M1034_g
+ N_A_27_47#_M1039_g N_A_27_47#_M1003_g N_A_27_47#_M1014_g N_A_27_47#_c_543_p
+ N_A_27_47#_c_289_n N_A_27_47#_c_290_n N_A_27_47#_c_304_n N_A_27_47#_c_416_p
+ N_A_27_47#_c_291_n N_A_27_47#_c_292_n N_A_27_47#_c_293_n N_A_27_47#_c_294_n
+ N_A_27_47#_c_295_n N_A_27_47#_c_296_n N_A_27_47#_c_308_n N_A_27_47#_c_297_n
+ N_A_27_47#_c_298_n N_A_27_47#_c_309_n N_A_27_47#_c_310_n N_A_27_47#_c_311_n
+ N_A_27_47#_c_312_n N_A_27_47#_c_313_n N_A_27_47#_c_299_n N_A_27_47#_c_315_n
+ N_A_27_47#_c_316_n N_A_27_47#_c_317_n N_A_27_47#_c_318_n N_A_27_47#_c_300_n
+ PM_SKY130_FD_SC_HD__DFSTP_4%A_27_47#
x_PM_SKY130_FD_SC_HD__DFSTP_4%D N_D_M1008_g N_D_M1028_g D D N_D_c_561_n
+ N_D_c_562_n PM_SKY130_FD_SC_HD__DFSTP_4%D
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_193_47# N_A_193_47#_M1022_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1009_g N_A_193_47#_c_599_n N_A_193_47#_c_600_n
+ N_A_193_47#_M1020_g N_A_193_47#_c_602_n N_A_193_47#_M1012_g
+ N_A_193_47#_c_604_n N_A_193_47#_M1030_g N_A_193_47#_c_605_n
+ N_A_193_47#_c_606_n N_A_193_47#_c_607_n N_A_193_47#_c_608_n
+ N_A_193_47#_c_609_n N_A_193_47#_c_610_n N_A_193_47#_c_611_n
+ N_A_193_47#_c_612_n N_A_193_47#_c_613_n N_A_193_47#_c_614_n
+ N_A_193_47#_c_615_n N_A_193_47#_c_616_n PM_SKY130_FD_SC_HD__DFSTP_4%A_193_47#
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_652_21# N_A_652_21#_M1005_d N_A_652_21#_M1033_d
+ N_A_652_21#_M1025_g N_A_652_21#_M1007_g N_A_652_21#_c_800_n
+ N_A_652_21#_c_884_p N_A_652_21#_c_801_n N_A_652_21#_c_795_n
+ N_A_652_21#_c_796_n N_A_652_21#_c_803_n N_A_652_21#_c_804_n
+ N_A_652_21#_c_805_n N_A_652_21#_c_797_n PM_SKY130_FD_SC_HD__DFSTP_4%A_652_21#
x_PM_SKY130_FD_SC_HD__DFSTP_4%SET_B N_SET_B_c_909_n N_SET_B_M1033_g
+ N_SET_B_M1002_g N_SET_B_M1021_g N_SET_B_M1001_g N_SET_B_c_913_n
+ N_SET_B_c_924_n N_SET_B_c_914_n N_SET_B_c_915_n SET_B N_SET_B_c_917_n
+ N_SET_B_c_918_n N_SET_B_c_919_n N_SET_B_c_920_n
+ PM_SKY130_FD_SC_HD__DFSTP_4%SET_B
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_476_47# N_A_476_47#_M1034_d N_A_476_47#_M1009_d
+ N_A_476_47#_c_1043_n N_A_476_47#_M1005_g N_A_476_47#_c_1044_n
+ N_A_476_47#_M1023_g N_A_476_47#_c_1045_n N_A_476_47#_M1017_g
+ N_A_476_47#_c_1046_n N_A_476_47#_M1024_g N_A_476_47#_c_1047_n
+ N_A_476_47#_c_1070_n N_A_476_47#_c_1075_n N_A_476_47#_c_1055_n
+ N_A_476_47#_c_1048_n N_A_476_47#_c_1049_n N_A_476_47#_c_1050_n
+ N_A_476_47#_c_1051_n N_A_476_47#_c_1052_n
+ PM_SKY130_FD_SC_HD__DFSTP_4%A_476_47#
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_1178_261# N_A_1178_261#_M1018_d
+ N_A_1178_261#_M1027_d N_A_1178_261#_M1015_g N_A_1178_261#_M1016_g
+ N_A_1178_261#_c_1201_n N_A_1178_261#_c_1206_n N_A_1178_261#_c_1207_n
+ N_A_1178_261#_c_1238_p N_A_1178_261#_c_1202_n N_A_1178_261#_c_1203_n
+ N_A_1178_261#_c_1209_n N_A_1178_261#_c_1210_n
+ PM_SKY130_FD_SC_HD__DFSTP_4%A_1178_261#
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_1028_413# N_A_1028_413#_M1012_d
+ N_A_1028_413#_M1003_d N_A_1028_413#_M1001_s N_A_1028_413#_M1018_g
+ N_A_1028_413#_M1027_g N_A_1028_413#_c_1281_n N_A_1028_413#_M1006_g
+ N_A_1028_413#_M1011_g N_A_1028_413#_c_1283_n N_A_1028_413#_c_1302_n
+ N_A_1028_413#_c_1294_n N_A_1028_413#_c_1310_n N_A_1028_413#_c_1284_n
+ N_A_1028_413#_c_1285_n N_A_1028_413#_c_1296_n N_A_1028_413#_c_1286_n
+ N_A_1028_413#_c_1297_n N_A_1028_413#_c_1298_n N_A_1028_413#_c_1384_n
+ N_A_1028_413#_c_1287_n N_A_1028_413#_c_1288_n N_A_1028_413#_c_1289_n
+ PM_SKY130_FD_SC_HD__DFSTP_4%A_1028_413#
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_1598_47# N_A_1598_47#_M1006_s
+ N_A_1598_47#_M1011_s N_A_1598_47#_M1026_g N_A_1598_47#_M1004_g
+ N_A_1598_47#_M1031_g N_A_1598_47#_M1010_g N_A_1598_47#_M1032_g
+ N_A_1598_47#_M1013_g N_A_1598_47#_M1037_g N_A_1598_47#_M1029_g
+ N_A_1598_47#_M1038_g N_A_1598_47#_M1035_g N_A_1598_47#_c_1452_n
+ N_A_1598_47#_c_1453_n N_A_1598_47#_c_1461_n N_A_1598_47#_c_1462_n
+ N_A_1598_47#_c_1454_n N_A_1598_47#_c_1455_n
+ PM_SKY130_FD_SC_HD__DFSTP_4%A_1598_47#
x_PM_SKY130_FD_SC_HD__DFSTP_4%VPWR N_VPWR_M1019_d N_VPWR_M1028_s N_VPWR_M1007_d
+ N_VPWR_M1023_d N_VPWR_M1015_d N_VPWR_M1001_d N_VPWR_M1011_d N_VPWR_M1010_d
+ N_VPWR_M1029_d N_VPWR_c_1569_n N_VPWR_c_1570_n N_VPWR_c_1571_n N_VPWR_c_1572_n
+ N_VPWR_c_1573_n N_VPWR_c_1574_n N_VPWR_c_1575_n N_VPWR_c_1576_n VPWR VPWR
+ N_VPWR_c_1577_n N_VPWR_c_1578_n N_VPWR_c_1579_n N_VPWR_c_1580_n
+ N_VPWR_c_1581_n N_VPWR_c_1582_n N_VPWR_c_1583_n N_VPWR_c_1584_n
+ N_VPWR_c_1585_n N_VPWR_c_1568_n N_VPWR_c_1587_n N_VPWR_c_1588_n
+ N_VPWR_c_1589_n N_VPWR_c_1590_n N_VPWR_c_1591_n N_VPWR_c_1592_n
+ N_VPWR_c_1593_n N_VPWR_c_1594_n N_VPWR_c_1595_n
+ PM_SKY130_FD_SC_HD__DFSTP_4%VPWR
x_PM_SKY130_FD_SC_HD__DFSTP_4%A_381_47# N_A_381_47#_M1008_d N_A_381_47#_M1028_d
+ N_A_381_47#_c_1763_n N_A_381_47#_c_1768_n N_A_381_47#_c_1764_n
+ N_A_381_47#_c_1770_n N_A_381_47#_c_1766_n N_A_381_47#_c_1772_n
+ N_A_381_47#_c_1773_n PM_SKY130_FD_SC_HD__DFSTP_4%A_381_47#
x_PM_SKY130_FD_SC_HD__DFSTP_4%Q N_Q_M1026_d N_Q_M1032_d N_Q_M1038_d N_Q_M1004_s
+ N_Q_M1013_s N_Q_M1035_s N_Q_c_1840_n N_Q_c_1829_n N_Q_c_1833_n N_Q_c_1834_n
+ N_Q_c_1895_p N_Q_c_1880_n N_Q_c_1856_n N_Q_c_1835_n N_Q_c_1830_n N_Q_c_1836_n
+ Q Q Q Q Q Q Q Q Q N_Q_c_1839_n PM_SKY130_FD_SC_HD__DFSTP_4%Q
x_PM_SKY130_FD_SC_HD__DFSTP_4%VGND N_VGND_M1036_d N_VGND_M1008_s N_VGND_M1025_d
+ N_VGND_M1024_s N_VGND_M1021_d N_VGND_M1006_d N_VGND_M1031_s N_VGND_M1037_s
+ N_VGND_c_1907_n N_VGND_c_1908_n N_VGND_c_1909_n N_VGND_c_1910_n
+ N_VGND_c_1911_n N_VGND_c_1912_n N_VGND_c_1913_n VGND VGND N_VGND_c_1914_n
+ N_VGND_c_1915_n N_VGND_c_1916_n N_VGND_c_1917_n N_VGND_c_1918_n
+ N_VGND_c_1919_n N_VGND_c_1920_n N_VGND_c_1921_n N_VGND_c_1922_n
+ N_VGND_c_1923_n N_VGND_c_1924_n N_VGND_c_1925_n N_VGND_c_1926_n
+ N_VGND_c_1927_n N_VGND_c_1928_n N_VGND_c_1929_n N_VGND_c_1930_n
+ N_VGND_c_1931_n PM_SKY130_FD_SC_HD__DFSTP_4%VGND
cc_1 VNB N_CLK_c_243_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_c_244_n 0.0229857f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK 0.0187424f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_c_246_n 0.01953f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_CLK_c_247_n 0.0141141f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_6 VNB N_A_27_47#_M1022_g 0.0364978f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_288_n 0.0180457f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_8 VNB N_A_27_47#_c_289_n 0.00174761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_290_n 0.00643757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_291_n 0.00246672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_292_n 0.00445416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_293_n 0.0327378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_294_n 0.00637933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_295_n 0.00847145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_296_n 0.00156937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_297_n 0.00506957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_298_n 0.0254428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_299_n 0.022701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_300_n 0.0159476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_M1008_g 0.0205663f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_21 VNB N_D_c_561_n 0.0258802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_D_c_562_n 0.00442451f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_23 VNB N_A_193_47#_c_599_n 0.0132632f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_24 VNB N_A_193_47#_c_600_n 0.00435992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_M1020_g 0.0199482f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_26 VNB N_A_193_47#_c_602_n 0.00803437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_M1012_g 0.0339782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_604_n 0.0100971f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_29 VNB N_A_193_47#_c_605_n 0.018279f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_30 VNB N_A_193_47#_c_606_n 0.0194566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_193_47#_c_607_n 0.00568843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_193_47#_c_608_n 0.00105673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_193_47#_c_609_n 0.0163665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_47#_c_610_n 0.00113053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_c_611_n 0.00189817f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_612_n 0.00500582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_193_47#_c_613_n 0.00145914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_614_n 0.00217053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_193_47#_c_615_n 0.0246637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_616_n 0.0161628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_652_21#_M1025_g 0.0422386f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_42 VNB N_A_652_21#_c_795_n 0.00136482f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_652_21#_c_796_n 0.00314488f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.19
cc_44 VNB N_A_652_21#_c_797_n 0.00513705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_SET_B_c_909_n 0.0308821f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_46 VNB N_SET_B_M1033_g 0.00706345f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_47 VNB N_SET_B_M1002_g 0.0179723f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_48 VNB N_SET_B_M1021_g 0.0183761f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_49 VNB N_SET_B_c_913_n 0.0075909f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_50 VNB N_SET_B_c_914_n 0.0252701f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_51 VNB N_SET_B_c_915_n 0.00436858f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_52 VNB SET_B 0.00646661f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_53 VNB N_SET_B_c_917_n 0.0137018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_918_n 0.00185354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_SET_B_c_919_n 3.85333e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_SET_B_c_920_n 0.00287603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_476_47#_c_1043_n 0.017726f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_58 VNB N_A_476_47#_c_1044_n 0.0138425f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_59 VNB N_A_476_47#_c_1045_n 0.0548714f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_476_47#_c_1046_n 0.0177765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_476_47#_c_1047_n 0.00507008f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_62 VNB N_A_476_47#_c_1048_n 0.00430167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_476_47#_c_1049_n 0.00446117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_476_47#_c_1050_n 0.00393532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_476_47#_c_1051_n 0.00107462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_476_47#_c_1052_n 0.0145441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1178_261#_M1016_g 0.0370862f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_68 VNB N_A_1178_261#_c_1201_n 0.00831402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1178_261#_c_1202_n 0.00717461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1178_261#_c_1203_n 0.00525762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1028_413#_M1018_g 0.0319034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1028_413#_c_1281_n 0.0390811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1028_413#_M1006_g 0.0419771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1028_413#_c_1283_n 0.00671176f $X=-0.19 $Y=-0.24 $X2=0.265
+ $Y2=1.19
cc_75 VNB N_A_1028_413#_c_1284_n 0.00499598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1028_413#_c_1285_n 0.0010444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1028_413#_c_1286_n 0.00897687f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1028_413#_c_1287_n 7.51809e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1028_413#_c_1288_n 0.012418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1028_413#_c_1289_n 0.00455313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1598_47#_M1026_g 0.018138f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_82 VNB N_A_1598_47#_M1004_g 4.83494e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_83 VNB N_A_1598_47#_M1031_g 0.017456f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_84 VNB N_A_1598_47#_M1010_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1598_47#_M1032_g 0.0172288f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_86 VNB N_A_1598_47#_M1013_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1598_47#_M1037_g 0.0172272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1598_47#_M1029_g 4.50048e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1598_47#_M1038_g 0.0218695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1598_47#_M1035_g 4.97409e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1598_47#_c_1452_n 0.00339441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_1598_47#_c_1453_n 0.0143242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_1598_47#_c_1454_n 3.08128e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_1598_47#_c_1455_n 0.0813174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VPWR_c_1568_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_381_47#_c_1763_n 0.00882912f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_97 VNB N_A_381_47#_c_1764_n 0.00229945f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_98 VNB N_Q_c_1829_n 0.00116361f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_99 VNB N_Q_c_1830_n 0.00116361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB Q 0.0201933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB Q 0.0307859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1907_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_103 VNB N_VGND_c_1908_n 0.00492922f $X=-0.19 $Y=-0.24 $X2=0.265 $Y2=1.53
cc_104 VNB N_VGND_c_1909_n 0.00404464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1910_n 0.0101869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1911_n 0.00254421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1912_n 0.00163878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1913_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1914_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1915_n 0.0164349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1916_n 0.0451324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1917_n 0.0192996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1918_n 0.0302303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1919_n 0.0149288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1920_n 0.0112161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1921_n 0.0164853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1922_n 0.517898f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1923_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1924_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1925_n 0.0056662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1926_n 0.00651127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1927_n 0.0402451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1928_n 0.0122102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1929_n 0.00427022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1930_n 0.00363423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1931_n 0.00436611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VPB N_CLK_c_248_n 0.0118724f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_128 VPB N_CLK_c_249_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_129 VPB N_CLK_c_250_n 0.0234494f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_130 VPB CLK 0.0178159f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_131 VPB N_CLK_c_246_n 0.0100888f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_132 VPB N_A_27_47#_M1000_g 0.0364742f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_133 VPB N_A_27_47#_M1039_g 0.021588f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_134 VPB N_A_27_47#_M1003_g 0.0202797f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_135 VPB N_A_27_47#_c_304_n 0.00131809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_291_n 0.0033408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_292_n 0.00245013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_27_47#_c_294_n 0.00546282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_27_47#_c_308_n 0.00355155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_309_n 0.0141666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_310_n 0.00223306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_311_n 0.0108096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_312_n 0.0015212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_313_n 0.00372072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_299_n 0.0115872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_315_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_316_n 0.00564526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_27_47#_c_317_n 0.0279259f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_318_n 0.00620409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_D_M1028_g 0.0293669f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_151 VPB N_D_c_561_n 0.00538482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_D_c_562_n 0.00459652f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_153 VPB N_A_193_47#_M1009_g 0.0465266f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_154 VPB N_A_193_47#_c_599_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_155 VPB N_A_193_47#_c_600_n 0.00328709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_193_47#_c_604_n 0.0110035f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_157 VPB N_A_193_47#_M1030_g 0.0394871f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_158 VPB N_A_193_47#_c_605_n 0.0125421f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_159 VPB N_A_193_47#_c_614_n 0.00217264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_193_47#_c_616_n 0.0183598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_652_21#_M1025_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_162 VPB N_A_652_21#_M1007_g 0.0208799f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_163 VPB N_A_652_21#_c_800_n 0.00189033f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_164 VPB N_A_652_21#_c_801_n 0.00247793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_652_21#_c_796_n 0.00270641f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.19
cc_166 VPB N_A_652_21#_c_803_n 0.00460198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_652_21#_c_804_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0.265 $Y2=1.53
cc_168 VPB N_A_652_21#_c_805_n 0.00112185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_SET_B_M1033_g 0.0474843f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_170 VPB N_SET_B_M1001_g 0.038305f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_171 VPB N_SET_B_c_913_n 0.0122551f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_172 VPB N_SET_B_c_924_n 0.00992356f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_173 VPB N_A_476_47#_M1023_g 0.0334449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_476_47#_M1017_g 0.0319093f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_175 VPB N_A_476_47#_c_1055_n 0.0121124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_476_47#_c_1049_n 0.00542515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_476_47#_c_1050_n 0.00271559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_476_47#_c_1051_n 0.00262972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_476_47#_c_1052_n 0.0306997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1178_261#_M1015_g 0.0268094f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_181 VPB N_A_1178_261#_c_1201_n 0.0286069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_1178_261#_c_1206_n 0.0164657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1178_261#_c_1207_n 0.0160465f $X=-0.19 $Y=1.305 $X2=0.245
+ $Y2=1.235
cc_184 VPB N_A_1178_261#_c_1202_n 0.0031237f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1178_261#_c_1209_n 0.0181025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1178_261#_c_1210_n 0.00940573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1028_413#_M1027_g 0.0263696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1028_413#_c_1281_n 0.02945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1028_413#_M1011_g 0.0408752f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.07
cc_190 VPB N_A_1028_413#_c_1283_n 0.00452788f $X=-0.19 $Y=1.305 $X2=0.265
+ $Y2=1.19
cc_191 VPB N_A_1028_413#_c_1294_n 0.00422026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1028_413#_c_1284_n 0.00190145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1028_413#_c_1296_n 0.0149976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1028_413#_c_1297_n 0.0037282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_1028_413#_c_1298_n 2.86428e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_1028_413#_c_1287_n 2.77041e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1028_413#_c_1288_n 0.00840405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1028_413#_c_1289_n 0.00450937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1598_47#_M1004_g 0.0203362f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_200 VPB N_A_1598_47#_M1010_g 0.0193938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1598_47#_M1013_g 0.0191708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_1598_47#_M1029_g 0.0191687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1598_47#_M1035_g 0.024213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1598_47#_c_1461_n 0.00606637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1598_47#_c_1462_n 0.00368113f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1569_n 0.00106376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1570_n 0.00578936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1571_n 0.0114969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1572_n 3.97306e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1573_n 0.00366994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1574_n 0.00282498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1575_n 0.00163878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1576_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1577_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1578_n 0.0163072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1579_n 0.0416374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1580_n 0.0307572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1581_n 0.01851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1582_n 0.0303512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1583_n 0.0154131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1584_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1585_n 0.0170749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1568_n 0.0678661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1587_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1588_n 0.00507833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1589_n 0.0091704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1590_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1591_n 0.011387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1592_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1593_n 0.00427244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1594_n 0.00363289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1595_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_381_47#_c_1763_n 0.0079947f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_234 VPB N_A_381_47#_c_1766_n 0.0018566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_Q_c_1833_n 0.00277073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_Q_c_1834_n 0.00201573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_Q_c_1835_n 0.00345381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_Q_c_1836_n 0.00136595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB Q 0.00856989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB Q 0.00951749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_Q_c_1839_n 0.0361798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 N_CLK_c_243_n N_A_27_47#_M1022_g 0.0200616f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_243 CLK N_A_27_47#_M1022_g 3.09846e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_244 N_CLK_c_247_n N_A_27_47#_M1022_g 0.00508029f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_245 N_CLK_c_250_n N_A_27_47#_M1000_g 0.0276478f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_246 CLK N_A_27_47#_M1000_g 5.73308e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_247 N_CLK_c_246_n N_A_27_47#_M1000_g 0.00530924f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_248 N_CLK_c_243_n N_A_27_47#_c_289_n 0.00684762f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_249 N_CLK_c_244_n N_A_27_47#_c_289_n 0.00787672f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_250 CLK N_A_27_47#_c_289_n 0.00736322f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_251 N_CLK_c_244_n N_A_27_47#_c_290_n 0.0059979f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_252 CLK N_A_27_47#_c_290_n 0.014414f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_253 N_CLK_c_246_n N_A_27_47#_c_290_n 3.2891e-19 $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_254 N_CLK_c_249_n N_A_27_47#_c_304_n 0.0128144f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_255 N_CLK_c_250_n N_A_27_47#_c_304_n 0.0013816f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_256 CLK N_A_27_47#_c_304_n 0.00728212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_257 N_CLK_c_244_n N_A_27_47#_c_291_n 0.00189711f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_258 N_CLK_c_250_n N_A_27_47#_c_291_n 0.00440146f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_259 CLK N_A_27_47#_c_291_n 0.0517133f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_260 N_CLK_c_246_n N_A_27_47#_c_291_n 9.99252e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_261 N_CLK_c_247_n N_A_27_47#_c_291_n 0.00246929f $X=0.245 $Y=1.07 $X2=0 $Y2=0
cc_262 N_CLK_c_249_n N_A_27_47#_c_308_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_263 N_CLK_c_250_n N_A_27_47#_c_308_n 0.00358837f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_264 CLK N_A_27_47#_c_308_n 0.0153363f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_265 N_CLK_c_246_n N_A_27_47#_c_308_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_266 N_CLK_c_249_n N_A_27_47#_c_310_n 0.00102822f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_267 CLK N_A_27_47#_c_299_n 0.00161876f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_268 N_CLK_c_246_n N_A_27_47#_c_299_n 0.0169694f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_269 N_CLK_c_249_n N_VPWR_c_1569_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_270 N_CLK_c_249_n N_VPWR_c_1577_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_271 N_CLK_c_249_n N_VPWR_c_1568_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_272 N_CLK_c_243_n N_VGND_c_1907_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_273 N_CLK_c_243_n N_VGND_c_1914_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_274 N_CLK_c_244_n N_VGND_c_1914_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_275 N_CLK_c_243_n N_VGND_c_1922_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_288_n N_D_M1008_g 0.0210908f $X=2.305 $Y=0.705 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_292_n N_D_M1008_g 0.00120175f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_316_n N_D_M1028_g 7.92917e-19 $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_292_n N_D_c_561_n 0.00106119f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_293_n N_D_c_561_n 0.00155965f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_292_n N_D_c_562_n 0.0453933f $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_293_n N_D_c_562_n 2.37218e-19 $X=2.435 $Y=0.87 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_309_n N_D_c_562_n 0.00575757f $X=2.385 $Y=1.87 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_316_n N_D_c_562_n 0.00408526f $X=2.765 $Y=1.74 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_309_n N_A_193_47#_M1000_d 6.81311e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_M1039_g N_A_193_47#_M1009_g 0.0191849f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_292_n N_A_193_47#_M1009_g 0.0053439f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_309_n N_A_193_47#_M1009_g 0.00702647f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_312_n N_A_193_47#_M1009_g 5.22576e-19 $X=2.675 $Y=1.87 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_315_n N_A_193_47#_M1009_g 0.0174486f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_316_n N_A_193_47#_M1009_g 0.010416f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_292_n N_A_193_47#_c_599_n 0.0101526f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_311_n N_A_193_47#_c_599_n 3.63007e-19 $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_315_n N_A_193_47#_c_599_n 0.0212215f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_316_n N_A_193_47#_c_599_n 0.00655916f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_292_n N_A_193_47#_c_600_n 0.00204176f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_293_n N_A_193_47#_c_600_n 0.0232669f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_288_n N_A_193_47#_M1020_g 0.0128045f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_292_n N_A_193_47#_M1020_g 4.48322e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_293_n N_A_193_47#_M1020_g 0.0214244f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_294_n N_A_193_47#_M1012_g 0.00402103f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_302 N_A_27_47#_c_295_n N_A_193_47#_M1012_g 0.0117214f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_297_n N_A_193_47#_M1012_g 0.00270619f $X=5.985 $Y=0.81 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_298_n N_A_193_47#_M1012_g 0.0209471f $X=5.985 $Y=0.93 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_300_n N_A_193_47#_M1012_g 0.0125268f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1003_g N_A_193_47#_M1030_g 0.0175645f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_294_n N_A_193_47#_M1030_g 0.00215568f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_308 N_A_27_47#_c_313_n N_A_193_47#_M1030_g 0.00434444f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_317_n N_A_193_47#_M1030_g 0.0159766f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_318_n N_A_193_47#_M1030_g 0.00180554f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_294_n N_A_193_47#_c_605_n 0.00355331f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_312 N_A_27_47#_c_295_n N_A_193_47#_c_605_n 0.00394592f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_313_n N_A_193_47#_c_605_n 5.11972e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_317_n N_A_193_47#_c_605_n 0.0106615f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_318_n N_A_193_47#_c_605_n 0.00101144f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_292_n N_A_193_47#_c_606_n 0.0173405f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_293_n N_A_193_47#_c_606_n 0.0059767f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_M1022_g N_A_193_47#_c_607_n 0.00656242f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_289_n N_A_193_47#_c_607_n 0.00216565f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_291_n N_A_193_47#_c_607_n 0.00510004f $X=0.755 $Y=1.235
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_292_n N_A_193_47#_c_608_n 0.00886175f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_294_n N_A_193_47#_c_609_n 0.0118781f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_295_n N_A_193_47#_c_609_n 0.00159218f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_313_n N_A_193_47#_c_609_n 9.05104e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_317_n N_A_193_47#_c_609_n 8.971e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_318_n N_A_193_47#_c_609_n 0.00270751f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_311_n N_A_193_47#_c_610_n 0.0945834f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_292_n N_A_193_47#_c_611_n 5.02791e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_288_n N_A_193_47#_c_612_n 5.21885e-19 $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_c_292_n N_A_193_47#_c_612_n 0.0209059f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_293_n N_A_193_47#_c_612_n 0.00155193f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_315_n N_A_193_47#_c_612_n 3.45191e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_316_n N_A_193_47#_c_612_n 0.00332918f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_294_n N_A_193_47#_c_613_n 0.00256294f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_295_n N_A_193_47#_c_613_n 0.0014885f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_313_n N_A_193_47#_c_613_n 0.0132733f $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_318_n N_A_193_47#_c_613_n 0.00178603f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_294_n N_A_193_47#_c_614_n 0.0285015f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_295_n N_A_193_47#_c_614_n 0.0123304f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_313_n N_A_193_47#_c_614_n 6.9568e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_317_n N_A_193_47#_c_614_n 6.19272e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_318_n N_A_193_47#_c_614_n 0.0119993f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_292_n N_A_193_47#_c_615_n 0.00673428f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_M1022_g N_A_193_47#_c_616_n 0.0272829f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_289_n N_A_193_47#_c_616_n 0.0118856f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_416_p N_A_193_47#_c_616_n 0.00826814f $X=0.725 $Y=1.795
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_c_291_n N_A_193_47#_c_616_n 0.0701221f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_348 N_A_27_47#_c_309_n N_A_193_47#_c_616_n 0.0247331f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_310_n N_A_193_47#_c_616_n 0.00238521f $X=0.845 $Y=1.87 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_292_n N_A_652_21#_M1025_g 5.35023e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_311_n N_A_652_21#_M1007_g 0.00197541f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_311_n N_A_652_21#_c_800_n 0.0147195f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_M1003_g N_A_652_21#_c_801_n 6.75516e-19 $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_311_n N_A_652_21#_c_801_n 0.021867f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_313_n N_A_652_21#_c_801_n 9.32161e-19 $X=5.29 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_318_n N_A_652_21#_c_801_n 0.0093814f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_294_n N_A_652_21#_c_796_n 0.041895f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_311_n N_A_652_21#_c_796_n 0.00686718f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_317_n N_A_652_21#_c_796_n 2.22171e-19 $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_318_n N_A_652_21#_c_796_n 0.0136142f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_311_n N_A_652_21#_c_803_n 0.0157473f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_M1039_g N_A_652_21#_c_804_n 0.0161874f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_311_n N_A_652_21#_c_804_n 0.00193898f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_315_n N_A_652_21#_c_804_n 0.00927772f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_311_n N_A_652_21#_c_805_n 0.00782494f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_294_n N_A_652_21#_c_797_n 0.0132853f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_296_n N_A_652_21#_c_797_n 0.0121054f $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_311_n N_SET_B_M1033_g 0.00205491f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_294_n N_SET_B_c_917_n 0.00399047f $X=4.965 $Y=1.655 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_295_n N_SET_B_c_917_n 0.0300923f $X=5.82 $Y=0.81 $X2=0 $Y2=0
cc_371 N_A_27_47#_c_296_n N_SET_B_c_917_n 0.00574094f $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_297_n N_SET_B_c_917_n 0.0167082f $X=5.985 $Y=0.81 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_294_n N_A_476_47#_c_1044_n 2.94773e-19 $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_311_n N_A_476_47#_M1023_g 0.00187886f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_294_n N_A_476_47#_c_1045_n 0.00469727f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_295_n N_A_476_47#_c_1045_n 0.0078216f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_296_n N_A_476_47#_c_1045_n 0.00630303f $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_317_n N_A_476_47#_c_1045_n 0.00228498f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_311_n N_A_476_47#_M1017_g 0.00301713f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_317_n N_A_476_47#_M1017_g 0.0626672f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_318_n N_A_476_47#_M1017_g 0.00172662f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_295_n N_A_476_47#_c_1046_n 0.00414107f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_M1039_g N_A_476_47#_c_1070_n 0.0090453f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_384 N_A_27_47#_c_311_n N_A_476_47#_c_1070_n 0.00517144f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_385 N_A_27_47#_c_312_n N_A_476_47#_c_1070_n 0.00306479f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_386 N_A_27_47#_c_315_n N_A_476_47#_c_1070_n 0.00186639f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_387 N_A_27_47#_c_316_n N_A_476_47#_c_1070_n 0.015267f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_292_n N_A_476_47#_c_1075_n 0.00676006f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_389 N_A_27_47#_c_293_n N_A_476_47#_c_1075_n 9.25786e-19 $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_M1039_g N_A_476_47#_c_1055_n 0.00650943f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_292_n N_A_476_47#_c_1055_n 0.00666284f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_392 N_A_27_47#_c_311_n N_A_476_47#_c_1055_n 0.013911f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_312_n N_A_476_47#_c_1055_n 0.00145075f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_394 N_A_27_47#_c_315_n N_A_476_47#_c_1055_n 0.00203066f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_c_316_n N_A_476_47#_c_1055_n 0.0283088f $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_311_n N_A_476_47#_c_1049_n 0.00472657f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_292_n N_A_476_47#_c_1050_n 0.007273f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_311_n N_A_476_47#_c_1050_n 0.00456576f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_399 N_A_27_47#_c_311_n N_A_476_47#_c_1051_n 0.00248872f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_294_n N_A_476_47#_c_1052_n 0.00640057f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_311_n N_A_476_47#_c_1052_n 0.00148193f $X=5.145 $Y=1.87
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_297_n N_A_1178_261#_M1016_g 8.41348e-19 $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_300_n N_A_1178_261#_M1016_g 0.0627906f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_297_n N_A_1178_261#_c_1201_n 3.96308e-19 $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_298_n N_A_1178_261#_c_1201_n 0.0149285f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_M1003_g N_A_1028_413#_c_1302_n 0.00493733f $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_313_n N_A_1028_413#_c_1302_n 0.00403604f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_317_n N_A_1028_413#_c_1302_n 9.00165e-19 $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_318_n N_A_1028_413#_c_1302_n 0.0148431f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_294_n N_A_1028_413#_c_1294_n 0.00537793f $X=4.965 $Y=1.655
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_313_n N_A_1028_413#_c_1294_n 0.00776519f $X=5.29 $Y=1.87
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_317_n N_A_1028_413#_c_1294_n 4.1977e-19 $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_318_n N_A_1028_413#_c_1294_n 0.0211547f $X=5.155 $Y=1.74
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_295_n N_A_1028_413#_c_1310_n 0.00680222f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_415 N_A_27_47#_c_297_n N_A_1028_413#_c_1310_n 0.0126727f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_298_n N_A_1028_413#_c_1310_n 5.72459e-19 $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_417 N_A_27_47#_c_300_n N_A_1028_413#_c_1310_n 0.00790984f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_418 N_A_27_47#_c_295_n N_A_1028_413#_c_1284_n 0.00259385f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_c_297_n N_A_1028_413#_c_1284_n 0.0183126f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_420 N_A_27_47#_c_298_n N_A_1028_413#_c_1284_n 0.00247612f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_c_295_n N_A_1028_413#_c_1285_n 0.00570635f $X=5.82 $Y=0.81
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_297_n N_A_1028_413#_c_1286_n 0.0218685f $X=5.985 $Y=0.81
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_298_n N_A_1028_413#_c_1286_n 0.00156489f $X=5.985 $Y=0.93
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_300_n N_A_1028_413#_c_1286_n 0.00248854f $X=5.985 $Y=0.765
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_M1003_g N_A_1028_413#_c_1298_n 0.0010081f $X=5.065 $Y=2.275
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_416_p N_VPWR_M1019_d 6.91013e-19 $X=0.725 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_427 N_A_27_47#_c_310_n N_VPWR_M1019_d 0.00191833f $X=0.845 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_428 N_A_27_47#_M1000_g N_VPWR_c_1569_n 0.00827983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_304_n N_VPWR_c_1569_n 0.00346402f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_416_p N_VPWR_c_1569_n 0.0133497f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_c_308_n N_VPWR_c_1569_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_310_n N_VPWR_c_1569_n 0.00355334f $X=0.845 $Y=1.87 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_M1000_g N_VPWR_c_1570_n 0.00190407f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_309_n N_VPWR_c_1570_n 0.00166908f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_M1003_g N_VPWR_c_1572_n 0.0019199f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_311_n N_VPWR_c_1572_n 0.001212f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_437 N_A_27_47#_c_304_n N_VPWR_c_1577_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_438 N_A_27_47#_c_308_n N_VPWR_c_1577_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_439 N_A_27_47#_M1000_g N_VPWR_c_1578_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_M1039_g N_VPWR_c_1579_n 0.00367119f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_M1003_g N_VPWR_c_1580_n 0.00427125f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_318_n N_VPWR_c_1580_n 0.0032218f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_M1000_g N_VPWR_c_1568_n 0.00534566f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_M1039_g N_VPWR_c_1568_n 0.00563088f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_M1003_g N_VPWR_c_1568_n 0.00577339f $X=5.065 $Y=2.275 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_c_304_n N_VPWR_c_1568_n 0.00397874f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_308_n N_VPWR_c_1568_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_309_n N_VPWR_c_1568_n 0.072227f $X=2.385 $Y=1.87 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_310_n N_VPWR_c_1568_n 0.0144765f $X=0.845 $Y=1.87 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_311_n N_VPWR_c_1568_n 0.111929f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_451 N_A_27_47#_c_312_n N_VPWR_c_1568_n 0.0160044f $X=2.675 $Y=1.87 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_313_n N_VPWR_c_1568_n 0.016077f $X=5.29 $Y=1.87 $X2=0 $Y2=0
cc_453 N_A_27_47#_c_316_n N_VPWR_c_1568_n 2.46058e-19 $X=2.765 $Y=1.74 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_318_n N_VPWR_c_1568_n 0.00246615f $X=5.155 $Y=1.74 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_311_n N_VPWR_c_1589_n 0.0014214f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_309_n N_A_381_47#_M1028_d 8.84929e-19 $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_288_n N_A_381_47#_c_1768_n 0.00223782f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_458 N_A_27_47#_c_292_n N_A_381_47#_c_1768_n 0.00713576f $X=2.435 $Y=0.87
+ $X2=0 $Y2=0
cc_459 N_A_27_47#_c_309_n N_A_381_47#_c_1770_n 0.019313f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_309_n N_A_381_47#_c_1766_n 0.0157335f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_288_n N_A_381_47#_c_1772_n 0.00399753f $X=2.305 $Y=0.705
+ $X2=0 $Y2=0
cc_462 N_A_27_47#_c_309_n N_A_381_47#_c_1773_n 0.0109514f $X=2.385 $Y=1.87 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_312_n N_A_381_47#_c_1773_n 0.00146426f $X=2.675 $Y=1.87
+ $X2=0 $Y2=0
cc_464 N_A_27_47#_c_316_n N_A_381_47#_c_1773_n 0.00827001f $X=2.765 $Y=1.74
+ $X2=0 $Y2=0
cc_465 N_A_27_47#_c_289_n N_VGND_M1036_d 0.00164712f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_466 N_A_27_47#_M1022_g N_VGND_c_1907_n 0.0078844f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_289_n N_VGND_c_1907_n 0.0170164f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_468 N_A_27_47#_c_299_n N_VGND_c_1907_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_M1022_g N_VGND_c_1908_n 0.00296522f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_288_n N_VGND_c_1908_n 0.00120909f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_295_n N_VGND_c_1910_n 0.0017326f $X=5.82 $Y=0.81 $X2=0 $Y2=0
cc_472 N_A_27_47#_c_296_n N_VGND_c_1910_n 0.0129707f $X=5.05 $Y=0.81 $X2=0 $Y2=0
cc_473 N_A_27_47#_c_543_p N_VGND_c_1914_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_289_n N_VGND_c_1914_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_M1022_g N_VGND_c_1915_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_288_n N_VGND_c_1916_n 0.00556304f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_292_n N_VGND_c_1916_n 0.00113905f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_293_n N_VGND_c_1916_n 2.48118e-19 $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_M1036_s N_VGND_c_1922_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_M1022_g N_VGND_c_1922_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_288_n N_VGND_c_1922_n 0.00678262f $X=2.305 $Y=0.705 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_543_p N_VGND_c_1922_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_289_n N_VGND_c_1922_n 0.00578908f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_c_292_n N_VGND_c_1922_n 0.00122477f $X=2.435 $Y=0.87 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_295_n N_VGND_c_1922_n 0.00615621f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_296_n N_VGND_c_1922_n 4.92512e-19 $X=5.05 $Y=0.81 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_c_300_n N_VGND_c_1922_n 0.00522127f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_295_n N_VGND_c_1927_n 0.00797153f $X=5.82 $Y=0.81 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_c_300_n N_VGND_c_1927_n 0.00368123f $X=5.985 $Y=0.765 $X2=0
+ $Y2=0
cc_490 N_D_M1028_g N_A_193_47#_c_600_n 0.0303627f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_491 N_D_c_561_n N_A_193_47#_c_600_n 0.00467503f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_492 N_D_c_562_n N_A_193_47#_c_600_n 0.00330794f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_493 N_D_M1008_g N_A_193_47#_c_606_n 0.00395556f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_494 N_D_c_561_n N_A_193_47#_c_606_n 8.88354e-19 $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_495 N_D_c_562_n N_A_193_47#_c_606_n 0.0127149f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_496 N_D_M1008_g N_A_193_47#_c_616_n 0.00372305f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_497 N_D_M1028_g N_A_193_47#_c_616_n 0.00471318f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_498 N_D_M1028_g N_VPWR_c_1570_n 0.0116766f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_499 N_D_M1028_g N_VPWR_c_1579_n 0.0035268f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_500 N_D_M1028_g N_VPWR_c_1568_n 0.00402871f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_501 N_D_M1008_g N_A_381_47#_c_1763_n 0.00557005f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_502 N_D_M1028_g N_A_381_47#_c_1763_n 0.0115166f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_503 N_D_c_561_n N_A_381_47#_c_1763_n 0.00753248f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_504 N_D_c_562_n N_A_381_47#_c_1763_n 0.0473419f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_505 N_D_M1008_g N_A_381_47#_c_1768_n 0.0126635f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_506 N_D_c_561_n N_A_381_47#_c_1768_n 0.0014463f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_507 N_D_c_562_n N_A_381_47#_c_1768_n 0.0217898f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_508 N_D_M1028_g N_A_381_47#_c_1770_n 0.011823f $X=1.83 $Y=2.065 $X2=0 $Y2=0
cc_509 N_D_c_562_n N_A_381_47#_c_1770_n 0.0109323f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_510 N_D_c_562_n N_A_381_47#_c_1773_n 0.0137404f $X=1.855 $Y=1.17 $X2=0 $Y2=0
cc_511 N_D_M1008_g N_VGND_c_1908_n 0.00942273f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_512 N_D_M1008_g N_VGND_c_1916_n 0.00339367f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_513 N_D_M1008_g N_VGND_c_1922_n 0.00393034f $X=1.83 $Y=0.555 $X2=0 $Y2=0
cc_514 N_A_193_47#_M1020_g N_A_652_21#_M1025_g 0.024565f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_515 N_A_193_47#_c_602_n N_A_652_21#_M1025_g 0.0114519f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_516 N_A_193_47#_c_609_n N_A_652_21#_M1025_g 9.99732e-19 $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_517 N_A_193_47#_c_611_n N_A_652_21#_M1025_g 0.00631121f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_518 N_A_193_47#_c_612_n N_A_652_21#_M1025_g 0.00191013f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_519 N_A_193_47#_c_615_n N_A_652_21#_M1025_g 0.0200607f $X=2.915 $Y=0.93 $X2=0
+ $Y2=0
cc_520 N_A_193_47#_c_609_n N_A_652_21#_c_800_n 5.47854e-19 $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_521 N_A_193_47#_c_609_n N_A_652_21#_c_801_n 0.00115455f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_522 N_A_193_47#_c_609_n N_A_652_21#_c_796_n 0.0140676f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_523 N_A_193_47#_c_609_n N_A_652_21#_c_803_n 8.37667e-19 $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_524 N_A_193_47#_c_609_n N_A_652_21#_c_797_n 0.00655125f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_525 N_A_193_47#_c_609_n N_SET_B_c_909_n 0.00381498f $X=5.165 $Y=1.19
+ $X2=-0.19 $Y2=-0.24
cc_526 N_A_193_47#_c_609_n N_SET_B_M1033_g 0.00121673f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_527 N_A_193_47#_c_609_n SET_B 0.00570533f $X=5.165 $Y=1.19 $X2=0 $Y2=0
cc_528 N_A_193_47#_M1012_g N_SET_B_c_917_n 0.00419104f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_529 N_A_193_47#_c_605_n N_SET_B_c_917_n 0.00120258f $X=5.47 $Y=1.26 $X2=0
+ $Y2=0
cc_530 N_A_193_47#_c_609_n N_SET_B_c_917_n 0.0878379f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_531 N_A_193_47#_c_613_n N_SET_B_c_917_n 0.02693f $X=5.31 $Y=1.19 $X2=0 $Y2=0
cc_532 N_A_193_47#_c_614_n N_SET_B_c_917_n 0.00112669f $X=5.31 $Y=1.19 $X2=0
+ $Y2=0
cc_533 N_A_193_47#_c_609_n N_SET_B_c_918_n 0.0263312f $X=5.165 $Y=1.19 $X2=0
+ $Y2=0
cc_534 N_A_193_47#_c_609_n N_A_476_47#_c_1044_n 0.00253485f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_535 N_A_193_47#_c_605_n N_A_476_47#_c_1045_n 0.00912806f $X=5.47 $Y=1.26
+ $X2=0 $Y2=0
cc_536 N_A_193_47#_c_609_n N_A_476_47#_c_1045_n 0.00101093f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_537 N_A_193_47#_c_614_n N_A_476_47#_c_1045_n 3.19592e-19 $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_538 N_A_193_47#_M1012_g N_A_476_47#_c_1046_n 0.0518139f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_539 N_A_193_47#_M1009_g N_A_476_47#_c_1070_n 0.00278769f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_540 N_A_193_47#_M1020_g N_A_476_47#_c_1075_n 0.008828f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_541 N_A_193_47#_c_606_n N_A_476_47#_c_1075_n 0.00573977f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_542 N_A_193_47#_c_611_n N_A_476_47#_c_1075_n 0.00194059f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_543 N_A_193_47#_c_612_n N_A_476_47#_c_1075_n 0.0194974f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_544 N_A_193_47#_c_615_n N_A_476_47#_c_1075_n 5.24271e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_545 N_A_193_47#_M1009_g N_A_476_47#_c_1055_n 8.73767e-19 $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_546 N_A_193_47#_c_610_n N_A_476_47#_c_1055_n 3.07745e-19 $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_547 N_A_193_47#_M1020_g N_A_476_47#_c_1048_n 0.00118778f $X=2.855 $Y=0.415
+ $X2=0 $Y2=0
cc_548 N_A_193_47#_c_602_n N_A_476_47#_c_1048_n 7.74259e-19 $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_549 N_A_193_47#_c_609_n N_A_476_47#_c_1048_n 0.0146154f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_550 N_A_193_47#_c_611_n N_A_476_47#_c_1048_n 0.0134967f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_551 N_A_193_47#_c_612_n N_A_476_47#_c_1048_n 0.0244992f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_552 N_A_193_47#_c_615_n N_A_476_47#_c_1048_n 7.73887e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_553 N_A_193_47#_c_609_n N_A_476_47#_c_1049_n 0.0232188f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_554 N_A_193_47#_c_602_n N_A_476_47#_c_1050_n 0.00262762f $X=2.855 $Y=1.245
+ $X2=0 $Y2=0
cc_555 N_A_193_47#_c_609_n N_A_476_47#_c_1050_n 0.0121342f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_556 N_A_193_47#_c_610_n N_A_476_47#_c_1050_n 0.00535278f $X=3.135 $Y=1.19
+ $X2=0 $Y2=0
cc_557 N_A_193_47#_c_612_n N_A_476_47#_c_1050_n 0.00527199f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_558 N_A_193_47#_c_615_n N_A_476_47#_c_1050_n 5.70501e-19 $X=2.915 $Y=0.93
+ $X2=0 $Y2=0
cc_559 N_A_193_47#_c_609_n N_A_476_47#_c_1051_n 0.00996075f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_560 N_A_193_47#_c_604_n N_A_476_47#_c_1052_n 5.76045e-19 $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_561 N_A_193_47#_c_605_n N_A_476_47#_c_1052_n 0.00482213f $X=5.47 $Y=1.26
+ $X2=0 $Y2=0
cc_562 N_A_193_47#_c_609_n N_A_476_47#_c_1052_n 0.00412912f $X=5.165 $Y=1.19
+ $X2=0 $Y2=0
cc_563 N_A_193_47#_M1012_g N_A_1178_261#_M1016_g 0.00243301f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_564 N_A_193_47#_c_604_n N_A_1178_261#_c_1201_n 0.0407126f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_565 N_A_193_47#_M1030_g N_A_1178_261#_c_1206_n 0.0407126f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_566 N_A_193_47#_M1030_g N_A_1028_413#_c_1302_n 0.00768489f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_567 N_A_193_47#_c_604_n N_A_1028_413#_c_1294_n 0.00103911f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_568 N_A_193_47#_M1030_g N_A_1028_413#_c_1294_n 0.0101662f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_569 N_A_193_47#_c_614_n N_A_1028_413#_c_1294_n 0.00496139f $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_570 N_A_193_47#_c_604_n N_A_1028_413#_c_1285_n 0.00827976f $X=5.605 $Y=1.455
+ $X2=0 $Y2=0
cc_571 N_A_193_47#_c_613_n N_A_1028_413#_c_1285_n 0.00200974f $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_572 N_A_193_47#_c_614_n N_A_1028_413#_c_1285_n 0.0123133f $X=5.31 $Y=1.19
+ $X2=0 $Y2=0
cc_573 N_A_193_47#_M1030_g N_A_1028_413#_c_1296_n 2.49577e-19 $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_574 N_A_193_47#_M1012_g N_A_1028_413#_c_1286_n 0.002035f $X=5.565 $Y=0.445
+ $X2=0 $Y2=0
cc_575 N_A_193_47#_M1030_g N_A_1028_413#_c_1298_n 0.011666f $X=5.605 $Y=2.275
+ $X2=0 $Y2=0
cc_576 N_A_193_47#_c_616_n N_VPWR_c_1569_n 0.0127357f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_577 N_A_193_47#_M1009_g N_VPWR_c_1570_n 0.00113058f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_578 N_A_193_47#_c_616_n N_VPWR_c_1570_n 0.0226552f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_579 N_A_193_47#_c_616_n N_VPWR_c_1578_n 0.015988f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_580 N_A_193_47#_M1009_g N_VPWR_c_1579_n 0.00541732f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_581 N_A_193_47#_M1030_g N_VPWR_c_1580_n 0.00369426f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_582 N_A_193_47#_M1009_g N_VPWR_c_1568_n 0.00628966f $X=2.315 $Y=2.275 $X2=0
+ $Y2=0
cc_583 N_A_193_47#_M1030_g N_VPWR_c_1568_n 0.00544628f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_584 N_A_193_47#_c_616_n N_VPWR_c_1568_n 0.00409094f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_585 N_A_193_47#_M1030_g N_VPWR_c_1591_n 0.00197636f $X=5.605 $Y=2.275 $X2=0
+ $Y2=0
cc_586 N_A_193_47#_c_606_n N_A_381_47#_M1008_d 4.25819e-19 $X=2.845 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_587 N_A_193_47#_c_606_n N_A_381_47#_c_1763_n 0.0148354f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_588 N_A_193_47#_c_607_n N_A_381_47#_c_1763_n 0.00135406f $X=1.295 $Y=0.85
+ $X2=0 $Y2=0
cc_589 N_A_193_47#_c_616_n N_A_381_47#_c_1763_n 0.0675462f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_590 N_A_193_47#_c_606_n N_A_381_47#_c_1768_n 0.0198802f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_591 N_A_193_47#_c_612_n N_A_381_47#_c_1768_n 0.00201969f $X=2.99 $Y=0.85
+ $X2=0 $Y2=0
cc_592 N_A_193_47#_c_606_n N_A_381_47#_c_1764_n 0.00435863f $X=2.845 $Y=0.85
+ $X2=0 $Y2=0
cc_593 N_A_193_47#_c_607_n N_A_381_47#_c_1764_n 0.00140429f $X=1.295 $Y=0.85
+ $X2=0 $Y2=0
cc_594 N_A_193_47#_c_616_n N_A_381_47#_c_1764_n 0.0138352f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_595 N_A_193_47#_c_616_n N_A_381_47#_c_1766_n 0.0114327f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_596 N_A_193_47#_M1009_g N_A_381_47#_c_1773_n 0.0102511f $X=2.315 $Y=2.275
+ $X2=0 $Y2=0
cc_597 N_A_193_47#_c_606_n N_VGND_c_1908_n 0.0012296f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_598 N_A_193_47#_c_616_n N_VGND_c_1908_n 0.00823827f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_599 N_A_193_47#_c_616_n N_VGND_c_1915_n 0.00978627f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_600 N_A_193_47#_M1020_g N_VGND_c_1916_n 0.00359964f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_601 N_A_193_47#_M1022_d N_VGND_c_1922_n 0.00324958f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_A_193_47#_M1020_g N_VGND_c_1922_n 0.0056346f $X=2.855 $Y=0.415 $X2=0
+ $Y2=0
cc_603 N_A_193_47#_M1012_g N_VGND_c_1922_n 0.00571363f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_604 N_A_193_47#_c_606_n N_VGND_c_1922_n 0.072327f $X=2.845 $Y=0.85 $X2=0
+ $Y2=0
cc_605 N_A_193_47#_c_607_n N_VGND_c_1922_n 0.0151383f $X=1.295 $Y=0.85 $X2=0
+ $Y2=0
cc_606 N_A_193_47#_c_611_n N_VGND_c_1922_n 0.0151785f $X=2.99 $Y=0.85 $X2=0
+ $Y2=0
cc_607 N_A_193_47#_c_616_n N_VGND_c_1922_n 0.00372614f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_608 N_A_193_47#_M1012_g N_VGND_c_1927_n 0.00437852f $X=5.565 $Y=0.445 $X2=0
+ $Y2=0
cc_609 N_A_193_47#_c_612_n A_586_47# 0.00109469f $X=2.99 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_610 N_A_652_21#_M1025_g N_SET_B_c_909_n 0.0189903f $X=3.335 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_611 N_A_652_21#_c_796_n N_SET_B_c_909_n 7.60504e-19 $X=4.625 $Y=1.835
+ $X2=-0.19 $Y2=-0.24
cc_612 N_A_652_21#_M1025_g N_SET_B_M1033_g 0.0137896f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_613 N_A_652_21#_M1007_g N_SET_B_M1033_g 0.0113783f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_614 N_A_652_21#_c_800_n N_SET_B_M1033_g 0.0139954f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_615 N_A_652_21#_c_803_n N_SET_B_M1033_g 0.00563707f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_616 N_A_652_21#_c_804_n N_SET_B_M1033_g 0.0201938f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_617 N_A_652_21#_M1025_g N_SET_B_M1002_g 0.0141659f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_618 N_A_652_21#_c_795_n N_SET_B_M1002_g 0.00124922f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_619 N_A_652_21#_c_797_n N_SET_B_M1002_g 3.79232e-19 $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_620 N_A_652_21#_M1025_g SET_B 0.00110794f $X=3.335 $Y=0.445 $X2=0 $Y2=0
cc_621 N_A_652_21#_c_797_n SET_B 0.0144281f $X=4.625 $Y=0.895 $X2=0 $Y2=0
cc_622 N_A_652_21#_c_795_n N_SET_B_c_917_n 9.52814e-19 $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_623 N_A_652_21#_c_797_n N_SET_B_c_917_n 0.0196649f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_624 N_A_652_21#_c_797_n N_SET_B_c_918_n 0.00250762f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_625 N_A_652_21#_c_795_n N_A_476_47#_c_1043_n 0.00809901f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_626 N_A_652_21#_c_797_n N_A_476_47#_c_1043_n 4.65467e-19 $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_627 N_A_652_21#_c_796_n N_A_476_47#_c_1044_n 0.00246574f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_628 N_A_652_21#_c_797_n N_A_476_47#_c_1044_n 0.0035345f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_629 N_A_652_21#_c_801_n N_A_476_47#_M1023_g 0.0138123f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_630 N_A_652_21#_c_796_n N_A_476_47#_M1023_g 0.00531645f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_631 N_A_652_21#_c_795_n N_A_476_47#_c_1045_n 0.00253676f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_632 N_A_652_21#_c_796_n N_A_476_47#_c_1045_n 2.06235e-19 $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_633 N_A_652_21#_c_797_n N_A_476_47#_c_1045_n 0.0148491f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_634 N_A_652_21#_c_801_n N_A_476_47#_M1017_g 0.00844681f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_635 N_A_652_21#_c_796_n N_A_476_47#_M1017_g 0.00507438f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_636 N_A_652_21#_c_795_n N_A_476_47#_c_1046_n 0.00422581f $X=4.475 $Y=0.46
+ $X2=0 $Y2=0
cc_637 N_A_652_21#_c_797_n N_A_476_47#_c_1047_n 0.00182302f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_638 N_A_652_21#_M1007_g N_A_476_47#_c_1070_n 0.00202046f $X=3.335 $Y=2.275
+ $X2=0 $Y2=0
cc_639 N_A_652_21#_M1025_g N_A_476_47#_c_1075_n 0.00854236f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_640 N_A_652_21#_M1025_g N_A_476_47#_c_1055_n 0.015293f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_641 N_A_652_21#_c_803_n N_A_476_47#_c_1055_n 0.0366983f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_642 N_A_652_21#_M1025_g N_A_476_47#_c_1048_n 0.0188229f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_643 N_A_652_21#_c_800_n N_A_476_47#_c_1049_n 0.00881126f $X=3.99 $Y=1.96
+ $X2=0 $Y2=0
cc_644 N_A_652_21#_c_805_n N_A_476_47#_c_1049_n 0.00337624f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_645 N_A_652_21#_M1025_g N_A_476_47#_c_1050_n 0.0109017f $X=3.335 $Y=0.445
+ $X2=0 $Y2=0
cc_646 N_A_652_21#_c_803_n N_A_476_47#_c_1050_n 0.0171213f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_647 N_A_652_21#_c_804_n N_A_476_47#_c_1050_n 0.0011995f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_648 N_A_652_21#_c_801_n N_A_476_47#_c_1051_n 0.0079382f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_649 N_A_652_21#_c_796_n N_A_476_47#_c_1051_n 0.0229291f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_650 N_A_652_21#_c_805_n N_A_476_47#_c_1051_n 0.00169427f $X=4.075 $Y=1.96
+ $X2=0 $Y2=0
cc_651 N_A_652_21#_c_797_n N_A_476_47#_c_1051_n 0.0037745f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_652 N_A_652_21#_c_801_n N_A_476_47#_c_1052_n 0.0029883f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_653 N_A_652_21#_c_796_n N_A_476_47#_c_1052_n 0.0130643f $X=4.625 $Y=1.835
+ $X2=0 $Y2=0
cc_654 N_A_652_21#_c_797_n N_A_476_47#_c_1052_n 0.00437877f $X=4.625 $Y=0.895
+ $X2=0 $Y2=0
cc_655 N_A_652_21#_c_800_n N_VPWR_M1007_d 0.00131929f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_656 N_A_652_21#_c_803_n N_VPWR_M1007_d 0.00154452f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_657 N_A_652_21#_c_801_n N_VPWR_M1023_d 0.00161389f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_658 N_A_652_21#_c_800_n N_VPWR_c_1571_n 0.00266175f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_659 N_A_652_21#_c_884_p N_VPWR_c_1571_n 0.0070924f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_660 N_A_652_21#_c_801_n N_VPWR_c_1571_n 0.00248431f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_661 N_A_652_21#_c_801_n N_VPWR_c_1572_n 0.0155298f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_662 N_A_652_21#_M1007_g N_VPWR_c_1579_n 0.00532975f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_663 N_A_652_21#_c_803_n N_VPWR_c_1579_n 0.00105935f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_664 N_A_652_21#_c_801_n N_VPWR_c_1580_n 8.80252e-19 $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_665 N_A_652_21#_M1033_d N_VPWR_c_1568_n 0.00202389f $X=3.94 $Y=2.065 $X2=0
+ $Y2=0
cc_666 N_A_652_21#_M1007_g N_VPWR_c_1568_n 0.0066225f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_667 N_A_652_21#_c_800_n N_VPWR_c_1568_n 0.00255051f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_668 N_A_652_21#_c_884_p N_VPWR_c_1568_n 0.00288476f $X=4.075 $Y=2.21 $X2=0
+ $Y2=0
cc_669 N_A_652_21#_c_801_n N_VPWR_c_1568_n 0.0034475f $X=4.54 $Y=1.96 $X2=0
+ $Y2=0
cc_670 N_A_652_21#_c_803_n N_VPWR_c_1568_n 0.00138626f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_671 N_A_652_21#_M1007_g N_VPWR_c_1589_n 0.00326498f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_672 N_A_652_21#_c_800_n N_VPWR_c_1589_n 0.0101842f $X=3.99 $Y=1.96 $X2=0
+ $Y2=0
cc_673 N_A_652_21#_c_803_n N_VPWR_c_1589_n 0.0109284f $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_674 N_A_652_21#_c_804_n N_VPWR_c_1589_n 6.81742e-19 $X=3.445 $Y=1.74 $X2=0
+ $Y2=0
cc_675 N_A_652_21#_M1025_g N_VGND_c_1909_n 0.0040279f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_676 N_A_652_21#_c_795_n N_VGND_c_1910_n 0.0192612f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_677 N_A_652_21#_M1025_g N_VGND_c_1916_n 0.0035977f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_678 N_A_652_21#_c_795_n N_VGND_c_1917_n 0.0118981f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_679 N_A_652_21#_c_797_n N_VGND_c_1917_n 0.00244068f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_680 N_A_652_21#_M1005_d N_VGND_c_1922_n 0.00186029f $X=4.34 $Y=0.235 $X2=0
+ $Y2=0
cc_681 N_A_652_21#_M1025_g N_VGND_c_1922_n 0.00580574f $X=3.335 $Y=0.445 $X2=0
+ $Y2=0
cc_682 N_A_652_21#_c_795_n N_VGND_c_1922_n 0.00426169f $X=4.475 $Y=0.46 $X2=0
+ $Y2=0
cc_683 N_A_652_21#_c_797_n N_VGND_c_1922_n 0.00183644f $X=4.625 $Y=0.895 $X2=0
+ $Y2=0
cc_684 N_SET_B_M1002_g N_A_476_47#_c_1043_n 0.0270653f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_909_n N_A_476_47#_c_1044_n 0.0146844f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_917_n N_A_476_47#_c_1044_n 8.12862e-19 $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_918_n N_A_476_47#_c_1044_n 7.28461e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_688 N_SET_B_M1033_g N_A_476_47#_M1023_g 0.0336841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_917_n N_A_476_47#_c_1045_n 0.00245454f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_909_n N_A_476_47#_c_1047_n 0.0270653f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_691 SET_B N_A_476_47#_c_1047_n 0.0021684f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_692 N_SET_B_c_917_n N_A_476_47#_c_1047_n 0.00277782f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_693 N_SET_B_c_918_n N_A_476_47#_c_1047_n 7.28461e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_909_n N_A_476_47#_c_1048_n 0.00218199f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_695 N_SET_B_M1033_g N_A_476_47#_c_1048_n 6.04572e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_696 N_SET_B_M1002_g N_A_476_47#_c_1048_n 0.00184201f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_697 SET_B N_A_476_47#_c_1048_n 0.0243988f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_698 N_SET_B_c_918_n N_A_476_47#_c_1048_n 0.00116251f $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_909_n N_A_476_47#_c_1049_n 0.00307815f $X=3.865 $Y=1.145 $X2=0
+ $Y2=0
cc_700 N_SET_B_M1033_g N_A_476_47#_c_1049_n 0.0103672f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_701 SET_B N_A_476_47#_c_1049_n 0.0263655f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_702 N_SET_B_c_917_n N_A_476_47#_c_1049_n 3.66303e-19 $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_918_n N_A_476_47#_c_1049_n 5.23607e-19 $X=4.055 $Y=0.85 $X2=0
+ $Y2=0
cc_704 N_SET_B_M1033_g N_A_476_47#_c_1050_n 5.20457e-19 $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_705 N_SET_B_M1033_g N_A_476_47#_c_1051_n 0.00354841f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_917_n N_A_476_47#_c_1051_n 0.00236582f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_707 N_SET_B_M1033_g N_A_476_47#_c_1052_n 0.0205296f $X=3.865 $Y=2.275 $X2=0
+ $Y2=0
cc_708 N_SET_B_M1021_g N_A_1178_261#_M1016_g 0.0658096f $X=6.765 $Y=0.445 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_913_n N_A_1178_261#_M1016_g 0.0116464f $X=6.895 $Y=1.535 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_915_n N_A_1178_261#_M1016_g 0.00104156f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_711 N_SET_B_M1001_g N_A_1178_261#_c_1206_n 0.00284189f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_712 N_SET_B_c_924_n N_A_1178_261#_c_1206_n 0.00234806f $X=6.895 $Y=1.685
+ $X2=0 $Y2=0
cc_713 N_SET_B_c_913_n N_A_1178_261#_c_1207_n 0.00234806f $X=6.895 $Y=1.535
+ $X2=0 $Y2=0
cc_714 N_SET_B_c_914_n N_A_1178_261#_c_1202_n 2.40292e-19 $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_915_n N_A_1178_261#_c_1202_n 0.00184604f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_919_n N_A_1178_261#_c_1202_n 0.00147872f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_717 N_SET_B_c_920_n N_A_1178_261#_c_1202_n 0.0116605f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_718 N_SET_B_M1001_g N_A_1178_261#_c_1209_n 0.00936381f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_719 N_SET_B_c_924_n N_A_1178_261#_c_1209_n 0.00778928f $X=6.895 $Y=1.685
+ $X2=0 $Y2=0
cc_720 N_SET_B_M1021_g N_A_1028_413#_M1018_g 0.0164357f $X=6.765 $Y=0.445 $X2=0
+ $Y2=0
cc_721 N_SET_B_c_914_n N_A_1028_413#_M1018_g 0.00943035f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_722 N_SET_B_c_915_n N_A_1028_413#_M1018_g 5.48549e-19 $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_920_n N_A_1028_413#_M1018_g 0.00790355f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_913_n N_A_1028_413#_M1027_g 0.00412516f $X=6.895 $Y=1.535 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_924_n N_A_1028_413#_M1027_g 0.0260901f $X=6.895 $Y=1.685 $X2=0
+ $Y2=0
cc_726 N_SET_B_c_917_n N_A_1028_413#_c_1310_n 0.00655755f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_727 N_SET_B_c_917_n N_A_1028_413#_c_1284_n 0.010616f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_728 N_SET_B_c_917_n N_A_1028_413#_c_1285_n 0.00391758f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_729 N_SET_B_M1001_g N_A_1028_413#_c_1296_n 0.00433068f $X=6.905 $Y=2.275
+ $X2=0 $Y2=0
cc_730 N_SET_B_M1021_g N_A_1028_413#_c_1286_n 0.00258467f $X=6.765 $Y=0.445
+ $X2=0 $Y2=0
cc_731 N_SET_B_c_913_n N_A_1028_413#_c_1286_n 0.00102632f $X=6.895 $Y=1.535
+ $X2=0 $Y2=0
cc_732 N_SET_B_c_914_n N_A_1028_413#_c_1286_n 0.00158445f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_915_n N_A_1028_413#_c_1286_n 0.0254752f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_734 N_SET_B_c_917_n N_A_1028_413#_c_1286_n 0.0180658f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_735 N_SET_B_c_919_n N_A_1028_413#_c_1286_n 3.39847e-19 $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_736 N_SET_B_c_913_n N_A_1028_413#_c_1287_n 6.19496e-19 $X=6.895 $Y=1.535
+ $X2=0 $Y2=0
cc_737 N_SET_B_c_919_n N_A_1028_413#_c_1287_n 8.97025e-19 $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_738 N_SET_B_c_920_n N_A_1028_413#_c_1287_n 0.0128812f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_739 N_SET_B_c_914_n N_A_1028_413#_c_1288_n 0.0218378f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_740 N_SET_B_c_920_n N_A_1028_413#_c_1288_n 0.00349124f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_741 N_SET_B_c_913_n N_A_1028_413#_c_1289_n 0.0101835f $X=6.895 $Y=1.535 $X2=0
+ $Y2=0
cc_742 N_SET_B_c_924_n N_A_1028_413#_c_1289_n 5.5231e-19 $X=6.895 $Y=1.685 $X2=0
+ $Y2=0
cc_743 N_SET_B_c_914_n N_A_1028_413#_c_1289_n 0.00347344f $X=6.825 $Y=0.98 $X2=0
+ $Y2=0
cc_744 N_SET_B_c_915_n N_A_1028_413#_c_1289_n 0.0229264f $X=6.99 $Y=0.9 $X2=0
+ $Y2=0
cc_745 N_SET_B_c_917_n N_A_1028_413#_c_1289_n 0.00838415f $X=6.985 $Y=0.85 $X2=0
+ $Y2=0
cc_746 N_SET_B_c_919_n N_A_1028_413#_c_1289_n 0.00102488f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_747 N_SET_B_c_920_n N_A_1028_413#_c_1289_n 0.00830557f $X=7.13 $Y=0.85 $X2=0
+ $Y2=0
cc_748 N_SET_B_M1033_g N_VPWR_c_1571_n 0.00368415f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_749 N_SET_B_M1033_g N_VPWR_c_1572_n 7.26951e-19 $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_750 N_SET_B_M1001_g N_VPWR_c_1573_n 0.00327827f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_751 N_SET_B_M1001_g N_VPWR_c_1581_n 0.00585385f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_752 N_SET_B_M1033_g N_VPWR_c_1568_n 0.00406312f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_753 N_SET_B_M1001_g N_VPWR_c_1568_n 0.0121898f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_754 N_SET_B_M1033_g N_VPWR_c_1589_n 0.00699603f $X=3.865 $Y=2.275 $X2=0 $Y2=0
cc_755 N_SET_B_M1001_g N_VPWR_c_1591_n 0.00306764f $X=6.905 $Y=2.275 $X2=0 $Y2=0
cc_756 N_SET_B_c_919_n N_VGND_M1021_d 0.00132095f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_757 N_SET_B_c_920_n N_VGND_M1021_d 9.16065e-19 $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_758 N_SET_B_c_909_n N_VGND_c_1909_n 0.00103531f $X=3.865 $Y=1.145 $X2=0 $Y2=0
cc_759 N_SET_B_M1002_g N_VGND_c_1909_n 0.0134999f $X=3.905 $Y=0.445 $X2=0 $Y2=0
cc_760 SET_B N_VGND_c_1909_n 0.0213368f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_761 N_SET_B_c_918_n N_VGND_c_1909_n 0.00267196f $X=4.055 $Y=0.85 $X2=0 $Y2=0
cc_762 N_SET_B_c_917_n N_VGND_c_1910_n 0.00564413f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_763 N_SET_B_c_915_n N_VGND_c_1922_n 0.00105154f $X=6.99 $Y=0.9 $X2=0 $Y2=0
cc_764 SET_B N_VGND_c_1922_n 9.94995e-19 $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_765 N_SET_B_c_917_n N_VGND_c_1922_n 0.134751f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_766 N_SET_B_c_918_n N_VGND_c_1922_n 0.0146581f $X=4.055 $Y=0.85 $X2=0 $Y2=0
cc_767 N_SET_B_c_919_n N_VGND_c_1922_n 0.0145559f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_768 N_SET_B_M1021_g N_VGND_c_1928_n 0.0199195f $X=6.765 $Y=0.445 $X2=0 $Y2=0
cc_769 N_SET_B_c_914_n N_VGND_c_1928_n 6.12458e-19 $X=6.825 $Y=0.98 $X2=0 $Y2=0
cc_770 N_SET_B_c_915_n N_VGND_c_1928_n 0.0401429f $X=6.99 $Y=0.9 $X2=0 $Y2=0
cc_771 N_SET_B_c_917_n N_VGND_c_1928_n 0.00146726f $X=6.985 $Y=0.85 $X2=0 $Y2=0
cc_772 N_SET_B_c_919_n N_VGND_c_1928_n 0.00339972f $X=7.13 $Y=0.85 $X2=0 $Y2=0
cc_773 N_A_476_47#_M1017_g N_A_1028_413#_c_1302_n 8.84083e-19 $X=4.705 $Y=2.275
+ $X2=0 $Y2=0
cc_774 N_A_476_47#_M1023_g N_VPWR_c_1571_n 0.00339367f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_775 N_A_476_47#_M1023_g N_VPWR_c_1572_n 0.00730335f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_776 N_A_476_47#_M1017_g N_VPWR_c_1572_n 0.00909428f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_777 N_A_476_47#_c_1070_n N_VPWR_c_1579_n 0.0377433f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_778 N_A_476_47#_M1017_g N_VPWR_c_1580_n 0.00414121f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_779 N_A_476_47#_M1009_d N_VPWR_c_1568_n 0.00172638f $X=2.39 $Y=2.065 $X2=0
+ $Y2=0
cc_780 N_A_476_47#_M1023_g N_VPWR_c_1568_n 0.00379591f $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_781 N_A_476_47#_M1017_g N_VPWR_c_1568_n 0.00402125f $X=4.705 $Y=2.275 $X2=0
+ $Y2=0
cc_782 N_A_476_47#_c_1070_n N_VPWR_c_1568_n 0.0132505f $X=3.02 $Y=2.335 $X2=0
+ $Y2=0
cc_783 N_A_476_47#_M1023_g N_VPWR_c_1589_n 7.14614e-19 $X=4.285 $Y=2.275 $X2=0
+ $Y2=0
cc_784 N_A_476_47#_c_1070_n N_A_381_47#_c_1773_n 0.0102747f $X=3.02 $Y=2.335
+ $X2=0 $Y2=0
cc_785 N_A_476_47#_c_1070_n A_562_413# 0.00859792f $X=3.02 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_786 N_A_476_47#_c_1055_n A_562_413# 0.00578953f $X=3.105 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_787 N_A_476_47#_c_1043_n N_VGND_c_1909_n 0.00301834f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_788 N_A_476_47#_c_1043_n N_VGND_c_1910_n 0.00375773f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_789 N_A_476_47#_c_1045_n N_VGND_c_1910_n 0.00681053f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_790 N_A_476_47#_c_1046_n N_VGND_c_1910_n 0.00458594f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_791 N_A_476_47#_c_1075_n N_VGND_c_1916_n 0.055608f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_792 N_A_476_47#_c_1043_n N_VGND_c_1917_n 0.00541969f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_793 N_A_476_47#_c_1045_n N_VGND_c_1917_n 0.00110285f $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_794 N_A_476_47#_M1034_d N_VGND_c_1922_n 0.00275359f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_795 N_A_476_47#_c_1043_n N_VGND_c_1922_n 0.00742824f $X=4.265 $Y=0.735 $X2=0
+ $Y2=0
cc_796 N_A_476_47#_c_1045_n N_VGND_c_1922_n 3.98471e-19 $X=5.13 $Y=0.825 $X2=0
+ $Y2=0
cc_797 N_A_476_47#_c_1046_n N_VGND_c_1922_n 0.00674913f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_798 N_A_476_47#_c_1075_n N_VGND_c_1922_n 0.0223868f $X=3.27 $Y=0.365 $X2=0
+ $Y2=0
cc_799 N_A_476_47#_c_1046_n N_VGND_c_1927_n 0.00437852f $X=5.205 $Y=0.735 $X2=0
+ $Y2=0
cc_800 N_A_476_47#_c_1075_n A_586_47# 0.00628999f $X=3.27 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_801 N_A_1178_261#_c_1202_n N_A_1028_413#_M1018_g 0.00949399f $X=7.745
+ $Y=1.575 $X2=0 $Y2=0
cc_802 N_A_1178_261#_c_1202_n N_A_1028_413#_M1027_g 0.0051921f $X=7.745 $Y=1.575
+ $X2=0 $Y2=0
cc_803 N_A_1178_261#_c_1209_n N_A_1028_413#_M1027_g 0.0145117f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_804 N_A_1178_261#_c_1202_n N_A_1028_413#_c_1281_n 0.0244516f $X=7.745
+ $Y=1.575 $X2=0 $Y2=0
cc_805 N_A_1178_261#_c_1203_n N_A_1028_413#_c_1281_n 0.00339526f $X=7.745
+ $Y=0.515 $X2=0 $Y2=0
cc_806 N_A_1178_261#_c_1210_n N_A_1028_413#_c_1281_n 0.00462612f $X=7.745
+ $Y=1.67 $X2=0 $Y2=0
cc_807 N_A_1178_261#_c_1202_n N_A_1028_413#_M1006_g 0.00182119f $X=7.745
+ $Y=1.575 $X2=0 $Y2=0
cc_808 N_A_1178_261#_c_1203_n N_A_1028_413#_M1006_g 6.42828e-19 $X=7.745
+ $Y=0.515 $X2=0 $Y2=0
cc_809 N_A_1178_261#_c_1238_p N_A_1028_413#_M1011_g 0.00122441f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_810 N_A_1178_261#_c_1202_n N_A_1028_413#_M1011_g 6.52815e-19 $X=7.745
+ $Y=1.575 $X2=0 $Y2=0
cc_811 N_A_1178_261#_c_1210_n N_A_1028_413#_M1011_g 9.12076e-19 $X=7.745 $Y=1.67
+ $X2=0 $Y2=0
cc_812 N_A_1178_261#_c_1201_n N_A_1028_413#_c_1294_n 0.00400927f $X=6.405
+ $Y=1.38 $X2=0 $Y2=0
cc_813 N_A_1178_261#_c_1209_n N_A_1028_413#_c_1294_n 0.0133834f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_814 N_A_1178_261#_M1016_g N_A_1028_413#_c_1310_n 0.00576956f $X=6.405
+ $Y=0.445 $X2=0 $Y2=0
cc_815 N_A_1178_261#_c_1201_n N_A_1028_413#_c_1284_n 0.0140658f $X=6.405 $Y=1.38
+ $X2=0 $Y2=0
cc_816 N_A_1178_261#_c_1209_n N_A_1028_413#_c_1284_n 0.0281674f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_817 N_A_1178_261#_M1015_g N_A_1028_413#_c_1296_n 0.0119267f $X=5.965 $Y=2.275
+ $X2=0 $Y2=0
cc_818 N_A_1178_261#_c_1206_n N_A_1028_413#_c_1296_n 0.00460004f $X=6.05
+ $Y=1.825 $X2=0 $Y2=0
cc_819 N_A_1178_261#_c_1209_n N_A_1028_413#_c_1296_n 0.0654175f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_820 N_A_1178_261#_M1016_g N_A_1028_413#_c_1286_n 0.0142383f $X=6.405 $Y=0.445
+ $X2=0 $Y2=0
cc_821 N_A_1178_261#_M1015_g N_A_1028_413#_c_1297_n 0.00296198f $X=5.965
+ $Y=2.275 $X2=0 $Y2=0
cc_822 N_A_1178_261#_M1015_g N_A_1028_413#_c_1298_n 0.00444241f $X=5.965
+ $Y=2.275 $X2=0 $Y2=0
cc_823 N_A_1178_261#_c_1206_n N_A_1028_413#_c_1298_n 0.00400927f $X=6.05
+ $Y=1.825 $X2=0 $Y2=0
cc_824 N_A_1178_261#_M1016_g N_A_1028_413#_c_1384_n 0.00331097f $X=6.405
+ $Y=0.445 $X2=0 $Y2=0
cc_825 N_A_1178_261#_c_1201_n N_A_1028_413#_c_1384_n 0.00412185f $X=6.405
+ $Y=1.38 $X2=0 $Y2=0
cc_826 N_A_1178_261#_c_1209_n N_A_1028_413#_c_1384_n 0.0136304f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_827 N_A_1178_261#_c_1202_n N_A_1028_413#_c_1287_n 0.0173655f $X=7.745
+ $Y=1.575 $X2=0 $Y2=0
cc_828 N_A_1178_261#_c_1209_n N_A_1028_413#_c_1288_n 0.0032134f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_829 N_A_1178_261#_c_1209_n N_A_1028_413#_c_1289_n 0.0708095f $X=7.51 $Y=1.67
+ $X2=0 $Y2=0
cc_830 N_A_1178_261#_c_1202_n N_A_1598_47#_c_1452_n 0.028344f $X=7.745 $Y=1.575
+ $X2=0 $Y2=0
cc_831 N_A_1178_261#_c_1203_n N_A_1598_47#_c_1452_n 0.0254195f $X=7.745 $Y=0.515
+ $X2=0 $Y2=0
cc_832 N_A_1178_261#_c_1238_p N_A_1598_47#_c_1461_n 0.0257383f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_833 N_A_1178_261#_c_1238_p N_A_1598_47#_c_1462_n 0.00670342f $X=7.595 $Y=1.87
+ $X2=0 $Y2=0
cc_834 N_A_1178_261#_c_1202_n N_A_1598_47#_c_1462_n 0.021487f $X=7.745 $Y=1.575
+ $X2=0 $Y2=0
cc_835 N_A_1178_261#_c_1210_n N_A_1598_47#_c_1462_n 0.0155746f $X=7.745 $Y=1.67
+ $X2=0 $Y2=0
cc_836 N_A_1178_261#_c_1202_n N_A_1598_47#_c_1454_n 0.0165785f $X=7.745 $Y=1.575
+ $X2=0 $Y2=0
cc_837 N_A_1178_261#_c_1209_n N_VPWR_M1001_d 0.00225674f $X=7.51 $Y=1.67 $X2=0
+ $Y2=0
cc_838 N_A_1178_261#_c_1209_n N_VPWR_c_1573_n 0.0195228f $X=7.51 $Y=1.67 $X2=0
+ $Y2=0
cc_839 N_A_1178_261#_M1015_g N_VPWR_c_1580_n 8.50188e-19 $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_840 N_A_1178_261#_c_1238_p N_VPWR_c_1582_n 0.00727431f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_841 N_A_1178_261#_M1027_d N_VPWR_c_1568_n 0.00535012f $X=7.46 $Y=1.645 $X2=0
+ $Y2=0
cc_842 N_A_1178_261#_M1015_g N_VPWR_c_1568_n 0.00145798f $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_843 N_A_1178_261#_c_1238_p N_VPWR_c_1568_n 0.00614354f $X=7.595 $Y=1.87 $X2=0
+ $Y2=0
cc_844 N_A_1178_261#_M1015_g N_VPWR_c_1591_n 0.0145664f $X=5.965 $Y=2.275 $X2=0
+ $Y2=0
cc_845 N_A_1178_261#_c_1203_n N_VGND_c_1918_n 0.0140151f $X=7.745 $Y=0.515 $X2=0
+ $Y2=0
cc_846 N_A_1178_261#_M1018_d N_VGND_c_1922_n 0.00391384f $X=7.46 $Y=0.235 $X2=0
+ $Y2=0
cc_847 N_A_1178_261#_M1016_g N_VGND_c_1922_n 0.00495706f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_848 N_A_1178_261#_c_1203_n N_VGND_c_1922_n 0.0121445f $X=7.745 $Y=0.515 $X2=0
+ $Y2=0
cc_849 N_A_1178_261#_M1016_g N_VGND_c_1927_n 0.00367922f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_850 N_A_1178_261#_M1016_g N_VGND_c_1928_n 0.00248483f $X=6.405 $Y=0.445 $X2=0
+ $Y2=0
cc_851 N_A_1028_413#_M1006_g N_A_1598_47#_M1026_g 0.0189726f $X=8.325 $Y=0.445
+ $X2=0 $Y2=0
cc_852 N_A_1028_413#_M1011_g N_A_1598_47#_M1004_g 0.0189726f $X=8.325 $Y=2.165
+ $X2=0 $Y2=0
cc_853 N_A_1028_413#_M1006_g N_A_1598_47#_c_1452_n 0.0198843f $X=8.325 $Y=0.445
+ $X2=0 $Y2=0
cc_854 N_A_1028_413#_M1006_g N_A_1598_47#_c_1453_n 0.00634889f $X=8.325 $Y=0.445
+ $X2=0 $Y2=0
cc_855 N_A_1028_413#_c_1283_n N_A_1598_47#_c_1453_n 0.00984432f $X=8.325 $Y=1.26
+ $X2=0 $Y2=0
cc_856 N_A_1028_413#_M1027_g N_A_1598_47#_c_1461_n 0.00145954f $X=7.385 $Y=2.065
+ $X2=0 $Y2=0
cc_857 N_A_1028_413#_c_1281_n N_A_1598_47#_c_1461_n 0.00240579f $X=8.25 $Y=1.26
+ $X2=0 $Y2=0
cc_858 N_A_1028_413#_M1011_g N_A_1598_47#_c_1461_n 0.0057641f $X=8.325 $Y=2.165
+ $X2=0 $Y2=0
cc_859 N_A_1028_413#_M1027_g N_A_1598_47#_c_1462_n 6.15526e-19 $X=7.385 $Y=2.065
+ $X2=0 $Y2=0
cc_860 N_A_1028_413#_c_1281_n N_A_1598_47#_c_1462_n 0.00836961f $X=8.25 $Y=1.26
+ $X2=0 $Y2=0
cc_861 N_A_1028_413#_M1011_g N_A_1598_47#_c_1462_n 0.0167403f $X=8.325 $Y=2.165
+ $X2=0 $Y2=0
cc_862 N_A_1028_413#_c_1283_n N_A_1598_47#_c_1462_n 0.00281021f $X=8.325 $Y=1.26
+ $X2=0 $Y2=0
cc_863 N_A_1028_413#_c_1281_n N_A_1598_47#_c_1454_n 0.00959921f $X=8.25 $Y=1.26
+ $X2=0 $Y2=0
cc_864 N_A_1028_413#_M1006_g N_A_1598_47#_c_1454_n 8.41951e-19 $X=8.325 $Y=0.445
+ $X2=0 $Y2=0
cc_865 N_A_1028_413#_c_1283_n N_A_1598_47#_c_1454_n 5.08488e-19 $X=8.325 $Y=1.26
+ $X2=0 $Y2=0
cc_866 N_A_1028_413#_c_1283_n N_A_1598_47#_c_1455_n 0.0189726f $X=8.325 $Y=1.26
+ $X2=0 $Y2=0
cc_867 N_A_1028_413#_c_1296_n N_VPWR_M1015_d 0.00216018f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_868 N_A_1028_413#_c_1302_n N_VPWR_c_1572_n 0.00557448f $X=5.57 $Y=2.29 $X2=0
+ $Y2=0
cc_869 N_A_1028_413#_M1027_g N_VPWR_c_1573_n 0.0153912f $X=7.385 $Y=2.065 $X2=0
+ $Y2=0
cc_870 N_A_1028_413#_c_1296_n N_VPWR_c_1573_n 0.00850121f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_871 N_A_1028_413#_M1011_g N_VPWR_c_1574_n 0.00609621f $X=8.325 $Y=2.165 $X2=0
+ $Y2=0
cc_872 N_A_1028_413#_c_1302_n N_VPWR_c_1580_n 0.0200526f $X=5.57 $Y=2.29 $X2=0
+ $Y2=0
cc_873 N_A_1028_413#_c_1296_n N_VPWR_c_1580_n 0.00267646f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_874 N_A_1028_413#_c_1298_n N_VPWR_c_1580_n 0.00720374f $X=5.655 $Y=2 $X2=0
+ $Y2=0
cc_875 N_A_1028_413#_c_1296_n N_VPWR_c_1581_n 0.0036467f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_876 N_A_1028_413#_c_1297_n N_VPWR_c_1581_n 0.0101929f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_877 N_A_1028_413#_M1027_g N_VPWR_c_1582_n 0.0046653f $X=7.385 $Y=2.065 $X2=0
+ $Y2=0
cc_878 N_A_1028_413#_M1011_g N_VPWR_c_1582_n 0.00542953f $X=8.325 $Y=2.165 $X2=0
+ $Y2=0
cc_879 N_A_1028_413#_M1003_d N_VPWR_c_1568_n 0.0026466f $X=5.14 $Y=2.065 $X2=0
+ $Y2=0
cc_880 N_A_1028_413#_M1001_s N_VPWR_c_1568_n 0.00394021f $X=6.57 $Y=2.065 $X2=0
+ $Y2=0
cc_881 N_A_1028_413#_M1027_g N_VPWR_c_1568_n 0.00934473f $X=7.385 $Y=2.065 $X2=0
+ $Y2=0
cc_882 N_A_1028_413#_M1011_g N_VPWR_c_1568_n 0.0110121f $X=8.325 $Y=2.165 $X2=0
+ $Y2=0
cc_883 N_A_1028_413#_c_1302_n N_VPWR_c_1568_n 0.00987026f $X=5.57 $Y=2.29 $X2=0
+ $Y2=0
cc_884 N_A_1028_413#_c_1296_n N_VPWR_c_1568_n 0.0124969f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_885 N_A_1028_413#_c_1297_n N_VPWR_c_1568_n 0.0086238f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_886 N_A_1028_413#_c_1298_n N_VPWR_c_1568_n 0.00578252f $X=5.655 $Y=2 $X2=0
+ $Y2=0
cc_887 N_A_1028_413#_c_1296_n N_VPWR_c_1591_n 0.0270337f $X=6.54 $Y=2 $X2=0
+ $Y2=0
cc_888 N_A_1028_413#_c_1297_n N_VPWR_c_1591_n 0.00887045f $X=6.695 $Y=2.21 $X2=0
+ $Y2=0
cc_889 N_A_1028_413#_c_1298_n N_VPWR_c_1591_n 0.0115187f $X=5.655 $Y=2 $X2=0
+ $Y2=0
cc_890 N_A_1028_413#_c_1296_n A_1136_413# 0.00166681f $X=6.54 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_891 N_A_1028_413#_c_1298_n A_1136_413# 0.00336335f $X=5.655 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_892 N_A_1028_413#_M1006_g N_VGND_c_1911_n 0.00587725f $X=8.325 $Y=0.445 $X2=0
+ $Y2=0
cc_893 N_A_1028_413#_M1018_g N_VGND_c_1918_n 0.00505556f $X=7.385 $Y=0.505 $X2=0
+ $Y2=0
cc_894 N_A_1028_413#_M1006_g N_VGND_c_1918_n 0.00544863f $X=8.325 $Y=0.445 $X2=0
+ $Y2=0
cc_895 N_A_1028_413#_M1012_d N_VGND_c_1922_n 0.00218745f $X=5.64 $Y=0.235 $X2=0
+ $Y2=0
cc_896 N_A_1028_413#_M1018_g N_VGND_c_1922_n 0.00991048f $X=7.385 $Y=0.505 $X2=0
+ $Y2=0
cc_897 N_A_1028_413#_M1006_g N_VGND_c_1922_n 0.0111099f $X=8.325 $Y=0.445 $X2=0
+ $Y2=0
cc_898 N_A_1028_413#_c_1310_n N_VGND_c_1922_n 0.0135115f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_899 N_A_1028_413#_c_1310_n N_VGND_c_1927_n 0.0361566f $X=6.32 $Y=0.39 $X2=0
+ $Y2=0
cc_900 N_A_1028_413#_M1018_g N_VGND_c_1928_n 0.0188993f $X=7.385 $Y=0.505 $X2=0
+ $Y2=0
cc_901 N_A_1028_413#_c_1287_n N_VGND_c_1928_n 2.67651e-19 $X=7.305 $Y=1.26 $X2=0
+ $Y2=0
cc_902 N_A_1028_413#_c_1310_n A_1224_47# 0.00244121f $X=6.32 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_903 N_A_1598_47#_c_1461_n N_VPWR_c_1573_n 0.00150514f $X=8.115 $Y=2 $X2=0
+ $Y2=0
cc_904 N_A_1598_47#_M1004_g N_VPWR_c_1574_n 0.0106489f $X=8.8 $Y=1.985 $X2=0
+ $Y2=0
cc_905 N_A_1598_47#_M1010_g N_VPWR_c_1574_n 7.45505e-19 $X=9.22 $Y=1.985 $X2=0
+ $Y2=0
cc_906 N_A_1598_47#_c_1453_n N_VPWR_c_1574_n 0.0089025f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_907 N_A_1598_47#_c_1462_n N_VPWR_c_1574_n 0.0431561f $X=8.115 $Y=1.915 $X2=0
+ $Y2=0
cc_908 N_A_1598_47#_M1010_g N_VPWR_c_1575_n 0.00262956f $X=9.22 $Y=1.985 $X2=0
+ $Y2=0
cc_909 N_A_1598_47#_M1013_g N_VPWR_c_1575_n 0.0134961f $X=9.64 $Y=1.985 $X2=0
+ $Y2=0
cc_910 N_A_1598_47#_M1029_g N_VPWR_c_1575_n 6.7514e-19 $X=10.06 $Y=1.985 $X2=0
+ $Y2=0
cc_911 N_A_1598_47#_M1013_g N_VPWR_c_1576_n 6.7947e-19 $X=9.64 $Y=1.985 $X2=0
+ $Y2=0
cc_912 N_A_1598_47#_M1029_g N_VPWR_c_1576_n 0.0114784f $X=10.06 $Y=1.985 $X2=0
+ $Y2=0
cc_913 N_A_1598_47#_M1035_g N_VPWR_c_1576_n 0.0134334f $X=10.48 $Y=1.985 $X2=0
+ $Y2=0
cc_914 N_A_1598_47#_c_1461_n N_VPWR_c_1582_n 0.0166647f $X=8.115 $Y=2 $X2=0
+ $Y2=0
cc_915 N_A_1598_47#_M1004_g N_VPWR_c_1583_n 0.00505556f $X=8.8 $Y=1.985 $X2=0
+ $Y2=0
cc_916 N_A_1598_47#_M1010_g N_VPWR_c_1583_n 0.0054895f $X=9.22 $Y=1.985 $X2=0
+ $Y2=0
cc_917 N_A_1598_47#_M1013_g N_VPWR_c_1584_n 0.0046653f $X=9.64 $Y=1.985 $X2=0
+ $Y2=0
cc_918 N_A_1598_47#_M1029_g N_VPWR_c_1584_n 0.0046653f $X=10.06 $Y=1.985 $X2=0
+ $Y2=0
cc_919 N_A_1598_47#_M1035_g N_VPWR_c_1585_n 0.0046653f $X=10.48 $Y=1.985 $X2=0
+ $Y2=0
cc_920 N_A_1598_47#_M1011_s N_VPWR_c_1568_n 0.00211564f $X=7.99 $Y=1.845 $X2=0
+ $Y2=0
cc_921 N_A_1598_47#_M1004_g N_VPWR_c_1568_n 0.00858194f $X=8.8 $Y=1.985 $X2=0
+ $Y2=0
cc_922 N_A_1598_47#_M1010_g N_VPWR_c_1568_n 0.00978844f $X=9.22 $Y=1.985 $X2=0
+ $Y2=0
cc_923 N_A_1598_47#_M1013_g N_VPWR_c_1568_n 0.00796766f $X=9.64 $Y=1.985 $X2=0
+ $Y2=0
cc_924 N_A_1598_47#_M1029_g N_VPWR_c_1568_n 0.00796766f $X=10.06 $Y=1.985 $X2=0
+ $Y2=0
cc_925 N_A_1598_47#_M1035_g N_VPWR_c_1568_n 0.00903731f $X=10.48 $Y=1.985 $X2=0
+ $Y2=0
cc_926 N_A_1598_47#_c_1461_n N_VPWR_c_1568_n 0.0121504f $X=8.115 $Y=2 $X2=0
+ $Y2=0
cc_927 N_A_1598_47#_M1031_g N_Q_c_1840_n 0.00871421f $X=9.22 $Y=0.56 $X2=0 $Y2=0
cc_928 N_A_1598_47#_M1032_g N_Q_c_1840_n 0.0103774f $X=9.64 $Y=0.56 $X2=0 $Y2=0
cc_929 N_A_1598_47#_c_1453_n N_Q_c_1840_n 0.0359313f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_930 N_A_1598_47#_c_1455_n N_Q_c_1840_n 0.0020061f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_931 N_A_1598_47#_M1031_g N_Q_c_1829_n 0.00126056f $X=9.22 $Y=0.56 $X2=0 $Y2=0
cc_932 N_A_1598_47#_c_1453_n N_Q_c_1829_n 0.016625f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_933 N_A_1598_47#_c_1455_n N_Q_c_1829_n 0.00207985f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_934 N_A_1598_47#_M1010_g N_Q_c_1833_n 0.0112131f $X=9.22 $Y=1.985 $X2=0 $Y2=0
cc_935 N_A_1598_47#_M1013_g N_Q_c_1833_n 0.0139621f $X=9.64 $Y=1.985 $X2=0 $Y2=0
cc_936 N_A_1598_47#_c_1453_n N_Q_c_1833_n 0.038022f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_937 N_A_1598_47#_c_1455_n N_Q_c_1833_n 0.00195136f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_938 N_A_1598_47#_M1004_g N_Q_c_1834_n 8.08741e-19 $X=8.8 $Y=1.985 $X2=0 $Y2=0
cc_939 N_A_1598_47#_M1010_g N_Q_c_1834_n 0.00214237f $X=9.22 $Y=1.985 $X2=0
+ $Y2=0
cc_940 N_A_1598_47#_c_1453_n N_Q_c_1834_n 0.0180277f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_941 N_A_1598_47#_c_1462_n N_Q_c_1834_n 0.002267f $X=8.115 $Y=1.915 $X2=0
+ $Y2=0
cc_942 N_A_1598_47#_c_1455_n N_Q_c_1834_n 0.00203971f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_943 N_A_1598_47#_M1037_g N_Q_c_1856_n 0.0104216f $X=10.06 $Y=0.56 $X2=0 $Y2=0
cc_944 N_A_1598_47#_M1038_g N_Q_c_1856_n 0.0110068f $X=10.48 $Y=0.56 $X2=0 $Y2=0
cc_945 N_A_1598_47#_c_1453_n N_Q_c_1856_n 0.037694f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_946 N_A_1598_47#_c_1455_n N_Q_c_1856_n 0.0020061f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_947 N_A_1598_47#_M1029_g N_Q_c_1835_n 0.0140063f $X=10.06 $Y=1.985 $X2=0
+ $Y2=0
cc_948 N_A_1598_47#_M1035_g N_Q_c_1835_n 0.0155339f $X=10.48 $Y=1.985 $X2=0
+ $Y2=0
cc_949 N_A_1598_47#_c_1453_n N_Q_c_1835_n 0.0396013f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_950 N_A_1598_47#_c_1455_n N_Q_c_1835_n 0.00195136f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_951 N_A_1598_47#_c_1453_n N_Q_c_1830_n 0.0129289f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_952 N_A_1598_47#_c_1455_n N_Q_c_1830_n 0.00207985f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_953 N_A_1598_47#_c_1453_n N_Q_c_1836_n 0.0125885f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_954 N_A_1598_47#_c_1455_n N_Q_c_1836_n 0.00203971f $X=10.48 $Y=1.16 $X2=0
+ $Y2=0
cc_955 N_A_1598_47#_M1031_g Q 0.00765112f $X=9.22 $Y=0.56 $X2=0 $Y2=0
cc_956 N_A_1598_47#_M1032_g Q 4.48464e-19 $X=9.64 $Y=0.56 $X2=0 $Y2=0
cc_957 N_A_1598_47#_M1010_g Q 0.0108942f $X=9.22 $Y=1.985 $X2=0 $Y2=0
cc_958 N_A_1598_47#_M1013_g Q 8.23709e-19 $X=9.64 $Y=1.985 $X2=0 $Y2=0
cc_959 N_A_1598_47#_M1038_g Q 0.00450247f $X=10.48 $Y=0.56 $X2=0 $Y2=0
cc_960 N_A_1598_47#_c_1453_n Q 0.0178088f $X=10.25 $Y=1.16 $X2=0 $Y2=0
cc_961 N_A_1598_47#_c_1455_n Q 0.00686754f $X=10.48 $Y=1.16 $X2=0 $Y2=0
cc_962 N_A_1598_47#_M1026_g N_VGND_c_1911_n 0.00731244f $X=8.8 $Y=0.56 $X2=0
+ $Y2=0
cc_963 N_A_1598_47#_M1031_g N_VGND_c_1911_n 6.95802e-19 $X=9.22 $Y=0.56 $X2=0
+ $Y2=0
cc_964 N_A_1598_47#_c_1452_n N_VGND_c_1911_n 0.0143899f $X=8.115 $Y=0.51 $X2=0
+ $Y2=0
cc_965 N_A_1598_47#_c_1453_n N_VGND_c_1911_n 0.00947484f $X=10.25 $Y=1.16 $X2=0
+ $Y2=0
cc_966 N_A_1598_47#_M1031_g N_VGND_c_1912_n 0.00144638f $X=9.22 $Y=0.56 $X2=0
+ $Y2=0
cc_967 N_A_1598_47#_M1032_g N_VGND_c_1912_n 0.00719509f $X=9.64 $Y=0.56 $X2=0
+ $Y2=0
cc_968 N_A_1598_47#_M1037_g N_VGND_c_1912_n 5.93299e-19 $X=10.06 $Y=0.56 $X2=0
+ $Y2=0
cc_969 N_A_1598_47#_M1032_g N_VGND_c_1913_n 5.98297e-19 $X=9.64 $Y=0.56 $X2=0
+ $Y2=0
cc_970 N_A_1598_47#_M1037_g N_VGND_c_1913_n 0.00755066f $X=10.06 $Y=0.56 $X2=0
+ $Y2=0
cc_971 N_A_1598_47#_M1038_g N_VGND_c_1913_n 0.00955696f $X=10.48 $Y=0.56 $X2=0
+ $Y2=0
cc_972 N_A_1598_47#_c_1452_n N_VGND_c_1918_n 0.00973496f $X=8.115 $Y=0.51 $X2=0
+ $Y2=0
cc_973 N_A_1598_47#_M1026_g N_VGND_c_1919_n 0.00505556f $X=8.8 $Y=0.56 $X2=0
+ $Y2=0
cc_974 N_A_1598_47#_M1031_g N_VGND_c_1919_n 0.00425202f $X=9.22 $Y=0.56 $X2=0
+ $Y2=0
cc_975 N_A_1598_47#_M1032_g N_VGND_c_1920_n 0.00348405f $X=9.64 $Y=0.56 $X2=0
+ $Y2=0
cc_976 N_A_1598_47#_M1037_g N_VGND_c_1920_n 0.00348405f $X=10.06 $Y=0.56 $X2=0
+ $Y2=0
cc_977 N_A_1598_47#_M1038_g N_VGND_c_1921_n 0.00348405f $X=10.48 $Y=0.56 $X2=0
+ $Y2=0
cc_978 N_A_1598_47#_M1006_s N_VGND_c_1922_n 0.00359633f $X=7.99 $Y=0.235 $X2=0
+ $Y2=0
cc_979 N_A_1598_47#_M1026_g N_VGND_c_1922_n 0.00858194f $X=8.8 $Y=0.56 $X2=0
+ $Y2=0
cc_980 N_A_1598_47#_M1031_g N_VGND_c_1922_n 0.00575022f $X=9.22 $Y=0.56 $X2=0
+ $Y2=0
cc_981 N_A_1598_47#_M1032_g N_VGND_c_1922_n 0.00414556f $X=9.64 $Y=0.56 $X2=0
+ $Y2=0
cc_982 N_A_1598_47#_M1037_g N_VGND_c_1922_n 0.00414556f $X=10.06 $Y=0.56 $X2=0
+ $Y2=0
cc_983 N_A_1598_47#_M1038_g N_VGND_c_1922_n 0.00521521f $X=10.48 $Y=0.56 $X2=0
+ $Y2=0
cc_984 N_A_1598_47#_c_1452_n N_VGND_c_1922_n 0.00895081f $X=8.115 $Y=0.51 $X2=0
+ $Y2=0
cc_985 N_VPWR_c_1568_n N_A_381_47#_M1028_d 0.00325229f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_986 N_VPWR_M1028_s N_A_381_47#_c_1763_n 0.00237137f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_987 N_VPWR_M1028_s N_A_381_47#_c_1770_n 0.00471078f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_988 N_VPWR_c_1570_n N_A_381_47#_c_1770_n 0.00880041f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_989 N_VPWR_c_1579_n N_A_381_47#_c_1770_n 0.0018545f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_990 N_VPWR_c_1568_n N_A_381_47#_c_1770_n 0.00198108f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_991 N_VPWR_M1028_s N_A_381_47#_c_1766_n 0.00187968f $X=1.495 $Y=1.645 $X2=0
+ $Y2=0
cc_992 N_VPWR_c_1570_n N_A_381_47#_c_1766_n 0.0114817f $X=1.62 $Y=2.22 $X2=0
+ $Y2=0
cc_993 N_VPWR_c_1578_n N_A_381_47#_c_1766_n 3.86777e-19 $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_994 N_VPWR_c_1568_n N_A_381_47#_c_1766_n 7.1462e-19 $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_995 N_VPWR_c_1579_n N_A_381_47#_c_1773_n 0.0115924f $X=3.43 $Y=2.72 $X2=0
+ $Y2=0
cc_996 N_VPWR_c_1568_n N_A_381_47#_c_1773_n 0.00307944f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_997 N_VPWR_c_1568_n A_562_413# 0.00355877f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_998 N_VPWR_c_1568_n A_956_413# 0.00250248f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_999 N_VPWR_c_1568_n A_1136_413# 0.00223276f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1000 N_VPWR_c_1568_n N_Q_M1004_s 0.00393857f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1001 N_VPWR_c_1568_n N_Q_M1013_s 0.00570907f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1002 N_VPWR_c_1568_n N_Q_M1035_s 0.00387172f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1003 N_VPWR_M1010_d N_Q_c_1833_n 0.00165831f $X=9.295 $Y=1.485 $X2=0 $Y2=0
cc_1004 N_VPWR_c_1575_n N_Q_c_1833_n 0.014901f $X=9.43 $Y=2.16 $X2=0 $Y2=0
cc_1005 N_VPWR_c_1584_n N_Q_c_1880_n 0.0113958f $X=10.105 $Y=2.72 $X2=0 $Y2=0
cc_1006 N_VPWR_c_1568_n N_Q_c_1880_n 0.00646998f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1007 N_VPWR_M1029_d N_Q_c_1835_n 0.00165831f $X=10.135 $Y=1.485 $X2=0 $Y2=0
cc_1008 N_VPWR_c_1576_n N_Q_c_1835_n 0.0171101f $X=10.27 $Y=2.02 $X2=0 $Y2=0
cc_1009 N_VPWR_c_1583_n Q 0.0148417f $X=9.34 $Y=2.72 $X2=0 $Y2=0
cc_1010 N_VPWR_c_1568_n Q 0.0092486f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1011 N_VPWR_c_1585_n N_Q_c_1839_n 0.0244536f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1012 N_VPWR_c_1568_n N_Q_c_1839_n 0.0134021f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_1013 N_A_381_47#_c_1763_n N_VGND_M1008_s 0.00105184f $X=1.515 $Y=1.795 $X2=0
+ $Y2=0
cc_1014 N_A_381_47#_c_1768_n N_VGND_M1008_s 0.00264874f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1015 N_A_381_47#_c_1764_n N_VGND_M1008_s 0.0019591f $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_1016 N_A_381_47#_c_1768_n N_VGND_c_1908_n 0.00883988f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1017 N_A_381_47#_c_1764_n N_VGND_c_1908_n 0.0114461f $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_1018 N_A_381_47#_c_1764_n N_VGND_c_1915_n 4.97798e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_1019 N_A_381_47#_c_1768_n N_VGND_c_1916_n 0.00245002f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1020 N_A_381_47#_c_1772_n N_VGND_c_1916_n 0.00861358f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1021 N_A_381_47#_M1008_d N_VGND_c_1922_n 0.00308719f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_1022 N_A_381_47#_c_1768_n N_VGND_c_1922_n 0.00232804f $X=1.955 $Y=0.73 $X2=0
+ $Y2=0
cc_1023 N_A_381_47#_c_1764_n N_VGND_c_1922_n 8.52239e-19 $X=1.6 $Y=0.73 $X2=0
+ $Y2=0
cc_1024 N_A_381_47#_c_1772_n N_VGND_c_1922_n 0.00295275f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_1025 N_Q_c_1840_n N_VGND_M1031_s 0.00306532f $X=9.765 $Y=0.8 $X2=0 $Y2=0
cc_1026 N_Q_c_1856_n N_VGND_M1037_s 0.00306532f $X=10.605 $Y=0.8 $X2=0 $Y2=0
cc_1027 N_Q_c_1840_n N_VGND_c_1912_n 0.014257f $X=9.765 $Y=0.8 $X2=0 $Y2=0
cc_1028 N_Q_c_1856_n N_VGND_c_1913_n 0.0163351f $X=10.605 $Y=0.8 $X2=0 $Y2=0
cc_1029 N_Q_c_1840_n N_VGND_c_1919_n 0.00205432f $X=9.765 $Y=0.8 $X2=0 $Y2=0
cc_1030 Q N_VGND_c_1919_n 0.013875f $X=8.94 $Y=0.425 $X2=0 $Y2=0
cc_1031 N_Q_c_1840_n N_VGND_c_1920_n 0.0020257f $X=9.765 $Y=0.8 $X2=0 $Y2=0
cc_1032 N_Q_c_1895_p N_VGND_c_1920_n 0.0106412f $X=9.85 $Y=0.715 $X2=0 $Y2=0
cc_1033 N_Q_c_1856_n N_VGND_c_1920_n 0.0020257f $X=10.605 $Y=0.8 $X2=0 $Y2=0
cc_1034 N_Q_c_1856_n N_VGND_c_1921_n 0.0020257f $X=10.605 $Y=0.8 $X2=0 $Y2=0
cc_1035 Q N_VGND_c_1921_n 0.022939f $X=10.725 $Y=0.425 $X2=0 $Y2=0
cc_1036 N_Q_M1026_d N_VGND_c_1922_n 0.0039413f $X=8.875 $Y=0.235 $X2=0 $Y2=0
cc_1037 N_Q_M1032_d N_VGND_c_1922_n 0.00263636f $X=9.715 $Y=0.235 $X2=0 $Y2=0
cc_1038 N_Q_M1038_d N_VGND_c_1922_n 0.00233692f $X=10.555 $Y=0.235 $X2=0 $Y2=0
cc_1039 N_Q_c_1840_n N_VGND_c_1922_n 0.00877041f $X=9.765 $Y=0.8 $X2=0 $Y2=0
cc_1040 N_Q_c_1895_p N_VGND_c_1922_n 0.00642326f $X=9.85 $Y=0.715 $X2=0 $Y2=0
cc_1041 N_Q_c_1856_n N_VGND_c_1922_n 0.00913773f $X=10.605 $Y=0.8 $X2=0 $Y2=0
cc_1042 Q N_VGND_c_1922_n 0.00918033f $X=8.94 $Y=0.425 $X2=0 $Y2=0
cc_1043 Q N_VGND_c_1922_n 0.0133273f $X=10.725 $Y=0.425 $X2=0 $Y2=0
cc_1044 N_VGND_c_1922_n A_586_47# 0.00231384f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1045 N_VGND_c_1922_n A_796_47# 0.00240916f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1046 N_VGND_c_1922_n A_1056_47# 0.00198596f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1047 N_VGND_c_1922_n A_1224_47# 0.00140476f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1048 N_VGND_c_1922_n A_1296_47# 0.00259801f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__clkdlybuf4s18_1.pex.spice
* Created: Tue Sep  1 19:00:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A 3 7 8 11 12 14
r31 11 14 54.9546 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.385 $Y=1.16
+ $X2=0.385 $Y2=1.375
r32 11 13 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.385 $Y=1.16
+ $X2=0.385 $Y2=1.025
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.16 $X2=0.385 $Y2=1.16
r34 8 12 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.385 $Y2=1.19
r35 7 14 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.375
r36 3 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_27_47# 1 2 9 13 15 16 19 23 25 26
+ 27 28 32
c65 32 0 1.1875e-19 $X=0.925 $Y=1.16
r66 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.16 $X2=0.925 $Y2=1.16
r67 30 32 8.09467 $w=4.93e-07 $l=3.35e-07 $layer=LI1_cond $X=0.967 $Y=1.495
+ $X2=0.967 $Y2=1.16
r68 29 32 6.64488 $w=4.93e-07 $l=2.75e-07 $layer=LI1_cond $X=0.967 $Y=0.885
+ $X2=0.967 $Y2=1.16
r69 27 30 9.18857 $w=1.7e-07 $l=2.86363e-07 $layer=LI1_cond $X=0.72 $Y=1.58
+ $X2=0.967 $Y2=1.495
r70 27 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=1.58
+ $X2=0.425 $Y2=1.58
r71 25 29 9.18857 $w=1.7e-07 $l=2.86363e-07 $layer=LI1_cond $X=0.72 $Y=0.8
+ $X2=0.967 $Y2=0.885
r72 25 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=0.8
+ $X2=0.425 $Y2=0.8
r73 21 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.425 $Y2=1.58
r74 21 23 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.26 $Y=1.665 $X2=0.26
+ $Y2=1.965
r75 17 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.425 $Y2=0.8
r76 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.26 $Y2=0.38
r77 15 33 50.2851 $w=3.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.23 $Y=1.2
+ $X2=0.925 $Y2=1.2
r78 15 16 3.56077 $w=3.5e-07 $l=9e-08 $layer=POLY_cond $X=1.23 $Y=1.2 $X2=1.32
+ $Y2=1.2
r79 11 16 34.0592 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.32 $Y=1.375
+ $X2=1.32 $Y2=1.2
r80 11 13 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=1.32 $Y=1.375 $X2=1.32
+ $Y2=2.075
r81 7 16 34.0592 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.32 $Y=1.025
+ $X2=1.32 $Y2=1.2
r82 7 9 180.75 $w=1.8e-07 $l=4.65e-07 $layer=POLY_cond $X=1.32 $Y=1.025 $X2=1.32
+ $Y2=0.56
r83 2 23 300 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.965
r84 1 19 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_282_47# 1 2 9 13 17 22 27 28 30 32
+ 33 34
c62 27 0 1.84838e-19 $X=2.52 $Y=1.16
r63 32 33 7.63251 $w=3.73e-07 $l=1.35e-07 $layer=LI1_cond $X=1.572 $Y=1.97
+ $X2=1.572 $Y2=1.835
r64 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.16 $X2=2.52 $Y2=1.16
r65 25 34 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=1.152
+ $X2=1.675 $Y2=1.152
r66 25 27 43.2261 $w=1.93e-07 $l=7.6e-07 $layer=LI1_cond $X=1.76 $Y=1.152
+ $X2=2.52 $Y2=1.152
r67 23 34 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.675 $Y=1.25
+ $X2=1.675 $Y2=1.152
r68 23 33 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.675 $Y=1.25
+ $X2=1.675 $Y2=1.835
r69 22 34 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.675 $Y=1.055
+ $X2=1.675 $Y2=1.152
r70 22 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.675 $Y=1.055
+ $X2=1.675 $Y2=0.825
r71 15 30 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=1.572 $Y=0.638
+ $X2=1.572 $Y2=0.825
r72 15 17 7.92881 $w=3.73e-07 $l=2.58e-07 $layer=LI1_cond $X=1.572 $Y=0.638
+ $X2=1.572 $Y2=0.38
r73 11 13 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=2.325 $Y=1.375
+ $X2=2.325 $Y2=2.075
r74 7 28 31.6967 $w=3.55e-07 $l=1.95e-07 $layer=POLY_cond $X=2.325 $Y=1.197
+ $X2=2.52 $Y2=1.197
r75 7 11 18.6398 $w=1.8e-07 $l=1.78e-07 $layer=POLY_cond $X=2.325 $Y=1.197
+ $X2=2.325 $Y2=1.375
r76 7 9 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=2.325 $Y=1.02
+ $X2=2.325 $Y2=0.56
r77 2 32 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.665 $X2=1.55 $Y2=1.97
r78 1 17 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_394_47# 1 2 9 13 16 20 22 23 24 25
+ 29 30 33
c66 30 0 1.84838e-19 $X=3.11 $Y=1.16
r67 30 33 57.9773 $w=3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.095 $Y=1.16
+ $X2=3.095 $Y2=1.375
r68 30 32 42.9806 $w=3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.095 $Y=1.16
+ $X2=3.095 $Y2=1.02
r69 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.16 $X2=3.11 $Y2=1.16
r70 27 29 8.8128 $w=3.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.025 $Y=1.42
+ $X2=3.025 $Y2=1.16
r71 26 29 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=3.025 $Y=0.885
+ $X2=3.025 $Y2=1.16
r72 24 27 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.855 $Y=1.505
+ $X2=3.025 $Y2=1.42
r73 24 25 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.855 $Y=1.505
+ $X2=2.26 $Y2=1.505
r74 22 26 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.855 $Y=0.8
+ $X2=3.025 $Y2=0.885
r75 22 23 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.855 $Y=0.8
+ $X2=2.26 $Y2=0.8
r76 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.095 $Y=1.59
+ $X2=2.26 $Y2=1.505
r77 18 20 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.095 $Y=1.59
+ $X2=2.095 $Y2=1.965
r78 14 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.095 $Y=0.715
+ $X2=2.26 $Y2=0.8
r79 14 16 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.095 $Y=0.715
+ $X2=2.095 $Y2=0.38
r80 13 33 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.17 $Y=1.985
+ $X2=3.17 $Y2=1.375
r81 9 32 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.17 $Y=0.445
+ $X2=3.17 $Y2=1.02
r82 2 20 300 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_PDIFF $count=2 $X=1.97
+ $Y=1.665 $X2=2.095 $Y2=1.965
r83 1 16 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.095 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
c41 1 0 1.1875e-19 $X=0.55 $Y=1.485
r42 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.76 $Y2=2.72
r51 25 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.76 $Y2=2.72
r53 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 16 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=2.72
+ $X2=2.875 $Y2=2.72
r58 15 33 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.04 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=2.72
+ $X2=2.875 $Y2=2.72
r60 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=2.635
+ $X2=2.875 $Y2=2.72
r61 11 13 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.875 $Y=2.635
+ $X2=2.875 $Y2=2
r62 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.635 $X2=0.76
+ $Y2=2.72
r63 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=2
r64 2 13 300 $w=1.7e-07 $l=6.04731e-07 $layer=licon1_PDIFF $count=2 $X=2.415
+ $Y=1.665 $X2=2.875 $Y2=2
r65 1 9 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.76 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%X 1 2 7 8 9 10 11 12 41 46
r16 30 46 2.33603 $w=3.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.405 $Y=1.945
+ $X2=3.405 $Y2=1.87
r17 21 41 2.24696 $w=2.25e-07 $l=1.45e-07 $layer=LI1_cond $X=3.477 $Y=0.545
+ $X2=3.477 $Y2=0.4
r18 11 46 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=3.405 $Y=1.865
+ $X2=3.405 $Y2=1.87
r19 11 44 5.02762 $w=3.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.405 $Y=1.865
+ $X2=3.405 $Y2=1.76
r20 11 12 8.09825 $w=3.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.405 $Y=1.95
+ $X2=3.405 $Y2=2.21
r21 11 30 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=3.405 $Y=1.95
+ $X2=3.405 $Y2=1.945
r22 10 44 11.7805 $w=2.23e-07 $l=2.3e-07 $layer=LI1_cond $X=3.477 $Y=1.53
+ $X2=3.477 $Y2=1.76
r23 9 10 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=3.477 $Y=1.19
+ $X2=3.477 $Y2=1.53
r24 8 9 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=3.477 $Y=0.85
+ $X2=3.477 $Y2=1.19
r25 7 41 1.07296 $w=2.88e-07 $l=2.7e-08 $layer=LI1_cond $X=3.45 $Y=0.4 $X2=3.477
+ $Y2=0.4
r26 7 37 2.58306 $w=2.88e-07 $l=6.5e-08 $layer=LI1_cond $X=3.45 $Y=0.4 $X2=3.385
+ $Y2=0.4
r27 7 8 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=3.477 $Y=0.57
+ $X2=3.477 $Y2=0.85
r28 7 21 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=3.477 $Y=0.57
+ $X2=3.477 $Y2=0.545
r29 2 11 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=3.245
+ $Y=1.485 $X2=3.385 $Y2=1.965
r30 1 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.385 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r46 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r48 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r49 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r50 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r51 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r52 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r53 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 25 37 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.752
+ $Y2=0
r55 25 27 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.15
+ $Y2=0
r56 20 37 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.752
+ $Y2=0
r57 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r58 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r59 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r60 16 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.53
+ $Y2=0
r61 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.875
+ $Y2=0
r62 15 33 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.45
+ $Y2=0
r63 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.875
+ $Y2=0
r64 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r65 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.38
r66 7 37 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0
r67 7 9 10.7927 $w=3.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0.38
r68 2 13 182 $w=1.7e-07 $l=5.27541e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.875 $Y2=0.38
r69 1 9 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.745 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__or4bb_2.pex.spice
* Created: Thu Aug 27 14:44:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4BB_2%C_N 3 7 8 9 13 14 15
c32 14 0 3.1948e-20 $X=0.515 $Y=1.16
c33 3 0 1.31674e-19 $X=0.47 $Y=2.26
r34 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r35 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r37 8 9 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.53
r38 8 14 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.16
r39 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.51 $Y=0.675
+ $X2=0.51 $Y2=0.995
r40 3 16 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.47 $Y=2.26
+ $X2=0.47 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%D_N 3 6 8 11 13
r37 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.16
+ $X2=1.035 $Y2=1.325
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.16
+ $X2=1.035 $Y2=0.995
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r40 8 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=1.035 $Y2=1.16
r41 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.955 $Y=1.695
+ $X2=0.955 $Y2=1.325
r42 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.955 $Y=0.675
+ $X2=0.955 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%A_206_93# 1 2 9 13 15 20 22 24 29 35
c71 22 0 1.56005e-19 $X=1.505 $Y=1.525
c72 20 0 1.87953e-19 $X=1.505 $Y=1.075
c73 15 0 1.31674e-19 $X=1.41 $Y=1.61
r74 34 35 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.895 $Y=1.16
+ $X2=1.915 $Y2=1.16
r75 30 34 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.67 $Y=1.16
+ $X2=1.895 $Y2=1.16
r76 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r77 26 29 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.16
+ $X2=1.67 $Y2=1.16
r78 24 25 17.5021 $w=2.37e-07 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=0.655
+ $X2=1.505 $Y2=0.655
r79 21 26 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=1.245
+ $X2=1.505 $Y2=1.16
r80 21 22 16.3445 $w=1.88e-07 $l=2.8e-07 $layer=LI1_cond $X=1.505 $Y=1.245
+ $X2=1.505 $Y2=1.525
r81 20 26 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=1.075
+ $X2=1.505 $Y2=1.16
r82 19 25 2.03416 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=1.505 $Y=0.825
+ $X2=1.505 $Y2=0.655
r83 19 20 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.505 $Y=0.825
+ $X2=1.505 $Y2=1.075
r84 15 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.41 $Y=1.61
+ $X2=1.505 $Y2=1.525
r85 15 17 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.41 $Y=1.61
+ $X2=1.165 $Y2=1.61
r86 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.325
+ $X2=1.915 $Y2=1.16
r87 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.915 $Y=1.325
+ $X2=1.915 $Y2=2.275
r88 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=1.16
r89 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=0.445
r90 2 17 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.61
r91 1 24 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.465 $X2=1.165 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%A_27_410# 1 2 9 13 16 19 21 24 25 26 29 30
+ 35 37
c88 30 0 3.1201e-19 $X=2.335 $Y=1.16
r89 32 35 3.93367 $w=3.73e-07 $l=1.28e-07 $layer=LI1_cond $X=0.172 $Y=0.637
+ $X2=0.3 $Y2=0.637
r90 30 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.16
+ $X2=2.335 $Y2=1.325
r91 30 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.16
+ $X2=2.335 $Y2=0.995
r92 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.335
+ $Y=1.16 $X2=2.335 $Y2=1.16
r93 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.335 $Y=1.415
+ $X2=2.335 $Y2=1.16
r94 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=1.5
+ $X2=2.335 $Y2=1.415
r95 25 26 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.25 $Y=1.5 $X2=1.94
+ $Y2=1.5
r96 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.855 $Y=1.585
+ $X2=1.94 $Y2=1.5
r97 23 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.855 $Y=1.585
+ $X2=1.855 $Y2=1.865
r98 22 37 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.95
+ $X2=0.215 $Y2=1.95
r99 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.77 $Y=1.95
+ $X2=1.855 $Y2=1.865
r100 21 22 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=1.77 $Y=1.95
+ $X2=0.345 $Y2=1.95
r101 17 37 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=1.95
r102 17 19 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=2.035
+ $X2=0.215 $Y2=2.29
r103 16 37 4.18896 $w=2.17e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.172 $Y=1.865
+ $X2=0.215 $Y2=1.95
r104 15 32 5.2298 $w=1.75e-07 $l=1.88e-07 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=0.637
r105 15 16 65.9117 $w=1.73e-07 $l=1.04e-06 $layer=LI1_cond $X=0.172 $Y=0.825
+ $X2=0.172 $Y2=1.865
r106 13 40 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.395 $Y=1.695
+ $X2=2.395 $Y2=1.325
r107 9 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.35 $Y=0.445
+ $X2=2.35 $Y2=0.995
r108 2 19 600 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.05 $X2=0.26 $Y2=2.29
r109 1 35 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.465 $X2=0.3 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%B 4 7 8 9 10 13
c43 13 0 1.28784e-20 $X=2.815 $Y=2.335
r44 13 15 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.815 $Y=2.335
+ $X2=2.815 $Y2=2.2
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.815
+ $Y=2.335 $X2=2.815 $Y2=2.335
r46 10 14 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.015 $Y=2.29 $X2=2.815
+ $Y2=2.29
r47 8 9 65.3429 $w=1.65e-07 $l=1.5e-07 $layer=POLY_cond $X=2.762 $Y=0.76
+ $X2=2.762 $Y2=0.91
r48 7 8 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.77 $Y=0.445 $X2=2.77
+ $Y2=0.76
r49 4 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.755 $Y=1.695
+ $X2=2.755 $Y2=2.2
r50 4 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.755 $Y=1.695
+ $X2=2.755 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%A 3 7 9 12 13
c42 7 0 1.96413e-19 $X=3.19 $Y=1.695
r43 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=1.16
+ $X2=3.175 $Y2=1.325
r44 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=1.16
+ $X2=3.175 $Y2=0.995
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.175
+ $Y=1.16 $X2=3.175 $Y2=1.16
r46 9 13 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.015 $Y=1.16
+ $X2=3.175 $Y2=1.16
r47 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.19 $Y=1.695
+ $X2=3.19 $Y2=1.325
r48 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.19 $Y=0.445
+ $X2=3.19 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%A_316_413# 1 2 3 10 12 15 17 19 22 24 30 33
+ 34 35 36 37 40 42 44 49 50 51 56 58 63
c128 56 0 1.14153e-19 $X=3.655 $Y=1.16
c129 49 0 1.06604e-19 $X=3.55 $Y=1.495
c130 42 0 2.82207e-20 $X=3.465 $Y=0.74
c131 36 0 1.96413e-19 $X=2.975 $Y=1.87
c132 33 0 1.28784e-20 $X=2.195 $Y=2.205
r133 62 63 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.68 $Y=1.16
+ $X2=4.1 $Y2=1.16
r134 57 62 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.655 $Y=1.16
+ $X2=3.68 $Y2=1.16
r135 56 59 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.602 $Y=1.16
+ $X2=3.602 $Y2=1.325
r136 56 58 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.602 $Y=1.16
+ $X2=3.602 $Y2=0.995
r137 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=1.16 $X2=3.655 $Y2=1.16
r138 51 53 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.06 $Y=1.58
+ $X2=3.06 $Y2=1.87
r139 49 59 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.55 $Y=1.495
+ $X2=3.55 $Y2=1.325
r140 46 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.55 $Y=0.825
+ $X2=3.55 $Y2=0.995
r141 45 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=1.58
+ $X2=3.06 $Y2=1.58
r142 44 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.465 $Y=1.58
+ $X2=3.55 $Y2=1.495
r143 44 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.465 $Y=1.58
+ $X2=3.145 $Y2=1.58
r144 43 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=0.74
+ $X2=2.98 $Y2=0.74
r145 42 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.465 $Y=0.74
+ $X2=3.55 $Y2=0.825
r146 42 43 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.465 $Y=0.74
+ $X2=3.065 $Y2=0.74
r147 38 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.655
+ $X2=2.98 $Y2=0.74
r148 38 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.98 $Y=0.655
+ $X2=2.98 $Y2=0.47
r149 36 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=1.87
+ $X2=3.06 $Y2=1.87
r150 36 37 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.975 $Y=1.87
+ $X2=2.28 $Y2=1.87
r151 34 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0.74
+ $X2=2.98 $Y2=0.74
r152 34 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.895 $Y=0.74
+ $X2=2.195 $Y2=0.74
r153 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.195 $Y=1.955
+ $X2=2.28 $Y2=1.87
r154 32 33 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.195 $Y=1.955
+ $X2=2.195 $Y2=2.205
r155 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=0.655
+ $X2=2.195 $Y2=0.74
r156 28 30 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.11 $Y=0.655
+ $X2=2.11 $Y2=0.47
r157 24 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=2.29
+ $X2=2.195 $Y2=2.205
r158 24 26 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.11 $Y=2.29
+ $X2=1.705 $Y2=2.29
r159 20 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.1 $Y=1.325
+ $X2=4.1 $Y2=1.16
r160 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.1 $Y=1.325
+ $X2=4.1 $Y2=1.985
r161 17 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.1 $Y=0.995
+ $X2=4.1 $Y2=1.16
r162 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.1 $Y=0.995
+ $X2=4.1 $Y2=0.56
r163 13 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.325
+ $X2=3.68 $Y2=1.16
r164 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.68 $Y=1.325
+ $X2=3.68 $Y2=1.985
r165 10 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=0.995
+ $X2=3.68 $Y2=1.16
r166 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.68 $Y=0.995
+ $X2=3.68 $Y2=0.56
r167 3 26 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=2.065 $X2=1.705 $Y2=2.29
r168 2 40 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=2.845
+ $Y=0.235 $X2=2.98 $Y2=0.47
r169 1 30 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.11 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%VPWR 1 2 3 12 16 18 20 24 26 31 39 45 48 52
c58 2 0 1.06604e-19 $X=3.265 $Y=1.485
r59 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r63 43 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r64 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 40 48 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.455 $Y2=2.72
r66 40 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 39 51 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.25 $Y=2.72
+ $X2=4.425 $Y2=2.72
r68 39 42 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.25 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 35 38 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r72 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 34 37 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r74 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r76 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r77 31 48 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.315 $Y=2.72
+ $X2=3.455 $Y2=2.72
r78 31 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.315 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r80 26 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r81 24 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r83 20 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.335 $Y=1.66
+ $X2=4.335 $Y2=2.34
r84 18 51 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.335 $Y=2.635
+ $X2=4.425 $Y2=2.72
r85 18 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.335 $Y=2.635
+ $X2=4.335 $Y2=2.34
r86 14 48 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=2.635
+ $X2=3.455 $Y2=2.72
r87 14 16 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.455 $Y=2.635
+ $X2=3.455 $Y2=2
r88 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r89 10 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.29
r90 3 23 400 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=1.485 $X2=4.335 $Y2=2.34
r91 3 20 400 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=1.485 $X2=4.335 $Y2=1.66
r92 2 16 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=1.485 $X2=3.465 $Y2=2
r93 1 12 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=0.545 $Y=2.05
+ $X2=0.68 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%X 1 2 12 14 15 16
r25 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=3.942 $Y=1.632
+ $X2=3.942 $Y2=1.845
r26 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=3.942 $Y=1.632
+ $X2=3.942 $Y2=1.495
r27 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=3.89 $Y=0.587
+ $X2=3.995 $Y2=0.587
r28 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.995 $Y=0.76
+ $X2=3.995 $Y2=0.587
r29 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.995 $Y=0.76
+ $X2=3.995 $Y2=1.495
r30 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=3.755
+ $Y=1.485 $X2=3.89 $Y2=1.845
r31 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=3.755
+ $Y=0.235 $X2=3.89 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR4BB_2%VGND 1 2 3 4 5 20 24 28 32 34 36 38 40 45 50
+ 55 61 64 67 70 74 76
c80 36 0 2.82207e-20 $X=4.335 $Y=0.39
r81 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r82 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r83 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r84 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r85 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r86 59 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r87 59 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r88 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r89 56 70 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.425
+ $Y2=0
r90 56 58 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.91
+ $Y2=0
r91 55 73 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.25 $Y=0 $X2=4.425
+ $Y2=0
r92 55 58 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.25 $Y=0 $X2=3.91
+ $Y2=0
r93 54 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r94 54 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r95 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r96 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.56
+ $Y2=0
r97 51 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.99
+ $Y2=0
r98 50 70 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.425
+ $Y2=0
r99 50 53 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=2.99
+ $Y2=0
r100 49 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r101 49 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r102 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r103 46 64 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.672
+ $Y2=0
r104 46 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.07
+ $Y2=0
r105 45 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.56
+ $Y2=0
r106 45 48 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=0
+ $X2=2.07 $Y2=0
r107 44 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r108 44 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r109 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r110 41 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.745
+ $Y2=0
r111 41 43 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.15
+ $Y2=0
r112 40 64 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.495 $Y=0
+ $X2=1.672 $Y2=0
r113 40 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.15
+ $Y2=0
r114 38 62 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r115 38 76 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r116 34 73 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.335 $Y=0.085
+ $X2=4.425 $Y2=0
r117 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.335 $Y=0.085
+ $X2=4.335 $Y2=0.39
r118 30 70 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.425 $Y2=0
r119 30 32 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.425 $Y2=0.4
r120 26 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r121 26 28 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.4
r122 22 64 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.672 $Y=0.085
+ $X2=1.672 $Y2=0
r123 22 24 10.2259 $w=3.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.672 $Y=0.085
+ $X2=1.672 $Y2=0.4
r124 18 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r125 18 20 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.66
r126 5 36 91 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_NDIFF $count=2 $X=4.175
+ $Y=0.235 $X2=4.335 $Y2=0.39
r127 4 32 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.235 $X2=3.45 $Y2=0.4
r128 3 28 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.56 $Y2=0.4
r129 2 24 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.685 $Y2=0.4
r130 1 20 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.465 $X2=0.745 $Y2=0.66
.ends


* File: sky130_fd_sc_hd__dlrtp_4.spice.SKY130_FD_SC_HD__DLRTP_4.pxi
* Created: Thu Aug 27 14:17:42 2020
* 
x_PM_SKY130_FD_SC_HD__DLRTP_4%GATE N_GATE_c_156_n N_GATE_c_151_n N_GATE_M1024_g
+ N_GATE_c_157_n N_GATE_M1011_g N_GATE_c_152_n N_GATE_c_158_n GATE GATE
+ N_GATE_c_154_n N_GATE_c_155_n PM_SKY130_FD_SC_HD__DLRTP_4%GATE
x_PM_SKY130_FD_SC_HD__DLRTP_4%A_27_47# N_A_27_47#_M1024_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1013_g N_A_27_47#_M1000_g N_A_27_47#_M1025_g N_A_27_47#_c_195_n
+ N_A_27_47#_c_196_n N_A_27_47#_M1019_g N_A_27_47#_c_207_n N_A_27_47#_c_330_p
+ N_A_27_47#_c_198_n N_A_27_47#_c_199_n N_A_27_47#_c_208_n N_A_27_47#_c_209_n
+ N_A_27_47#_c_200_n N_A_27_47#_c_201_n N_A_27_47#_c_211_n N_A_27_47#_c_212_n
+ N_A_27_47#_c_213_n N_A_27_47#_c_214_n N_A_27_47#_c_215_n N_A_27_47#_c_216_n
+ N_A_27_47#_c_202_n PM_SKY130_FD_SC_HD__DLRTP_4%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRTP_4%D N_D_M1022_g N_D_M1016_g D N_D_c_341_n
+ N_D_c_342_n PM_SKY130_FD_SC_HD__DLRTP_4%D
x_PM_SKY130_FD_SC_HD__DLRTP_4%A_300_47# N_A_300_47#_M1022_s N_A_300_47#_M1016_s
+ N_A_300_47#_M1005_g N_A_300_47#_M1012_g N_A_300_47#_c_387_n
+ N_A_300_47#_c_380_n N_A_300_47#_c_388_n N_A_300_47#_c_389_n
+ N_A_300_47#_c_381_n N_A_300_47#_c_382_n N_A_300_47#_c_383_n
+ N_A_300_47#_c_384_n N_A_300_47#_c_385_n PM_SKY130_FD_SC_HD__DLRTP_4%A_300_47#
x_PM_SKY130_FD_SC_HD__DLRTP_4%A_193_47# N_A_193_47#_M1013_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1008_g N_A_193_47#_M1004_g N_A_193_47#_c_464_n
+ N_A_193_47#_c_471_n N_A_193_47#_c_465_n N_A_193_47#_c_466_n
+ N_A_193_47#_c_472_n N_A_193_47#_c_473_n N_A_193_47#_c_474_n
+ N_A_193_47#_c_475_n N_A_193_47#_c_467_n N_A_193_47#_c_476_n
+ N_A_193_47#_c_477_n N_A_193_47#_c_468_n PM_SKY130_FD_SC_HD__DLRTP_4%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRTP_4%A_725_21# N_A_725_21#_M1003_s N_A_725_21#_M1001_d
+ N_A_725_21#_M1009_g N_A_725_21#_M1006_g N_A_725_21#_c_587_n
+ N_A_725_21#_M1007_g N_A_725_21#_M1002_g N_A_725_21#_c_588_n
+ N_A_725_21#_M1017_g N_A_725_21#_M1014_g N_A_725_21#_c_589_n
+ N_A_725_21#_M1018_g N_A_725_21#_M1015_g N_A_725_21#_c_590_n
+ N_A_725_21#_M1020_g N_A_725_21#_M1023_g N_A_725_21#_c_601_n
+ N_A_725_21#_c_602_n N_A_725_21#_c_591_n N_A_725_21#_c_611_p
+ N_A_725_21#_c_592_n N_A_725_21#_c_667_p N_A_725_21#_c_635_p
+ N_A_725_21#_c_593_n N_A_725_21#_c_640_p N_A_725_21#_c_594_n
+ PM_SKY130_FD_SC_HD__DLRTP_4%A_725_21#
x_PM_SKY130_FD_SC_HD__DLRTP_4%A_562_413# N_A_562_413#_M1008_d
+ N_A_562_413#_M1025_d N_A_562_413#_M1003_g N_A_562_413#_M1001_g
+ N_A_562_413#_c_739_n N_A_562_413#_c_740_n N_A_562_413#_c_747_n
+ N_A_562_413#_c_748_n N_A_562_413#_c_741_n N_A_562_413#_c_742_n
+ N_A_562_413#_c_745_n N_A_562_413#_c_743_n
+ PM_SKY130_FD_SC_HD__DLRTP_4%A_562_413#
x_PM_SKY130_FD_SC_HD__DLRTP_4%RESET_B N_RESET_B_c_821_n N_RESET_B_M1021_g
+ N_RESET_B_M1010_g RESET_B N_RESET_B_c_822_n N_RESET_B_c_823_n
+ PM_SKY130_FD_SC_HD__DLRTP_4%RESET_B
x_PM_SKY130_FD_SC_HD__DLRTP_4%VPWR N_VPWR_M1011_d N_VPWR_M1016_d N_VPWR_M1006_d
+ N_VPWR_M1001_s N_VPWR_M1010_d N_VPWR_M1014_d N_VPWR_M1023_d N_VPWR_c_862_n
+ N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_865_n N_VPWR_c_866_n N_VPWR_c_867_n
+ N_VPWR_c_868_n N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_871_n VPWR
+ N_VPWR_c_872_n N_VPWR_c_873_n N_VPWR_c_874_n N_VPWR_c_875_n N_VPWR_c_876_n
+ N_VPWR_c_877_n N_VPWR_c_878_n N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n
+ N_VPWR_c_882_n N_VPWR_c_861_n PM_SKY130_FD_SC_HD__DLRTP_4%VPWR
x_PM_SKY130_FD_SC_HD__DLRTP_4%Q N_Q_M1007_s N_Q_M1018_s N_Q_M1002_s N_Q_M1015_s
+ N_Q_c_991_n N_Q_c_988_n N_Q_c_997_n N_Q_c_1001_n N_Q_c_989_n N_Q_c_986_n Q Q Q
+ Q N_Q_c_1015_n N_Q_c_1018_n PM_SKY130_FD_SC_HD__DLRTP_4%Q
x_PM_SKY130_FD_SC_HD__DLRTP_4%VGND N_VGND_M1024_d N_VGND_M1022_d N_VGND_M1009_d
+ N_VGND_M1021_d N_VGND_M1017_d N_VGND_M1020_d N_VGND_c_1046_n N_VGND_c_1047_n
+ N_VGND_c_1048_n N_VGND_c_1049_n N_VGND_c_1050_n N_VGND_c_1051_n
+ N_VGND_c_1052_n N_VGND_c_1053_n VGND N_VGND_c_1054_n N_VGND_c_1055_n
+ N_VGND_c_1056_n N_VGND_c_1057_n N_VGND_c_1058_n N_VGND_c_1059_n
+ N_VGND_c_1060_n N_VGND_c_1061_n N_VGND_c_1062_n N_VGND_c_1063_n
+ N_VGND_c_1064_n PM_SKY130_FD_SC_HD__DLRTP_4%VGND
cc_1 VNB N_GATE_c_151_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_c_152_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_c_154_n 0.0212744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_c_155_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1013_g 0.0398153f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_195_n 0.0133385f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_c_196_n 0.00520223f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_9 VNB N_A_27_47#_M1019_g 0.0464035f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_10 VNB N_A_27_47#_c_198_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_199_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_200_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_201_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_202_n 0.0230796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_D_M1022_g 0.0259137f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_16 VNB N_D_M1016_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_17 VNB N_D_c_341_n 0.00410732f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_18 VNB N_D_c_342_n 0.0422167f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_19 VNB N_A_300_47#_M1012_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_300_47#_c_380_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_300_47#_c_381_n 0.00496114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_300_47#_c_382_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_23 VNB N_A_300_47#_c_383_n 0.00266162f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_24 VNB N_A_300_47#_c_384_n 0.0274388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_300_47#_c_385_n 0.01709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_c_464_n 0.0141407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_465_n 0.0271289f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_28 VNB N_A_193_47#_c_466_n 0.00381134f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_29 VNB N_A_193_47#_c_467_n 0.0176114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_468_n 0.00469707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_725_21#_M1009_g 0.0513173f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_32 VNB N_A_725_21#_c_587_n 0.016009f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_33 VNB N_A_725_21#_c_588_n 0.0155423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_725_21#_c_589_n 0.0152501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_725_21#_c_590_n 0.0190067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_725_21#_c_591_n 0.00462291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_725_21#_c_592_n 0.0032549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_725_21#_c_593_n 0.00188136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_725_21#_c_594_n 0.0773531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_562_413#_M1003_g 0.0239034f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_41 VNB N_A_562_413#_M1001_g 4.92816e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_42 VNB N_A_562_413#_c_739_n 0.0496142f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_43 VNB N_A_562_413#_c_740_n 0.00703905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_562_413#_c_741_n 0.00738412f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_45 VNB N_A_562_413#_c_742_n 0.0118425f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_46 VNB N_A_562_413#_c_743_n 0.0105408f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_47 VNB N_RESET_B_c_821_n 0.0167184f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_48 VNB N_RESET_B_c_822_n 0.0200549f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_49 VNB N_RESET_B_c_823_n 0.00294307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VPWR_c_861_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_Q_c_986_n 6.78457e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB Q 0.0246209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1046_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1047_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_55 VNB N_VGND_c_1048_n 0.00598407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1049_n 0.00278314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1050_n 0.0177881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1051_n 0.00223657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1052_n 0.0100504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1053_n 0.0171925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1054_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1055_n 0.0273338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1056_n 0.0412073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1057_n 0.0261275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1058_n 0.0131639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1059_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1060_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1061_n 0.00507544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1062_n 0.00523213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1063_n 0.00380306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1064_n 0.372537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VPB N_GATE_c_156_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_73 VPB N_GATE_c_157_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_74 VPB N_GATE_c_158_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_75 VPB GATE 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_76 VPB N_GATE_c_154_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_77 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_78 VPB N_A_27_47#_M1025_g 0.0320638f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_79 VPB N_A_27_47#_c_195_n 0.0174243f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_80 VPB N_A_27_47#_c_196_n 0.00955572f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_81 VPB N_A_27_47#_c_207_n 0.0121291f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_82 VPB N_A_27_47#_c_208_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_209_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_200_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_211_n 0.0226938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_212_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_47#_c_213_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_47#_c_214_n 0.00344459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_27_47#_c_215_n 0.00529835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_27_47#_c_216_n 0.00947367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_27_47#_c_202_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_D_M1016_g 0.0462632f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_93 VPB N_D_c_341_n 0.00235173f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_94 VPB N_A_300_47#_M1012_g 0.0366983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_300_47#_c_387_n 0.00718148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_300_47#_c_388_n 0.00409088f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_97 VPB N_A_300_47#_c_389_n 0.00291454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_300_47#_c_382_n 0.00355393f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_99 VPB N_A_193_47#_M1004_g 0.0212488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_193_47#_c_464_n 0.00807078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_193_47#_c_471_n 0.00294853f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_102 VPB N_A_193_47#_c_472_n 0.00925296f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_103 VPB N_A_193_47#_c_473_n 0.00238933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_193_47#_c_474_n 0.00716976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_193_47#_c_475_n 0.00258599f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_193_47#_c_476_n 0.00920811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_193_47#_c_477_n 0.0330434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_193_47#_c_468_n 0.00264136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_725_21#_M1009_g 0.019403f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_110 VPB N_A_725_21#_M1006_g 0.0275278f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_111 VPB N_A_725_21#_M1002_g 0.0180708f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_112 VPB N_A_725_21#_M1014_g 0.0184109f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_113 VPB N_A_725_21#_M1015_g 0.0187462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_725_21#_M1023_g 0.025555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_725_21#_c_601_n 0.00678489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_725_21#_c_602_n 0.0414704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_725_21#_c_593_n 0.00274615f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_725_21#_c_594_n 0.0157737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_562_413#_M1001_g 0.0266617f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_120 VPB N_A_562_413#_c_745_n 0.00556334f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_121 VPB N_A_562_413#_c_743_n 0.00397469f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_122 VPB N_RESET_B_M1010_g 0.0195786f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_123 VPB N_RESET_B_c_822_n 0.00406869f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_124 VPB N_RESET_B_c_823_n 0.00291233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_862_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_126 VPB N_VPWR_c_863_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_127 VPB N_VPWR_c_864_n 0.00761302f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_865_n 0.00598254f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_866_n 0.00111373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_867_n 3.28374e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_868_n 0.0167807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_869_n 0.00169029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_870_n 0.0100504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_871_n 0.0418135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_872_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_873_n 0.0296723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_874_n 0.0416819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_875_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_876_n 0.0131639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_877_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_878_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_879_n 0.00555175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_880_n 0.00417584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_881_n 0.00490136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_882_n 0.00380306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_861_n 0.0577381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_Q_c_988_n 0.00278502f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_148 VPB N_Q_c_989_n 9.5962e-19 $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_149 VPB Q 0.00375704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 N_GATE_c_151_n N_A_27_47#_M1013_g 0.0187834f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_151 N_GATE_c_155_n N_A_27_47#_M1013_g 0.0041981f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_152 N_GATE_c_158_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_153 N_GATE_c_154_n N_A_27_47#_M1000_g 0.00527228f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_154 N_GATE_c_151_n N_A_27_47#_c_198_n 0.00663556f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_155 N_GATE_c_152_n N_A_27_47#_c_198_n 0.0105293f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_156 N_GATE_c_152_n N_A_27_47#_c_199_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_157 GATE N_A_27_47#_c_199_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_158 N_GATE_c_154_n N_A_27_47#_c_199_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_159 N_GATE_c_157_n N_A_27_47#_c_208_n 0.0135489f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_160 N_GATE_c_158_n N_A_27_47#_c_208_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_161 N_GATE_c_157_n N_A_27_47#_c_209_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_162 N_GATE_c_158_n N_A_27_47#_c_209_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_163 GATE N_A_27_47#_c_209_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_164 N_GATE_c_154_n N_A_27_47#_c_209_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_165 N_GATE_c_154_n N_A_27_47#_c_200_n 0.00319708f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_166 N_GATE_c_152_n N_A_27_47#_c_201_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_167 GATE N_A_27_47#_c_201_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_168 N_GATE_c_155_n N_A_27_47#_c_201_n 0.0015185f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_169 N_GATE_c_156_n N_A_27_47#_c_212_n 0.0033897f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_170 N_GATE_c_158_n N_A_27_47#_c_212_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_171 GATE N_A_27_47#_c_212_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_172 N_GATE_c_156_n N_A_27_47#_c_213_n 7.60515e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_173 N_GATE_c_158_n N_A_27_47#_c_213_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_174 GATE N_A_27_47#_c_202_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_175 N_GATE_c_154_n N_A_27_47#_c_202_n 0.0165992f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_176 N_GATE_c_157_n N_VPWR_c_862_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_177 N_GATE_c_157_n N_VPWR_c_872_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_178 N_GATE_c_157_n N_VPWR_c_861_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_179 N_GATE_c_151_n N_VGND_c_1046_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_180 N_GATE_c_151_n N_VGND_c_1054_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_181 N_GATE_c_152_n N_VGND_c_1054_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_182 N_GATE_c_151_n N_VGND_c_1064_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_211_n N_D_M1016_g 0.00583826f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_211_n N_D_c_341_n 0.0087134f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1013_g N_D_c_342_n 0.00512711f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A_27_47#_M1025_g N_A_300_47#_M1012_g 0.0356141f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_196_n N_A_300_47#_M1012_g 0.0248435f $X=2.81 $Y=1.32 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_211_n N_A_300_47#_M1012_g 0.00493352f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_214_n N_A_300_47#_M1012_g 0.00140912f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_215_n N_A_300_47#_M1012_g 0.00239179f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_211_n N_A_300_47#_c_388_n 0.0116439f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_214_n N_A_300_47#_c_388_n 0.00130924f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_215_n N_A_300_47#_c_388_n 0.00675603f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_211_n N_A_300_47#_c_389_n 0.0115282f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_211_n N_A_300_47#_c_381_n 0.00675641f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_211_n N_A_300_47#_c_382_n 0.0108494f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_214_n N_A_300_47#_c_382_n 0.00124596f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_215_n N_A_300_47#_c_382_n 0.00570493f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_211_n N_A_300_47#_c_384_n 0.00107604f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_M1025_g N_A_193_47#_M1004_g 0.0144372f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_M1013_g N_A_193_47#_c_464_n 0.00780615f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_198_n N_A_193_47#_c_464_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_200_n N_A_193_47#_c_464_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_201_n N_A_193_47#_c_464_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_211_n N_A_193_47#_c_464_n 0.0184751f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_212_n N_A_193_47#_c_464_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_213_n N_A_193_47#_c_464_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_208_n N_A_193_47#_c_471_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_211_n N_A_193_47#_c_471_n 0.00195186f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_202_n N_A_193_47#_c_471_n 0.00780615f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_196_n N_A_193_47#_c_465_n 0.0188813f $X=2.81 $Y=1.32 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_M1019_g N_A_193_47#_c_465_n 0.0192792f $X=3.225 $Y=0.415 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_215_n N_A_193_47#_c_465_n 4.13927e-19 $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_195_n N_A_193_47#_c_466_n 7.03475e-19 $X=3.15 $Y=1.32 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_196_n N_A_193_47#_c_466_n 0.00136198f $X=2.81 $Y=1.32 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_M1019_g N_A_193_47#_c_466_n 0.00256371f $X=3.225 $Y=0.415
+ $X2=0 $Y2=0
cc_217 N_A_27_47#_c_215_n N_A_193_47#_c_466_n 0.00180905f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_M1025_g N_A_193_47#_c_472_n 0.00772267f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_219 N_A_27_47#_c_195_n N_A_193_47#_c_472_n 0.00118095f $X=3.15 $Y=1.32 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_207_n N_A_193_47#_c_472_n 0.00185018f $X=2.675 $Y=1.685
+ $X2=0 $Y2=0
cc_221 N_A_27_47#_c_211_n N_A_193_47#_c_472_n 0.0875256f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_214_n N_A_193_47#_c_472_n 0.0266068f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_215_n N_A_193_47#_c_472_n 0.00879532f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_M1000_g N_A_193_47#_c_473_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_208_n N_A_193_47#_c_473_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_211_n N_A_193_47#_c_473_n 0.0259095f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_213_n N_A_193_47#_c_473_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1000_g N_A_193_47#_c_474_n 0.00780615f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_M1025_g N_A_193_47#_c_475_n 0.00151176f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_230 N_A_27_47#_c_195_n N_A_193_47#_c_475_n 0.00114785f $X=3.15 $Y=1.32 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1019_g N_A_193_47#_c_467_n 0.0126141f $X=3.225 $Y=0.415 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_195_n N_A_193_47#_c_476_n 0.00413065f $X=3.15 $Y=1.32 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_207_n N_A_193_47#_c_476_n 0.0051426f $X=2.675 $Y=1.685 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_195_n N_A_193_47#_c_477_n 0.0185785f $X=3.15 $Y=1.32 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_207_n N_A_193_47#_c_477_n 0.016673f $X=2.675 $Y=1.685 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_195_n N_A_193_47#_c_468_n 0.0129153f $X=3.15 $Y=1.32 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1019_g N_A_193_47#_c_468_n 0.0049729f $X=3.225 $Y=0.415 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_214_n N_A_193_47#_c_468_n 0.00148697f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_215_n N_A_193_47#_c_468_n 0.0232128f $X=2.56 $Y=1.53 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_216_n N_A_193_47#_c_468_n 0.0051426f $X=2.675 $Y=1.52 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_M1019_g N_A_725_21#_M1009_g 0.0429816f $X=3.225 $Y=0.415 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1019_g N_A_562_413#_c_747_n 0.0125275f $X=3.225 $Y=0.415
+ $X2=0 $Y2=0
cc_243 N_A_27_47#_M1025_g N_A_562_413#_c_748_n 0.00281839f $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_244 N_A_27_47#_M1019_g N_A_562_413#_c_741_n 0.00562201f $X=3.225 $Y=0.415
+ $X2=0 $Y2=0
cc_245 N_A_27_47#_M1019_g N_A_562_413#_c_742_n 0.00348305f $X=3.225 $Y=0.415
+ $X2=0 $Y2=0
cc_246 N_A_27_47#_M1025_g N_A_562_413#_c_745_n 9.31897e-19 $X=2.735 $Y=2.275
+ $X2=0 $Y2=0
cc_247 N_A_27_47#_c_195_n N_A_562_413#_c_745_n 6.71539e-19 $X=3.15 $Y=1.32 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_208_n N_VPWR_M1011_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_249 N_A_27_47#_M1000_g N_VPWR_c_862_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_208_n N_VPWR_c_862_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_209_n N_VPWR_c_862_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_212_n N_VPWR_c_862_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1025_g N_VPWR_c_863_n 0.00404706f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_211_n N_VPWR_c_863_n 0.0019389f $X=2.415 $Y=1.53 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_208_n N_VPWR_c_872_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_209_n N_VPWR_c_872_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_257 N_A_27_47#_M1000_g N_VPWR_c_873_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1025_g N_VPWR_c_874_n 0.00585385f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1000_g N_VPWR_c_861_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1025_g N_VPWR_c_861_n 0.00704377f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_208_n N_VPWR_c_861_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_209_n N_VPWR_c_861_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_198_n N_VGND_M1024_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_264 N_A_27_47#_M1013_g N_VGND_c_1046_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_198_n N_VGND_c_1046_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_200_n N_VGND_c_1046_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_202_n N_VGND_c_1046_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1019_g N_VGND_c_1048_n 0.0017297f $X=3.225 $Y=0.415 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_330_p N_VGND_c_1054_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_198_n N_VGND_c_1054_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1013_g N_VGND_c_1055_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1019_g N_VGND_c_1056_n 0.0037981f $X=3.225 $Y=0.415 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1024_s N_VGND_c_1064_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1013_g N_VGND_c_1064_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1019_g N_VGND_c_1064_n 0.00555936f $X=3.225 $Y=0.415 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_330_p N_VGND_c_1064_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_198_n N_VGND_c_1064_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_278 N_D_c_342_n N_A_300_47#_M1012_g 0.03863f $X=1.835 $Y=1.04 $X2=0 $Y2=0
cc_279 N_D_M1016_g N_A_300_47#_c_387_n 0.012851f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_280 N_D_M1022_g N_A_300_47#_c_380_n 0.0144498f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_281 N_D_c_341_n N_A_300_47#_c_380_n 0.00627239f $X=1.63 $Y=1.04 $X2=0 $Y2=0
cc_282 N_D_c_342_n N_A_300_47#_c_380_n 0.00123166f $X=1.835 $Y=1.04 $X2=0 $Y2=0
cc_283 N_D_M1016_g N_A_300_47#_c_388_n 0.00794545f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_284 N_D_M1016_g N_A_300_47#_c_389_n 0.00412429f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_285 N_D_c_341_n N_A_300_47#_c_389_n 0.0229667f $X=1.63 $Y=1.04 $X2=0 $Y2=0
cc_286 N_D_c_342_n N_A_300_47#_c_389_n 0.00131849f $X=1.835 $Y=1.04 $X2=0 $Y2=0
cc_287 N_D_M1022_g N_A_300_47#_c_381_n 0.00563568f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_288 N_D_c_341_n N_A_300_47#_c_381_n 0.0107593f $X=1.63 $Y=1.04 $X2=0 $Y2=0
cc_289 N_D_c_341_n N_A_300_47#_c_382_n 0.0164827f $X=1.63 $Y=1.04 $X2=0 $Y2=0
cc_290 N_D_c_342_n N_A_300_47#_c_382_n 0.00552652f $X=1.835 $Y=1.04 $X2=0 $Y2=0
cc_291 N_D_M1022_g N_A_300_47#_c_383_n 0.00120855f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_292 N_D_c_341_n N_A_300_47#_c_383_n 0.0138491f $X=1.63 $Y=1.04 $X2=0 $Y2=0
cc_293 N_D_c_342_n N_A_300_47#_c_383_n 0.0042466f $X=1.835 $Y=1.04 $X2=0 $Y2=0
cc_294 N_D_M1022_g N_A_300_47#_c_384_n 0.0197208f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_295 N_D_M1022_g N_A_300_47#_c_385_n 0.015283f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_296 N_D_M1022_g N_A_193_47#_c_464_n 0.00202363f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_297 N_D_M1016_g N_A_193_47#_c_464_n 0.00457813f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_298 N_D_c_341_n N_A_193_47#_c_464_n 0.0207394f $X=1.63 $Y=1.04 $X2=0 $Y2=0
cc_299 N_D_c_342_n N_A_193_47#_c_464_n 0.00255999f $X=1.835 $Y=1.04 $X2=0 $Y2=0
cc_300 N_D_M1016_g N_A_193_47#_c_471_n 0.00135447f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_301 N_D_M1016_g N_A_193_47#_c_472_n 0.00294239f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_302 N_D_M1016_g N_VPWR_c_863_n 0.00304701f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_303 N_D_M1016_g N_VPWR_c_873_n 0.00543342f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_304 N_D_M1016_g N_VPWR_c_861_n 0.00734866f $X=1.835 $Y=2.165 $X2=0 $Y2=0
cc_305 N_D_M1022_g N_VGND_c_1047_n 0.0110406f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_306 N_D_M1022_g N_VGND_c_1055_n 0.00337001f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_307 N_D_M1022_g N_VGND_c_1064_n 0.0053254f $X=1.835 $Y=0.445 $X2=0 $Y2=0
cc_308 N_D_c_342_n N_VGND_c_1064_n 0.00103829f $X=1.835 $Y=1.04 $X2=0 $Y2=0
cc_309 N_A_300_47#_c_387_n N_A_193_47#_c_464_n 0.00107843f $X=1.625 $Y=1.99
+ $X2=0 $Y2=0
cc_310 N_A_300_47#_c_389_n N_A_193_47#_c_464_n 0.00845026f $X=1.79 $Y=1.58 $X2=0
+ $Y2=0
cc_311 N_A_300_47#_c_383_n N_A_193_47#_c_464_n 0.018988f $X=1.625 $Y=0.51 $X2=0
+ $Y2=0
cc_312 N_A_300_47#_c_387_n N_A_193_47#_c_471_n 0.0462772f $X=1.625 $Y=1.99 $X2=0
+ $Y2=0
cc_313 N_A_300_47#_c_381_n N_A_193_47#_c_465_n 9.56555e-19 $X=2.06 $Y=1.095
+ $X2=0 $Y2=0
cc_314 N_A_300_47#_c_384_n N_A_193_47#_c_465_n 0.0117556f $X=2.26 $Y=0.93 $X2=0
+ $Y2=0
cc_315 N_A_300_47#_c_385_n N_A_193_47#_c_465_n 0.00200147f $X=2.26 $Y=0.765
+ $X2=0 $Y2=0
cc_316 N_A_300_47#_c_381_n N_A_193_47#_c_466_n 0.0129081f $X=2.06 $Y=1.095 $X2=0
+ $Y2=0
cc_317 N_A_300_47#_c_384_n N_A_193_47#_c_466_n 9.50608e-19 $X=2.26 $Y=0.93 $X2=0
+ $Y2=0
cc_318 N_A_300_47#_c_385_n N_A_193_47#_c_466_n 2.04855e-19 $X=2.26 $Y=0.765
+ $X2=0 $Y2=0
cc_319 N_A_300_47#_M1012_g N_A_193_47#_c_472_n 0.00365242f $X=2.255 $Y=2.165
+ $X2=0 $Y2=0
cc_320 N_A_300_47#_c_387_n N_A_193_47#_c_472_n 0.0227796f $X=1.625 $Y=1.99 $X2=0
+ $Y2=0
cc_321 N_A_300_47#_c_388_n N_A_193_47#_c_472_n 0.00551435f $X=1.975 $Y=1.58
+ $X2=0 $Y2=0
cc_322 N_A_300_47#_c_387_n N_A_193_47#_c_473_n 0.00272304f $X=1.625 $Y=1.99
+ $X2=0 $Y2=0
cc_323 N_A_300_47#_c_385_n N_A_193_47#_c_467_n 0.0197936f $X=2.26 $Y=0.765 $X2=0
+ $Y2=0
cc_324 N_A_300_47#_M1012_g N_A_193_47#_c_468_n 0.00370009f $X=2.255 $Y=2.165
+ $X2=0 $Y2=0
cc_325 N_A_300_47#_c_381_n N_A_193_47#_c_468_n 0.00178567f $X=2.06 $Y=1.095
+ $X2=0 $Y2=0
cc_326 N_A_300_47#_c_384_n N_A_193_47#_c_468_n 9.9633e-19 $X=2.26 $Y=0.93 $X2=0
+ $Y2=0
cc_327 N_A_300_47#_c_385_n N_A_562_413#_c_747_n 6.54613e-19 $X=2.26 $Y=0.765
+ $X2=0 $Y2=0
cc_328 N_A_300_47#_M1012_g N_VPWR_c_863_n 0.0238376f $X=2.255 $Y=2.165 $X2=0
+ $Y2=0
cc_329 N_A_300_47#_c_387_n N_VPWR_c_863_n 0.0232987f $X=1.625 $Y=1.99 $X2=0
+ $Y2=0
cc_330 N_A_300_47#_c_388_n N_VPWR_c_863_n 0.013562f $X=1.975 $Y=1.58 $X2=0 $Y2=0
cc_331 N_A_300_47#_c_387_n N_VPWR_c_873_n 0.0159418f $X=1.625 $Y=1.99 $X2=0
+ $Y2=0
cc_332 N_A_300_47#_M1012_g N_VPWR_c_874_n 0.00212864f $X=2.255 $Y=2.165 $X2=0
+ $Y2=0
cc_333 N_A_300_47#_M1016_s N_VPWR_c_861_n 0.00174533f $X=1.5 $Y=1.845 $X2=0
+ $Y2=0
cc_334 N_A_300_47#_M1012_g N_VPWR_c_861_n 0.00262666f $X=2.255 $Y=2.165 $X2=0
+ $Y2=0
cc_335 N_A_300_47#_c_387_n N_VPWR_c_861_n 0.00576627f $X=1.625 $Y=1.99 $X2=0
+ $Y2=0
cc_336 N_A_300_47#_c_381_n N_VGND_M1022_d 0.00156939f $X=2.06 $Y=1.095 $X2=0
+ $Y2=0
cc_337 N_A_300_47#_c_380_n N_VGND_c_1047_n 0.00259081f $X=1.975 $Y=0.7 $X2=0
+ $Y2=0
cc_338 N_A_300_47#_c_381_n N_VGND_c_1047_n 0.0141976f $X=2.06 $Y=1.095 $X2=0
+ $Y2=0
cc_339 N_A_300_47#_c_385_n N_VGND_c_1047_n 0.00964732f $X=2.26 $Y=0.765 $X2=0
+ $Y2=0
cc_340 N_A_300_47#_c_380_n N_VGND_c_1055_n 0.00255672f $X=1.975 $Y=0.7 $X2=0
+ $Y2=0
cc_341 N_A_300_47#_c_383_n N_VGND_c_1055_n 0.00711582f $X=1.625 $Y=0.51 $X2=0
+ $Y2=0
cc_342 N_A_300_47#_c_384_n N_VGND_c_1056_n 9.84895e-19 $X=2.26 $Y=0.93 $X2=0
+ $Y2=0
cc_343 N_A_300_47#_c_385_n N_VGND_c_1056_n 0.0046653f $X=2.26 $Y=0.765 $X2=0
+ $Y2=0
cc_344 N_A_300_47#_M1022_s N_VGND_c_1064_n 0.00283248f $X=1.5 $Y=0.235 $X2=0
+ $Y2=0
cc_345 N_A_300_47#_c_380_n N_VGND_c_1064_n 0.00473142f $X=1.975 $Y=0.7 $X2=0
+ $Y2=0
cc_346 N_A_300_47#_c_381_n N_VGND_c_1064_n 0.00552372f $X=2.06 $Y=1.095 $X2=0
+ $Y2=0
cc_347 N_A_300_47#_c_383_n N_VGND_c_1064_n 0.00607883f $X=1.625 $Y=0.51 $X2=0
+ $Y2=0
cc_348 N_A_300_47#_c_384_n N_VGND_c_1064_n 0.00117722f $X=2.26 $Y=0.93 $X2=0
+ $Y2=0
cc_349 N_A_300_47#_c_385_n N_VGND_c_1064_n 0.00454932f $X=2.26 $Y=0.765 $X2=0
+ $Y2=0
cc_350 N_A_193_47#_c_468_n N_A_725_21#_M1009_g 9.55756e-19 $X=3.1 $Y=1.575 $X2=0
+ $Y2=0
cc_351 N_A_193_47#_M1004_g N_A_725_21#_M1006_g 0.0313447f $X=3.34 $Y=2.275 $X2=0
+ $Y2=0
cc_352 N_A_193_47#_c_476_n N_A_725_21#_c_602_n 4.66982e-19 $X=3.185 $Y=1.74
+ $X2=0 $Y2=0
cc_353 N_A_193_47#_c_477_n N_A_725_21#_c_602_n 0.0313447f $X=3.34 $Y=1.74 $X2=0
+ $Y2=0
cc_354 N_A_193_47#_c_465_n N_A_562_413#_c_747_n 0.00144439f $X=2.805 $Y=0.87
+ $X2=0 $Y2=0
cc_355 N_A_193_47#_c_466_n N_A_562_413#_c_747_n 0.0162478f $X=3.015 $Y=0.87
+ $X2=0 $Y2=0
cc_356 N_A_193_47#_c_467_n N_A_562_413#_c_747_n 0.00412044f $X=2.805 $Y=0.705
+ $X2=0 $Y2=0
cc_357 N_A_193_47#_M1004_g N_A_562_413#_c_748_n 0.0116262f $X=3.34 $Y=2.275
+ $X2=0 $Y2=0
cc_358 N_A_193_47#_c_475_n N_A_562_413#_c_748_n 0.00179474f $X=3.02 $Y=1.87
+ $X2=0 $Y2=0
cc_359 N_A_193_47#_c_476_n N_A_562_413#_c_748_n 0.0149106f $X=3.185 $Y=1.74
+ $X2=0 $Y2=0
cc_360 N_A_193_47#_c_477_n N_A_562_413#_c_748_n 0.00111122f $X=3.34 $Y=1.74
+ $X2=0 $Y2=0
cc_361 N_A_193_47#_c_466_n N_A_562_413#_c_741_n 0.0184898f $X=3.015 $Y=0.87
+ $X2=0 $Y2=0
cc_362 N_A_193_47#_c_466_n N_A_562_413#_c_742_n 0.0027819f $X=3.015 $Y=0.87
+ $X2=0 $Y2=0
cc_363 N_A_193_47#_c_477_n N_A_562_413#_c_742_n 0.00291146f $X=3.34 $Y=1.74
+ $X2=0 $Y2=0
cc_364 N_A_193_47#_c_468_n N_A_562_413#_c_742_n 0.0160678f $X=3.1 $Y=1.575 $X2=0
+ $Y2=0
cc_365 N_A_193_47#_c_475_n N_A_562_413#_c_745_n 0.0013063f $X=3.02 $Y=1.87 $X2=0
+ $Y2=0
cc_366 N_A_193_47#_c_476_n N_A_562_413#_c_745_n 0.0251673f $X=3.185 $Y=1.74
+ $X2=0 $Y2=0
cc_367 N_A_193_47#_c_477_n N_A_562_413#_c_745_n 0.00856317f $X=3.34 $Y=1.74
+ $X2=0 $Y2=0
cc_368 N_A_193_47#_c_468_n N_A_562_413#_c_745_n 0.0103836f $X=3.1 $Y=1.575 $X2=0
+ $Y2=0
cc_369 N_A_193_47#_c_472_n N_VPWR_M1016_d 6.81311e-19 $X=2.875 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_474_n N_VPWR_c_862_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_c_472_n N_VPWR_c_863_n 0.0184727f $X=2.875 $Y=1.87 $X2=0
+ $Y2=0
cc_372 N_A_193_47#_c_475_n N_VPWR_c_863_n 9.60836e-19 $X=3.02 $Y=1.87 $X2=0
+ $Y2=0
cc_373 N_A_193_47#_c_476_n N_VPWR_c_863_n 0.00218529f $X=3.185 $Y=1.74 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_474_n N_VPWR_c_873_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_375 N_A_193_47#_M1004_g N_VPWR_c_874_n 0.00366111f $X=3.34 $Y=2.275 $X2=0
+ $Y2=0
cc_376 N_A_193_47#_M1004_g N_VPWR_c_861_n 0.00549379f $X=3.34 $Y=2.275 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_c_472_n N_VPWR_c_861_n 0.0755222f $X=2.875 $Y=1.87 $X2=0
+ $Y2=0
cc_378 N_A_193_47#_c_473_n N_VPWR_c_861_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_379 N_A_193_47#_c_474_n N_VPWR_c_861_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_380 N_A_193_47#_c_475_n N_VPWR_c_861_n 0.0149279f $X=3.02 $Y=1.87 $X2=0 $Y2=0
cc_381 N_A_193_47#_c_472_n A_466_369# 0.00388705f $X=2.875 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_193_47#_c_467_n N_VGND_c_1047_n 0.00174223f $X=2.805 $Y=0.705 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_c_464_n N_VGND_c_1055_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_384 N_A_193_47#_c_465_n N_VGND_c_1056_n 9.43262e-19 $X=2.805 $Y=0.87 $X2=0
+ $Y2=0
cc_385 N_A_193_47#_c_466_n N_VGND_c_1056_n 0.00182549f $X=3.015 $Y=0.87 $X2=0
+ $Y2=0
cc_386 N_A_193_47#_c_467_n N_VGND_c_1056_n 0.00425892f $X=2.805 $Y=0.705 $X2=0
+ $Y2=0
cc_387 N_A_193_47#_M1013_d N_VGND_c_1064_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_388 N_A_193_47#_c_464_n N_VGND_c_1064_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_389 N_A_193_47#_c_465_n N_VGND_c_1064_n 0.00121904f $X=2.805 $Y=0.87 $X2=0
+ $Y2=0
cc_390 N_A_193_47#_c_466_n N_VGND_c_1064_n 0.00328555f $X=3.015 $Y=0.87 $X2=0
+ $Y2=0
cc_391 N_A_193_47#_c_467_n N_VGND_c_1064_n 0.00628992f $X=2.805 $Y=0.705 $X2=0
+ $Y2=0
cc_392 N_A_725_21#_c_591_n N_A_562_413#_M1003_g 0.00734947f $X=4.43 $Y=0.4 $X2=0
+ $Y2=0
cc_393 N_A_725_21#_c_611_p N_A_562_413#_M1003_g 0.00820318f $X=5.455 $Y=0.74
+ $X2=0 $Y2=0
cc_394 N_A_725_21#_c_592_n N_A_562_413#_M1003_g 8.67038e-19 $X=4.595 $Y=0.74
+ $X2=0 $Y2=0
cc_395 N_A_725_21#_c_601_n N_A_562_413#_M1001_g 0.0167742f $X=4.755 $Y=1.7 $X2=0
+ $Y2=0
cc_396 N_A_725_21#_c_602_n N_A_562_413#_M1001_g 0.00640354f $X=3.93 $Y=1.7 $X2=0
+ $Y2=0
cc_397 N_A_725_21#_M1009_g N_A_562_413#_c_739_n 0.0175191f $X=3.7 $Y=0.445 $X2=0
+ $Y2=0
cc_398 N_A_725_21#_c_601_n N_A_562_413#_c_739_n 0.0113698f $X=4.755 $Y=1.7 $X2=0
+ $Y2=0
cc_399 N_A_725_21#_c_602_n N_A_562_413#_c_739_n 0.00424117f $X=3.93 $Y=1.7 $X2=0
+ $Y2=0
cc_400 N_A_725_21#_c_592_n N_A_562_413#_c_739_n 0.0100964f $X=4.595 $Y=0.74
+ $X2=0 $Y2=0
cc_401 N_A_725_21#_M1009_g N_A_562_413#_c_747_n 0.00158904f $X=3.7 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_725_21#_M1006_g N_A_562_413#_c_748_n 0.00369776f $X=3.7 $Y=2.275
+ $X2=0 $Y2=0
cc_403 N_A_725_21#_M1009_g N_A_562_413#_c_741_n 0.010318f $X=3.7 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_A_725_21#_M1009_g N_A_562_413#_c_742_n 0.00570022f $X=3.7 $Y=0.445
+ $X2=0 $Y2=0
cc_405 N_A_725_21#_M1009_g N_A_562_413#_c_745_n 0.0114233f $X=3.7 $Y=0.445 $X2=0
+ $Y2=0
cc_406 N_A_725_21#_M1006_g N_A_562_413#_c_745_n 0.0143765f $X=3.7 $Y=2.275 $X2=0
+ $Y2=0
cc_407 N_A_725_21#_c_601_n N_A_562_413#_c_745_n 0.0249855f $X=4.755 $Y=1.7 $X2=0
+ $Y2=0
cc_408 N_A_725_21#_c_602_n N_A_562_413#_c_745_n 0.00797618f $X=3.93 $Y=1.7 $X2=0
+ $Y2=0
cc_409 N_A_725_21#_M1009_g N_A_562_413#_c_743_n 0.0180695f $X=3.7 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_725_21#_c_601_n N_A_562_413#_c_743_n 0.0284222f $X=4.755 $Y=1.7 $X2=0
+ $Y2=0
cc_411 N_A_725_21#_c_602_n N_A_562_413#_c_743_n 0.0059817f $X=3.93 $Y=1.7 $X2=0
+ $Y2=0
cc_412 N_A_725_21#_c_587_n N_RESET_B_c_821_n 0.0209688f $X=5.54 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_413 N_A_725_21#_c_591_n N_RESET_B_c_821_n 0.00151117f $X=4.43 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_414 N_A_725_21#_c_611_p N_RESET_B_c_821_n 0.0117213f $X=5.455 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_415 N_A_725_21#_c_593_n N_RESET_B_c_821_n 0.00210354f $X=5.54 $Y=1.16
+ $X2=-0.19 $Y2=-0.24
cc_416 N_A_725_21#_M1002_g N_RESET_B_M1010_g 0.0221909f $X=5.54 $Y=1.985 $X2=0
+ $Y2=0
cc_417 N_A_725_21#_c_635_p N_RESET_B_M1010_g 0.0131717f $X=5.455 $Y=1.62 $X2=0
+ $Y2=0
cc_418 N_A_725_21#_c_593_n N_RESET_B_M1010_g 0.00295902f $X=5.54 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A_725_21#_c_611_p N_RESET_B_c_822_n 0.0024858f $X=5.455 $Y=0.74 $X2=0
+ $Y2=0
cc_420 N_A_725_21#_c_635_p N_RESET_B_c_822_n 0.00121226f $X=5.455 $Y=1.62 $X2=0
+ $Y2=0
cc_421 N_A_725_21#_c_593_n N_RESET_B_c_822_n 0.00107425f $X=5.54 $Y=1.16 $X2=0
+ $Y2=0
cc_422 N_A_725_21#_c_640_p N_RESET_B_c_822_n 3.98165e-19 $X=4.85 $Y=1.755 $X2=0
+ $Y2=0
cc_423 N_A_725_21#_c_594_n N_RESET_B_c_822_n 0.0214597f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_424 N_A_725_21#_c_601_n N_RESET_B_c_823_n 0.0131995f $X=4.755 $Y=1.7 $X2=0
+ $Y2=0
cc_425 N_A_725_21#_c_611_p N_RESET_B_c_823_n 0.0362828f $X=5.455 $Y=0.74 $X2=0
+ $Y2=0
cc_426 N_A_725_21#_c_592_n N_RESET_B_c_823_n 0.00496106f $X=4.595 $Y=0.74 $X2=0
+ $Y2=0
cc_427 N_A_725_21#_c_635_p N_RESET_B_c_823_n 0.0106304f $X=5.455 $Y=1.62 $X2=0
+ $Y2=0
cc_428 N_A_725_21#_c_593_n N_RESET_B_c_823_n 0.0153384f $X=5.54 $Y=1.16 $X2=0
+ $Y2=0
cc_429 N_A_725_21#_c_640_p N_RESET_B_c_823_n 0.0127431f $X=4.85 $Y=1.755 $X2=0
+ $Y2=0
cc_430 N_A_725_21#_c_594_n N_RESET_B_c_823_n 0.0012594f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_431 N_A_725_21#_c_601_n N_VPWR_M1001_s 0.00675912f $X=4.755 $Y=1.7 $X2=0
+ $Y2=0
cc_432 N_A_725_21#_c_635_p N_VPWR_M1010_d 0.0103088f $X=5.455 $Y=1.62 $X2=0
+ $Y2=0
cc_433 N_A_725_21#_M1006_g N_VPWR_c_864_n 0.0045387f $X=3.7 $Y=2.275 $X2=0 $Y2=0
cc_434 N_A_725_21#_c_601_n N_VPWR_c_864_n 0.0157229f $X=4.755 $Y=1.7 $X2=0 $Y2=0
cc_435 N_A_725_21#_c_602_n N_VPWR_c_864_n 0.00522755f $X=3.93 $Y=1.7 $X2=0 $Y2=0
cc_436 N_A_725_21#_c_601_n N_VPWR_c_866_n 0.0123588f $X=4.755 $Y=1.7 $X2=0 $Y2=0
cc_437 N_A_725_21#_M1002_g N_VPWR_c_867_n 0.0106906f $X=5.54 $Y=1.985 $X2=0
+ $Y2=0
cc_438 N_A_725_21#_M1014_g N_VPWR_c_867_n 7.54305e-19 $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_439 N_A_725_21#_c_635_p N_VPWR_c_867_n 0.0205447f $X=5.455 $Y=1.62 $X2=0
+ $Y2=0
cc_440 N_A_725_21#_M1002_g N_VPWR_c_868_n 0.00505556f $X=5.54 $Y=1.985 $X2=0
+ $Y2=0
cc_441 N_A_725_21#_M1014_g N_VPWR_c_868_n 0.00518588f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_442 N_A_725_21#_M1014_g N_VPWR_c_869_n 0.00456367f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_443 N_A_725_21#_M1015_g N_VPWR_c_869_n 0.0165681f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_444 N_A_725_21#_M1023_g N_VPWR_c_869_n 7.29212e-19 $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_445 N_A_725_21#_c_594_n N_VPWR_c_869_n 0.00244604f $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_446 N_A_725_21#_M1015_g N_VPWR_c_871_n 6.78711e-19 $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_447 N_A_725_21#_M1023_g N_VPWR_c_871_n 0.0147395f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_448 N_A_725_21#_M1006_g N_VPWR_c_874_n 0.00541489f $X=3.7 $Y=2.275 $X2=0
+ $Y2=0
cc_449 N_A_725_21#_c_667_p N_VPWR_c_875_n 0.0121054f $X=4.85 $Y=2.27 $X2=0 $Y2=0
cc_450 N_A_725_21#_M1015_g N_VPWR_c_876_n 0.00388479f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_451 N_A_725_21#_M1023_g N_VPWR_c_876_n 0.00505556f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_452 N_A_725_21#_M1001_d N_VPWR_c_861_n 0.00385995f $X=4.715 $Y=1.485 $X2=0
+ $Y2=0
cc_453 N_A_725_21#_M1006_g N_VPWR_c_861_n 0.0106979f $X=3.7 $Y=2.275 $X2=0 $Y2=0
cc_454 N_A_725_21#_M1002_g N_VPWR_c_861_n 0.00859622f $X=5.54 $Y=1.985 $X2=0
+ $Y2=0
cc_455 N_A_725_21#_M1014_g N_VPWR_c_861_n 0.00911393f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_456 N_A_725_21#_M1015_g N_VPWR_c_861_n 0.00676354f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_457 N_A_725_21#_M1023_g N_VPWR_c_861_n 0.00860861f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_458 N_A_725_21#_c_601_n N_VPWR_c_861_n 0.0142526f $X=4.755 $Y=1.7 $X2=0 $Y2=0
cc_459 N_A_725_21#_c_602_n N_VPWR_c_861_n 0.00110429f $X=3.93 $Y=1.7 $X2=0 $Y2=0
cc_460 N_A_725_21#_c_667_p N_VPWR_c_861_n 0.00724021f $X=4.85 $Y=2.27 $X2=0
+ $Y2=0
cc_461 N_A_725_21#_c_587_n N_Q_c_991_n 0.00361433f $X=5.54 $Y=0.995 $X2=0 $Y2=0
cc_462 N_A_725_21#_c_588_n N_Q_c_991_n 0.00646762f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_463 N_A_725_21#_c_589_n N_Q_c_991_n 5.83114e-19 $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_464 N_A_725_21#_M1015_g N_Q_c_988_n 0.00608036f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_465 N_A_725_21#_M1023_g N_Q_c_988_n 0.00538211f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_466 N_A_725_21#_c_594_n N_Q_c_988_n 0.00382365f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_467 N_A_725_21#_c_587_n N_Q_c_997_n 0.00201876f $X=5.54 $Y=0.995 $X2=0 $Y2=0
cc_468 N_A_725_21#_c_588_n N_Q_c_997_n 0.00314065f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_469 N_A_725_21#_c_611_p N_Q_c_997_n 3.33421e-19 $X=5.455 $Y=0.74 $X2=0 $Y2=0
cc_470 N_A_725_21#_c_594_n N_Q_c_997_n 0.00253843f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_471 N_A_725_21#_M1002_g N_Q_c_1001_n 0.00306727f $X=5.54 $Y=1.985 $X2=0 $Y2=0
cc_472 N_A_725_21#_M1014_g N_Q_c_1001_n 0.00305099f $X=5.995 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_A_725_21#_c_594_n N_Q_c_1001_n 0.00262533f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_474 N_A_725_21#_M1002_g N_Q_c_989_n 0.00470014f $X=5.54 $Y=1.985 $X2=0 $Y2=0
cc_475 N_A_725_21#_M1014_g N_Q_c_989_n 0.0118076f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_476 N_A_725_21#_M1015_g N_Q_c_989_n 5.15734e-19 $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_477 N_A_725_21#_c_593_n N_Q_c_989_n 0.0137852f $X=5.54 $Y=1.16 $X2=0 $Y2=0
cc_478 N_A_725_21#_c_587_n N_Q_c_986_n 9.2199e-19 $X=5.54 $Y=0.995 $X2=0 $Y2=0
cc_479 N_A_725_21#_c_588_n N_Q_c_986_n 0.00265448f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_480 N_A_725_21#_c_593_n N_Q_c_986_n 0.0370808f $X=5.54 $Y=1.16 $X2=0 $Y2=0
cc_481 N_A_725_21#_c_594_n N_Q_c_986_n 0.0115123f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_482 N_A_725_21#_M1014_g Q 0.00636811f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_483 N_A_725_21#_c_590_n Q 0.0143541f $X=6.89 $Y=0.995 $X2=0 $Y2=0
cc_484 N_A_725_21#_c_594_n Q 0.031228f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_485 N_A_725_21#_c_588_n N_Q_c_1015_n 0.00759671f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_486 N_A_725_21#_c_589_n N_Q_c_1015_n 0.0121098f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_487 N_A_725_21#_c_594_n N_Q_c_1015_n 0.0409199f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_488 N_A_725_21#_c_589_n N_Q_c_1018_n 0.00289643f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_489 N_A_725_21#_c_594_n N_Q_c_1018_n 5.29963e-19 $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_490 N_A_725_21#_c_611_p N_VGND_M1021_d 0.0102296f $X=5.455 $Y=0.74 $X2=0
+ $Y2=0
cc_491 N_A_725_21#_M1009_g N_VGND_c_1048_n 0.0115145f $X=3.7 $Y=0.445 $X2=0
+ $Y2=0
cc_492 N_A_725_21#_c_591_n N_VGND_c_1048_n 0.0211756f $X=4.43 $Y=0.4 $X2=0 $Y2=0
cc_493 N_A_725_21#_c_587_n N_VGND_c_1049_n 0.00312335f $X=5.54 $Y=0.995 $X2=0
+ $Y2=0
cc_494 N_A_725_21#_c_591_n N_VGND_c_1049_n 0.0071136f $X=4.43 $Y=0.4 $X2=0 $Y2=0
cc_495 N_A_725_21#_c_611_p N_VGND_c_1049_n 0.0189838f $X=5.455 $Y=0.74 $X2=0
+ $Y2=0
cc_496 N_A_725_21#_c_587_n N_VGND_c_1050_n 0.00425543f $X=5.54 $Y=0.995 $X2=0
+ $Y2=0
cc_497 N_A_725_21#_c_588_n N_VGND_c_1050_n 0.00517132f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_498 N_A_725_21#_c_611_p N_VGND_c_1050_n 0.00258263f $X=5.455 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_725_21#_c_588_n N_VGND_c_1051_n 0.00428312f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_500 N_A_725_21#_c_589_n N_VGND_c_1051_n 0.00929972f $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_501 N_A_725_21#_c_590_n N_VGND_c_1051_n 5.95615e-19 $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_A_725_21#_c_594_n N_VGND_c_1051_n 4.93017e-19 $X=6.89 $Y=1.16 $X2=0
+ $Y2=0
cc_503 N_A_725_21#_c_589_n N_VGND_c_1053_n 5.57058e-19 $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_725_21#_c_590_n N_VGND_c_1053_n 0.00897931f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_A_725_21#_M1009_g N_VGND_c_1056_n 0.0046653f $X=3.7 $Y=0.445 $X2=0
+ $Y2=0
cc_506 N_A_725_21#_c_591_n N_VGND_c_1057_n 0.0207942f $X=4.43 $Y=0.4 $X2=0 $Y2=0
cc_507 N_A_725_21#_c_611_p N_VGND_c_1057_n 0.00732922f $X=5.455 $Y=0.74 $X2=0
+ $Y2=0
cc_508 N_A_725_21#_c_589_n N_VGND_c_1058_n 0.00388479f $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_509 N_A_725_21#_c_590_n N_VGND_c_1058_n 0.00505556f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_510 N_A_725_21#_M1003_s N_VGND_c_1064_n 0.00209319f $X=4.305 $Y=0.235 $X2=0
+ $Y2=0
cc_511 N_A_725_21#_M1009_g N_VGND_c_1064_n 0.00813035f $X=3.7 $Y=0.445 $X2=0
+ $Y2=0
cc_512 N_A_725_21#_c_587_n N_VGND_c_1064_n 0.00585509f $X=5.54 $Y=0.995 $X2=0
+ $Y2=0
cc_513 N_A_725_21#_c_588_n N_VGND_c_1064_n 0.00586927f $X=5.995 $Y=0.995 $X2=0
+ $Y2=0
cc_514 N_A_725_21#_c_589_n N_VGND_c_1064_n 0.00373675f $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_515 N_A_725_21#_c_590_n N_VGND_c_1064_n 0.00465936f $X=6.89 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_A_725_21#_c_591_n N_VGND_c_1064_n 0.0123694f $X=4.43 $Y=0.4 $X2=0 $Y2=0
cc_517 N_A_725_21#_c_611_p N_VGND_c_1064_n 0.0186317f $X=5.455 $Y=0.74 $X2=0
+ $Y2=0
cc_518 N_A_725_21#_c_611_p A_943_47# 0.00441372f $X=5.455 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_519 N_A_562_413#_M1003_g N_RESET_B_c_821_n 0.0424142f $X=4.64 $Y=0.56
+ $X2=-0.19 $Y2=-0.24
cc_520 N_A_562_413#_M1001_g N_RESET_B_M1010_g 0.0244798f $X=4.64 $Y=1.985 $X2=0
+ $Y2=0
cc_521 N_A_562_413#_M1003_g N_RESET_B_c_822_n 0.0213898f $X=4.64 $Y=0.56 $X2=0
+ $Y2=0
cc_522 N_A_562_413#_M1003_g N_RESET_B_c_823_n 0.0031862f $X=4.64 $Y=0.56 $X2=0
+ $Y2=0
cc_523 N_A_562_413#_M1001_g N_RESET_B_c_823_n 0.00343566f $X=4.64 $Y=1.985 $X2=0
+ $Y2=0
cc_524 N_A_562_413#_c_739_n N_RESET_B_c_823_n 0.00821388f $X=4.565 $Y=1.16 $X2=0
+ $Y2=0
cc_525 N_A_562_413#_c_740_n N_RESET_B_c_823_n 0.00629189f $X=4.64 $Y=1.16 $X2=0
+ $Y2=0
cc_526 N_A_562_413#_c_743_n N_RESET_B_c_823_n 0.0195733f $X=4.15 $Y=1.16 $X2=0
+ $Y2=0
cc_527 N_A_562_413#_c_748_n N_VPWR_c_863_n 0.00489615f $X=3.485 $Y=2.34 $X2=0
+ $Y2=0
cc_528 N_A_562_413#_M1001_g N_VPWR_c_864_n 0.00105344f $X=4.64 $Y=1.985 $X2=0
+ $Y2=0
cc_529 N_A_562_413#_M1001_g N_VPWR_c_866_n 0.00859497f $X=4.64 $Y=1.985 $X2=0
+ $Y2=0
cc_530 N_A_562_413#_M1001_g N_VPWR_c_867_n 6.54137e-19 $X=4.64 $Y=1.985 $X2=0
+ $Y2=0
cc_531 N_A_562_413#_c_748_n N_VPWR_c_874_n 0.0343719f $X=3.485 $Y=2.34 $X2=0
+ $Y2=0
cc_532 N_A_562_413#_M1001_g N_VPWR_c_875_n 0.00505556f $X=4.64 $Y=1.985 $X2=0
+ $Y2=0
cc_533 N_A_562_413#_M1025_d N_VPWR_c_861_n 0.00383902f $X=2.81 $Y=2.065 $X2=0
+ $Y2=0
cc_534 N_A_562_413#_M1001_g N_VPWR_c_861_n 0.00477699f $X=4.64 $Y=1.985 $X2=0
+ $Y2=0
cc_535 N_A_562_413#_c_748_n N_VPWR_c_861_n 0.0212261f $X=3.485 $Y=2.34 $X2=0
+ $Y2=0
cc_536 N_A_562_413#_c_748_n A_683_413# 0.00145479f $X=3.485 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_537 N_A_562_413#_c_745_n A_683_413# 0.00208506f $X=3.57 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_538 N_A_562_413#_c_747_n N_VGND_c_1047_n 0.00209539f $X=3.335 $Y=0.45 $X2=0
+ $Y2=0
cc_539 N_A_562_413#_M1003_g N_VGND_c_1048_n 0.00234993f $X=4.64 $Y=0.56 $X2=0
+ $Y2=0
cc_540 N_A_562_413#_c_739_n N_VGND_c_1048_n 5.64862e-19 $X=4.565 $Y=1.16 $X2=0
+ $Y2=0
cc_541 N_A_562_413#_c_747_n N_VGND_c_1048_n 0.010424f $X=3.335 $Y=0.45 $X2=0
+ $Y2=0
cc_542 N_A_562_413#_c_743_n N_VGND_c_1048_n 0.0123605f $X=4.15 $Y=1.16 $X2=0
+ $Y2=0
cc_543 N_A_562_413#_M1003_g N_VGND_c_1049_n 0.00183303f $X=4.64 $Y=0.56 $X2=0
+ $Y2=0
cc_544 N_A_562_413#_c_747_n N_VGND_c_1056_n 0.0221606f $X=3.335 $Y=0.45 $X2=0
+ $Y2=0
cc_545 N_A_562_413#_M1003_g N_VGND_c_1057_n 0.00415469f $X=4.64 $Y=0.56 $X2=0
+ $Y2=0
cc_546 N_A_562_413#_M1008_d N_VGND_c_1064_n 0.00237979f $X=2.87 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_A_562_413#_M1003_g N_VGND_c_1064_n 0.00709954f $X=4.64 $Y=0.56 $X2=0
+ $Y2=0
cc_548 N_A_562_413#_c_747_n N_VGND_c_1064_n 0.0222941f $X=3.335 $Y=0.45 $X2=0
+ $Y2=0
cc_549 N_A_562_413#_c_747_n A_660_47# 0.00365607f $X=3.335 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_550 N_A_562_413#_c_741_n A_660_47# 0.00149829f $X=3.42 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_551 N_RESET_B_M1010_g N_VPWR_c_866_n 5.74285e-19 $X=5.06 $Y=1.985 $X2=0 $Y2=0
cc_552 N_RESET_B_M1010_g N_VPWR_c_867_n 0.0100483f $X=5.06 $Y=1.985 $X2=0 $Y2=0
cc_553 N_RESET_B_M1010_g N_VPWR_c_875_n 0.00505556f $X=5.06 $Y=1.985 $X2=0 $Y2=0
cc_554 N_RESET_B_M1010_g N_VPWR_c_861_n 0.00861019f $X=5.06 $Y=1.985 $X2=0 $Y2=0
cc_555 N_RESET_B_c_821_n N_VGND_c_1049_n 0.00994415f $X=5.06 $Y=0.995 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_821_n N_VGND_c_1057_n 0.00327422f $X=5.06 $Y=0.995 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_821_n N_VGND_c_1064_n 0.00391018f $X=5.06 $Y=0.995 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_861_n A_466_369# 0.00476473f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_559 N_VPWR_c_861_n A_683_413# 0.00170472f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_560 N_VPWR_c_861_n N_Q_M1002_s 0.00468958f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_561 N_VPWR_c_861_n N_Q_M1015_s 0.00629193f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_562 N_VPWR_c_869_n N_Q_c_988_n 0.0713882f $X=6.22 $Y=1.66 $X2=0 $Y2=0
cc_563 N_VPWR_c_876_n N_Q_c_988_n 0.0133661f $X=6.945 $Y=2.72 $X2=0 $Y2=0
cc_564 N_VPWR_c_861_n N_Q_c_988_n 0.00762533f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_565 N_VPWR_c_867_n N_Q_c_1001_n 0.0410574f $X=5.3 $Y=2.02 $X2=0 $Y2=0
cc_566 N_VPWR_c_869_n N_Q_c_989_n 0.0722051f $X=6.22 $Y=1.66 $X2=0 $Y2=0
cc_567 N_VPWR_c_868_n Q 0.0177053f $X=6.135 $Y=2.72 $X2=0 $Y2=0
cc_568 N_VPWR_c_861_n Q 0.0106089f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_569 N_VPWR_c_871_n Q 0.0269253f $X=7.1 $Y=1.66 $X2=0 $Y2=0
cc_570 N_VPWR_c_869_n N_Q_c_1015_n 0.0202473f $X=6.22 $Y=1.66 $X2=0 $Y2=0
cc_571 N_Q_c_1015_n N_VGND_M1017_d 0.00194737f $X=6.575 $Y=1.045 $X2=0 $Y2=0
cc_572 Q N_VGND_M1020_d 0.00272121f $X=7.095 $Y=0.765 $X2=0 $Y2=0
cc_573 N_Q_c_997_n N_VGND_c_1050_n 0.019461f $X=5.88 $Y=0.37 $X2=0 $Y2=0
cc_574 N_Q_c_991_n N_VGND_c_1051_n 0.00800894f $X=5.88 $Y=0.765 $X2=0 $Y2=0
cc_575 N_Q_c_997_n N_VGND_c_1051_n 0.0176123f $X=5.88 $Y=0.37 $X2=0 $Y2=0
cc_576 N_Q_c_1015_n N_VGND_c_1051_n 0.0178223f $X=6.575 $Y=1.045 $X2=0 $Y2=0
cc_577 N_Q_c_1018_n N_VGND_c_1051_n 0.0250227f $X=6.66 $Y=0.49 $X2=0 $Y2=0
cc_578 Q N_VGND_c_1053_n 0.0232877f $X=7.095 $Y=0.765 $X2=0 $Y2=0
cc_579 N_Q_c_1018_n N_VGND_c_1058_n 0.0131012f $X=6.66 $Y=0.49 $X2=0 $Y2=0
cc_580 N_Q_M1007_s N_VGND_c_1064_n 0.00243335f $X=5.615 $Y=0.235 $X2=0 $Y2=0
cc_581 N_Q_M1018_s N_VGND_c_1064_n 0.00311299f $X=6.505 $Y=0.235 $X2=0 $Y2=0
cc_582 N_Q_c_997_n N_VGND_c_1064_n 0.0129403f $X=5.88 $Y=0.37 $X2=0 $Y2=0
cc_583 Q N_VGND_c_1064_n 0.00129832f $X=7.095 $Y=0.765 $X2=0 $Y2=0
cc_584 N_Q_c_1015_n N_VGND_c_1064_n 0.0194974f $X=6.575 $Y=1.045 $X2=0 $Y2=0
cc_585 N_Q_c_1018_n N_VGND_c_1064_n 0.00756902f $X=6.66 $Y=0.49 $X2=0 $Y2=0
cc_586 N_VGND_c_1064_n A_466_47# 0.0139156f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_587 N_VGND_c_1064_n A_660_47# 0.00687059f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_588 N_VGND_c_1064_n A_943_47# 0.00323135f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__sdfxtp_1.spice
* Created: Thu Aug 27 14:47:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdfxtp_1.pex.spice"
.subckt sky130_fd_sc_hd__sdfxtp_1  VNB VPB CLK SCE D SCD VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SCD	SCD
* D	D
* SCE	SCE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1029 N_VGND_M1029_d N_CLK_M1029_g N_A_27_47#_M1029_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_193_47#_M1015_d N_A_27_47#_M1015_g N_VGND_M1029_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_SCE_M1031_g N_A_299_47#_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0714 AS=0.1176 PD=0.76 PS=1.4 NRD=17.136 NRS=2.856 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1013 A_483_47# N_A_299_47#_M1013_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0714 PD=0.66 PS=0.76 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1014 N_A_556_369#_M1014_d N_D_M1014_g A_483_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0504 PD=0.75 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1025 A_657_47# N_SCE_M1025_g N_A_556_369#_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0483 AS=0.0693 PD=0.65 PS=0.75 NRD=17.136 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_SCD_M1011_g A_657_47# VNB NSHORT L=0.15 W=0.42 AD=0.1302
+ AS=0.0483 PD=1.46 PS=0.65 NRD=12.852 NRS=17.136 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_A_933_413#_M1030_d N_A_27_47#_M1030_g N_A_556_369#_M1030_s VNB NSHORT
+ L=0.15 W=0.36 AD=0.0594 AS=0.099 PD=0.69 PS=1.27 NRD=18.324 NRS=3.324 M=1
+ R=2.4 SA=75000.2 SB=75003.4 A=0.054 P=1.02 MULT=1
MM1027 A_1030_47# N_A_193_47#_M1027_g N_A_933_413#_M1030_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0634154 AS=0.0594 PD=0.701538 PS=0.69 NRD=40.38 NRS=0 M=1 R=2.4
+ SA=75000.7 SB=75002.9 A=0.054 P=1.02 MULT=1
MM1007 N_VGND_M1007_d N_A_1092_183#_M1007_g A_1030_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.118313 AS=0.0739846 PD=0.966792 PS=0.818462 NRD=47.136 NRS=34.608 M=1
+ R=2.8 SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1016 N_A_1092_183#_M1016_d N_A_933_413#_M1016_g N_VGND_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.126592 AS=0.180287 PD=1.2736 PS=1.47321 NRD=4.68 NRS=25.308
+ M=1 R=4.26667 SA=75001.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1002 N_A_1349_413#_M1002_d N_A_193_47#_M1002_g N_A_1092_183#_M1016_d VNB
+ NSHORT L=0.15 W=0.36 AD=0.0657 AS=0.071208 PD=0.725 PS=0.7164 NRD=26.664
+ NRS=16.656 M=1 R=2.4 SA=75002.4 SB=75001.2 A=0.054 P=1.02 MULT=1
MM1003 A_1478_47# N_A_27_47#_M1003_g N_A_1349_413#_M1002_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0657 PD=0.687692 PS=0.725 NRD=38.076 NRS=1.656 M=1
+ R=2.4 SA=75002.9 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1017 N_VGND_M1017_d N_A_1520_315#_M1017_g A_1478_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_1349_413#_M1004_g N_A_1520_315#_M1004_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.099125 AS=0.169 PD=0.955 PS=1.82 NRD=2.76 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1000 N_Q_M1000_d N_A_1520_315#_M1000_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.099125 PD=1.82 PS=0.955 NRD=0 NRS=1.836 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_CLK_M1005_g N_A_27_47#_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1028 N_A_193_47#_M1028_d N_A_27_47#_M1028_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1018_d N_SCE_M1018_g N_A_299_47#_M1018_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.088 AS=0.1664 PD=0.915 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1010 A_467_369# N_SCE_M1010_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0944 AS=0.088 PD=0.935 PS=0.915 NRD=28.4665 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1021 N_A_556_369#_M1021_d N_D_M1021_g A_467_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.0944 PD=0.91 PS=0.935 NRD=0 NRS=28.4665 M=1 R=4.26667
+ SA=75001.1 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 A_640_369# N_A_299_47#_M1012_g N_A_556_369#_M1021_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0864 PD=0.96 PS=0.91 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_SCD_M1009_g A_640_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1728 AS=0.1024 PD=1.82 PS=0.96 NRD=1.5366 NRS=32.308 M=1 R=4.26667
+ SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_933_413#_M1023_d N_A_193_47#_M1023_g N_A_556_369#_M1023_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06615 AS=0.1281 PD=0.735 PS=1.45 NRD=9.3772 NRS=18.7544 M=1
+ R=2.8 SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1006 A_1026_413# N_A_27_47#_M1006_g N_A_933_413#_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0693 AS=0.06615 PD=0.75 PS=0.735 NRD=51.5943 NRS=7.0329 M=1 R=2.8
+ SA=75000.7 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_A_1092_183#_M1022_g A_1026_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.128423 AS=0.0693 PD=0.904615 PS=0.75 NRD=111.384 NRS=51.5943 M=1
+ R=2.8 SA=75001.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1008 N_A_1092_183#_M1008_d N_A_933_413#_M1008_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.15 W=0.75 AD=0.140385 AS=0.229327 PD=1.37821 PS=1.61538 NRD=0 NRS=0 M=1
+ R=5 SA=75001.2 SB=75001.1 A=0.1125 P=1.8 MULT=1
MM1026 N_A_1349_413#_M1026_d N_A_27_47#_M1026_g N_A_1092_183#_M1008_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0567 AS=0.0786154 PD=0.69 PS=0.771795 NRD=0
+ NRS=23.443 M=1 R=2.8 SA=75002.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1019 A_1433_413# N_A_193_47#_M1019_g N_A_1349_413#_M1026_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09135 AS=0.0567 PD=0.855 PS=0.69 NRD=76.2193 NRS=0 M=1 R=2.8
+ SA=75002.7 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_1520_315#_M1001_g A_1433_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1575 AS=0.09135 PD=1.59 PS=0.855 NRD=49.25 NRS=76.2193 M=1 R=2.8
+ SA=75003.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_1349_413#_M1020_g N_A_1520_315#_M1020_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.1525 AS=0.26 PD=1.305 PS=2.52 NRD=2.9353 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1024 N_Q_M1024_d N_A_1520_315#_M1024_g N_VPWR_M1020_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1525 PD=2.52 PS=1.305 NRD=0 NRS=1.9503 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_110 VNB 0 8.70797e-20 $X=0.145 $Y=-0.085
c_215 VPB 0 1.42307e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__sdfxtp_1.pxi.spice"
*
.ends
*
*

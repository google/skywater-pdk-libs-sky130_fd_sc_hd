* File: sky130_fd_sc_hd__a31oi_1.spice
* Created: Thu Aug 27 14:04:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a31oi_1.spice.pex"
.subckt sky130_fd_sc_hd__a31oi_1  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1007 A_109_47# N_A3_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.169 PD=0.86 PS=1.82 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.5
+ A=0.0975 P=1.6 MULT=1
MM1003 A_181_47# N_A2_M1003_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.118625
+ AS=0.06825 PD=1.015 PS=0.86 NRD=23.532 NRS=9.228 M=1 R=4.33333 SA=75000.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A1_M1004_g A_181_47# VNB NSHORT L=0.15 W=0.65 AD=0.105625
+ AS=0.118625 PD=0.975 PS=1.015 NRD=0 NRS=23.532 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.105625 PD=1.84 PS=0.975 NRD=0.912 NRS=9.228 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_109_297#_M1006_d N_A3_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_109_297#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.135 PD=1.305 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 N_A_109_297#_M1005_d N_A1_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1625 AS=0.1525 PD=1.325 PS=1.305 NRD=0 NRS=5.8903 M=1 R=6.66667
+ SA=75001.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_109_297#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.1625 PD=2.54 PS=1.325 NRD=0.9653 NRS=9.8303 M=1 R=6.66667
+ SA=75001.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__a31oi_1.spice.SKY130_FD_SC_HD__A31OI_1.pxi"
*
.ends
*
*

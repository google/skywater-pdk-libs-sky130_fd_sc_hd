* File: sky130_fd_sc_hd__clkdlybuf4s25_1.pxi.spice
* Created: Tue Sep  1 19:00:51 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A N_A_M1001_g N_A_M1004_g A N_A_c_65_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_27_47# N_A_27_47#_M1001_s
+ N_A_27_47#_M1004_s N_A_27_47#_M1005_g N_A_27_47#_M1007_g N_A_27_47#_c_98_n
+ N_A_27_47#_c_104_n N_A_27_47#_c_99_n N_A_27_47#_c_100_n N_A_27_47#_c_105_n
+ N_A_27_47#_c_106_n N_A_27_47#_c_101_n N_A_27_47#_c_107_n N_A_27_47#_c_102_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_244_47# N_A_244_47#_M1005_d
+ N_A_244_47#_M1007_d N_A_244_47#_M1002_g N_A_244_47#_M1000_g
+ N_A_244_47#_c_167_n N_A_244_47#_c_168_n N_A_244_47#_c_169_n
+ N_A_244_47#_c_170_n N_A_244_47#_c_174_n N_A_244_47#_c_171_n
+ N_A_244_47#_c_172_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_244_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_355_47# N_A_355_47#_M1002_s
+ N_A_355_47#_M1000_s N_A_355_47#_M1006_g N_A_355_47#_M1003_g
+ N_A_355_47#_c_242_n N_A_355_47#_c_243_n N_A_355_47#_c_232_n
+ N_A_355_47#_c_233_n N_A_355_47#_c_237_n N_A_355_47#_c_238_n
+ N_A_355_47#_c_234_n N_A_355_47#_c_240_n N_A_355_47#_c_235_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%A_355_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%VPWR N_VPWR_M1004_d N_VPWR_M1000_d
+ N_VPWR_c_311_n N_VPWR_c_312_n VPWR N_VPWR_c_313_n N_VPWR_c_314_n
+ N_VPWR_c_315_n N_VPWR_c_310_n N_VPWR_c_317_n N_VPWR_c_318_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%X N_X_M1006_d N_X_M1003_d X X X X X X X X
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%VGND N_VGND_M1001_d N_VGND_M1002_d
+ N_VGND_c_373_n VGND N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S25_1%VGND
cc_1 VNB N_A_M1001_g 0.0394167f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.445
cc_2 VNB A 0.00938906f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_65_n 0.0328953f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_4 VNB N_A_27_47#_M1005_g 0.0283759f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_47#_M1007_g 6.23468e-19 $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_6 VNB N_A_27_47#_c_98_n 0.0193059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_99_n 0.00236293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_100_n 0.00990326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_101_n 0.00308192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_102_n 0.0341907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_244_47#_M1002_g 0.0302179f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_12 VNB N_A_244_47#_M1000_g 7.21333e-19 $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_13 VNB N_A_244_47#_c_167_n 0.00473673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_244_47#_c_168_n 0.00835538f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_244_47#_c_169_n 0.0535809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_244_47#_c_170_n 0.00882648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_244_47#_c_171_n 0.00117137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_244_47#_c_172_n 0.00211047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_355_47#_M1006_g 0.0370131f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_A_355_47#_c_232_n 0.00325488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_355_47#_c_233_n 0.00151839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_355_47#_c_234_n 0.0105541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_355_47#_c_235_n 0.0263801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_310_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 0.0165088f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.985
cc_26 VNB X 0.0390164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_373_n 0.00558575f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_28 VNB N_VGND_c_374_n 0.0168024f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_29 VNB N_VGND_c_375_n 0.0231521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_376_n 0.206746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_377_n 0.00631673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_378_n 0.0332818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_379_n 0.0144583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_M1004_g 0.0291685f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_35 VPB A 0.00348705f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_36 VPB N_A_c_65_n 0.00714927f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_37 VPB N_A_27_47#_M1007_g 0.0437201f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_38 VPB N_A_27_47#_c_104_n 0.0319414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_105_n 0.00298872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_106_n 0.00770758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_107_n 0.00177659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_244_47#_M1000_g 0.047741f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_43 VPB N_A_244_47#_c_174_n 0.00978325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_244_47#_c_171_n 0.0101433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_355_47#_M1003_g 0.0251646f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_46 VPB N_A_355_47#_c_237_n 0.0072151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_355_47#_c_238_n 0.00316189f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_355_47#_c_234_n 0.00369559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_355_47#_c_240_n 0.00315466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_355_47#_c_235_n 0.00497508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_311_n 0.00554519f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_52 VPB N_VPWR_c_312_n 0.00422131f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_53 VPB N_VPWR_c_313_n 0.0178727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_314_n 0.0338362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_315_n 0.023341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_310_n 0.0508921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_317_n 0.00622207f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_318_n 0.0103166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB X 0.0138609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB X 0.0116399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 0.0260894f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 N_A_M1001_g N_A_27_47#_M1005_g 0.0191f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_63 N_A_c_65_n N_A_27_47#_M1007_g 0.0315386f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_M1001_g N_A_27_47#_c_98_n 0.0083825f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_65 N_A_M1004_g N_A_27_47#_c_104_n 0.0130364f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1001_g N_A_27_47#_c_99_n 0.0114536f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_67 A N_A_27_47#_c_99_n 0.00519649f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_M1001_g N_A_27_47#_c_100_n 0.00355291f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_69 A N_A_27_47#_c_100_n 0.0270132f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_65_n N_A_27_47#_c_100_n 0.00608644f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_A_27_47#_c_105_n 0.0126616f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_72 A N_A_27_47#_c_105_n 0.00380172f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_A_27_47#_c_106_n 0.00423547f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_74 A N_A_27_47#_c_106_n 0.0266346f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_65_n N_A_27_47#_c_106_n 0.00173603f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_A_27_47#_c_101_n 0.00624254f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_77 A N_A_27_47#_c_101_n 0.0181868f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_78 A N_A_27_47#_c_107_n 0.00186331f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_c_65_n N_A_27_47#_c_107_n 0.0048828f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_65_n N_A_27_47#_c_102_n 0.0160041f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_M1001_g N_A_244_47#_c_170_n 7.61571e-19 $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_M1004_g N_A_244_47#_c_174_n 3.10665e-19 $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_M1004_g N_VPWR_c_311_n 0.00704462f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1004_g N_VPWR_c_313_n 0.0054895f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1004_g N_VPWR_c_310_n 0.0110689f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1001_g N_VGND_c_373_n 0.00323908f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_VGND_c_374_n 0.00438006f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_M1001_g N_VGND_c_376_n 0.00709551f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_27_47#_M1005_g N_A_244_47#_c_167_n 0.00422729f $X=1.095 $Y=0.56 $X2=0
+ $Y2=0
cc_90 N_A_27_47#_c_101_n N_A_244_47#_c_167_n 0.00822194f $X=0.83 $Y=1.295 $X2=0
+ $Y2=0
cc_91 N_A_27_47#_c_102_n N_A_244_47#_c_169_n 0.00461614f $X=1.095 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_M1005_g N_A_244_47#_c_170_n 0.0197049f $X=1.095 $Y=0.56 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_c_101_n N_A_244_47#_c_170_n 0.00983042f $X=0.83 $Y=1.295 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_M1007_g N_A_244_47#_c_174_n 0.0121322f $X=1.095 $Y=2.075 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_105_n N_A_244_47#_c_171_n 0.00635339f $X=0.655 $Y=1.575 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_c_101_n N_A_244_47#_c_171_n 0.00194246f $X=0.83 $Y=1.295 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_107_n N_A_244_47#_c_171_n 0.00689186f $X=0.83 $Y=1.49 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_c_102_n N_A_244_47#_c_171_n 0.0128123f $X=1.095 $Y=1.16 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_101_n N_A_244_47#_c_172_n 0.00854995f $X=0.83 $Y=1.295 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_102_n N_A_244_47#_c_172_n 0.00202606f $X=1.095 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_M1005_g N_A_355_47#_c_242_n 8.06133e-19 $X=1.095 $Y=0.56 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_M1007_g N_A_355_47#_c_243_n 7.6947e-19 $X=1.095 $Y=2.075 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_M1005_g N_A_355_47#_c_233_n 4.04566e-19 $X=1.095 $Y=0.56 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_105_n N_VPWR_M1004_d 0.00338617f $X=0.655 $Y=1.575 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_27_47#_M1007_g N_VPWR_c_311_n 0.00757328f $X=1.095 $Y=2.075 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_105_n N_VPWR_c_311_n 0.0273849f $X=0.655 $Y=1.575 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_102_n N_VPWR_c_311_n 5.35972e-19 $X=1.095 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_c_104_n N_VPWR_c_313_n 0.0221174f $X=0.265 $Y=1.995 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_M1007_g N_VPWR_c_314_n 0.00939206f $X=1.095 $Y=2.075 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_M1004_s N_VPWR_c_310_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_M1007_g N_VPWR_c_310_n 0.0176049f $X=1.095 $Y=2.075 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_c_104_n N_VPWR_c_310_n 0.0130273f $X=0.265 $Y=1.995 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_101_n N_VGND_M1001_d 0.00302667f $X=0.83 $Y=1.295 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_27_47#_M1005_g N_VGND_c_373_n 0.00709904f $X=1.095 $Y=0.56 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_99_n N_VGND_c_373_n 0.00448114f $X=0.655 $Y=0.82 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_101_n N_VGND_c_373_n 0.0220299f $X=0.83 $Y=1.295 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_102_n N_VGND_c_373_n 5.61301e-19 $X=1.095 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_c_98_n N_VGND_c_374_n 0.0206917f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_99_n N_VGND_c_374_n 0.00226107f $X=0.655 $Y=0.82 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1001_s N_VGND_c_376_n 0.00217517f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_M1005_g N_VGND_c_376_n 0.0158083f $X=1.095 $Y=0.56 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_98_n N_VGND_c_376_n 0.0123339f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_99_n N_VGND_c_376_n 0.00396529f $X=0.655 $Y=0.82 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_101_n N_VGND_c_376_n 0.00359769f $X=0.83 $Y=1.295 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_M1005_g N_VGND_c_378_n 0.00874704f $X=1.095 $Y=0.56 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_c_101_n N_VGND_c_378_n 9.77487e-19 $X=0.83 $Y=1.295 $X2=0
+ $Y2=0
cc_127 N_A_244_47#_M1002_g N_A_355_47#_M1006_g 0.0134495f $X=2.165 $Y=0.56 $X2=0
+ $Y2=0
cc_128 N_A_244_47#_M1000_g N_A_355_47#_M1003_g 0.0181181f $X=2.165 $Y=2.075
+ $X2=0 $Y2=0
cc_129 N_A_244_47#_M1002_g N_A_355_47#_c_242_n 0.0148195f $X=2.165 $Y=0.56 $X2=0
+ $Y2=0
cc_130 N_A_244_47#_c_170_n N_A_355_47#_c_242_n 0.0395108f $X=1.36 $Y=0.4 $X2=0
+ $Y2=0
cc_131 N_A_244_47#_M1000_g N_A_355_47#_c_243_n 0.0195096f $X=2.165 $Y=2.075
+ $X2=0 $Y2=0
cc_132 N_A_244_47#_c_171_n N_A_355_47#_c_243_n 0.0648823f $X=1.42 $Y=1.79 $X2=0
+ $Y2=0
cc_133 N_A_244_47#_M1002_g N_A_355_47#_c_232_n 0.0147913f $X=2.165 $Y=0.56 $X2=0
+ $Y2=0
cc_134 N_A_244_47#_c_168_n N_A_355_47#_c_232_n 0.024568f $X=2.255 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_244_47#_c_169_n N_A_355_47#_c_232_n 0.00296734f $X=2.255 $Y=1.16
+ $X2=0 $Y2=0
cc_136 N_A_244_47#_M1002_g N_A_355_47#_c_233_n 0.00395296f $X=2.165 $Y=0.56
+ $X2=0 $Y2=0
cc_137 N_A_244_47#_c_168_n N_A_355_47#_c_233_n 0.0199832f $X=2.255 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_244_47#_c_169_n N_A_355_47#_c_233_n 0.00531537f $X=2.255 $Y=1.16
+ $X2=0 $Y2=0
cc_139 N_A_244_47#_c_170_n N_A_355_47#_c_233_n 0.0148182f $X=1.36 $Y=0.4 $X2=0
+ $Y2=0
cc_140 N_A_244_47#_M1000_g N_A_355_47#_c_237_n 0.0185718f $X=2.165 $Y=2.075
+ $X2=0 $Y2=0
cc_141 N_A_244_47#_c_168_n N_A_355_47#_c_237_n 0.0184842f $X=2.255 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_244_47#_c_169_n N_A_355_47#_c_237_n 0.00280725f $X=2.255 $Y=1.16
+ $X2=0 $Y2=0
cc_143 N_A_244_47#_M1000_g N_A_355_47#_c_238_n 0.00402784f $X=2.165 $Y=2.075
+ $X2=0 $Y2=0
cc_144 N_A_244_47#_c_168_n N_A_355_47#_c_238_n 0.0152539f $X=2.255 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_244_47#_c_169_n N_A_355_47#_c_238_n 0.0050987f $X=2.255 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_244_47#_c_171_n N_A_355_47#_c_238_n 0.0143863f $X=1.42 $Y=1.79 $X2=0
+ $Y2=0
cc_147 N_A_244_47#_M1002_g N_A_355_47#_c_234_n 0.00259068f $X=2.165 $Y=0.56
+ $X2=0 $Y2=0
cc_148 N_A_244_47#_M1000_g N_A_355_47#_c_234_n 7.03652e-19 $X=2.165 $Y=2.075
+ $X2=0 $Y2=0
cc_149 N_A_244_47#_c_168_n N_A_355_47#_c_234_n 0.014622f $X=2.255 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_244_47#_c_169_n N_A_355_47#_c_234_n 0.00334716f $X=2.255 $Y=1.16
+ $X2=0 $Y2=0
cc_151 N_A_244_47#_M1000_g N_A_355_47#_c_240_n 0.00348724f $X=2.165 $Y=2.075
+ $X2=0 $Y2=0
cc_152 N_A_244_47#_M1002_g N_A_355_47#_c_235_n 5.65741e-19 $X=2.165 $Y=0.56
+ $X2=0 $Y2=0
cc_153 N_A_244_47#_M1000_g N_A_355_47#_c_235_n 5.65741e-19 $X=2.165 $Y=2.075
+ $X2=0 $Y2=0
cc_154 N_A_244_47#_c_169_n N_A_355_47#_c_235_n 0.00873969f $X=2.255 $Y=1.16
+ $X2=0 $Y2=0
cc_155 N_A_244_47#_M1000_g N_VPWR_c_312_n 0.0329643f $X=2.165 $Y=2.075 $X2=0
+ $Y2=0
cc_156 N_A_244_47#_M1000_g N_VPWR_c_314_n 0.00722788f $X=2.165 $Y=2.075 $X2=0
+ $Y2=0
cc_157 N_A_244_47#_c_174_n N_VPWR_c_314_n 0.0296441f $X=1.36 $Y=1.995 $X2=0
+ $Y2=0
cc_158 N_A_244_47#_M1007_d N_VPWR_c_310_n 0.00213418f $X=1.22 $Y=1.665 $X2=0
+ $Y2=0
cc_159 N_A_244_47#_M1000_g N_VPWR_c_310_n 0.0129983f $X=2.165 $Y=2.075 $X2=0
+ $Y2=0
cc_160 N_A_244_47#_c_174_n N_VPWR_c_310_n 0.017069f $X=1.36 $Y=1.995 $X2=0 $Y2=0
cc_161 N_A_244_47#_c_170_n N_VGND_c_373_n 0.0175745f $X=1.36 $Y=0.4 $X2=0 $Y2=0
cc_162 N_A_244_47#_M1005_d N_VGND_c_376_n 0.00213418f $X=1.22 $Y=0.235 $X2=0
+ $Y2=0
cc_163 N_A_244_47#_M1002_g N_VGND_c_376_n 0.0077411f $X=2.165 $Y=0.56 $X2=0
+ $Y2=0
cc_164 N_A_244_47#_c_170_n N_VGND_c_376_n 0.0177132f $X=1.36 $Y=0.4 $X2=0 $Y2=0
cc_165 N_A_244_47#_M1002_g N_VGND_c_378_n 0.00572733f $X=2.165 $Y=0.56 $X2=0
+ $Y2=0
cc_166 N_A_244_47#_c_170_n N_VGND_c_378_n 0.0308657f $X=1.36 $Y=0.4 $X2=0 $Y2=0
cc_167 N_A_244_47#_M1002_g N_VGND_c_379_n 0.0204027f $X=2.165 $Y=0.56 $X2=0
+ $Y2=0
cc_168 N_A_355_47#_c_237_n N_VPWR_M1000_d 0.00484989f $X=2.595 $Y=1.58 $X2=0
+ $Y2=0
cc_169 N_A_355_47#_M1003_g N_VPWR_c_312_n 0.00867095f $X=2.975 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_355_47#_c_243_n N_VPWR_c_312_n 0.0486212f $X=1.9 $Y=1.96 $X2=0 $Y2=0
cc_171 N_A_355_47#_c_237_n N_VPWR_c_312_n 0.0420202f $X=2.595 $Y=1.58 $X2=0
+ $Y2=0
cc_172 N_A_355_47#_c_234_n N_VPWR_c_312_n 0.00282779f $X=2.68 $Y=1.325 $X2=0
+ $Y2=0
cc_173 N_A_355_47#_c_235_n N_VPWR_c_312_n 4.21248e-19 $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_174 N_A_355_47#_c_243_n N_VPWR_c_314_n 0.0153696f $X=1.9 $Y=1.96 $X2=0 $Y2=0
cc_175 N_A_355_47#_M1003_g N_VPWR_c_315_n 0.00564131f $X=2.975 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_355_47#_M1000_s N_VPWR_c_310_n 0.00355752f $X=1.775 $Y=1.665 $X2=0
+ $Y2=0
cc_177 N_A_355_47#_M1003_g N_VPWR_c_310_n 0.01194f $X=2.975 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_355_47#_c_243_n N_VPWR_c_310_n 0.00936871f $X=1.9 $Y=1.96 $X2=0 $Y2=0
cc_179 N_A_355_47#_M1006_g X 0.00906555f $X=2.975 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A_355_47#_c_234_n X 0.00149519f $X=2.68 $Y=1.325 $X2=0 $Y2=0
cc_181 N_A_355_47#_M1006_g X 0.0118614f $X=2.975 $Y=0.445 $X2=0 $Y2=0
cc_182 N_A_355_47#_M1003_g X 0.00548454f $X=2.975 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_355_47#_c_237_n X 0.00282048f $X=2.595 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A_355_47#_c_234_n X 0.0368768f $X=2.68 $Y=1.325 $X2=0 $Y2=0
cc_185 N_A_355_47#_c_240_n X 0.00666717f $X=2.68 $Y=1.495 $X2=0 $Y2=0
cc_186 N_A_355_47#_M1003_g X 0.0138754f $X=2.975 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_355_47#_c_237_n X 0.00600589f $X=2.595 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A_355_47#_c_234_n X 8.51344e-19 $X=2.68 $Y=1.325 $X2=0 $Y2=0
cc_189 N_A_355_47#_M1003_g X 0.00659964f $X=2.975 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_355_47#_c_232_n N_VGND_M1002_d 0.00359381f $X=2.595 $Y=0.82 $X2=0
+ $Y2=0
cc_191 N_A_355_47#_c_234_n N_VGND_M1002_d 0.00457774f $X=2.68 $Y=1.325 $X2=0
+ $Y2=0
cc_192 N_A_355_47#_M1006_g N_VGND_c_375_n 0.005323f $X=2.975 $Y=0.445 $X2=0
+ $Y2=0
cc_193 N_A_355_47#_M1002_s N_VGND_c_376_n 0.00355752f $X=1.775 $Y=0.235 $X2=0
+ $Y2=0
cc_194 N_A_355_47#_M1006_g N_VGND_c_376_n 0.0111608f $X=2.975 $Y=0.445 $X2=0
+ $Y2=0
cc_195 N_A_355_47#_c_242_n N_VGND_c_376_n 0.00935749f $X=1.9 $Y=0.42 $X2=0 $Y2=0
cc_196 N_A_355_47#_c_232_n N_VGND_c_376_n 0.00502649f $X=2.595 $Y=0.82 $X2=0
+ $Y2=0
cc_197 N_A_355_47#_c_234_n N_VGND_c_376_n 7.24644e-19 $X=2.68 $Y=1.325 $X2=0
+ $Y2=0
cc_198 N_A_355_47#_c_242_n N_VGND_c_378_n 0.0153256f $X=1.9 $Y=0.42 $X2=0 $Y2=0
cc_199 N_A_355_47#_c_232_n N_VGND_c_378_n 0.00228044f $X=2.595 $Y=0.82 $X2=0
+ $Y2=0
cc_200 N_A_355_47#_M1006_g N_VGND_c_379_n 0.006114f $X=2.975 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_355_47#_c_242_n N_VGND_c_379_n 0.0233972f $X=1.9 $Y=0.42 $X2=0 $Y2=0
cc_202 N_A_355_47#_c_232_n N_VGND_c_379_n 0.02298f $X=2.595 $Y=0.82 $X2=0 $Y2=0
cc_203 N_A_355_47#_c_234_n N_VGND_c_379_n 0.0182037f $X=2.68 $Y=1.325 $X2=0
+ $Y2=0
cc_204 N_A_355_47#_c_235_n N_VGND_c_379_n 4.33043e-19 $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_310_n N_X_M1003_d 0.00401972f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_206 N_VPWR_c_315_n X 0.0372578f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_207 N_VPWR_c_310_n X 0.0213531f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_208 X N_VGND_c_375_n 0.0370374f $X=3.36 $Y=0.425 $X2=0 $Y2=0
cc_209 N_X_M1006_d N_VGND_c_376_n 0.00402019f $X=3.05 $Y=0.235 $X2=0 $Y2=0
cc_210 X N_VGND_c_376_n 0.0217739f $X=3.36 $Y=0.425 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_8.pex.spice
* Created: Tue Sep  1 19:10:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%A 3 5 7 10 12 14 15 16 24
c43 15 0 1.46759e-19 $X=0.23 $Y=0.85
r44 23 24 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.155
+ $X2=0.905 $Y2=1.155
r45 20 23 21.5061 $w=5.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.155
+ $X2=0.475 $Y2=1.155
r46 16 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r47 15 16 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=0.242 $Y=0.85
+ $X2=0.242 $Y2=1.16
r48 12 24 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.155
r49 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.985
r50 8 24 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=1.155
r51 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=0.445
r52 5 23 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.155
r53 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.985
r54 1 23 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=1.155
r55 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%A_110_47# 1 2 9 13 17 21 25 29
+ 33 37 41 45 49 53 57 61 63 65 69 73 77 84 87
r170 84 85 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.245
+ $Y=1.16 $X2=3.245 $Y2=1.16
r171 81 84 78.3661 $w=2.48e-07 $l=1.7e-06 $layer=LI1_cond $X=1.545 $Y=1.2
+ $X2=3.245 $Y2=1.2
r172 81 82 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.545
+ $Y=1.16 $X2=1.545 $Y2=1.16
r173 79 87 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=1.2
+ $X2=0.695 $Y2=1.2
r174 79 81 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=0.82 $Y=1.2
+ $X2=1.545 $Y2=1.2
r175 75 87 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.695 $Y2=1.2
r176 75 77 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.695 $Y2=1.69
r177 71 87 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.075
+ $X2=0.695 $Y2=1.2
r178 71 73 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=0.695 $Y=1.075
+ $X2=0.695 $Y2=0.445
r179 67 69 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.345 $Y=1.325
+ $X2=4.345 $Y2=1.985
r180 63 67 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=4.345 $Y=1.137
+ $X2=4.345 $Y2=1.325
r181 63 65 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.345 $Y=0.95
+ $X2=4.345 $Y2=0.445
r182 59 61 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.915 $Y=1.325
+ $X2=3.915 $Y2=1.985
r183 55 63 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=4.345 $Y2=1.137
r184 55 59 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=3.915 $Y2=1.325
r185 55 57 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.915 $Y=0.95
+ $X2=3.915 $Y2=0.445
r186 51 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.485 $Y=1.325
+ $X2=3.485 $Y2=1.985
r187 47 55 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.915 $Y2=1.137
r188 47 51 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.485 $Y2=1.325
r189 47 85 35.5938 $w=3.75e-07 $l=2.4e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.245 $Y2=1.137
r190 47 49 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.485 $Y=0.95
+ $X2=3.485 $Y2=0.445
r191 43 45 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.055 $Y=1.325
+ $X2=3.055 $Y2=1.985
r192 39 85 28.1785 $w=3.75e-07 $l=1.9e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.245 $Y2=1.137
r193 39 43 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.055 $Y2=1.325
r194 39 41 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.055 $Y=0.95
+ $X2=3.055 $Y2=0.445
r195 35 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.625 $Y=1.325
+ $X2=2.625 $Y2=1.985
r196 31 39 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=3.055 $Y2=1.137
r197 31 35 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=2.625 $Y2=1.325
r198 31 33 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.625 $Y=0.95
+ $X2=2.625 $Y2=0.445
r199 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.195 $Y=1.325
+ $X2=2.195 $Y2=1.985
r200 23 31 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.625 $Y2=1.137
r201 23 27 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.195 $Y2=1.325
r202 23 25 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.195 $Y=0.95
+ $X2=2.195 $Y2=0.445
r203 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=1.325
+ $X2=1.765 $Y2=1.985
r204 15 23 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=1.765 $Y=1.137
+ $X2=2.195 $Y2=1.137
r205 15 19 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=1.765 $Y=1.137
+ $X2=1.765 $Y2=1.325
r206 15 82 32.6277 $w=3.75e-07 $l=2.2e-07 $layer=POLY_cond $X=1.765 $Y=1.137
+ $X2=1.545 $Y2=1.137
r207 15 17 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.765 $Y=0.95
+ $X2=1.765 $Y2=0.445
r208 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=1.985
r209 7 82 31.1446 $w=3.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.335 $Y=1.137
+ $X2=1.545 $Y2=1.137
r210 7 11 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=1.335 $Y=1.137
+ $X2=1.335 $Y2=1.325
r211 7 9 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.335 $Y=0.95
+ $X2=1.335 $Y2=0.445
r212 2 77 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.69
r213 1 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%KAPWR 1 2 3 4 5 6 20 34 35 38
+ 39 40 43 44 45 48 49 50 52 53 54 56 59 66
c108 52 0 1.98896e-19 $X=4.565 $Y=2.21
c109 45 0 1.77237e-19 $X=2.97 $Y=2.21
c110 6 0 4.2343e-20 $X=4.42 $Y=1.485
c111 5 0 1.26035e-19 $X=3.56 $Y=1.485
r112 59 62 20.3142 $w=2.93e-07 $l=5.2e-07 $layer=LI1_cond $X=0.242 $Y=1.69
+ $X2=0.242 $Y2=2.21
r113 56 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=2.21
+ $X2=0.26 $Y2=2.21
r114 52 54 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=4.565 $Y=2.21
+ $X2=4.42 $Y2=2.21
r115 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.565 $Y=2.21
+ $X2=4.565 $Y2=2.21
r116 50 54 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=3.85 $Y=2.24
+ $X2=4.42 $Y2=2.24
r117 47 50 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.705 $Y=2.21
+ $X2=3.85 $Y2=2.21
r118 47 49 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=3.705 $Y=2.21
+ $X2=3.56 $Y2=2.21
r119 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.705 $Y=2.21
+ $X2=3.705 $Y2=2.21
r120 45 49 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=2.97 $Y=2.24
+ $X2=3.56 $Y2=2.24
r121 42 45 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.825 $Y=2.21
+ $X2=2.97 $Y2=2.21
r122 42 44 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=2.825 $Y=2.21
+ $X2=2.68 $Y2=2.21
r123 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.825 $Y=2.21
+ $X2=2.825 $Y2=2.21
r124 40 44 0.429825 $w=2e-07 $l=5.6e-07 $layer=MET1_cond $X=2.12 $Y=2.24
+ $X2=2.68 $Y2=2.24
r125 37 40 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=2.12 $Y2=2.21
r126 37 39 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.975 $Y=2.21
+ $X2=1.83 $Y2=2.21
r127 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.975 $Y=2.21
+ $X2=1.975 $Y2=2.21
r128 35 39 0.433663 $w=2e-07 $l=5.65e-07 $layer=MET1_cond $X=1.265 $Y=2.24
+ $X2=1.83 $Y2=2.24
r129 33 66 23.0489 $w=2.58e-07 $l=5.2e-07 $layer=LI1_cond $X=1.12 $Y=2.21
+ $X2=1.12 $Y2=1.69
r130 32 35 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.12 $Y=2.21
+ $X2=1.265 $Y2=2.21
r131 32 34 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.12 $Y=2.21
+ $X2=0.975 $Y2=2.21
r132 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=2.21
+ $X2=1.12 $Y2=2.21
r133 20 56 0.0777288 $w=2.51e-07 $l=1.59295e-07 $layer=MET1_cond $X=0.405
+ $Y=2.24 $X2=0.26 $Y2=2.21
r134 20 34 0.437501 $w=2e-07 $l=5.7e-07 $layer=MET1_cond $X=0.405 $Y=2.24
+ $X2=0.975 $Y2=2.24
r135 6 53 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.485 $X2=4.56 $Y2=2.22
r136 5 48 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.485 $X2=3.7 $Y2=2.22
r137 4 43 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.485 $X2=2.84 $Y2=2.22
r138 3 38 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.485 $X2=1.98 $Y2=2.22
r139 2 66 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=1.69
r140 1 59 300 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.69
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%X 1 2 3 4 5 6 7 8 27 31 32 33
+ 37 41 43 47 51 53 57 62 63 65 66 68 69 70 71
c153 69 0 1.68378e-19 $X=4.37 $Y=0.85
r154 71 86 2.23356 $w=6.15e-07 $l=1.2e-07 $layer=LI1_cond $X=4.245 $Y=1.615
+ $X2=4.245 $Y2=1.495
r155 71 86 0.314433 $w=9.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.245 $Y=1.47
+ $X2=4.245 $Y2=1.495
r156 70 71 3.52165 $w=9.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.245 $Y=1.19
+ $X2=4.245 $Y2=1.47
r157 69 85 1.61223 $w=6.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.82
+ $X2=4.245 $Y2=0.905
r158 69 70 3.39588 $w=9.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.245 $Y=0.92
+ $X2=4.245 $Y2=1.19
r159 69 85 0.18866 $w=9.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.245 $Y=0.92
+ $X2=4.245 $Y2=0.905
r160 55 69 1.61223 $w=6.15e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.245 $Y2=0.82
r161 55 57 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.445
r162 54 68 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=1.615
+ $X2=3.27 $Y2=1.615
r163 53 71 4.87019 $w=2.4e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=1.615
+ $X2=4.245 $Y2=1.615
r164 53 54 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=1.615
+ $X2=3.4 $Y2=1.615
r165 52 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=0.82 $X2=3.27
+ $Y2=0.82
r166 51 69 6.19726 $w=1.7e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=0.82
+ $X2=4.245 $Y2=0.82
r167 51 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=0.82
+ $X2=3.4 $Y2=0.82
r168 45 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.82
r169 45 47 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.445
r170 44 65 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=1.615
+ $X2=2.41 $Y2=1.615
r171 43 68 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=3.27 $Y2=1.615
r172 43 44 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=2.54 $Y2=1.615
r173 42 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=0.82
+ $X2=2.41 $Y2=0.82
r174 41 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=0.82
+ $X2=3.27 $Y2=0.82
r175 41 42 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=0.82 $X2=2.54
+ $Y2=0.82
r176 35 63 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.82
r177 35 37 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.445
r178 34 62 3.55196 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=1.55 $Y2=1.615
r179 33 65 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=1.615
+ $X2=2.41 $Y2=1.615
r180 33 34 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=1.615
+ $X2=1.68 $Y2=1.615
r181 31 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=0.82
+ $X2=2.41 $Y2=0.82
r182 31 32 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=0.82 $X2=1.68
+ $Y2=0.82
r183 25 32 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.68 $Y2=0.82
r184 25 27 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.55 $Y2=0.445
r185 8 71 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.485 $X2=4.13 $Y2=1.69
r186 7 68 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=1.485 $X2=3.27 $Y2=1.69
r187 6 65 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.485 $X2=2.41 $Y2=1.69
r188 5 62 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.485 $X2=1.55 $Y2=1.69
r189 4 57 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.445
r190 3 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.445
r191 2 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.445
r192 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%VGND 1 2 3 4 5 6 19 21 25 29 33
+ 37 41 44 45 47 48 50 51 53 54 55 57 76 77 83
c84 57 0 1.46759e-19 $X=0.99 $Y=0
r85 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r86 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r87 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r88 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r89 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r90 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r91 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r92 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r93 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r94 65 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r95 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r96 62 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.12
+ $Y2=0
r97 62 64 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.61
+ $Y2=0
r98 61 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r99 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r100 58 80 3.93884 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r101 58 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.69
+ $Y2=0
r102 57 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.12
+ $Y2=0
r103 57 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.69
+ $Y2=0
r104 55 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r105 55 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r106 53 73 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.37
+ $Y2=0
r107 53 54 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.58
+ $Y2=0
r108 52 76 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.83
+ $Y2=0
r109 52 54 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.58
+ $Y2=0
r110 50 70 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.45
+ $Y2=0
r111 50 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.7
+ $Y2=0
r112 49 73 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.37
+ $Y2=0
r113 49 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.7
+ $Y2=0
r114 47 67 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.53
+ $Y2=0
r115 47 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.84
+ $Y2=0
r116 46 70 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=3.45
+ $Y2=0
r117 46 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.84
+ $Y2=0
r118 44 64 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.61
+ $Y2=0
r119 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.98
+ $Y2=0
r120 43 67 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.53
+ $Y2=0
r121 43 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.98
+ $Y2=0
r122 39 54 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r123 39 41 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.4
r124 35 51 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r125 35 37 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.4
r126 31 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r127 31 33 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.4
r128 27 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r129 27 29 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.4
r130 23 83 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r131 23 25 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.445
r132 19 80 3.17127 $w=2.45e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.195 $Y2=0
r133 19 21 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.267 $Y2=0.38
r134 6 41 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.235 $X2=4.565 $Y2=0.4
r135 5 37 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.4
r136 4 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.4
r137 3 29 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.4
r138 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.445
r139 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_8%VPWR 1 8 9
c67 8 0 3.76133e-19 $X=4.83 $Y=2.72
r68 8 9 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r69 4 8 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=4.83
+ $Y2=2.72
r70 1 9 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=4.83
+ $Y2=2.72
r71 1 4 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
.ends


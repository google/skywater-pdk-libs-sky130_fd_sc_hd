* File: sky130_fd_sc_hd__nand4bb_1.spice.pex
* Created: Thu Aug 27 14:30:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%B_N 3 6 8 9 13 14 15
c29 15 0 6.81442e-20 $X=0.562 $Y=0.995
r30 13 16 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=1.325
r31 13 15 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=0.995
r32 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r33 8 9 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.53
r34 8 14 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.16
r35 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r36 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%D 3 6 8 11 13
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.16
+ $X2=1.105 $Y2=1.325
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.16
+ $X2=1.105 $Y2=0.995
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=1.16 $X2=1.135 $Y2=1.16
r37 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.015 $Y=1.985
+ $X2=1.015 $Y2=1.325
r38 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.015 $Y=0.56
+ $X2=1.015 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%C 3 6 8 9 13 15
r36 13 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.16
+ $X2=1.625 $Y2=1.325
r37 13 15 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.16
+ $X2=1.625 $Y2=0.995
r38 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.16 $X2=1.635 $Y2=1.16
r39 8 9 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=1.61 $Y=0.85 $X2=1.61
+ $Y2=1.16
r40 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.555 $Y=1.985
+ $X2=1.555 $Y2=1.325
r41 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.555 $Y=0.56
+ $X2=1.555 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%A_27_93# 1 2 9 12 16 19 20 21 24 25 28 33
+ 34 37
c82 21 0 6.81442e-20 $X=1.27 $Y=0.46
r83 33 34 12.0264 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=0.255 $Y=2.34
+ $X2=0.255 $Y2=2.065
r84 31 34 73.5169 $w=1.73e-07 $l=1.16e-06 $layer=LI1_cond $X=0.172 $Y=0.905
+ $X2=0.172 $Y2=2.065
r85 30 31 5.92518 $w=3.38e-07 $l=9.5e-08 $layer=LI1_cond $X=0.255 $Y=0.81
+ $X2=0.255 $Y2=0.905
r86 28 30 6.77908 $w=3.38e-07 $l=2e-07 $layer=LI1_cond $X=0.255 $Y=0.61
+ $X2=0.255 $Y2=0.81
r87 25 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.16
+ $X2=2.115 $Y2=1.325
r88 25 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.16
+ $X2=2.115 $Y2=0.995
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=1.16 $X2=2.115 $Y2=1.16
r90 22 24 24.901 $w=2.78e-07 $l=6.05e-07 $layer=LI1_cond $X=2.11 $Y=0.555
+ $X2=2.11 $Y2=1.16
r91 20 22 7.1467 $w=1.9e-07 $l=1.81384e-07 $layer=LI1_cond $X=1.97 $Y=0.46
+ $X2=2.11 $Y2=0.555
r92 20 21 40.8612 $w=1.88e-07 $l=7e-07 $layer=LI1_cond $X=1.97 $Y=0.46 $X2=1.27
+ $Y2=0.46
r93 18 21 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.27 $Y2=0.46
r94 18 19 9.33971 $w=1.88e-07 $l=1.6e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.175 $Y2=0.715
r95 17 30 4.14298 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=0.425 $Y=0.81
+ $X2=0.255 $Y2=0.81
r96 16 19 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=1.08 $Y=0.81
+ $X2=1.175 $Y2=0.715
r97 16 17 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=1.08 $Y=0.81
+ $X2=0.425 $Y2=0.81
r98 12 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.055 $Y=1.985
+ $X2=2.055 $Y2=1.325
r99 9 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.055 $Y=0.56
+ $X2=2.055 $Y2=0.995
r100 2 33 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.34
r101 1 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%A_496_21# 1 2 7 9 12 15 18 19 21 22 25 28
+ 32 34
r66 30 32 5.2456 $w=2.88e-07 $l=1.32e-07 $layer=LI1_cond $X=3.8 $Y=0.4 $X2=3.932
+ $Y2=0.4
r67 28 34 2.86771 $w=3.32e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.932 $Y=1.835
+ $X2=3.845 $Y2=1.92
r68 27 32 1.74699 $w=2.45e-07 $l=1.45e-07 $layer=LI1_cond $X=3.932 $Y=0.545
+ $X2=3.932 $Y2=0.4
r69 27 28 60.6797 $w=2.43e-07 $l=1.29e-06 $layer=LI1_cond $X=3.932 $Y=0.545
+ $X2=3.932 $Y2=1.835
r70 23 34 2.86771 $w=3.32e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=2.005
+ $X2=3.845 $Y2=1.92
r71 23 25 9.19211 $w=4.18e-07 $l=3.35e-07 $layer=LI1_cond $X=3.845 $Y=2.005
+ $X2=3.845 $Y2=2.34
r72 21 34 3.83825 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.635 $Y=1.92
+ $X2=3.845 $Y2=1.92
r73 21 22 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.635 $Y=1.92
+ $X2=3.09 $Y2=1.92
r74 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.925
+ $Y=1.16 $X2=2.925 $Y2=1.16
r75 16 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.965 $Y=1.835
+ $X2=3.09 $Y2=1.92
r76 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.965 $Y=1.835
+ $X2=2.965 $Y2=1.16
r77 14 19 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=2.63 $Y=1.16
+ $X2=2.925 $Y2=1.16
r78 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.63 $Y=1.16
+ $X2=2.555 $Y2=1.16
r79 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.555 $Y=1.325
+ $X2=2.555 $Y2=1.16
r80 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.555 $Y=1.325
+ $X2=2.555 $Y2=1.985
r81 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.555 $Y=0.995
+ $X2=2.555 $Y2=1.16
r82 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.555 $Y=0.995
+ $X2=2.555 $Y2=0.56
r83 2 25 600 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=2.065 $X2=3.8 $Y2=2.34
r84 1 30 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.8 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%A_N 3 7 9 10 11 16
r33 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.155
+ $X2=3.555 $Y2=1.32
r34 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.155
+ $X2=3.555 $Y2=0.99
r35 10 11 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=3.515 $Y=1.155
+ $X2=3.515 $Y2=1.53
r36 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.555
+ $Y=1.155 $X2=3.555 $Y2=1.155
r37 9 10 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=3.515 $Y=0.85
+ $X2=3.515 $Y2=1.155
r38 7 19 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=3.495 $Y=2.275
+ $X2=3.495 $Y2=1.32
r39 3 18 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.495 $Y=0.445
+ $X2=3.495 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%VPWR 1 2 3 4 15 19 22 23 24 26 41 42 45 49
+ 55
r55 54 55 10.3517 $w=6.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=2.49
+ $X2=3.45 $Y2=2.49
r56 51 54 5.60068 $w=6.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=2.49
+ $X2=3.285 $Y2=2.49
r57 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 48 51 4.27171 $w=6.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.765 $Y=2.49
+ $X2=2.99 $Y2=2.49
r59 48 49 8.83288 $w=6.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=2.49
+ $X2=2.68 $Y2=2.49
r60 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 42 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 41 55 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r63 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r65 37 49 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=2.72 $X2=2.68
+ $Y2=2.72
r66 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r67 34 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r68 34 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r70 31 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.76 $Y2=2.72
r71 31 33 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.76 $Y2=2.72
r73 26 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 24 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r76 22 33 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.64 $Y=2.72 $X2=1.61
+ $Y2=2.72
r77 22 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=2.72
+ $X2=1.805 $Y2=2.72
r78 21 37 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.97 $Y=2.72
+ $X2=2.53 $Y2=2.72
r79 21 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=2.72
+ $X2=1.805 $Y2=2.72
r80 17 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=2.635
+ $X2=1.805 $Y2=2.72
r81 17 19 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.805 $Y=2.635
+ $X2=1.805 $Y2=2
r82 13 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=2.72
r83 13 15 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=1.92
r84 4 54 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=2.065 $X2=3.285 $Y2=2.34
r85 3 48 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.485 $X2=2.765 $Y2=2.34
r86 2 19 300 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=2 $X=1.63
+ $Y=1.485 $X2=1.805 $Y2=2
r87 1 15 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=2.065 $X2=0.76 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%Y 1 2 3 10 12 14 18 22 23 24 25 35 41
r42 35 46 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.545 $Y=0.85
+ $X2=2.545 $Y2=0.825
r43 25 33 3.24686 $w=2.9e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.405 $Y=1.58
+ $X2=2.545 $Y2=1.495
r44 25 33 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.545 $Y=1.47
+ $X2=2.545 $Y2=1.495
r45 24 25 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.545 $Y=1.19
+ $X2=2.545 $Y2=1.47
r46 23 46 3.81656 $w=5.08e-07 $l=3e-08 $layer=LI1_cond $X=2.675 $Y=0.795
+ $X2=2.675 $Y2=0.825
r47 23 24 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=2.545 $Y=0.88
+ $X2=2.545 $Y2=1.19
r48 23 35 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=2.545 $Y=0.88
+ $X2=2.545 $Y2=0.85
r49 22 23 6.68397 $w=5.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.675 $Y=0.51
+ $X2=2.675 $Y2=0.795
r50 22 41 3.04883 $w=5.08e-07 $l=1.3e-07 $layer=LI1_cond $X=2.675 $Y=0.51
+ $X2=2.675 $Y2=0.38
r51 16 25 3.24686 $w=2.9e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.305 $Y=1.665
+ $X2=2.405 $Y2=1.58
r52 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.305 $Y=1.665
+ $X2=2.305 $Y2=2.34
r53 15 21 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=1.58
+ $X2=1.285 $Y2=1.58
r54 14 25 3.3199 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=2.14 $Y=1.58
+ $X2=2.405 $Y2=1.58
r55 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.14 $Y=1.58 $X2=1.45
+ $Y2=1.58
r56 10 21 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.665
+ $X2=1.285 $Y2=1.58
r57 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.285 $Y=1.665
+ $X2=1.285 $Y2=2.34
r58 3 25 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.485 $X2=2.305 $Y2=1.66
r59 3 18 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.485 $X2=2.305 $Y2=2.34
r60 2 21 400 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.485 $X2=1.285 $Y2=1.66
r61 2 12 400 $w=1.7e-07 $l=9.47497e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.485 $X2=1.285 $Y2=2.34
r62 1 41 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.63
+ $Y=0.235 $X2=2.765 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4BB_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r48 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r49 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r50 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r51 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 28 31 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r53 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r54 27 30 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r55 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r56 25 37 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.747
+ $Y2=0
r57 25 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.15
+ $Y2=0
r58 20 37 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.747
+ $Y2=0
r59 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r60 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r61 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r62 16 30 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.99
+ $Y2=0
r63 16 17 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.275
+ $Y2=0
r64 15 33 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r65 15 17 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.275
+ $Y2=0
r66 11 17 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=0.085
+ $X2=3.275 $Y2=0
r67 11 13 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.275 $Y=0.085
+ $X2=3.275 $Y2=0.38
r68 7 37 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0
r69 7 9 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0.38
r70 2 13 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.16
+ $Y=0.235 $X2=3.285 $Y2=0.38
r71 1 9 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.745 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__and3b_2.spice
* Created: Thu Aug 27 14:08:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and3b_2.pex.spice"
.subckt sky130_fd_sc_hd__and3b_2  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1005 N_A_109_53#_M1005_d N_A_N_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.1092 PD=1.4 PS=1.36 NRD=4.284 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_301_53# N_A_109_53#_M1002_g N_A_215_311#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1003 A_373_53# N_B_M1003_g A_301_53# VNB NSHORT L=0.15 W=0.42 AD=0.05355
+ AS=0.0441 PD=0.675 PS=0.63 NRD=20.712 NRS=14.28 M=1 R=2.8 SA=75000.5
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g A_373_53# VNB NSHORT L=0.15 W=0.42
+ AD=0.0998187 AS=0.05355 PD=0.859626 PS=0.675 NRD=47.136 NRS=20.712 M=1 R=2.8
+ SA=75000.9 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_215_311#_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.154481 PD=0.92 PS=1.33037 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1009_d N_A_215_311#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_109_53#_M1006_d N_A_N_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_109_53#_M1010_g N_A_215_311#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_215_311#_M1007_d N_B_M1007_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.074375 AS=0.0567 PD=0.815 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_C_M1008_g N_A_215_311#_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.074375 PD=0.789718 PS=0.815 NRD=70.4866 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1008_d N_A_215_311#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.205282 AS=0.135 PD=1.88028 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_215_311#_M1001_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__and3b_2.pxi.spice"
*
.ends
*
*

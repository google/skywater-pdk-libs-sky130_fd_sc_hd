* File: sky130_fd_sc_hd__and2b_4.spice.pex
* Created: Thu Aug 27 14:07:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND2B_4%A_33_199# 1 2 9 12 15 16 17 19 20 25 26 32
+ 35
r70 31 33 0.698946 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=3.44 $Y=1.695
+ $X2=3.44 $Y2=1.7
r71 31 32 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=1.695
+ $X2=3.44 $Y2=1.53
r72 26 36 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.355 $Y=1.16
+ $X2=0.355 $Y2=1.325
r73 26 35 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.355 $Y=1.16
+ $X2=0.355 $Y2=0.995
r74 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.16 $X2=0.34 $Y2=1.16
r75 22 25 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.25 $Y=1.16 $X2=0.34
+ $Y2=1.16
r76 20 29 10.7156 $w=1.91e-07 $l=1.76125e-07 $layer=LI1_cond $X=3.46 $Y=0.845
+ $X2=3.437 $Y2=0.68
r77 20 32 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.46 $Y=0.845
+ $X2=3.46 $Y2=1.53
r78 19 33 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.42 $Y=1.915
+ $X2=3.42 $Y2=1.7
r79 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=2
+ $X2=3.42 $Y2=1.915
r80 16 17 195.722 $w=1.68e-07 $l=3e-06 $layer=LI1_cond $X=3.335 $Y=2 $X2=0.335
+ $Y2=2
r81 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.25 $Y=1.915
+ $X2=0.335 $Y2=2
r82 14 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.25 $Y=1.325
+ $X2=0.25 $Y2=1.16
r83 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.25 $Y=1.325
+ $X2=0.25 $Y2=1.915
r84 12 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r85 9 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
r86 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.485 $X2=3.42 $Y2=1.695
r87 1 29 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.465 $X2=3.415 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_4%B 3 6 8 11 12 13
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r37 8 12 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.89 $Y2=1.16
r38 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r39 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r40 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.84 $Y=0.56 $X2=0.84
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_4%A_27_47# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 37 39 40 41 46 47 52 65
r114 64 65 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.28 $Y=1.16
+ $X2=2.7 $Y2=1.16
r115 63 64 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.27 $Y=1.16 $X2=2.28
+ $Y2=1.16
r116 60 61 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.84 $Y=1.16 $X2=1.86
+ $Y2=1.16
r117 53 63 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.175 $Y=1.16
+ $X2=2.27 $Y2=1.16
r118 53 61 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.175 $Y=1.16
+ $X2=1.86 $Y2=1.16
r119 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.175
+ $Y=1.16 $X2=2.175 $Y2=1.16
r120 50 60 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=1.495 $Y=1.16
+ $X2=1.84 $Y2=1.16
r121 50 57 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.495 $Y=1.16
+ $X2=1.41 $Y2=1.16
r122 49 52 21.7684 $w=3.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.495 $Y=1.175
+ $X2=2.175 $Y2=1.175
r123 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.495
+ $Y=1.16 $X2=1.495 $Y2=1.16
r124 47 49 4.48172 $w=3.58e-07 $l=1.4e-07 $layer=LI1_cond $X=1.355 $Y=1.175
+ $X2=1.495 $Y2=1.175
r125 46 47 10.4571 $w=2.1e-07 $l=1.88786e-07 $layer=LI1_cond $X=1.25 $Y=0.995
+ $X2=1.232 $Y2=1.175
r126 45 46 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=1.25 $Y=0.805
+ $X2=1.25 $Y2=0.995
r127 41 47 26.7324 $w=2.04e-07 $l=4.47e-07 $layer=LI1_cond $X=1.232 $Y=1.622
+ $X2=1.232 $Y2=1.175
r128 41 43 20.2266 $w=2.43e-07 $l=4.3e-07 $layer=LI1_cond $X=1.11 $Y=1.622
+ $X2=0.68 $Y2=1.622
r129 39 45 6.83868 $w=1.9e-07 $l=1.44914e-07 $layer=LI1_cond $X=1.145 $Y=0.71
+ $X2=1.25 $Y2=0.805
r130 39 40 42.0287 $w=1.88e-07 $l=7.2e-07 $layer=LI1_cond $X=1.145 $Y=0.71
+ $X2=0.425 $Y2=0.71
r131 35 40 7.51555 $w=1.9e-07 $l=2.102e-07 $layer=LI1_cond $X=0.257 $Y=0.615
+ $X2=0.425 $Y2=0.71
r132 35 37 8.0843 $w=3.33e-07 $l=2.35e-07 $layer=LI1_cond $X=0.257 $Y=0.615
+ $X2=0.257 $Y2=0.38
r133 31 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.16
r134 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.985
r135 28 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=1.16
r136 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=0.56
r137 24 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.325
+ $X2=2.28 $Y2=1.16
r138 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.28 $Y=1.325
+ $X2=2.28 $Y2=1.985
r139 21 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.27 $Y2=1.16
r140 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.27 $Y2=0.56
r141 17 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.325
+ $X2=1.86 $Y2=1.16
r142 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.86 $Y=1.325
+ $X2=1.86 $Y2=1.985
r143 14 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=0.995
+ $X2=1.84 $Y2=1.16
r144 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.84 $Y=0.995
+ $X2=1.84 $Y2=0.56
r145 10 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r146 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.985
r147 7 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r148 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r149 2 43 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r150 1 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_4%A_N 3 6 12 15 16 17
c35 17 0 1.4468e-19 $X=3.132 $Y=0.995
c36 16 0 1.19177e-19 $X=3.12 $Y=1.16
c37 6 0 3.45336e-19 $X=3.205 $Y=1.695
r38 15 18 51.062 $w=2.95e-07 $l=1.8e-07 $layer=POLY_cond $X=3.132 $Y=1.16
+ $X2=3.132 $Y2=1.34
r39 15 17 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=3.132 $Y=1.16
+ $X2=3.132 $Y2=0.995
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.16 $X2=3.12 $Y2=1.16
r41 12 16 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=3.052 $Y=1.19
+ $X2=3.052 $Y2=1.16
r42 6 18 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=3.205 $Y=1.695
+ $X2=3.205 $Y2=1.34
r43 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.205 $Y=0.675
+ $X2=3.205 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_4%VPWR 1 2 3 4 13 15 19 23 27 29 31 36 41 48
+ 49 55 58 61
r60 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r61 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 49 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r65 46 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=2.91 $Y2=2.72
r66 46 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 45 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r68 45 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r69 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 42 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r71 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 41 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.91 $Y2=2.72
r73 41 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.53 $Y2=2.72
r74 40 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r75 40 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 37 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=2.72
+ $X2=1.155 $Y2=2.72
r78 37 39 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.32 $Y=2.72
+ $X2=1.61 $Y2=2.72
r79 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 36 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.905 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 35 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r82 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 32 52 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r84 32 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r85 31 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=2.72
+ $X2=1.155 $Y2=2.72
r86 31 34 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=0.69
+ $Y2=2.72
r87 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 29 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 25 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=2.635
+ $X2=2.91 $Y2=2.72
r90 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.91 $Y=2.635
+ $X2=2.91 $Y2=2.36
r91 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.635
+ $X2=2.07 $Y2=2.72
r92 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.07 $Y=2.635
+ $X2=2.07 $Y2=2.36
r93 17 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.635
+ $X2=1.155 $Y2=2.72
r94 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.155 $Y=2.635
+ $X2=1.155 $Y2=2.36
r95 13 52 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r96 13 15 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r97 4 27 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.485 $X2=2.91 $Y2=2.36
r98 3 23 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.485 $X2=2.07 $Y2=2.36
r99 2 19 600 $w=1.7e-07 $l=9.65337e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.155 $Y2=2.36
r100 1 15 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_4%X 1 2 3 4 13 18 23 26 30 32
c43 32 0 3.11092e-19 $X=2.525 $Y=0.85
c44 23 0 1.78923e-19 $X=2.585 $Y=1.535
r45 30 32 0.993485 $w=2.88e-07 $l=2.5e-08 $layer=LI1_cond $X=2.585 $Y=0.825
+ $X2=2.585 $Y2=0.85
r46 26 30 2.95929 $w=2.9e-07 $l=1.05e-07 $layer=LI1_cond $X=2.585 $Y=0.72
+ $X2=2.585 $Y2=0.825
r47 26 32 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=2.585 $Y=0.88
+ $X2=2.585 $Y2=0.85
r48 23 26 26.0293 $w=2.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.585 $Y=1.535
+ $X2=2.585 $Y2=0.88
r49 23 25 2.95929 $w=2.9e-07 $l=1.05e-07 $layer=LI1_cond $X=2.585 $Y=1.535
+ $X2=2.585 $Y2=1.64
r50 21 26 31.5451 $w=2.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.715 $Y=0.72
+ $X2=2.44 $Y2=0.72
r51 20 21 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=1.62 $Y=0.72
+ $X2=1.715 $Y2=0.72
r52 18 20 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=1.62 $Y=0.66 $X2=1.62
+ $Y2=0.72
r53 13 25 4.08664 $w=2.1e-07 $l=1.45e-07 $layer=LI1_cond $X=2.44 $Y=1.64
+ $X2=2.585 $Y2=1.64
r54 13 15 41.7229 $w=2.08e-07 $l=7.9e-07 $layer=LI1_cond $X=2.44 $Y=1.64
+ $X2=1.65 $Y2=1.64
r55 4 25 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.355
+ $Y=1.485 $X2=2.49 $Y2=1.62
r56 3 15 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.65 $Y2=1.62
r57 2 26 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.235 $X2=2.485 $Y2=0.74
r58 1 18 182 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_4%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r62 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r63 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r64 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r65 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r66 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r67 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=0 $X2=2.91
+ $Y2=0
r68 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.075 $Y=0 $X2=3.45
+ $Y2=0
r69 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r70 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r71 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r72 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.05
+ $Y2=0
r73 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.53
+ $Y2=0
r74 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.91
+ $Y2=0
r75 34 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.53
+ $Y2=0
r76 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r77 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r78 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r79 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r80 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.61
+ $Y2=0
r81 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.05
+ $Y2=0
r82 29 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=1.61
+ $Y2=0
r83 27 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r84 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r85 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r86 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.69
+ $Y2=0
r87 22 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r88 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0
r89 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0.36
r90 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0
r91 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0.36
r92 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r93 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r94 3 20 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.235 $X2=2.91 $Y2=0.36
r95 2 16 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.235 $X2=2.05 $Y2=0.36
r96 1 12 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.915
+ $Y=0.235 $X2=1.12 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__dlrbp_1.spice.SKY130_FD_SC_HD__DLRBP_1.pxi
* Created: Thu Aug 27 14:16:53 2020
* 
x_PM_SKY130_FD_SC_HD__DLRBP_1%GATE N_GATE_c_155_n N_GATE_c_150_n N_GATE_M1021_g
+ N_GATE_c_156_n N_GATE_M1007_g N_GATE_c_151_n N_GATE_c_157_n GATE GATE
+ N_GATE_c_153_n N_GATE_c_154_n PM_SKY130_FD_SC_HD__DLRBP_1%GATE
x_PM_SKY130_FD_SC_HD__DLRBP_1%A_27_47# N_A_27_47#_M1021_s N_A_27_47#_M1007_s
+ N_A_27_47#_M1010_g N_A_27_47#_M1000_g N_A_27_47#_M1001_g N_A_27_47#_c_194_n
+ N_A_27_47#_c_195_n N_A_27_47#_M1011_g N_A_27_47#_c_207_n N_A_27_47#_c_197_n
+ N_A_27_47#_c_198_n N_A_27_47#_c_199_n N_A_27_47#_c_208_n N_A_27_47#_c_209_n
+ N_A_27_47#_c_200_n N_A_27_47#_c_201_n N_A_27_47#_c_211_n N_A_27_47#_c_212_n
+ N_A_27_47#_c_213_n N_A_27_47#_c_214_n N_A_27_47#_c_215_n N_A_27_47#_c_216_n
+ N_A_27_47#_c_202_n PM_SKY130_FD_SC_HD__DLRBP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRBP_1%D N_D_M1003_g N_D_M1017_g D N_D_c_341_n
+ N_D_c_342_n PM_SKY130_FD_SC_HD__DLRBP_1%D
x_PM_SKY130_FD_SC_HD__DLRBP_1%A_299_47# N_A_299_47#_M1003_s N_A_299_47#_M1017_s
+ N_A_299_47#_M1006_g N_A_299_47#_M1012_g N_A_299_47#_c_387_n
+ N_A_299_47#_c_380_n N_A_299_47#_c_388_n N_A_299_47#_c_389_n
+ N_A_299_47#_c_381_n N_A_299_47#_c_382_n N_A_299_47#_c_383_n
+ N_A_299_47#_c_384_n N_A_299_47#_c_385_n PM_SKY130_FD_SC_HD__DLRBP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__DLRBP_1%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_c_463_n N_A_193_47#_M1018_g N_A_193_47#_M1022_g
+ N_A_193_47#_c_464_n N_A_193_47#_c_465_n N_A_193_47#_c_466_n
+ N_A_193_47#_c_470_n N_A_193_47#_c_471_n N_A_193_47#_c_472_n
+ N_A_193_47#_c_473_n N_A_193_47#_c_474_n N_A_193_47#_c_475_n
+ N_A_193_47#_c_476_n PM_SKY130_FD_SC_HD__DLRBP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRBP_1%A_711_307# N_A_711_307#_M1015_s
+ N_A_711_307#_M1013_d N_A_711_307#_M1009_g N_A_711_307#_M1023_g
+ N_A_711_307#_c_581_n N_A_711_307#_M1008_g N_A_711_307#_M1004_g
+ N_A_711_307#_c_582_n N_A_711_307#_c_583_n N_A_711_307#_M1002_g
+ N_A_711_307#_M1016_g N_A_711_307#_c_585_n N_A_711_307#_c_596_n
+ N_A_711_307#_c_597_n N_A_711_307#_c_586_n N_A_711_307#_c_607_p
+ N_A_711_307#_c_587_n N_A_711_307#_c_606_p N_A_711_307#_c_622_p
+ N_A_711_307#_c_588_n N_A_711_307#_c_630_p
+ PM_SKY130_FD_SC_HD__DLRBP_1%A_711_307#
x_PM_SKY130_FD_SC_HD__DLRBP_1%A_560_47# N_A_560_47#_M1018_d N_A_560_47#_M1001_d
+ N_A_560_47#_M1013_g N_A_560_47#_c_694_n N_A_560_47#_M1015_g
+ N_A_560_47#_c_695_n N_A_560_47#_c_696_n N_A_560_47#_c_705_n
+ N_A_560_47#_c_706_n N_A_560_47#_c_697_n N_A_560_47#_c_703_n
+ N_A_560_47#_c_698_n N_A_560_47#_c_699_n PM_SKY130_FD_SC_HD__DLRBP_1%A_560_47#
x_PM_SKY130_FD_SC_HD__DLRBP_1%RESET_B N_RESET_B_M1020_g N_RESET_B_M1005_g
+ RESET_B RESET_B N_RESET_B_c_775_n N_RESET_B_c_776_n RESET_B
+ PM_SKY130_FD_SC_HD__DLRBP_1%RESET_B
x_PM_SKY130_FD_SC_HD__DLRBP_1%A_1308_47# N_A_1308_47#_M1002_s
+ N_A_1308_47#_M1016_s N_A_1308_47#_M1019_g N_A_1308_47#_M1014_g
+ N_A_1308_47#_c_810_n N_A_1308_47#_c_815_n N_A_1308_47#_c_811_n
+ N_A_1308_47#_c_812_n N_A_1308_47#_c_823_n N_A_1308_47#_c_813_n
+ PM_SKY130_FD_SC_HD__DLRBP_1%A_1308_47#
x_PM_SKY130_FD_SC_HD__DLRBP_1%VPWR N_VPWR_M1007_d N_VPWR_M1017_d N_VPWR_M1009_d
+ N_VPWR_M1013_s N_VPWR_M1005_d N_VPWR_M1016_d N_VPWR_c_851_n N_VPWR_c_852_n
+ N_VPWR_c_853_n VPWR N_VPWR_c_854_n N_VPWR_c_855_n N_VPWR_c_856_n
+ N_VPWR_c_857_n N_VPWR_c_858_n N_VPWR_c_850_n N_VPWR_c_860_n N_VPWR_c_861_n
+ N_VPWR_c_862_n N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_865_n
+ PM_SKY130_FD_SC_HD__DLRBP_1%VPWR
x_PM_SKY130_FD_SC_HD__DLRBP_1%Q N_Q_M1008_d N_Q_M1004_d Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HD__DLRBP_1%Q
x_PM_SKY130_FD_SC_HD__DLRBP_1%Q_N N_Q_N_M1019_d N_Q_N_M1014_d Q_N Q_N Q_N
+ N_Q_N_c_982_n Q_N PM_SKY130_FD_SC_HD__DLRBP_1%Q_N
x_PM_SKY130_FD_SC_HD__DLRBP_1%VGND N_VGND_M1021_d N_VGND_M1003_d N_VGND_M1023_d
+ N_VGND_M1020_d N_VGND_M1002_d N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n
+ N_VGND_c_997_n VGND N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n
+ N_VGND_c_1001_n N_VGND_c_1002_n N_VGND_c_1003_n N_VGND_c_1004_n
+ N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n N_VGND_c_1008_n
+ N_VGND_c_1009_n PM_SKY130_FD_SC_HD__DLRBP_1%VGND
cc_1 VNB N_GATE_c_150_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_c_151_n 0.023495f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE 0.0127963f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_GATE_c_153_n 0.0210526f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_GATE_c_154_n 0.0148348f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1010_g 0.0398194f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_194_n 0.0131032f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_27_47#_c_195_n 0.00481214f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_9 VNB N_A_27_47#_M1011_g 0.0469778f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_10 VNB N_A_27_47#_c_197_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_198_n 0.00225297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_199_n 0.00790266f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_200_n 7.88168e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_201_n 0.00420082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_202_n 0.0231108f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1003_g 0.0258946f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_17 VNB N_D_M1017_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_341_n 0.00407935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_19 VNB N_D_c_342_n 0.0421617f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_20 VNB N_A_299_47#_M1012_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_299_47#_c_380_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_381_n 0.00503217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_47#_c_382_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_24 VNB N_A_299_47#_c_383_n 0.00265154f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_25 VNB N_A_299_47#_c_384_n 0.0267054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_299_47#_c_385_n 0.0166855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_463_n 0.0471774f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_28 VNB N_A_193_47#_c_464_n 0.0140955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_c_465_n 0.00526473f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_193_47#_c_466_n 0.00419558f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_31 VNB N_A_711_307#_M1023_g 0.050595f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_32 VNB N_A_711_307#_c_581_n 0.0211172f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_33 VNB N_A_711_307#_c_582_n 0.047203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_711_307#_c_583_n 0.0255903f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_35 VNB N_A_711_307#_M1002_g 0.0357177f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_36 VNB N_A_711_307#_c_585_n 0.00829564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_711_307#_c_586_n 0.00482174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_711_307#_c_587_n 0.00345373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_711_307#_c_588_n 0.00147514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_560_47#_c_694_n 0.0224584f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_41 VNB N_A_560_47#_c_695_n 0.0402072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_560_47#_c_696_n 0.00895781f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_43 VNB N_A_560_47#_c_697_n 0.00752442f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_44 VNB N_A_560_47#_c_698_n 0.00338161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_560_47#_c_699_n 0.0110123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB RESET_B 0.00718508f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_47 VNB N_RESET_B_c_775_n 0.020948f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_48 VNB N_RESET_B_c_776_n 0.0192541f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_49 VNB N_A_1308_47#_c_810_n 0.00275283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1308_47#_c_811_n 0.00397886f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_51 VNB N_A_1308_47#_c_812_n 0.0260627f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_52 VNB N_A_1308_47#_c_813_n 0.0197073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VPWR_c_850_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB Q 0.0095977f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_55 VNB Q_N 0.0303491f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_56 VNB N_Q_N_c_982_n 0.0133709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_994_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_995_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_996_n 0.00603643f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_60 VNB N_VGND_c_997_n 0.00276055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_998_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_999_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1000_n 0.0410013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1001_n 0.0279074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1002_n 0.0150402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1003_n 0.39647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1004_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1005_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1006_n 0.00517156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1007_n 0.0270084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1008_n 0.0147422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1009_n 0.00506835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VPB N_GATE_c_155_n 0.0129163f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_74 VPB N_GATE_c_156_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_75 VPB N_GATE_c_157_n 0.02422f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_76 VPB GATE 0.0127706f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_77 VPB N_GATE_c_153_n 0.0106946f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_78 VPB N_A_27_47#_M1000_g 0.039528f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_79 VPB N_A_27_47#_M1001_g 0.0300673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_80 VPB N_A_27_47#_c_194_n 0.0172883f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_81 VPB N_A_27_47#_c_195_n 0.00790086f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_82 VPB N_A_27_47#_c_207_n 0.0121288f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_83 VPB N_A_27_47#_c_208_n 0.00126297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_209_n 0.0300458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_200_n 6.03631e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_211_n 0.0224566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_47#_c_212_n 0.00377566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_47#_c_213_n 0.00547825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_27_47#_c_214_n 0.00344459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_27_47#_c_215_n 0.00529835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_27_47#_c_216_n 0.00947367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_27_47#_c_202_n 0.0116052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_D_M1017_g 0.0462501f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_94 VPB N_D_c_341_n 0.00235013f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_95 VPB N_A_299_47#_M1012_g 0.0366983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_299_47#_c_387_n 0.00712099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_299_47#_c_388_n 0.00409088f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_98 VPB N_A_299_47#_c_389_n 0.00290124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_299_47#_c_382_n 0.00355393f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_100 VPB N_A_193_47#_M1022_g 0.0205785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_193_47#_c_464_n 0.00804665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_193_47#_c_466_n 0.00254097f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_103 VPB N_A_193_47#_c_470_n 0.00293933f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_104 VPB N_A_193_47#_c_471_n 0.00861819f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_105 VPB N_A_193_47#_c_472_n 0.00238602f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.19
cc_106 VPB N_A_193_47#_c_473_n 0.00711634f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.53
cc_107 VPB N_A_193_47#_c_474_n 0.00247667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_193_47#_c_475_n 0.0268882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_193_47#_c_476_n 0.00796076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_711_307#_M1009_g 0.0291104f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_111 VPB N_A_711_307#_M1023_g 0.0183372f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_112 VPB N_A_711_307#_M1004_g 0.0241438f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_113 VPB N_A_711_307#_c_582_n 0.0229504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_711_307#_c_583_n 0.00708238f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_115 VPB N_A_711_307#_M1016_g 0.0474763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_711_307#_c_585_n 5.25028e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_711_307#_c_596_n 0.00457073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_711_307#_c_597_n 0.047134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_711_307#_c_588_n 0.00214566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_560_47#_M1013_g 0.0257812f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_121 VPB N_A_560_47#_c_695_n 0.0145744f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_560_47#_c_696_n 9.45393e-19 $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_123 VPB N_A_560_47#_c_703_n 0.00880117f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_124 VPB N_A_560_47#_c_698_n 0.00182699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_RESET_B_M1005_g 0.0227316f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_126 VPB RESET_B 0.00478222f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_127 VPB N_RESET_B_c_775_n 0.00410784f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_128 VPB N_A_1308_47#_M1014_g 0.0226364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_1308_47#_c_815_n 0.00435864f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_130 VPB N_A_1308_47#_c_811_n 0.00470632f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_131 VPB N_A_1308_47#_c_812_n 0.00693673f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_132 VPB N_VPWR_c_851_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_852_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_134 VPB N_VPWR_c_853_n 0.00289402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_854_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_855_n 0.0295132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_856_n 0.013238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_857_n 0.0288197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_858_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_850_n 0.0597909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_860_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_861_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_862_n 0.0387638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_863_n 0.0273201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_864_n 0.0146748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_865_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB Q 0.0146865f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_148 VPB Q_N 0.0458373f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_149 N_GATE_c_150_n N_A_27_47#_M1010_g 0.0187874f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_150 N_GATE_c_154_n N_A_27_47#_M1010_g 0.00412893f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_151 N_GATE_c_157_n N_A_27_47#_M1000_g 0.0260433f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_152 N_GATE_c_153_n N_A_27_47#_M1000_g 0.00519338f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_153 N_GATE_c_150_n N_A_27_47#_c_198_n 0.00674622f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_154 N_GATE_c_151_n N_A_27_47#_c_198_n 0.0104954f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_155 N_GATE_c_151_n N_A_27_47#_c_199_n 0.00711144f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_156 GATE N_A_27_47#_c_199_n 0.0198215f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_157 N_GATE_c_153_n N_A_27_47#_c_199_n 7.3212e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_158 N_GATE_c_156_n N_A_27_47#_c_208_n 0.0135762f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_159 N_GATE_c_157_n N_A_27_47#_c_208_n 0.00216816f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_160 N_GATE_c_156_n N_A_27_47#_c_209_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_161 N_GATE_c_157_n N_A_27_47#_c_209_n 0.00423203f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_162 GATE N_A_27_47#_c_209_n 0.0217264f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_163 N_GATE_c_153_n N_A_27_47#_c_209_n 5.66731e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_164 N_GATE_c_153_n N_A_27_47#_c_200_n 0.00319971f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_165 N_GATE_c_151_n N_A_27_47#_c_201_n 0.00179459f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_166 GATE N_A_27_47#_c_201_n 0.0283946f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_167 N_GATE_c_154_n N_A_27_47#_c_201_n 0.00151497f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_168 N_GATE_c_155_n N_A_27_47#_c_212_n 0.00338266f $X=0.3 $Y=1.59 $X2=0 $Y2=0
cc_169 N_GATE_c_157_n N_A_27_47#_c_212_n 0.00102651f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_170 GATE N_A_27_47#_c_212_n 0.00651178f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_171 N_GATE_c_155_n N_A_27_47#_c_213_n 7.61436e-19 $X=0.3 $Y=1.59 $X2=0 $Y2=0
cc_172 N_GATE_c_157_n N_A_27_47#_c_213_n 0.00428034f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_173 GATE N_A_27_47#_c_202_n 9.15599e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_174 N_GATE_c_153_n N_A_27_47#_c_202_n 0.0161155f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_175 N_GATE_c_156_n N_VPWR_c_851_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_176 N_GATE_c_156_n N_VPWR_c_854_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_177 N_GATE_c_156_n N_VPWR_c_850_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_178 N_GATE_c_150_n N_VGND_c_994_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_179 N_GATE_c_150_n N_VGND_c_998_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_180 N_GATE_c_151_n N_VGND_c_998_n 4.87495e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_181 N_GATE_c_150_n N_VGND_c_1003_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_211_n N_D_M1017_g 0.00583826f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_211_n N_D_c_341_n 0.0087134f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1010_g N_D_c_342_n 0.00520956f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1001_g N_A_299_47#_M1012_g 0.0353942f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_195_n N_A_299_47#_M1012_g 0.0248407f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_211_n N_A_299_47#_M1012_g 0.00493352f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_214_n N_A_299_47#_M1012_g 0.00140912f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_215_n N_A_299_47#_M1012_g 0.00239179f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_211_n N_A_299_47#_c_388_n 0.0116439f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_214_n N_A_299_47#_c_388_n 0.00130924f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_215_n N_A_299_47#_c_388_n 0.00675603f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_211_n N_A_299_47#_c_389_n 0.0115067f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_211_n N_A_299_47#_c_381_n 0.00675641f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_211_n N_A_299_47#_c_382_n 0.0108494f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_214_n N_A_299_47#_c_382_n 0.00124596f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_215_n N_A_299_47#_c_382_n 0.00570493f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_211_n N_A_299_47#_c_384_n 0.00107604f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_195_n N_A_193_47#_c_463_n 0.0207633f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_M1011_g N_A_193_47#_c_463_n 0.0365214f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_215_n N_A_193_47#_c_463_n 5.58399e-19 $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_M1001_g N_A_193_47#_M1022_g 0.019647f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_M1010_g N_A_193_47#_c_464_n 0.00779983f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_198_n N_A_193_47#_c_464_n 0.0100297f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_200_n N_A_193_47#_c_464_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_201_n N_A_193_47#_c_464_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_211_n N_A_193_47#_c_464_n 0.0184539f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_212_n N_A_193_47#_c_464_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_213_n N_A_193_47#_c_464_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_195_n N_A_193_47#_c_465_n 0.00183728f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_M1011_g N_A_193_47#_c_465_n 0.00221014f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_212 N_A_27_47#_c_214_n N_A_193_47#_c_465_n 5.91364e-19 $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_215_n N_A_193_47#_c_465_n 0.00623896f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_194_n N_A_193_47#_c_466_n 0.0133727f $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_M1011_g N_A_193_47#_c_466_n 0.0049549f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_214_n N_A_193_47#_c_466_n 0.00101104f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_215_n N_A_193_47#_c_466_n 0.0151027f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_216_n N_A_193_47#_c_466_n 0.00406305f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_208_n N_A_193_47#_c_470_n 0.00294892f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_211_n N_A_193_47#_c_470_n 0.00195186f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_202_n N_A_193_47#_c_470_n 0.00779983f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_M1001_g N_A_193_47#_c_471_n 0.00736818f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_194_n N_A_193_47#_c_471_n 0.00108869f $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_207_n N_A_193_47#_c_471_n 0.00185018f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_211_n N_A_193_47#_c_471_n 0.0871075f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_214_n N_A_193_47#_c_471_n 0.0266068f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_215_n N_A_193_47#_c_471_n 0.00864674f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1000_g N_A_193_47#_c_472_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_208_n N_A_193_47#_c_472_n 0.00551586f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_211_n N_A_193_47#_c_472_n 0.0259095f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_213_n N_A_193_47#_c_472_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1000_g N_A_193_47#_c_473_n 0.00779983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_M1001_g N_A_193_47#_c_474_n 0.00145643f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_194_n N_A_193_47#_c_474_n 0.00123942f $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_194_n N_A_193_47#_c_475_n 0.0180829f $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_207_n N_A_193_47#_c_475_n 0.0166555f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_194_n N_A_193_47#_c_476_n 0.00400792f $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_207_n N_A_193_47#_c_476_n 0.00597161f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_214_n N_A_193_47#_c_476_n 4.76211e-19 $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_215_n N_A_193_47#_c_476_n 0.00815409f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_M1011_g N_A_711_307#_M1023_g 0.0425818f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_242 N_A_27_47#_M1001_g N_A_560_47#_c_705_n 0.0049672f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_M1011_g N_A_560_47#_c_706_n 0.0149072f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1011_g N_A_560_47#_c_697_n 0.00652775f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_245 N_A_27_47#_c_194_n N_A_560_47#_c_703_n 6.91978e-19 $X=3.14 $Y=1.32 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_M1011_g N_A_560_47#_c_699_n 0.00346936f $X=3.215 $Y=0.415
+ $X2=0 $Y2=0
cc_247 N_A_27_47#_c_208_n N_VPWR_M1007_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_248 N_A_27_47#_M1000_g N_VPWR_c_851_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_208_n N_VPWR_c_851_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_209_n N_VPWR_c_851_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_212_n N_VPWR_c_851_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_252 N_A_27_47#_M1001_g N_VPWR_c_852_n 0.00401328f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_211_n N_VPWR_c_852_n 0.0019389f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_208_n N_VPWR_c_854_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_209_n N_VPWR_c_854_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_256 N_A_27_47#_M1000_g N_VPWR_c_855_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1000_g N_VPWR_c_850_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1001_g N_VPWR_c_850_n 0.00611433f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_208_n N_VPWR_c_850_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_209_n N_VPWR_c_850_n 0.00993215f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_261 N_A_27_47#_M1001_g N_VPWR_c_862_n 0.00497675f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_198_n N_VGND_M1021_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_263 N_A_27_47#_M1010_g N_VGND_c_994_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_198_n N_VGND_c_994_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_200_n N_VGND_c_994_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_202_n N_VGND_c_994_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_M1011_g N_VGND_c_996_n 0.00172953f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_197_n N_VGND_c_998_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_198_n N_VGND_c_998_n 0.00243651f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_270 N_A_27_47#_M1010_g N_VGND_c_999_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_271 N_A_27_47#_M1011_g N_VGND_c_1000_n 0.0037981f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1021_s N_VGND_c_1003_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1010_g N_VGND_c_1003_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1011_g N_VGND_c_1003_n 0.00570274f $X=3.215 $Y=0.415 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_197_n N_VGND_c_1003_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_198_n N_VGND_c_1003_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_277 N_D_c_342_n N_A_299_47#_M1012_g 0.03863f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_278 N_D_M1017_g N_A_299_47#_c_387_n 0.012851f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_279 N_D_M1003_g N_A_299_47#_c_380_n 0.0144406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_280 N_D_c_341_n N_A_299_47#_c_380_n 0.00627239f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_281 N_D_c_342_n N_A_299_47#_c_380_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_282 N_D_M1017_g N_A_299_47#_c_388_n 0.00794545f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_283 N_D_M1017_g N_A_299_47#_c_389_n 0.00412429f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_284 N_D_c_341_n N_A_299_47#_c_389_n 0.0229667f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_285 N_D_c_342_n N_A_299_47#_c_389_n 0.00131849f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_286 N_D_M1003_g N_A_299_47#_c_381_n 0.00563568f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_287 N_D_c_341_n N_A_299_47#_c_381_n 0.0107593f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_288 N_D_c_341_n N_A_299_47#_c_382_n 0.0164827f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_289 N_D_c_342_n N_A_299_47#_c_382_n 0.00552652f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_290 N_D_M1003_g N_A_299_47#_c_383_n 0.00120855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_291 N_D_c_341_n N_A_299_47#_c_383_n 0.0138491f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_292 N_D_c_342_n N_A_299_47#_c_383_n 0.0042466f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_293 N_D_M1003_g N_A_299_47#_c_384_n 0.0197189f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_294 N_D_M1003_g N_A_299_47#_c_385_n 0.015283f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_295 N_D_M1003_g N_A_193_47#_c_464_n 0.00203374f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_296 N_D_M1017_g N_A_193_47#_c_464_n 0.00459933f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_297 N_D_c_341_n N_A_193_47#_c_464_n 0.0209974f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_298 N_D_c_342_n N_A_193_47#_c_464_n 0.00256393f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_299 N_D_M1017_g N_A_193_47#_c_470_n 0.00134564f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_300 N_D_M1017_g N_A_193_47#_c_471_n 0.00294239f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_301 N_D_M1017_g N_VPWR_c_852_n 0.00304701f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_302 N_D_M1017_g N_VPWR_c_855_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_303 N_D_M1017_g N_VPWR_c_850_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_304 N_D_M1003_g N_VGND_c_995_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_305 N_D_M1003_g N_VGND_c_999_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_306 N_D_M1003_g N_VGND_c_1003_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_307 N_D_c_342_n N_VGND_c_1003_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_308 N_A_299_47#_c_381_n N_A_193_47#_c_463_n 3.13306e-19 $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_309 N_A_299_47#_c_384_n N_A_193_47#_c_463_n 0.0167604f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_310 N_A_299_47#_c_385_n N_A_193_47#_c_463_n 0.0264449f $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_311 N_A_299_47#_c_387_n N_A_193_47#_c_464_n 0.0010921f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_312 N_A_299_47#_c_389_n N_A_193_47#_c_464_n 0.00859001f $X=1.785 $Y=1.58
+ $X2=0 $Y2=0
cc_313 N_A_299_47#_c_383_n N_A_193_47#_c_464_n 0.0191833f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_314 N_A_299_47#_c_381_n N_A_193_47#_c_465_n 0.0150553f $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_315 N_A_299_47#_c_384_n N_A_193_47#_c_465_n 9.34289e-19 $X=2.255 $Y=0.93
+ $X2=0 $Y2=0
cc_316 N_A_299_47#_M1012_g N_A_193_47#_c_466_n 0.00370009f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_317 N_A_299_47#_c_381_n N_A_193_47#_c_466_n 0.00176972f $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_318 N_A_299_47#_c_384_n N_A_193_47#_c_466_n 9.9292e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_319 N_A_299_47#_c_387_n N_A_193_47#_c_470_n 0.0471072f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_320 N_A_299_47#_M1012_g N_A_193_47#_c_471_n 0.00365242f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_321 N_A_299_47#_c_387_n N_A_193_47#_c_471_n 0.022748f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_322 N_A_299_47#_c_388_n N_A_193_47#_c_471_n 0.00551435f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_323 N_A_299_47#_c_387_n N_A_193_47#_c_472_n 0.00273055f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_324 N_A_299_47#_M1012_g N_A_560_47#_c_705_n 5.24267e-19 $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_325 N_A_299_47#_c_385_n N_A_560_47#_c_706_n 6.66135e-19 $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_326 N_A_299_47#_M1012_g N_VPWR_c_852_n 0.0234054f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_327 N_A_299_47#_c_387_n N_VPWR_c_852_n 0.0232987f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_328 N_A_299_47#_c_388_n N_VPWR_c_852_n 0.013562f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_329 N_A_299_47#_c_387_n N_VPWR_c_855_n 0.0159418f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_330 N_A_299_47#_M1017_s N_VPWR_c_850_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_331 N_A_299_47#_M1012_g N_VPWR_c_850_n 0.00262666f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_332 N_A_299_47#_c_387_n N_VPWR_c_850_n 0.00576627f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_333 N_A_299_47#_M1012_g N_VPWR_c_862_n 0.00212864f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_334 N_A_299_47#_c_381_n N_VGND_M1003_d 0.00156939f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_380_n N_VGND_c_995_n 0.00259081f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_336 N_A_299_47#_c_381_n N_VGND_c_995_n 0.0141976f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_337 N_A_299_47#_c_385_n N_VGND_c_995_n 0.00941159f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_380_n N_VGND_c_999_n 0.00255672f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_339 N_A_299_47#_c_383_n N_VGND_c_999_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_340 N_A_299_47#_c_384_n N_VGND_c_1000_n 9.84895e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_341 N_A_299_47#_c_385_n N_VGND_c_1000_n 0.0046653f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_342 N_A_299_47#_M1003_s N_VGND_c_1003_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_343 N_A_299_47#_c_380_n N_VGND_c_1003_n 0.00473142f $X=1.97 $Y=0.7 $X2=0
+ $Y2=0
cc_344 N_A_299_47#_c_381_n N_VGND_c_1003_n 0.00552372f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_345 N_A_299_47#_c_383_n N_VGND_c_1003_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_c_384_n N_VGND_c_1003_n 0.00117722f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_347 N_A_299_47#_c_385_n N_VGND_c_1003_n 0.00440683f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_348 N_A_193_47#_M1022_g N_A_711_307#_M1009_g 0.0263455f $X=3.15 $Y=2.275
+ $X2=0 $Y2=0
cc_349 N_A_193_47#_c_476_n N_A_711_307#_M1009_g 2.15098e-19 $X=3.18 $Y=1.74
+ $X2=0 $Y2=0
cc_350 N_A_193_47#_c_475_n N_A_711_307#_c_597_n 0.0167148f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_351 N_A_193_47#_c_476_n N_A_711_307#_c_597_n 3.98623e-19 $X=3.18 $Y=1.74
+ $X2=0 $Y2=0
cc_352 N_A_193_47#_M1022_g N_A_560_47#_c_705_n 0.00894354f $X=3.15 $Y=2.275
+ $X2=0 $Y2=0
cc_353 N_A_193_47#_c_471_n N_A_560_47#_c_705_n 0.00268701f $X=2.865 $Y=1.87
+ $X2=0 $Y2=0
cc_354 N_A_193_47#_c_474_n N_A_560_47#_c_705_n 0.00279139f $X=3.01 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_193_47#_c_476_n N_A_560_47#_c_705_n 0.0121101f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_356 N_A_193_47#_c_463_n N_A_560_47#_c_706_n 0.00702246f $X=2.725 $Y=0.705
+ $X2=0 $Y2=0
cc_357 N_A_193_47#_c_465_n N_A_560_47#_c_706_n 0.0167325f $X=2.925 $Y=0.9 $X2=0
+ $Y2=0
cc_358 N_A_193_47#_c_465_n N_A_560_47#_c_697_n 0.0150278f $X=2.925 $Y=0.9 $X2=0
+ $Y2=0
cc_359 N_A_193_47#_M1022_g N_A_560_47#_c_703_n 0.00376601f $X=3.15 $Y=2.275
+ $X2=0 $Y2=0
cc_360 N_A_193_47#_c_466_n N_A_560_47#_c_703_n 0.0113318f $X=3.01 $Y=1.575 $X2=0
+ $Y2=0
cc_361 N_A_193_47#_c_474_n N_A_560_47#_c_703_n 0.00283423f $X=3.01 $Y=1.87 $X2=0
+ $Y2=0
cc_362 N_A_193_47#_c_475_n N_A_560_47#_c_703_n 0.00425391f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_363 N_A_193_47#_c_476_n N_A_560_47#_c_703_n 0.0275893f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_364 N_A_193_47#_c_465_n N_A_560_47#_c_699_n 0.00291029f $X=2.925 $Y=0.9 $X2=0
+ $Y2=0
cc_365 N_A_193_47#_c_466_n N_A_560_47#_c_699_n 0.0167234f $X=3.01 $Y=1.575 $X2=0
+ $Y2=0
cc_366 N_A_193_47#_c_475_n N_A_560_47#_c_699_n 4.91178e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_367 N_A_193_47#_c_471_n N_VPWR_M1017_d 6.81311e-19 $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_368 N_A_193_47#_c_473_n N_VPWR_c_851_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_193_47#_c_471_n N_VPWR_c_852_n 0.0184713f $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_474_n N_VPWR_c_852_n 9.65502e-19 $X=3.01 $Y=1.87 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_c_476_n N_VPWR_c_852_n 0.00216873f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_372 N_A_193_47#_c_473_n N_VPWR_c_855_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_373 N_A_193_47#_M1022_g N_VPWR_c_850_n 0.00538581f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_471_n N_VPWR_c_850_n 0.0747938f $X=2.865 $Y=1.87 $X2=0
+ $Y2=0
cc_375 N_A_193_47#_c_472_n N_VPWR_c_850_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_376 N_A_193_47#_c_473_n N_VPWR_c_850_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_c_474_n N_VPWR_c_850_n 0.0148714f $X=3.01 $Y=1.87 $X2=0 $Y2=0
cc_378 N_A_193_47#_M1022_g N_VPWR_c_862_n 0.00366111f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_471_n A_465_369# 0.00388705f $X=2.865 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_380 N_A_193_47#_c_463_n N_VGND_c_995_n 0.0018389f $X=2.725 $Y=0.705 $X2=0
+ $Y2=0
cc_381 N_A_193_47#_c_464_n N_VGND_c_999_n 0.00732874f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_382 N_A_193_47#_c_463_n N_VGND_c_1000_n 0.00629197f $X=2.725 $Y=0.705 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_M1010_d N_VGND_c_1003_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_384 N_A_193_47#_c_463_n N_VGND_c_1003_n 0.00753081f $X=2.725 $Y=0.705 $X2=0
+ $Y2=0
cc_385 N_A_193_47#_c_464_n N_VGND_c_1003_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_386 N_A_193_47#_c_465_n N_VGND_c_1003_n 0.00570891f $X=2.925 $Y=0.9 $X2=0
+ $Y2=0
cc_387 N_A_711_307#_c_596_n N_A_560_47#_M1013_g 0.0164134f $X=4.78 $Y=1.7 $X2=0
+ $Y2=0
cc_388 N_A_711_307#_c_597_n N_A_560_47#_M1013_g 0.00687993f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_389 N_A_711_307#_c_606_p N_A_560_47#_M1013_g 0.00649326f $X=4.865 $Y=2.27
+ $X2=0 $Y2=0
cc_390 N_A_711_307#_c_607_p N_A_560_47#_c_694_n 0.0113641f $X=5.655 $Y=0.74
+ $X2=0 $Y2=0
cc_391 N_A_711_307#_M1023_g N_A_560_47#_c_695_n 0.0208156f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_392 N_A_711_307#_c_596_n N_A_560_47#_c_695_n 0.0148917f $X=4.78 $Y=1.7 $X2=0
+ $Y2=0
cc_393 N_A_711_307#_c_597_n N_A_560_47#_c_695_n 0.00487525f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_394 N_A_711_307#_c_587_n N_A_560_47#_c_695_n 0.0110111f $X=4.54 $Y=0.74 $X2=0
+ $Y2=0
cc_395 N_A_711_307#_M1023_g N_A_560_47#_c_706_n 0.00160708f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_396 N_A_711_307#_M1023_g N_A_560_47#_c_697_n 0.0103832f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_397 N_A_711_307#_M1009_g N_A_560_47#_c_703_n 0.0213969f $X=3.63 $Y=2.275
+ $X2=0 $Y2=0
cc_398 N_A_711_307#_M1023_g N_A_560_47#_c_703_n 0.00748409f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_399 N_A_711_307#_c_596_n N_A_560_47#_c_703_n 0.0192637f $X=4.78 $Y=1.7 $X2=0
+ $Y2=0
cc_400 N_A_711_307#_c_597_n N_A_560_47#_c_703_n 0.0103945f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_401 N_A_711_307#_M1023_g N_A_560_47#_c_698_n 0.0244837f $X=3.69 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_711_307#_c_596_n N_A_560_47#_c_698_n 0.02399f $X=4.78 $Y=1.7 $X2=0
+ $Y2=0
cc_403 N_A_711_307#_c_597_n N_A_560_47#_c_698_n 0.0067022f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_404 N_A_711_307#_M1004_g N_RESET_B_M1005_g 0.00675716f $X=5.935 $Y=1.985
+ $X2=0 $Y2=0
cc_405 N_A_711_307#_c_622_p N_RESET_B_M1005_g 0.0164645f $X=5.655 $Y=1.65 $X2=0
+ $Y2=0
cc_406 N_A_711_307#_c_588_n N_RESET_B_M1005_g 0.00360226f $X=5.805 $Y=1.16 $X2=0
+ $Y2=0
cc_407 N_A_711_307#_c_583_n RESET_B 0.00338448f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_408 N_A_711_307#_c_596_n RESET_B 0.0177238f $X=4.78 $Y=1.7 $X2=0 $Y2=0
cc_409 N_A_711_307#_c_607_p RESET_B 0.0604948f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_410 N_A_711_307#_c_587_n RESET_B 0.00545394f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_411 N_A_711_307#_c_622_p RESET_B 0.0283296f $X=5.655 $Y=1.65 $X2=0 $Y2=0
cc_412 N_A_711_307#_c_588_n RESET_B 0.0222979f $X=5.805 $Y=1.16 $X2=0 $Y2=0
cc_413 N_A_711_307#_c_630_p RESET_B 0.0122277f $X=4.865 $Y=1.755 $X2=0 $Y2=0
cc_414 N_A_711_307#_c_583_n N_RESET_B_c_775_n 0.00715465f $X=6.01 $Y=1.16 $X2=0
+ $Y2=0
cc_415 N_A_711_307#_c_607_p N_RESET_B_c_775_n 0.0017807f $X=5.655 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A_711_307#_c_588_n N_RESET_B_c_775_n 2.97021e-19 $X=5.805 $Y=1.16 $X2=0
+ $Y2=0
cc_417 N_A_711_307#_c_630_p N_RESET_B_c_775_n 7.74669e-19 $X=4.865 $Y=1.755
+ $X2=0 $Y2=0
cc_418 N_A_711_307#_c_581_n N_RESET_B_c_776_n 0.0066515f $X=5.935 $Y=0.995 $X2=0
+ $Y2=0
cc_419 N_A_711_307#_c_607_p N_RESET_B_c_776_n 0.0131853f $X=5.655 $Y=0.74 $X2=0
+ $Y2=0
cc_420 N_A_711_307#_c_588_n N_RESET_B_c_776_n 0.00291283f $X=5.805 $Y=1.16 $X2=0
+ $Y2=0
cc_421 N_A_711_307#_M1016_g N_A_1308_47#_M1014_g 0.0227021f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_422 N_A_711_307#_M1002_g N_A_1308_47#_c_810_n 0.0183974f $X=6.875 $Y=0.445
+ $X2=0 $Y2=0
cc_423 N_A_711_307#_M1016_g N_A_1308_47#_c_815_n 0.0307383f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_424 N_A_711_307#_c_585_n N_A_1308_47#_c_811_n 0.018261f $X=6.875 $Y=1.16
+ $X2=0 $Y2=0
cc_425 N_A_711_307#_c_585_n N_A_1308_47#_c_812_n 0.0197483f $X=6.875 $Y=1.16
+ $X2=0 $Y2=0
cc_426 N_A_711_307#_c_582_n N_A_1308_47#_c_823_n 0.0179878f $X=6.8 $Y=1.16 $X2=0
+ $Y2=0
cc_427 N_A_711_307#_c_585_n N_A_1308_47#_c_823_n 0.00223011f $X=6.875 $Y=1.16
+ $X2=0 $Y2=0
cc_428 N_A_711_307#_M1002_g N_A_1308_47#_c_813_n 0.0200172f $X=6.875 $Y=0.445
+ $X2=0 $Y2=0
cc_429 N_A_711_307#_c_596_n N_VPWR_M1013_s 0.00663785f $X=4.78 $Y=1.7 $X2=0
+ $Y2=0
cc_430 N_A_711_307#_c_622_p N_VPWR_M1005_d 0.0221843f $X=5.655 $Y=1.65 $X2=0
+ $Y2=0
cc_431 N_A_711_307#_c_588_n N_VPWR_M1005_d 8.26946e-19 $X=5.805 $Y=1.16 $X2=0
+ $Y2=0
cc_432 N_A_711_307#_M1016_g N_VPWR_c_853_n 0.00537515f $X=6.875 $Y=2.165 $X2=0
+ $Y2=0
cc_433 N_A_711_307#_c_606_p N_VPWR_c_856_n 0.00972841f $X=4.865 $Y=2.27 $X2=0
+ $Y2=0
cc_434 N_A_711_307#_M1004_g N_VPWR_c_857_n 0.00468308f $X=5.935 $Y=1.985 $X2=0
+ $Y2=0
cc_435 N_A_711_307#_M1016_g N_VPWR_c_857_n 0.00541359f $X=6.875 $Y=2.165 $X2=0
+ $Y2=0
cc_436 N_A_711_307#_M1013_d N_VPWR_c_850_n 0.00490525f $X=4.69 $Y=1.485 $X2=0
+ $Y2=0
cc_437 N_A_711_307#_M1009_g N_VPWR_c_850_n 0.0103589f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_438 N_A_711_307#_M1004_g N_VPWR_c_850_n 0.00921791f $X=5.935 $Y=1.985 $X2=0
+ $Y2=0
cc_439 N_A_711_307#_M1016_g N_VPWR_c_850_n 0.0110992f $X=6.875 $Y=2.165 $X2=0
+ $Y2=0
cc_440 N_A_711_307#_c_596_n N_VPWR_c_850_n 0.00903489f $X=4.78 $Y=1.7 $X2=0
+ $Y2=0
cc_441 N_A_711_307#_c_597_n N_VPWR_c_850_n 0.00123717f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_442 N_A_711_307#_c_606_p N_VPWR_c_850_n 0.00637538f $X=4.865 $Y=2.27 $X2=0
+ $Y2=0
cc_443 N_A_711_307#_M1009_g N_VPWR_c_862_n 0.00520872f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_444 N_A_711_307#_M1009_g N_VPWR_c_863_n 0.00483063f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_445 N_A_711_307#_c_596_n N_VPWR_c_863_n 0.0390798f $X=4.78 $Y=1.7 $X2=0 $Y2=0
cc_446 N_A_711_307#_c_597_n N_VPWR_c_863_n 0.00807403f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_447 N_A_711_307#_c_606_p N_VPWR_c_863_n 0.0215518f $X=4.865 $Y=2.27 $X2=0
+ $Y2=0
cc_448 N_A_711_307#_M1004_g N_VPWR_c_864_n 0.0131127f $X=5.935 $Y=1.985 $X2=0
+ $Y2=0
cc_449 N_A_711_307#_c_583_n N_VPWR_c_864_n 5.88929e-19 $X=6.01 $Y=1.16 $X2=0
+ $Y2=0
cc_450 N_A_711_307#_c_622_p N_VPWR_c_864_n 0.055093f $X=5.655 $Y=1.65 $X2=0
+ $Y2=0
cc_451 N_A_711_307#_c_581_n Q 0.00708343f $X=5.935 $Y=0.995 $X2=0 $Y2=0
cc_452 N_A_711_307#_M1004_g Q 0.00898269f $X=5.935 $Y=1.985 $X2=0 $Y2=0
cc_453 N_A_711_307#_c_582_n Q 0.0353039f $X=6.8 $Y=1.16 $X2=0 $Y2=0
cc_454 N_A_711_307#_M1002_g Q 0.00240253f $X=6.875 $Y=0.445 $X2=0 $Y2=0
cc_455 N_A_711_307#_M1016_g Q 0.00408436f $X=6.875 $Y=2.165 $X2=0 $Y2=0
cc_456 N_A_711_307#_c_588_n Q 0.0488918f $X=5.805 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_711_307#_c_607_p N_VGND_M1020_d 0.0200993f $X=5.655 $Y=0.74 $X2=0
+ $Y2=0
cc_458 N_A_711_307#_c_588_n N_VGND_M1020_d 9.49324e-19 $X=5.805 $Y=1.16 $X2=0
+ $Y2=0
cc_459 N_A_711_307#_M1023_g N_VGND_c_996_n 0.0115105f $X=3.69 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_A_711_307#_c_586_n N_VGND_c_996_n 0.0227609f $X=4.39 $Y=0.655 $X2=0
+ $Y2=0
cc_461 N_A_711_307#_M1002_g N_VGND_c_997_n 0.00310635f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_462 N_A_711_307#_M1023_g N_VGND_c_1000_n 0.0046653f $X=3.69 $Y=0.445 $X2=0
+ $Y2=0
cc_463 N_A_711_307#_c_581_n N_VGND_c_1001_n 0.0046653f $X=5.935 $Y=0.995 $X2=0
+ $Y2=0
cc_464 N_A_711_307#_M1002_g N_VGND_c_1001_n 0.00579312f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_465 N_A_711_307#_M1015_s N_VGND_c_1003_n 0.00215226f $X=4.295 $Y=0.235 $X2=0
+ $Y2=0
cc_466 N_A_711_307#_M1023_g N_VGND_c_1003_n 0.00813035f $X=3.69 $Y=0.445 $X2=0
+ $Y2=0
cc_467 N_A_711_307#_c_581_n N_VGND_c_1003_n 0.00929621f $X=5.935 $Y=0.995 $X2=0
+ $Y2=0
cc_468 N_A_711_307#_M1002_g N_VGND_c_1003_n 0.0118997f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_469 N_A_711_307#_c_586_n N_VGND_c_1003_n 0.011424f $X=4.39 $Y=0.655 $X2=0
+ $Y2=0
cc_470 N_A_711_307#_c_607_p N_VGND_c_1003_n 0.0182342f $X=5.655 $Y=0.74 $X2=0
+ $Y2=0
cc_471 N_A_711_307#_c_586_n N_VGND_c_1007_n 0.0193675f $X=4.39 $Y=0.655 $X2=0
+ $Y2=0
cc_472 N_A_711_307#_c_607_p N_VGND_c_1007_n 0.00843435f $X=5.655 $Y=0.74 $X2=0
+ $Y2=0
cc_473 N_A_711_307#_c_581_n N_VGND_c_1008_n 0.00985451f $X=5.935 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_711_307#_c_583_n N_VGND_c_1008_n 6.83192e-19 $X=6.01 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_A_711_307#_c_607_p N_VGND_c_1008_n 0.0510955f $X=5.655 $Y=0.74 $X2=0
+ $Y2=0
cc_476 N_A_711_307#_c_607_p A_941_47# 0.0050941f $X=5.655 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_477 N_A_560_47#_M1013_g N_RESET_B_M1005_g 0.0210644f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_478 N_A_560_47#_c_695_n RESET_B 0.00935533f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_479 N_A_560_47#_c_696_n RESET_B 0.0127404f $X=4.622 $Y=1.16 $X2=0 $Y2=0
cc_480 N_A_560_47#_c_698_n RESET_B 0.02034f $X=4.115 $Y=1.16 $X2=0 $Y2=0
cc_481 N_A_560_47#_c_696_n N_RESET_B_c_775_n 0.0215022f $X=4.622 $Y=1.16 $X2=0
+ $Y2=0
cc_482 N_A_560_47#_c_694_n N_RESET_B_c_776_n 0.0386574f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_560_47#_c_705_n N_VPWR_c_852_n 0.00578043f $X=3.27 $Y=2.34 $X2=0
+ $Y2=0
cc_484 N_A_560_47#_M1013_g N_VPWR_c_856_n 0.00388479f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_A_560_47#_M1001_d N_VPWR_c_850_n 0.00173718f $X=2.805 $Y=2.065 $X2=0
+ $Y2=0
cc_486 N_A_560_47#_M1013_g N_VPWR_c_850_n 0.00389183f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_487 N_A_560_47#_c_705_n N_VPWR_c_850_n 0.0100566f $X=3.27 $Y=2.34 $X2=0 $Y2=0
cc_488 N_A_560_47#_c_703_n N_VPWR_c_850_n 0.0121128f $X=3.52 $Y=1.96 $X2=0 $Y2=0
cc_489 N_A_560_47#_c_705_n N_VPWR_c_862_n 0.0226583f $X=3.27 $Y=2.34 $X2=0 $Y2=0
cc_490 N_A_560_47#_c_703_n N_VPWR_c_862_n 0.0156263f $X=3.52 $Y=1.96 $X2=0 $Y2=0
cc_491 N_A_560_47#_M1013_g N_VPWR_c_863_n 0.0117394f $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_492 N_A_560_47#_M1013_g N_VPWR_c_864_n 6.44953e-19 $X=4.615 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_A_560_47#_c_703_n A_645_413# 0.0058803f $X=3.52 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_494 N_A_560_47#_c_706_n N_VGND_c_995_n 0.00233913f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_495 N_A_560_47#_c_694_n N_VGND_c_996_n 0.00298695f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_496 N_A_560_47#_c_695_n N_VGND_c_996_n 0.00169847f $X=4.54 $Y=1.16 $X2=0
+ $Y2=0
cc_497 N_A_560_47#_c_706_n N_VGND_c_996_n 0.01063f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_498 N_A_560_47#_c_698_n N_VGND_c_996_n 0.0122055f $X=4.115 $Y=1.16 $X2=0
+ $Y2=0
cc_499 N_A_560_47#_c_706_n N_VGND_c_1000_n 0.0247905f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_500 N_A_560_47#_M1018_d N_VGND_c_1003_n 0.00288975f $X=2.8 $Y=0.235 $X2=0
+ $Y2=0
cc_501 N_A_560_47#_c_694_n N_VGND_c_1003_n 0.00739361f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_A_560_47#_c_706_n N_VGND_c_1003_n 0.0247067f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_503 N_A_560_47#_c_694_n N_VGND_c_1007_n 0.00428022f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_560_47#_c_694_n N_VGND_c_1008_n 0.00186338f $X=4.63 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_A_560_47#_c_706_n A_658_47# 0.0038256f $X=3.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_506 N_A_560_47#_c_697_n A_658_47# 0.00152789f $X=3.415 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_507 N_RESET_B_M1005_g N_VPWR_c_856_n 0.00468308f $X=5.075 $Y=1.985 $X2=0
+ $Y2=0
cc_508 N_RESET_B_M1005_g N_VPWR_c_850_n 0.00809505f $X=5.075 $Y=1.985 $X2=0
+ $Y2=0
cc_509 N_RESET_B_M1005_g N_VPWR_c_863_n 6.32662e-19 $X=5.075 $Y=1.985 $X2=0
+ $Y2=0
cc_510 N_RESET_B_M1005_g N_VPWR_c_864_n 0.0114795f $X=5.075 $Y=1.985 $X2=0 $Y2=0
cc_511 N_RESET_B_c_776_n N_VGND_c_1003_n 0.00410127f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_512 N_RESET_B_c_776_n N_VGND_c_1007_n 0.00341689f $X=5.05 $Y=0.995 $X2=0
+ $Y2=0
cc_513 N_RESET_B_c_776_n N_VGND_c_1008_n 0.0112079f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_514 N_A_1308_47#_M1014_g N_VPWR_c_853_n 0.0132029f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_515 N_A_1308_47#_c_815_n N_VPWR_c_853_n 0.0454653f $X=6.665 $Y=2.165 $X2=0
+ $Y2=0
cc_516 N_A_1308_47#_c_811_n N_VPWR_c_853_n 0.00978365f $X=7.31 $Y=1.16 $X2=0
+ $Y2=0
cc_517 N_A_1308_47#_c_812_n N_VPWR_c_853_n 0.00160788f $X=7.31 $Y=1.16 $X2=0
+ $Y2=0
cc_518 N_A_1308_47#_c_815_n N_VPWR_c_857_n 0.0153916f $X=6.665 $Y=2.165 $X2=0
+ $Y2=0
cc_519 N_A_1308_47#_M1014_g N_VPWR_c_858_n 0.0046653f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_520 N_A_1308_47#_M1016_s N_VPWR_c_850_n 0.00352456f $X=6.54 $Y=1.845 $X2=0
+ $Y2=0
cc_521 N_A_1308_47#_M1014_g N_VPWR_c_850_n 0.008846f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_522 N_A_1308_47#_c_815_n N_VPWR_c_850_n 0.00941829f $X=6.665 $Y=2.165 $X2=0
+ $Y2=0
cc_523 N_A_1308_47#_c_810_n Q 0.0595519f $X=6.665 $Y=0.51 $X2=0 $Y2=0
cc_524 N_A_1308_47#_c_815_n Q 0.0924595f $X=6.665 $Y=2.165 $X2=0 $Y2=0
cc_525 N_A_1308_47#_c_823_n Q 0.0264547f $X=6.705 $Y=1.16 $X2=0 $Y2=0
cc_526 N_A_1308_47#_M1014_g Q_N 0.0158846f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_527 N_A_1308_47#_c_811_n Q_N 0.0262099f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_528 N_A_1308_47#_c_812_n Q_N 0.00800507f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_529 N_A_1308_47#_c_813_n Q_N 0.0136059f $X=7.325 $Y=0.995 $X2=0 $Y2=0
cc_530 N_A_1308_47#_c_811_n N_VGND_c_997_n 0.0100674f $X=7.31 $Y=1.16 $X2=0
+ $Y2=0
cc_531 N_A_1308_47#_c_812_n N_VGND_c_997_n 0.00156823f $X=7.31 $Y=1.16 $X2=0
+ $Y2=0
cc_532 N_A_1308_47#_c_813_n N_VGND_c_997_n 0.00870521f $X=7.325 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_A_1308_47#_c_810_n N_VGND_c_1001_n 0.0136871f $X=6.665 $Y=0.51 $X2=0
+ $Y2=0
cc_534 N_A_1308_47#_c_813_n N_VGND_c_1002_n 0.0046653f $X=7.325 $Y=0.995 $X2=0
+ $Y2=0
cc_535 N_A_1308_47#_M1002_s N_VGND_c_1003_n 0.00352456f $X=6.54 $Y=0.235 $X2=0
+ $Y2=0
cc_536 N_A_1308_47#_c_810_n N_VGND_c_1003_n 0.00856983f $X=6.665 $Y=0.51 $X2=0
+ $Y2=0
cc_537 N_A_1308_47#_c_813_n N_VGND_c_1003_n 0.008846f $X=7.325 $Y=0.995 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_850_n A_465_369# 0.00476473f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_539 N_VPWR_c_850_n A_645_413# 0.00267862f $X=7.59 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_540 N_VPWR_c_850_n N_Q_M1004_d 0.00382897f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_541 N_VPWR_c_857_n Q 0.0244536f $X=7.01 $Y=2.72 $X2=0 $Y2=0
cc_542 N_VPWR_c_850_n Q 0.0134021f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_543 N_VPWR_c_850_n N_Q_N_M1014_d 0.00382897f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_544 N_VPWR_c_858_n Q_N 0.018001f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_545 N_VPWR_c_850_n Q_N 0.00993603f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_546 Q N_VGND_c_1001_n 0.0244536f $X=6.1 $Y=0.425 $X2=0 $Y2=0
cc_547 N_Q_M1008_d N_VGND_c_1003_n 0.00387172f $X=6.01 $Y=0.235 $X2=0 $Y2=0
cc_548 Q N_VGND_c_1003_n 0.0134021f $X=6.1 $Y=0.425 $X2=0 $Y2=0
cc_549 N_Q_N_c_982_n N_VGND_c_1002_n 0.0171222f $X=7.65 $Y=0.425 $X2=0 $Y2=0
cc_550 N_Q_N_M1019_d N_VGND_c_1003_n 0.00379446f $X=7.425 $Y=0.235 $X2=0 $Y2=0
cc_551 N_Q_N_c_982_n N_VGND_c_1003_n 0.00983509f $X=7.65 $Y=0.425 $X2=0 $Y2=0
cc_552 N_VGND_c_1003_n A_465_47# 0.0108492f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_553 N_VGND_c_1003_n A_658_47# 0.00669936f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24
cc_554 N_VGND_c_1003_n A_941_47# 0.00353055f $X=7.59 $Y=0 $X2=-0.19 $Y2=-0.24

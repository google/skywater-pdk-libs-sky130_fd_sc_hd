* File: sky130_fd_sc_hd__or4bb_4.spice
* Created: Thu Aug 27 14:44:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or4bb_4.spice.pex"
.subckt sky130_fd_sc_hd__or4bb_4  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_C_N_M1014_g N_A_27_410#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.1092 PD=0.715 PS=1.36 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_A_205_93#_M1016_d N_D_N_M1016_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.06195 PD=1.36 PS=0.715 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_315_380#_M1004_d N_A_205_93#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1235 AS=0.169 PD=1.03 PS=1.82 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_27_410#_M1007_g N_A_315_380#_M1004_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=0 NRS=4.608 M=1 R=4.33333
+ SA=75000.7 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_315_380#_M1005_d N_B_M1005_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_A_315_380#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.08775 PD=1.03 PS=0.92 NRD=17.532 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1008_d N_A_315_380#_M1008_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75002.1
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1008_d N_A_315_380#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1012 N_X_M1012_d N_A_315_380#_M1012_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1012_d N_A_315_380#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1017 N_VPWR_M1017_d N_C_N_M1017_g N_A_27_410#_M1017_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.122612 AS=0.1092 PD=1.32 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_205_93#_M1018_d N_D_N_M1018_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.11295 AS=0.122612 PD=1.4 PS=1.32 NRD=0 NRS=111.128 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_397_297# N_A_205_93#_M1002_g N_A_315_380#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.18 AS=0.257925 PD=1.36 PS=2.52 NRD=24.6053 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1003 A_499_297# N_A_27_410#_M1003_g A_397_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.18 PD=1.27 PS=1.36 NRD=15.7403 NRS=24.6053 M=1 R=6.66667 SA=75000.7
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1000 A_583_297# N_B_M1000_g A_499_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A_M1019_g A_583_297# VPB PHIGHVT L=0.15 W=1 AD=0.19
+ AS=0.135 PD=1.38 PS=1.27 NRD=9.8303 NRS=15.7403 M=1 R=6.66667 SA=75001.5
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_315_380#_M1001_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.19 PD=1.27 PS=1.38 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.1
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1006 N_X_M1001_d N_A_315_380#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1010_d N_A_315_380#_M1010_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_X_M1010_d N_A_315_380#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__or4bb_4.spice.SKY130_FD_SC_HD__OR4BB_4.pxi"
*
.ends
*
*

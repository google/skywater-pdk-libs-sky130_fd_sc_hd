* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
M1000 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=8.224e+11p pd=6.71e+06u as=1.134e+11p ps=1.38e+06u
M1001 a_228_47# a_27_47# VPWR VPB phighvt w=820000u l=150000u
+  ad=3.116e+11p pd=2.4e+06u as=1.5189e+12p ps=9.27e+06u
M1002 VPWR a_362_333# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1003 a_228_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=2.6325e+11p pd=2.11e+06u as=0p ps=0u
M1004 VPWR a_228_47# a_362_333# VPB phighvt w=820000u l=150000u
+  ad=0p pd=0u as=2.173e+11p ps=2.17e+06u
M1005 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 X a_362_333# VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1007 X a_362_333# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_362_333# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_228_47# a_362_333# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
.ends

* File: sky130_fd_sc_hd__a22o_2.spice
* Created: Thu Aug 27 14:02:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a22o_2.spice.pex"
.subckt sky130_fd_sc_hd__a22o_2  VNB VPB B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1011 A_109_47# N_B2_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65 AD=0.07475
+ AS=0.169 PD=0.88 PS=1.82 NRD=11.076 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1000 N_A_27_297#_M1000_d N_B1_M1000_g A_109_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.07475 PD=1.82 PS=0.88 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 A_381_47# N_A1_M1001_g N_A_27_297#_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.169 PD=0.98 PS=1.82 NRD=20.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g A_381_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.102375 AS=0.10725 PD=0.965 PS=0.98 NRD=0 NRS=20.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_27_297#_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.102375 PD=0.92 PS=0.965 NRD=0 NRS=7.38 M=1 R=4.33333
+ SA=75001.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1007_d N_A_27_297#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1755 PD=0.92 PS=1.84 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_109_297#_M1008_d N_B2_M1008_g N_A_27_297#_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_27_297#_M1002_d N_B1_M1002_g N_A_109_297#_M1008_d VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1010 N_A_109_297#_M1010_d N_A1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.26 PD=1.33 PS=2.52 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_109_297#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1575 AS=0.165 PD=1.315 PS=1.33 NRD=7.8603 NRS=5.8903 M=1 R=6.66667
+ SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1005_d N_A_27_297#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1575 AS=0.135 PD=1.315 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_27_297#_M1004_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.135 PD=2.54 PS=1.27 NRD=0.9653 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__a22o_2.spice.SKY130_FD_SC_HD__A22O_2.pxi"
*
.ends
*
*

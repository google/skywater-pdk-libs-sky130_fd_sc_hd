* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
M1000 VGND a_283_47# a_390_47# VNB nshort w=650000u l=500000u
+  ad=5.686e+11p pd=5.6e+06u as=1.69e+11p ps=1.82e+06u
M1001 X a_390_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
M1002 a_283_47# a_27_47# VGND VNB nshort w=650000u l=500000u
+  ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1003 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1004 VPWR a_390_47# X VPB phighvt w=1e+06u l=150000u
+  ad=1.0458e+12p pd=8.16e+06u as=2.75e+11p ps=2.55e+06u
M1005 VGND a_390_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 VPWR a_283_47# a_390_47# VPB phighvt w=820000u l=500000u
+  ad=0p pd=0u as=2.132e+11p ps=2.16e+06u
M1008 a_283_47# a_27_47# VPWR VPB phighvt w=820000u l=500000u
+  ad=2.173e+11p pd=2.17e+06u as=0p ps=0u
M1009 X a_390_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

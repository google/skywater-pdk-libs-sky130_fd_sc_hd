* File: sky130_fd_sc_hd__nand4bb_2.spice
* Created: Tue Sep  1 19:17:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand4bb_2.pex.spice"
.subckt sky130_fd_sc_hd__nand4bb_2  VNB VPB B_N A_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* A_N	A_N
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_B_N_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1006 N_A_193_47#_M1006_d N_A_N_M1006_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1974 AS=0.0567 PD=1.78 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_A_193_47#_M1009_g N_A_341_47#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1009_d N_A_193_47#_M1015_g N_A_341_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1014 N_A_591_47#_M1014_d N_A_27_47#_M1014_g N_A_341_47#_M1015_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_A_591_47#_M1014_d N_A_27_47#_M1018_g N_A_341_47#_M1018_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_591_47#_M1010_d N_C_M1010_g N_A_781_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1016 N_A_591_47#_M1010_d N_C_M1016_g N_A_781_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1003 N_A_781_47#_M1016_s N_D_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_A_781_47#_M1007_d N_D_M1007_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_B_N_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1019 N_A_193_47#_M1019_d N_A_N_M1019_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1974 AS=0.0567 PD=1.78 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_193_47#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A_193_47#_M1008_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1008_d N_A_27_47#_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_27_47#_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.395 AS=0.135 PD=1.79 PS=1.27 NRD=14.7553 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1001_d N_C_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.395
+ AS=0.135 PD=1.79 PS=1.27 NRD=14.7553 NRS=0 M=1 R=6.66667 SA=75002.4 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_C_M1013_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1002 N_Y_M1002_d N_D_M1002_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1002_d N_D_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.6 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__nand4bb_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a21bo_4.pex.spice
* Created: Tue Sep  1 18:51:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21BO_4%B1_N 3 6 8 11 13
c32 11 0 9.79304e-20 $X=0.665 $Y=1.16
r33 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.16
+ $X2=0.665 $Y2=1.325
r34 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.16
+ $X2=0.665 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.665
+ $Y=1.16 $X2=0.665 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.67 $Y=1.985
+ $X2=0.67 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.67 $Y=0.56 $X2=0.67
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%A_205_21# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 38 44 45 49 53 55 58 59 63 67
c139 55 0 4.87616e-20 $X=4.685 $Y=0.755
r140 75 76 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.96 $Y=1.16
+ $X2=2.39 $Y2=1.16
r141 71 73 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.1 $Y=1.16
+ $X2=1.53 $Y2=1.16
r142 67 69 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.825 $Y=0.57
+ $X2=4.825 $Y2=0.755
r143 61 63 17.1785 $w=1.83e-07 $l=2.85e-07 $layer=LI1_cond $X=2.725 $Y=0.707
+ $X2=3.01 $Y2=0.707
r144 59 76 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.445 $Y=1.16
+ $X2=2.39 $Y2=1.16
r145 58 60 14.1743 $w=2.41e-07 $l=2.8e-07 $layer=LI1_cond $X=2.445 $Y=1.16
+ $X2=2.725 $Y2=1.16
r146 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.445
+ $Y=1.16 $X2=2.445 $Y2=1.16
r147 56 65 3.05 $w=1.7e-07 $l=9.80051e-08 $layer=LI1_cond $X=3.645 $Y=0.755
+ $X2=3.56 $Y2=0.727
r148 55 69 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.685 $Y=0.755
+ $X2=4.825 $Y2=0.755
r149 55 56 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.685 $Y=0.755
+ $X2=3.645 $Y2=0.755
r150 51 65 3.05 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.56 $Y=0.84 $X2=3.56
+ $Y2=0.727
r151 51 53 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.56 $Y=0.84
+ $X2=3.56 $Y2=1.62
r152 47 65 3.05 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.56 $Y=0.615 $X2=3.56
+ $Y2=0.727
r153 47 49 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.56 $Y=0.615
+ $X2=3.56 $Y2=0.42
r154 45 65 3.05 $w=1.7e-07 $l=9.75705e-08 $layer=LI1_cond $X=3.475 $Y=0.7
+ $X2=3.56 $Y2=0.727
r155 45 63 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.475 $Y=0.7
+ $X2=3.01 $Y2=0.7
r156 44 60 2.78154 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0.995
+ $X2=2.725 $Y2=1.16
r157 43 61 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=2.725 $Y=0.8
+ $X2=2.725 $Y2=0.707
r158 43 44 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.725 $Y=0.8
+ $X2=2.725 $Y2=0.995
r159 41 75 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.765 $Y=1.16
+ $X2=1.96 $Y2=1.16
r160 41 73 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.765 $Y=1.16
+ $X2=1.53 $Y2=1.16
r161 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.16 $X2=1.765 $Y2=1.16
r162 38 58 3.86752 $w=3.3e-07 $l=8e-08 $layer=LI1_cond $X=2.365 $Y=1.16
+ $X2=2.445 $Y2=1.16
r163 38 40 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=2.365 $Y=1.16
+ $X2=1.765 $Y2=1.16
r164 34 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=1.325
+ $X2=2.39 $Y2=1.16
r165 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.39 $Y=1.325
+ $X2=2.39 $Y2=1.985
r166 31 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=0.995
+ $X2=2.39 $Y2=1.16
r167 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.39 $Y=0.995
+ $X2=2.39 $Y2=0.56
r168 27 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.325
+ $X2=1.96 $Y2=1.16
r169 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.96 $Y=1.325
+ $X2=1.96 $Y2=1.985
r170 24 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=0.995
+ $X2=1.96 $Y2=1.16
r171 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.96 $Y=0.995
+ $X2=1.96 $Y2=0.56
r172 20 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.53 $Y=1.325
+ $X2=1.53 $Y2=1.16
r173 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.53 $Y=1.325
+ $X2=1.53 $Y2=1.985
r174 17 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=1.16
r175 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=0.56
r176 13 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.325
+ $X2=1.1 $Y2=1.16
r177 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.1 $Y=1.325
+ $X2=1.1 $Y2=1.985
r178 10 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=0.995
+ $X2=1.1 $Y2=1.16
r179 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.1 $Y=0.995
+ $X2=1.1 $Y2=0.56
r180 3 53 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.56 $Y2=1.62
r181 2 67 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.235 $X2=4.82 $Y2=0.57
r182 1 65 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.425
+ $Y=0.235 $X2=3.56 $Y2=0.76
r183 1 49 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.425
+ $Y=0.235 $X2=3.56 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%A_42_47# 1 2 7 9 12 14 16 19 22 23 26 27 29
+ 33 38 48
c104 38 0 9.79304e-20 $X=0.335 $Y=2.02
r105 47 48 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.35 $Y=1.16
+ $X2=3.77 $Y2=1.16
r106 38 40 7.57428 $w=4.51e-07 $l=2.8e-07 $layer=LI1_cond $X=0.335 $Y=2.02
+ $X2=0.335 $Y2=2.3
r107 37 38 1.62306 $w=4.51e-07 $l=6e-08 $layer=LI1_cond $X=0.335 $Y=1.96
+ $X2=0.335 $Y2=2.02
r108 33 35 15.3925 $w=4.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.322 $Y=0.36
+ $X2=0.322 $Y2=0.84
r109 30 47 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=3.22 $Y=1.16
+ $X2=3.35 $Y2=1.16
r110 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.16 $X2=3.22 $Y2=1.16
r111 27 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.15 $Y=1.44
+ $X2=2.785 $Y2=1.44
r112 27 29 7.24924 $w=3.08e-07 $l=1.95e-07 $layer=LI1_cond $X=3.15 $Y=1.355
+ $X2=3.15 $Y2=1.16
r113 25 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.525
+ $X2=2.785 $Y2=1.44
r114 25 26 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.785 $Y=1.525
+ $X2=2.785 $Y2=1.935
r115 24 38 6.51405 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.565 $Y=2.02
+ $X2=0.335 $Y2=2.02
r116 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.7 $Y=2.02
+ $X2=2.785 $Y2=1.935
r117 23 24 139.289 $w=1.68e-07 $l=2.135e-06 $layer=LI1_cond $X=2.7 $Y=2.02
+ $X2=0.565 $Y2=2.02
r118 22 37 7.52558 $w=4.51e-07 $l=2.1609e-07 $layer=LI1_cond $X=0.217 $Y=1.795
+ $X2=0.335 $Y2=1.96
r119 22 35 48.9148 $w=2.23e-07 $l=9.55e-07 $layer=LI1_cond $X=0.217 $Y=1.795
+ $X2=0.217 $Y2=0.84
r120 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.77 $Y=1.325
+ $X2=3.77 $Y2=1.16
r121 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.77 $Y=1.325
+ $X2=3.77 $Y2=1.985
r122 14 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.77 $Y=0.995
+ $X2=3.77 $Y2=1.16
r123 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.77 $Y=0.995
+ $X2=3.77 $Y2=0.56
r124 10 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.325
+ $X2=3.35 $Y2=1.16
r125 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.35 $Y=1.325
+ $X2=3.35 $Y2=1.985
r126 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=0.995
+ $X2=3.35 $Y2=1.16
r127 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.35 $Y=0.995
+ $X2=3.35 $Y2=0.56
r128 2 40 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.485 $X2=0.455 $Y2=2.3
r129 2 37 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.485 $X2=0.455 $Y2=1.96
r130 1 33 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.235 $X2=0.375 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%A2 3 7 10 13 16 17 19 20 24 26 28 30 35 37
+ 39 42
c79 30 0 9.49649e-20 $X=5.22 $Y=1.445
c80 24 0 1.1533e-19 $X=4.19 $Y=1.16
c81 13 0 2.74367e-20 $X=5.45 $Y=1.985
c82 3 0 2.98924e-20 $X=4.19 $Y=1.985
r83 39 42 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.305 $Y=1.595
+ $X2=5.305 $Y2=1.53
r84 30 39 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.305 $Y=1.68
+ $X2=5.305 $Y2=1.595
r85 30 42 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.305 $Y=1.52
+ $X2=5.305 $Y2=1.53
r86 29 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.305 $Y=1.29
+ $X2=5.305 $Y2=1.52
r87 28 30 46.8468 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=4.42 $Y=1.68 $X2=5.22
+ $Y2=1.68
r88 24 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.16
+ $X2=4.19 $Y2=0.995
r89 23 26 6.17535 $w=2.63e-07 $l=1.42e-07 $layer=LI1_cond $X=4.19 $Y=1.142
+ $X2=4.332 $Y2=1.142
r90 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=1.16 $X2=4.19 $Y2=1.16
r91 20 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.51 $Y=1.16
+ $X2=5.51 $Y2=1.325
r92 20 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.51 $Y=1.16
+ $X2=5.51 $Y2=0.995
r93 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.51
+ $Y=1.16 $X2=5.51 $Y2=1.16
r94 17 29 7.04737 $w=2.35e-07 $l=1.54771e-07 $layer=LI1_cond $X=5.39 $Y=1.172
+ $X2=5.305 $Y2=1.29
r95 17 19 5.88482 $w=2.33e-07 $l=1.2e-07 $layer=LI1_cond $X=5.39 $Y=1.172
+ $X2=5.51 $Y2=1.172
r96 16 28 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=4.332 $Y=1.595
+ $X2=4.42 $Y2=1.68
r97 15 26 3.18883 $w=1.75e-07 $l=1.33e-07 $layer=LI1_cond $X=4.332 $Y=1.275
+ $X2=4.332 $Y2=1.142
r98 15 16 20.2805 $w=1.73e-07 $l=3.2e-07 $layer=LI1_cond $X=4.332 $Y=1.275
+ $X2=4.332 $Y2=1.595
r99 13 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.45 $Y=1.985
+ $X2=5.45 $Y2=1.325
r100 10 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.45 $Y=0.56
+ $X2=5.45 $Y2=0.995
r101 7 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.23 $Y=0.56
+ $X2=4.23 $Y2=0.995
r102 1 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.325
+ $X2=4.19 $Y2=1.16
r103 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.19 $Y=1.325
+ $X2=4.19 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%A1 1 3 6 8 10 13 15 22
c45 15 0 5.7329e-20 $X=4.845 $Y=1.19
c46 8 0 4.87616e-20 $X=5.03 $Y=0.995
r47 20 22 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=5.03 $Y2=1.16
r48 17 20 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.61 $Y=1.16 $X2=4.79
+ $Y2=1.16
r49 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.79
+ $Y=1.16 $X2=4.79 $Y2=1.16
r50 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.03 $Y=1.325
+ $X2=5.03 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.03 $Y=1.325
+ $X2=5.03 $Y2=1.985
r52 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.03 $Y=0.995
+ $X2=5.03 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.03 $Y=0.995
+ $X2=5.03 $Y2=0.56
r54 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.61 $Y=1.325
+ $X2=4.61 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.61 $Y=1.325 $X2=4.61
+ $Y2=1.985
r56 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.61 $Y=0.995
+ $X2=4.61 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.61 $Y=0.995 $X2=4.61
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%VPWR 1 2 3 4 5 18 20 24 28 32 36 38 39 40 46
+ 51 59 66 67 70 73 76 79
r102 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r103 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r104 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r106 67 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r107 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r108 64 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.405 $Y=2.72
+ $X2=5.24 $Y2=2.72
r109 64 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.405 $Y=2.72
+ $X2=5.75 $Y2=2.72
r110 63 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r111 63 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r112 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r113 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.4 $Y2=2.72
r114 60 62 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.83 $Y2=2.72
r115 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=2.72
+ $X2=5.24 $Y2=2.72
r116 59 62 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.075 $Y=2.72
+ $X2=4.83 $Y2=2.72
r117 58 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r118 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r120 55 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r121 54 57 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r122 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r123 52 73 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.77 $Y=2.72
+ $X2=2.602 $Y2=2.72
r124 52 54 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.77 $Y=2.72
+ $X2=2.99 $Y2=2.72
r125 51 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.235 $Y=2.72
+ $X2=4.4 $Y2=2.72
r126 51 57 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.235 $Y=2.72
+ $X2=3.91 $Y2=2.72
r127 50 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r128 50 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r129 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r130 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=1.745 $Y2=2.72
r131 47 49 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=2.07 $Y2=2.72
r132 46 73 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.602 $Y2=2.72
r133 46 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 44 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r135 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 40 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r137 38 43 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=2.72 $X2=0.69
+ $Y2=2.72
r138 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=2.72
+ $X2=0.885 $Y2=2.72
r139 34 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=2.635
+ $X2=5.24 $Y2=2.72
r140 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.24 $Y=2.635
+ $X2=5.24 $Y2=2.36
r141 30 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=2.635 $X2=4.4
+ $Y2=2.72
r142 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.4 $Y=2.635
+ $X2=4.4 $Y2=2.36
r143 26 73 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.602 $Y=2.635
+ $X2=2.602 $Y2=2.72
r144 26 28 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=2.602 $Y=2.635
+ $X2=2.602 $Y2=2.36
r145 22 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=2.635
+ $X2=1.745 $Y2=2.72
r146 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.745 $Y=2.635
+ $X2=1.745 $Y2=2.36
r147 21 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.05 $Y=2.72
+ $X2=0.885 $Y2=2.72
r148 20 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=2.72
+ $X2=1.745 $Y2=2.72
r149 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.58 $Y=2.72
+ $X2=1.05 $Y2=2.72
r150 16 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=2.635
+ $X2=0.885 $Y2=2.72
r151 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.885 $Y=2.635
+ $X2=0.885 $Y2=2.36
r152 5 36 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=5.105
+ $Y=1.485 $X2=5.24 $Y2=2.36
r153 4 32 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.485 $X2=4.4 $Y2=2.36
r154 3 28 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.6 $Y2=2.36
r155 2 24 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.485 $X2=1.745 $Y2=2.36
r156 1 18 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.745
+ $Y=1.485 $X2=0.885 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%X 1 2 3 4 13 17 20 24 27 33
r45 30 33 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.315 $Y=1.68
+ $X2=2.175 $Y2=1.68
r46 24 27 3.18761 $w=2.33e-07 $l=6.5e-08 $layer=LI1_cond $X=1.117 $Y=1.595
+ $X2=1.117 $Y2=1.53
r47 20 24 2.95087 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.117 $Y=1.68
+ $X2=1.117 $Y2=1.595
r48 20 30 4.81805 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=1.235 $Y=1.68
+ $X2=1.315 $Y2=1.68
r49 20 27 0.490401 $w=2.33e-07 $l=1e-08 $layer=LI1_cond $X=1.117 $Y=1.52
+ $X2=1.117 $Y2=1.53
r50 19 20 36.0445 $w=2.33e-07 $l=7.35e-07 $layer=LI1_cond $X=1.117 $Y=0.785
+ $X2=1.117 $Y2=1.52
r51 15 17 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.315 $Y=0.7
+ $X2=2.175 $Y2=0.7
r52 13 19 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=1.235 $Y=0.7
+ $X2=1.117 $Y2=0.785
r53 13 15 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.235 $Y=0.7 $X2=1.315
+ $Y2=0.7
r54 4 33 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=1.485 $X2=2.175 $Y2=1.68
r55 3 30 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.485 $X2=1.315 $Y2=1.68
r56 2 17 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.235 $X2=2.175 $Y2=0.7
r57 1 15 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.315 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%A_603_297# 1 2 3 4 15 17 18 21 23 29 32
c53 23 0 1.1533e-19 $X=5.57 $Y=2.02
r54 32 33 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.975 $Y=2.02
+ $X2=3.975 $Y2=2.295
r55 27 29 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=5.697 $Y=1.935
+ $X2=5.697 $Y2=1.63
r56 24 32 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.065 $Y=2.02 $X2=3.975
+ $Y2=2.02
r57 24 26 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.065 $Y=2.02
+ $X2=4.82 $Y2=2.02
r58 23 27 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.57 $Y=2.02
+ $X2=5.697 $Y2=1.935
r59 23 26 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.57 $Y=2.02
+ $X2=4.82 $Y2=2.02
r60 19 32 5.23737 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=1.935
+ $X2=3.975 $Y2=2.02
r61 19 21 20.0253 $w=1.78e-07 $l=3.25e-07 $layer=LI1_cond $X=3.975 $Y=1.935
+ $X2=3.975 $Y2=1.61
r62 17 33 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.885 $Y=2.295
+ $X2=3.975 $Y2=2.295
r63 17 18 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.885 $Y=2.295
+ $X2=3.225 $Y2=2.295
r64 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.14 $Y=2.21
+ $X2=3.225 $Y2=2.295
r65 13 15 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.14 $Y=2.21
+ $X2=3.14 $Y2=1.86
r66 4 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.525
+ $Y=1.485 $X2=5.66 $Y2=1.63
r67 3 26 600 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=1 $X=4.685
+ $Y=1.485 $X2=4.82 $Y2=2.02
r68 2 32 600 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.485 $X2=3.98 $Y2=2.055
r69 2 21 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.485 $X2=3.98 $Y2=1.61
r70 1 15 300 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=2 $X=3.015
+ $Y=1.485 $X2=3.14 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_HD__A21BO_4%VGND 1 2 3 4 5 18 20 24 28 32 34 36 38 39 40
+ 46 55 60 66 68 72
r91 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r92 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r93 65 66 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=0.18
+ $X2=3.285 $Y2=0.18
r94 63 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r95 62 65 2.93378 $w=5.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.99 $Y=0.18
+ $X2=3.12 $Y2=0.18
r96 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r97 59 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r98 58 62 10.3811 $w=5.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=0.18
+ $X2=2.99 $Y2=0.18
r99 58 60 6.31924 $w=5.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.53 $Y=0.18
+ $X2=2.515 $Y2=0.18
r100 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r101 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r102 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r103 53 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r104 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r105 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r106 50 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r107 49 52 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r108 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r109 47 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.02
+ $Y2=0
r110 47 49 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=4.37 $Y2=0
r111 46 71 4.21407 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=5.545 $Y=0
+ $X2=5.762 $Y2=0
r112 46 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=0
+ $X2=5.29 $Y2=0
r113 44 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r114 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r115 40 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r116 38 43 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.69
+ $Y2=0
r117 38 39 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.88
+ $Y2=0
r118 34 71 3.14599 $w=2.8e-07 $l=1.17346e-07 $layer=LI1_cond $X=5.685 $Y=0.085
+ $X2=5.762 $Y2=0
r119 34 36 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.685 $Y=0.085
+ $X2=5.685 $Y2=0.38
r120 30 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r121 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.36
r122 28 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=4.02
+ $Y2=0
r123 28 66 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=3.285 $Y2=0
r124 27 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=1.745
+ $Y2=0
r125 27 60 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.91 $Y=0
+ $X2=2.515 $Y2=0
r126 22 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=0.085
+ $X2=1.745 $Y2=0
r127 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.745 $Y=0.085
+ $X2=1.745 $Y2=0.36
r128 21 39 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=0.88
+ $Y2=0
r129 20 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=1.745
+ $Y2=0
r130 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=1.05
+ $Y2=0
r131 16 39 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=0.085
+ $X2=0.88 $Y2=0
r132 16 18 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=0.88 $Y=0.085
+ $X2=0.88 $Y2=0.36
r133 5 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.525
+ $Y=0.235 $X2=5.66 $Y2=0.38
r134 4 32 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.235 $X2=4.02 $Y2=0.36
r135 3 65 91 $w=1.7e-07 $l=7.14773e-07 $layer=licon1_NDIFF $count=2 $X=2.465
+ $Y=0.235 $X2=3.12 $Y2=0.36
r136 2 24 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.235 $X2=1.745 $Y2=0.36
r137 1 18 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.745
+ $Y=0.235 $X2=0.885 $Y2=0.36
.ends


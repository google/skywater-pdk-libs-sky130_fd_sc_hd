* File: sky130_fd_sc_hd__a211oi_4.spice
* Created: Tue Sep  1 18:51:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a211oi_4.pex.spice"
.subckt sky130_fd_sc_hd__a211oi_4  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_109_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75006.6 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A2_M1018_g N_A_109_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75006.2 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1018_d N_A2_M1025_g N_A_109_47#_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75005.8 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_A1_M1013_g N_A_109_47#_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1013_d N_A1_M1014_g N_A_109_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1020_d N_A1_M1020_g N_A_109_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1024 N_Y_M1020_d N_A1_M1024_g N_A_109_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1030 N_VGND_M1030_d N_A2_M1030_g N_A_109_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.08775 PD=0.985 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1002_d N_B1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.091 PD=0.985 PS=0.93 NRD=7.38 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1023_d N_B1_M1023_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.091 PD=0.925 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1023_d N_C1_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.08775 PD=0.925 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1021 N_Y_M1021_d N_C1_M1021_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1027 N_Y_M1021_d N_C1_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1031 N_Y_M1031_d N_C1_M1031_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.08775 PD=0.93 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75006.1 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1026 N_Y_M1031_d N_B1_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.1885 PD=0.93 PS=1.88 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75006.6 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75006.6 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1001_d N_A2_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75006.2 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A2_M1019_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75005.8 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1019_d N_A1_M1000_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1004_d N_A1_M1022_g N_A_27_297#_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1028 N_VPWR_M1028_d N_A1_M1028_g N_A_27_297#_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1029 N_VPWR_M1028_d N_A2_M1029_g N_A_27_297#_M1029_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1011 N_A_27_297#_M1029_s N_B1_M1011_g N_A_781_297#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1016 N_A_27_297#_M1016_d N_B1_M1016_g N_A_781_297#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1007 N_A_27_297#_M1016_d N_B1_M1007_g A_949_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.15 PD=1.27 PS=1.3 NRD=0 NRS=18.6953 M=1 R=6.66667 SA=75004.4
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1010 A_949_297# N_C1_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.15
+ AS=0.14 PD=1.3 PS=1.28 NRD=18.6953 NRS=0 M=1 R=6.66667 SA=75004.8 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1005 N_A_781_297#_M1005_d N_C1_M1005_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.3
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1017 N_A_781_297#_M1005_d N_C1_M1017_g N_Y_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=3.9203 M=1 R=6.66667 SA=75005.7
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1008 A_1301_297# N_C1_M1008_g N_Y_M1017_s VPB PHIGHVT L=0.15 W=1 AD=0.155
+ AS=0.15 PD=1.31 PS=1.3 NRD=19.6803 NRS=0 M=1 R=6.66667 SA=75006.1 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1012 N_A_27_297#_M1012_d N_B1_M1012_g A_1301_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.155 PD=2.52 PS=1.31 NRD=0 NRS=19.6803 M=1 R=6.66667 SA=75006.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=12.4227 P=18.69
*
.include "sky130_fd_sc_hd__a211oi_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nor3_2.pex.spice
* Created: Thu Aug 27 14:32:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR3_2%A 1 3 6 8 10 13 15 16 24
r40 22 24 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=0.645 $Y=1.16
+ $X2=0.91 $Y2=1.16
r41 19 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.645 $Y2=1.16
r42 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r43 15 16 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.645 $Y2=1.18
r44 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r45 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r46 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r47 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r48 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r49 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r50 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_2%B 1 3 6 8 10 13 15 16 24
r47 22 24 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.525 $Y=1.16
+ $X2=1.75 $Y2=1.16
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.16 $X2=1.525 $Y2=1.16
r49 19 22 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.525 $Y2=1.16
r50 15 16 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=2.075 $Y2=1.18
r51 15 23 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=1.615 $Y=1.18
+ $X2=1.525 $Y2=1.18
r52 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r54 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r56 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325 $X2=1.33
+ $Y2=1.985
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995 $X2=1.33
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_2%C 1 3 6 8 10 13 15 16 24 25 27
c46 16 0 8.40227e-20 $X=2.47 $Y=1.445
r47 23 25 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.8 $Y=1.16 $X2=3.13
+ $Y2=1.16
r48 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=1.16 $X2=2.8 $Y2=1.16
r49 20 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.71 $Y=1.16 $X2=2.8
+ $Y2=1.16
r50 16 27 10.6547 $w=2.63e-07 $l=2.45e-07 $layer=LI1_cond $X=2.507 $Y=1.53
+ $X2=2.507 $Y2=1.285
r51 15 27 3.06002 $w=2.65e-07 $l=1.05e-07 $layer=LI1_cond $X=2.507 $Y=1.18
+ $X2=2.507 $Y2=1.285
r52 15 24 7.14137 $w=3.78e-07 $l=1.6e-07 $layer=LI1_cond $X=2.64 $Y=1.18 $X2=2.8
+ $Y2=1.18
r53 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.13 $Y=1.325
+ $X2=3.13 $Y2=1.16
r54 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.13 $Y=1.325
+ $X2=3.13 $Y2=1.985
r55 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.13 $Y=0.995
+ $X2=3.13 $Y2=1.16
r56 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.13 $Y=0.995
+ $X2=3.13 $Y2=0.56
r57 4 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.325
+ $X2=2.71 $Y2=1.16
r58 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.71 $Y=1.325 $X2=2.71
+ $Y2=1.985
r59 1 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=0.995
+ $X2=2.71 $Y2=1.16
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.71 $Y=0.995 $X2=2.71
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_2%A_27_297# 1 2 3 10 12 14 18 20 27 29
r35 21 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=1.54
+ $X2=1.12 $Y2=1.54
r36 20 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.96 $Y2=1.54
r37 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.245 $Y2=1.54
r38 16 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=1.54
r39 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=2.3
r40 15 25 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r41 14 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=1.12 $Y2=1.54
r42 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=0.405 $Y2=1.54
r43 10 25 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r44 10 12 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r45 3 29 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r46 2 27 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r47 2 18 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r48 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r49 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_2%VPWR 1 6 8 10 20 21 24
r41 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 20 21 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r43 18 21 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 17 20 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 17 18 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 15 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r48 15 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 10 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r50 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r53 4 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r54 4 6 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=1.96
r55 1 6 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_2%A_281_297# 1 2 3 12 14 15 18 20 24 26
c31 20 0 8.40227e-20 $X=3.215 $Y=2.38
r32 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.34 $Y=2.295
+ $X2=3.34 $Y2=1.96
r33 21 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.625 $Y=2.38
+ $X2=2.52 $Y2=2.38
r34 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.215 $Y=2.38
+ $X2=3.34 $Y2=2.295
r35 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.215 $Y=2.38
+ $X2=2.625 $Y2=2.38
r36 16 26 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.295
+ $X2=2.52 $Y2=2.38
r37 16 18 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.52 $Y=2.295
+ $X2=2.52 $Y2=1.96
r38 14 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.415 $Y=2.38
+ $X2=2.52 $Y2=2.38
r39 14 15 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.415 $Y=2.38
+ $X2=1.665 $Y2=2.38
r40 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.54 $Y=2.295
+ $X2=1.665 $Y2=2.38
r41 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=2.295
+ $X2=1.54 $Y2=1.96
r42 3 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.205
+ $Y=1.485 $X2=3.34 $Y2=1.96
r43 2 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=2.375
+ $Y=1.485 $X2=2.5 $Y2=1.96
r44 1 12 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_2%Y 1 2 3 4 15 17 18 21 23 27 31 34 36 42
r75 39 42 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.365 $Y=1.54
+ $X2=2.92 $Y2=1.54
r76 36 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.475 $Y=1.54
+ $X2=3.365 $Y2=1.54
r77 36 39 0.130009 $w=4.58e-07 $l=5e-09 $layer=LI1_cond $X=3.365 $Y=1.45
+ $X2=3.365 $Y2=1.455
r78 34 36 14.1709 $w=4.58e-07 $l=5.45e-07 $layer=LI1_cond $X=3.365 $Y=0.905
+ $X2=3.365 $Y2=1.45
r79 25 34 27.4192 $w=1.78e-07 $l=4.45e-07 $layer=LI1_cond $X=2.92 $Y=0.815
+ $X2=3.365 $Y2=0.815
r80 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.92 $Y=0.725
+ $X2=2.92 $Y2=0.39
r81 24 31 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r82 23 25 10.1667 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0.815
+ $X2=2.92 $Y2=0.815
r83 23 24 64.697 $w=1.78e-07 $l=1.05e-06 $layer=LI1_cond $X=2.755 $Y=0.815
+ $X2=1.705 $Y2=0.815
r84 19 31 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725 $X2=1.54
+ $Y2=0.815
r85 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r86 17 31 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r87 17 18 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r88 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r89 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725 $X2=0.7
+ $Y2=0.39
r90 4 42 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.785
+ $Y=1.485 $X2=2.92 $Y2=1.62
r91 3 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.785
+ $Y=0.235 $X2=2.92 $Y2=0.39
r92 2 21 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r93 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_2%VGND 1 2 3 4 5 16 18 22 24 26 29 30 31 41 51
+ 57 60
r55 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r56 56 57 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=0.235
+ $X2=2.585 $Y2=0.235
r57 53 56 8.03615 $w=6.38e-07 $l=4.3e-07 $layer=LI1_cond $X=2.07 $Y=0.235
+ $X2=2.5 $Y2=0.235
r58 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r59 50 53 2.05576 $w=6.38e-07 $l=1.1e-07 $layer=LI1_cond $X=1.96 $Y=0.235
+ $X2=2.07 $Y2=0.235
r60 50 51 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.235
+ $X2=1.875 $Y2=0.235
r61 45 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r62 45 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r63 44 57 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=2.585
+ $Y2=0
r64 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r65 41 59 4.33193 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.467
+ $Y2=0
r66 41 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r67 40 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r68 39 51 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.875
+ $Y2=0
r69 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r70 36 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r71 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 33 47 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r73 33 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r74 31 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r75 31 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 29 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r77 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r78 28 39 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.61
+ $Y2=0
r79 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r80 24 59 3.10591 $w=2.9e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.4 $Y=0.085
+ $X2=3.467 $Y2=0
r81 24 26 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.4 $Y=0.085
+ $X2=3.4 $Y2=0.39
r82 20 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r83 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r84 16 47 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r85 16 18 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r86 5 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.34 $Y2=0.39
r87 4 56 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.235 $X2=2.5 $Y2=0.39
r88 3 50 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r89 2 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r90 1 18 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


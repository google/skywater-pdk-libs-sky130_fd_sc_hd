* File: sky130_fd_sc_hd__dlrbp_2.spice.pex
* Created: Thu Aug 27 14:17:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRBP_2%GATE 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.235 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%A_27_47# 1 2 9 13 17 19 20 23 27 30 34 35 36
+ 41 44 46 49 50 53 56 57 60 64
c147 57 0 1.8552e-19 $X=2.555 $Y=1.53
c148 13 0 2.6965e-20 $X=0.89 $Y=2.135
c149 9 0 2.6965e-20 $X=0.89 $Y=0.445
r150 57 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r151 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.53
+ $X2=2.555 $Y2=1.53
r152 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r153 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r154 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.53
+ $X2=2.555 $Y2=1.53
r155 49 50 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.41 $Y=1.53
+ $X2=0.84 $Y2=1.53
r156 48 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r157 47 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r158 45 64 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r159 44 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r160 44 46 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r161 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r162 38 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r163 37 41 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r164 36 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r165 36 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r166 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r167 34 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r168 28 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r169 28 30 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r170 26 60 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r171 26 27 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r172 25 60 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r173 21 23 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.22 $Y=1.245
+ $X2=3.22 $Y2=0.415
r174 20 25 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r175 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=3.22 $Y2=1.245
r176 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=2.805 $Y2=1.32
r177 17 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.73 $Y=2.275
+ $X2=2.73 $Y2=1.685
r178 11 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r179 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r180 7 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r181 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r182 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r183 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%A_299_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c86 32 0 1.12109e-19 $X=2.255 $Y=0.93
c87 18 0 7.13094e-20 $X=1.97 $Y=0.7
r88 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=1.095
r89 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=0.765
r90 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r91 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r92 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.155 $Y2=0.93
r93 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.055 $Y2=1.495
r94 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=2.055 $Y2=1.495
r95 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=1.785 $Y2=1.58
r96 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r97 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=2.155 $Y2=0.93
r98 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=1.705 $Y2=0.7
r99 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r100 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r101 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=2.165
+ $X2=2.25 $Y2=1.095
r102 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.765
r103 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r104 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%A_193_47# 1 2 9 12 16 19 20 24 26 28 29 32
+ 35 39 42 43
c125 42 0 2.54761e-19 $X=3.18 $Y=1.74
c126 19 0 2.83694e-19 $X=3.01 $Y=1.575
r127 42 45 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.18 $Y2=1.875
r128 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r129 35 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.87
+ $X2=3.015 $Y2=1.87
r130 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r131 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r132 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.87
+ $X2=3.015 $Y2=1.87
r133 28 29 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=2.87 $Y=1.87
+ $X2=1.3 $Y2=1.87
r134 24 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=0.87
+ $X2=2.8 $Y2=0.705
r135 23 26 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=0.87
+ $X2=3.01 $Y2=0.87
r136 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=0.87 $X2=2.8 $Y2=0.87
r137 20 32 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r138 20 21 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r139 19 43 8.96365 $w=3.1e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.01 $Y=1.575
+ $X2=3.095 $Y2=1.74
r140 18 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=0.87
r141 18 19 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=1.575
r142 16 21 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r143 12 45 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.15 $Y=2.275
+ $X2=3.15 $Y2=1.875
r144 9 39 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.79 $Y=0.415
+ $X2=2.79 $Y2=0.705
r145 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r146 1 16 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%A_711_307# 1 2 9 13 15 17 20 22 24 27 29 30
+ 33 37 39 40 43 45 49 51 56 58 63 65 67
c146 65 0 1.13195e-19 $X=5.535 $Y=1.16
c147 43 0 1.91094e-19 $X=3.925 $Y=1.7
c148 39 0 1.02435e-19 $X=6.915 $Y=1.16
c149 30 0 2.69497e-19 $X=6.05 $Y=1.16
c150 13 0 2.1991e-19 $X=3.695 $Y=0.445
r151 69 71 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.63 $Y=1.7
+ $X2=3.695 $Y2=1.7
r152 66 76 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=5.535 $Y=1.16
+ $X2=5.975 $Y2=1.16
r153 65 68 7.88116 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.47 $Y=1.16
+ $X2=5.47 $Y2=1.325
r154 65 67 7.88116 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.47 $Y=1.16
+ $X2=5.47 $Y2=0.995
r155 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.535
+ $Y=1.16 $X2=5.535 $Y2=1.16
r156 58 60 6.14636 $w=2.98e-07 $l=1.6e-07 $layer=LI1_cond $X=4.42 $Y=0.58
+ $X2=4.42 $Y2=0.74
r157 56 68 12.2584 $w=1.88e-07 $l=2.1e-07 $layer=LI1_cond $X=5.415 $Y=1.535
+ $X2=5.415 $Y2=1.325
r158 53 67 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5.415 $Y=0.825
+ $X2=5.415 $Y2=0.995
r159 52 63 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.94 $Y=1.62
+ $X2=4.855 $Y2=1.7
r160 51 56 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.32 $Y=1.62
+ $X2=5.415 $Y2=1.535
r161 51 52 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.32 $Y=1.62
+ $X2=4.94 $Y2=1.62
r162 47 63 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=1.865
+ $X2=4.855 $Y2=1.7
r163 47 49 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.855 $Y=1.865
+ $X2=4.855 $Y2=2.27
r164 46 60 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.57 $Y=0.74 $X2=4.42
+ $Y2=0.74
r165 45 53 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.32 $Y=0.74
+ $X2=5.415 $Y2=0.825
r166 45 46 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.32 $Y=0.74
+ $X2=4.57 $Y2=0.74
r167 43 71 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.695 $Y2=1.7
r168 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r169 40 63 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=1.7
+ $X2=4.855 $Y2=1.7
r170 40 42 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=4.77 $Y=1.7
+ $X2=3.925 $Y2=1.7
r171 35 39 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.915 $Y=1.325
+ $X2=6.915 $Y2=1.16
r172 35 37 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.915 $Y=1.325
+ $X2=6.915 $Y2=2.165
r173 31 39 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.915 $Y=0.995
+ $X2=6.915 $Y2=1.16
r174 31 33 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.915 $Y=0.995
+ $X2=6.915 $Y2=0.445
r175 30 76 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.05 $Y=1.16
+ $X2=5.975 $Y2=1.16
r176 29 39 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.84 $Y=1.16
+ $X2=6.915 $Y2=1.16
r177 29 30 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=6.84 $Y=1.16
+ $X2=6.05 $Y2=1.16
r178 25 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.975 $Y=1.325
+ $X2=5.975 $Y2=1.16
r179 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.975 $Y=1.325
+ $X2=5.975 $Y2=1.985
r180 22 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.975 $Y=0.995
+ $X2=5.975 $Y2=1.16
r181 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.975 $Y=0.995
+ $X2=5.975 $Y2=0.56
r182 18 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.325
+ $X2=5.535 $Y2=1.16
r183 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.535 $Y=1.325
+ $X2=5.535 $Y2=1.985
r184 15 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=0.995
+ $X2=5.535 $Y2=1.16
r185 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.535 $Y=0.995
+ $X2=5.535 $Y2=0.56
r186 11 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=1.7
r187 11 13 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=0.445
r188 7 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=1.7
r189 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.63 $Y=1.865
+ $X2=3.63 $Y2=2.275
r190 2 63 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.855 $Y2=1.755
r191 2 49 600 $w=1.7e-07 $l=8.5443e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.855 $Y2=2.27
r192 1 58 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.235 $X2=4.425 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%A_561_413# 1 2 7 9 12 14 15 16 20 25 27 30
+ 34
c82 34 0 1.54137e-19 $X=3.33 $Y=0.995
c83 16 0 2.87957e-19 $X=3.27 $Y=2.34
r84 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.16 $X2=4.115 $Y2=1.16
r85 28 34 0.89609 $w=3.3e-07 $l=3.47851e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=3.33 $Y2=0.995
r86 28 30 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=4.115 $Y2=1.16
r87 27 33 18.4264 $w=2.8e-07 $l=4.19452e-07 $layer=LI1_cond $X=3.52 $Y=1.96
+ $X2=3.437 $Y2=2.34
r88 26 34 8.61065 $w=1.7e-07 $l=4.14246e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.33 $Y2=0.995
r89 26 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.96
r90 25 34 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=0.995
+ $X2=3.33 $Y2=0.995
r91 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=0.995
r92 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r93 20 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.005 $Y2=0.45
r94 16 33 3.65648 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.27 $Y=2.34
+ $X2=3.437 $Y2=2.34
r95 16 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.27 $Y=2.34
+ $X2=2.94 $Y2=2.34
r96 14 31 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.115 $Y2=1.16
r97 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.635 $Y2=1.16
r98 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=1.325
+ $X2=4.635 $Y2=1.16
r99 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.635 $Y=1.325
+ $X2=4.635 $Y2=1.985
r100 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=0.995
+ $X2=4.635 $Y2=1.16
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.635 $Y=0.995
+ $X2=4.635 $Y2=0.56
r102 2 18 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.065 $X2=2.94 $Y2=2.34
r103 1 22 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3.005 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%RESET_B 3 6 8 11 12 13
c37 12 0 1.27311e-19 $X=5.055 $Y=1.16
r38 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.16
+ $X2=5.055 $Y2=1.325
r39 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.16
+ $X2=5.055 $Y2=0.995
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.16 $X2=5.055 $Y2=1.16
r41 8 12 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.885 $Y=1.16
+ $X2=5.055 $Y2=1.16
r42 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.065 $Y=1.985
+ $X2=5.065 $Y2=1.325
r43 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.065 $Y=0.56
+ $X2=5.065 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%A_1316_47# 1 2 7 9 12 14 16 20 24 28 32 35
r69 33 37 8.25342 $w=2.92e-07 $l=5e-08 $layer=POLY_cond $X=7.34 $Y=1.16 $X2=7.39
+ $Y2=1.16
r70 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.16 $X2=7.34 $Y2=1.16
r71 30 35 1.36975 $w=3.3e-07 $l=1.68e-07 $layer=LI1_cond $X=6.87 $Y=1.16
+ $X2=6.702 $Y2=1.16
r72 30 32 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=6.87 $Y=1.16
+ $X2=7.34 $Y2=1.16
r73 26 35 5.13366 $w=3.32e-07 $l=1.65e-07 $layer=LI1_cond $X=6.702 $Y=1.325
+ $X2=6.702 $Y2=1.16
r74 26 28 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=6.702 $Y=1.325
+ $X2=6.702 $Y2=2
r75 22 35 5.13366 $w=3.32e-07 $l=1.65997e-07 $layer=LI1_cond $X=6.7 $Y=0.995
+ $X2=6.702 $Y2=1.16
r76 22 24 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=6.7 $Y=0.995
+ $X2=6.7 $Y2=0.51
r77 14 37 69.3288 $w=2.92e-07 $l=4.2e-07 $layer=POLY_cond $X=7.81 $Y=1.16
+ $X2=7.39 $Y2=1.16
r78 14 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.81 $Y=1.295
+ $X2=7.81 $Y2=1.985
r79 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.81 $Y=1.025
+ $X2=7.81 $Y2=0.56
r80 10 37 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=1.325
+ $X2=7.39 $Y2=1.16
r81 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.39 $Y=1.325
+ $X2=7.39 $Y2=1.985
r82 7 37 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=0.995
+ $X2=7.39 $Y2=1.16
r83 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.39 $Y=0.995 $X2=7.39
+ $Y2=0.56
r84 2 28 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=6.58
+ $Y=1.845 $X2=6.705 $Y2=2
r85 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.235 $X2=6.705 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 45 47 51
+ 53 58 71 76 81 86 92 95 99 105 107 110 113 117
c129 35 0 1.30285e-19 $X=5.275 $Y=2.02
r130 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r131 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r132 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r133 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 104 105 10.7902 $w=6.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.425 $Y=2.47
+ $X2=4.6 $Y2=2.47
r135 101 104 0.981855 $w=6.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.37 $Y=2.47
+ $X2=4.425 $Y2=2.47
r136 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r137 98 101 9.46152 $w=6.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.84 $Y=2.47
+ $X2=4.37 $Y2=2.47
r138 98 99 9.18355 $w=6.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=2.47
+ $X2=3.755 $Y2=2.47
r139 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r140 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r141 90 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r142 90 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r143 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r144 87 113 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.192 $Y2=2.72
r145 87 89 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.59 $Y2=2.72
r146 86 116 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=7.935 $Y=2.72
+ $X2=8.107 $Y2=2.72
r147 86 89 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=2.72
+ $X2=7.59 $Y2=2.72
r148 85 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r149 85 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r150 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r151 82 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.23 $Y2=2.72
r152 82 84 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.67 $Y2=2.72
r153 81 113 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.045 $Y=2.72
+ $X2=7.192 $Y2=2.72
r154 81 84 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.045 $Y=2.72
+ $X2=6.67 $Y2=2.72
r155 80 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r156 80 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r157 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r158 77 107 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.49 $Y=2.72
+ $X2=5.3 $Y2=2.72
r159 77 79 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.49 $Y=2.72
+ $X2=5.75 $Y2=2.72
r160 76 110 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.1 $Y=2.72
+ $X2=6.23 $Y2=2.72
r161 76 79 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.1 $Y=2.72
+ $X2=5.75 $Y2=2.72
r162 75 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r163 75 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r164 74 105 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=4.6 $Y2=2.72
r165 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r166 71 107 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.11 $Y=2.72
+ $X2=5.3 $Y2=2.72
r167 71 74 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.11 $Y=2.72
+ $X2=4.83 $Y2=2.72
r168 70 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r169 69 99 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.755 $Y2=2.72
r170 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r171 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r172 67 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r173 66 69 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r174 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r175 64 95 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r176 64 66 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r177 62 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r178 62 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r179 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r180 59 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r181 59 61 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r182 58 95 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r183 58 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r184 53 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r185 53 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r186 51 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r187 51 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r188 47 50 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=8.065 $Y=1.66
+ $X2=8.065 $Y2=2.34
r189 45 116 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=8.065 $Y=2.635
+ $X2=8.107 $Y2=2.72
r190 45 50 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=8.065 $Y=2.635
+ $X2=8.065 $Y2=2.34
r191 41 113 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.192 $Y=2.635
+ $X2=7.192 $Y2=2.72
r192 41 43 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=7.192 $Y=2.635
+ $X2=7.192 $Y2=2
r193 37 110 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.23 $Y=2.635
+ $X2=6.23 $Y2=2.72
r194 37 39 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=6.23 $Y=2.635
+ $X2=6.23 $Y2=2
r195 33 107 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.72
r196 33 35 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.02
r197 29 95 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r198 29 31 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r199 25 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r200 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r201 8 50 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=2.34
r202 8 47 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=1.66
r203 7 43 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=6.99
+ $Y=1.845 $X2=7.175 $Y2=2
r204 6 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.05
+ $Y=1.485 $X2=6.185 $Y2=2
r205 5 35 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=5.14
+ $Y=1.485 $X2=5.275 $Y2=2.02
r206 4 104 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.485 $X2=4.425 $Y2=2.34
r207 3 98 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.705
+ $Y=2.065 $X2=3.84 $Y2=2.3
r208 2 31 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r209 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%Q 1 2 7 10 11 12 13 14 24
r39 14 18 18.2037 $w=5.28e-07 $l=6.39922e-07 $layer=LI1_cond $X=6.02 $Y=1.19
+ $X2=5.765 $Y2=0.665
r40 13 24 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.805 $Y=2.21
+ $X2=5.805 $Y2=1.96
r41 12 18 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.765 $Y=0.51
+ $X2=5.765 $Y2=0.665
r42 11 24 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=5.805 $Y=1.66
+ $X2=5.805 $Y2=1.96
r43 10 11 7.03284 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=5.872 $Y=1.495
+ $X2=5.872 $Y2=1.66
r44 7 14 5.90853 $w=5.28e-07 $l=1.75442e-07 $layer=LI1_cond $X=5.927 $Y=1.325
+ $X2=6.02 $Y2=1.19
r45 7 10 7.12419 $w=2.73e-07 $l=1.7e-07 $layer=LI1_cond $X=5.927 $Y=1.325
+ $X2=5.927 $Y2=1.495
r46 2 24 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=5.61
+ $Y=1.485 $X2=5.765 $Y2=1.96
r47 1 12 182 $w=1.7e-07 $l=4.15331e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.235 $X2=5.765 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%Q_N 1 2 8 12 13 14 16 17 18 19 20 36
c29 16 0 2.65541e-19 $X=7.68 $Y=1.19
c30 8 0 1.13751e-20 $X=7.68 $Y=1.055
r31 20 36 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=8.08 $Y=1.19 $X2=8.05
+ $Y2=1.19
r32 18 19 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=7.64 $Y=1.82
+ $X2=7.64 $Y2=2.21
r33 15 36 12.1647 $w=2.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.765 $Y=1.19
+ $X2=8.05 $Y2=1.19
r34 15 16 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.765 $Y=1.19
+ $X2=7.68 $Y2=1.19
r35 13 18 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.64 $Y=1.73 $X2=7.64
+ $Y2=1.82
r36 13 14 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.64 $Y=1.73
+ $X2=7.64 $Y2=1.605
r37 11 17 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=7.64 $Y=0.7 $X2=7.64
+ $Y2=0.51
r38 11 12 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.64 $Y=0.7
+ $X2=7.64 $Y2=0.825
r39 9 16 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.68 $Y=1.325
+ $X2=7.68 $Y2=1.19
r40 9 14 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.68 $Y=1.325
+ $X2=7.68 $Y2=1.605
r41 8 16 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.68 $Y=1.055
+ $X2=7.68 $Y2=1.19
r42 8 12 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.68 $Y=1.055
+ $X2=7.68 $Y2=0.825
r43 2 18 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=7.465
+ $Y=1.485 $X2=7.6 $Y2=1.82
r44 1 17 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=7.465
+ $Y=0.235 $X2=7.6 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 50 52 57 62 70 75 80 85 91 94 97 100 103 106 110
c138 110 0 2.71124e-20 $X=8.05 $Y=0
c139 36 0 1.39212e-19 $X=5.275 $Y=0.36
c140 2 0 7.13094e-20 $X=1.905 $Y=0.235
r141 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r142 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r143 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r144 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r145 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r146 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r147 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r148 89 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r149 89 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r150 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r151 86 106 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.34 $Y=0
+ $X2=7.187 $Y2=0
r152 86 88 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.34 $Y=0 $X2=7.59
+ $Y2=0
r153 85 109 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=7.935 $Y=0
+ $X2=8.107 $Y2=0
r154 85 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=0 $X2=7.59
+ $Y2=0
r155 84 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r156 84 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r157 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r158 81 103 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.19
+ $Y2=0
r159 81 83 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.67
+ $Y2=0
r160 80 106 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.035 $Y=0
+ $X2=7.187 $Y2=0
r161 80 83 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.035 $Y=0
+ $X2=6.67 $Y2=0
r162 79 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r163 79 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r164 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r165 76 100 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.49 $Y=0 $X2=5.3
+ $Y2=0
r166 76 78 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.49 $Y=0 $X2=5.75
+ $Y2=0
r167 75 103 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.02 $Y=0 $X2=6.19
+ $Y2=0
r168 75 78 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.02 $Y=0 $X2=5.75
+ $Y2=0
r169 74 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r170 74 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r171 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r172 71 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.905
+ $Y2=0
r173 71 73 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.83
+ $Y2=0
r174 70 100 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=5.3
+ $Y2=0
r175 70 73 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=4.83
+ $Y2=0
r176 69 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r177 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r178 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r179 66 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r180 65 68 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r181 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r182 63 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r183 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r184 62 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.905
+ $Y2=0
r185 62 68 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.45
+ $Y2=0
r186 61 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r187 61 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r188 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r189 58 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r190 58 60 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r191 57 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r192 57 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r193 52 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r194 52 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r195 50 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r196 50 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r197 46 109 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=8.065 $Y=0.085
+ $X2=8.107 $Y2=0
r198 46 48 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=8.065 $Y=0.085
+ $X2=8.065 $Y2=0.38
r199 42 106 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.187 $Y=0.085
+ $X2=7.187 $Y2=0
r200 42 44 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=7.187 $Y=0.085
+ $X2=7.187 $Y2=0.38
r201 38 103 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0
r202 38 40 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0.38
r203 34 100 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0
r204 34 36 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0.36
r205 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0
r206 30 32 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0.445
r207 26 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r208 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r209 22 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r210 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r211 7 48 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.38
r212 6 44 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.99
+ $Y=0.235 $X2=7.175 $Y2=0.38
r213 5 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.05
+ $Y=0.235 $X2=6.185 $Y2=0.38
r214 4 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.14
+ $Y=0.235 $X2=5.275 $Y2=0.36
r215 3 32 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.235 $X2=3.905 $Y2=0.445
r216 2 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r217 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__dlclkp_4.pex.spice
* Created: Tue Sep  1 19:04:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%CLK 4 5 7 8 10 13 15 17 20 24 26 27 30 31
+ 37 41 43 46 47
c131 46 0 9.51314e-20 $X=5.575 $Y=1.16
c132 37 0 6.14555e-20 $X=5.315 $Y=1.19
c133 26 0 6.52821e-20 $X=0.235 $Y=1.19
c134 20 0 2.71124e-20 $X=0.47 $Y=0.805
c135 15 0 1.57241e-19 $X=5.575 $Y=0.995
r136 46 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.16
+ $X2=5.575 $Y2=1.325
r137 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.575
+ $Y=1.16 $X2=5.575 $Y2=1.16
r138 41 44 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r139 41 43 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r140 38 47 11.0976 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.315 $Y=1.19
+ $X2=5.575 $Y2=1.19
r141 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.315 $Y=1.19
+ $X2=5.315 $Y2=1.19
r142 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.38 $Y=1.19
+ $X2=0.235 $Y2=1.19
r143 30 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.17 $Y=1.19
+ $X2=5.315 $Y2=1.19
r144 30 31 5.92821 $w=1.4e-07 $l=4.79e-06 $layer=MET1_cond $X=5.17 $Y=1.19
+ $X2=0.38 $Y2=1.19
r145 26 27 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.21 $Y=1.19
+ $X2=0.21 $Y2=1.53
r146 26 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r147 26 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=1.19
+ $X2=0.235 $Y2=1.19
r148 22 24 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r149 18 20 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r150 15 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=0.995
+ $X2=5.575 $Y2=1.16
r151 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.575 $Y=0.995
+ $X2=5.575 $Y2=0.56
r152 13 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.515 $Y=1.985
+ $X2=5.515 $Y2=1.325
r153 8 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=1.665
r154 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r155 5 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.47 $Y2=0.805
r156 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r157 4 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r158 4 44 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r159 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r160 1 43 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%A_27_47# 1 2 9 13 17 20 24 28 29 30 35 36
+ 39 41 43 45 49 51 54 57 58 64 69 72 76 81
c191 76 0 7.61476e-20 $X=2.85 $Y=1.74
c192 51 0 2.78233e-20 $X=2.65 $Y=0.87
c193 35 0 1.2348e-19 $X=0.695 $Y=1.795
c194 30 0 3.29888e-20 $X=0.61 $Y=1.88
c195 13 0 2.69707e-20 $X=0.89 $Y=2.135
c196 9 0 3.83113e-20 $X=0.89 $Y=0.445
r197 65 81 5.07737 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=1.905
+ $X2=1.695 $Y2=1.905
r198 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.87
+ $X2=1.61 $Y2=1.87
r199 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.87
+ $X2=0.695 $Y2=1.87
r200 58 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.87
+ $X2=0.695 $Y2=1.87
r201 57 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.465 $Y=1.87
+ $X2=1.61 $Y2=1.87
r202 57 58 0.773513 $w=1.4e-07 $l=6.25e-07 $layer=MET1_cond $X=1.465 $Y=1.87
+ $X2=0.84 $Y2=1.87
r203 55 76 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.76 $Y=1.74 $X2=2.85
+ $Y2=1.74
r204 54 56 7.87097 $w=3.1e-07 $l=2e-07 $layer=LI1_cond $X=2.675 $Y=1.74
+ $X2=2.675 $Y2=1.94
r205 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=1.74 $X2=2.76 $Y2=1.74
r206 49 72 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.377 $Y=0.87
+ $X2=2.377 $Y2=0.705
r207 48 51 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.38 $Y=0.87
+ $X2=2.65 $Y2=0.87
r208 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=0.87 $X2=2.38 $Y2=0.87
r209 44 69 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r210 43 46 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r211 43 45 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r212 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r213 39 54 8.96365 $w=3.1e-07 $l=1.77059e-07 $layer=LI1_cond $X=2.65 $Y=1.575
+ $X2=2.675 $Y2=1.74
r214 38 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=1.035
+ $X2=2.65 $Y2=0.87
r215 38 39 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.65 $Y=1.035
+ $X2=2.65 $Y2=1.575
r216 36 56 4.25403 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.505 $Y=1.94
+ $X2=2.675 $Y2=1.94
r217 36 81 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.505 $Y=1.94
+ $X2=1.695 $Y2=1.94
r218 35 61 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.88
r219 35 46 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.4
r220 32 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r221 31 41 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r222 30 61 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.88
r223 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r224 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r225 28 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r226 22 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r227 22 24 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r228 18 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.85 $Y=1.875
+ $X2=2.85 $Y2=1.74
r229 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.85 $Y=1.875
+ $X2=2.85 $Y2=2.275
r230 17 72 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.365 $Y=0.415
+ $X2=2.365 $Y2=0.705
r231 11 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r232 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r233 7 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r234 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r235 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r236 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%GATE 1 3 4 6 8 12
r44 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.785
+ $Y=0.93 $X2=1.785 $Y2=0.93
r45 8 12 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.615 $Y=0.89
+ $X2=1.785 $Y2=0.89
r46 4 11 38.5938 $w=3.29e-07 $l=1.86145e-07 $layer=POLY_cond $X=1.83 $Y=1.095
+ $X2=1.785 $Y2=0.93
r47 4 6 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.83 $Y=1.095 $X2=1.83
+ $Y2=2.165
r48 1 11 39.3263 $w=3.29e-07 $l=1.91181e-07 $layer=POLY_cond $X=1.83 $Y=0.76
+ $X2=1.785 $Y2=0.93
r49 1 3 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.83 $Y=0.76 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%A_193_47# 1 2 9 11 12 15 19 22 26 30 32 33
+ 34
c96 32 0 7.61476e-20 $X=2.25 $Y=1.52
r97 32 34 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.25 $Y=1.52
+ $X2=2.045 $Y2=1.52
r98 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.52 $X2=2.25 $Y2=1.52
r99 29 30 1.57103 $w=2.3e-07 $l=1.33e-07 $layer=LI1_cond $X=1.28 $Y=1.47
+ $X2=1.147 $Y2=1.47
r100 29 34 38.3313 $w=2.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.28 $Y=1.47
+ $X2=2.045 $Y2=1.47
r101 24 30 4.89986 $w=2.45e-07 $l=1.24599e-07 $layer=LI1_cond $X=1.127 $Y=1.585
+ $X2=1.147 $Y2=1.47
r102 24 26 19.2074 $w=2.23e-07 $l=3.75e-07 $layer=LI1_cond $X=1.127 $Y=1.585
+ $X2=1.127 $Y2=1.96
r103 20 30 4.89986 $w=2.45e-07 $l=1.15e-07 $layer=LI1_cond $X=1.147 $Y=1.355
+ $X2=1.147 $Y2=1.47
r104 20 22 36.7477 $w=2.63e-07 $l=8.45e-07 $layer=LI1_cond $X=1.147 $Y=1.355
+ $X2=1.147 $Y2=0.51
r105 18 33 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.25 $Y=1.55 $X2=2.25
+ $Y2=1.52
r106 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.55
+ $X2=2.25 $Y2=1.685
r107 17 33 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.25 $Y=1.395
+ $X2=2.25 $Y2=1.52
r108 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.8 $Y=1.245
+ $X2=2.8 $Y2=0.415
r109 12 17 29.8935 $w=1.5e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.385 $Y=1.32
+ $X2=2.25 $Y2=1.395
r110 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.725 $Y=1.32
+ $X2=2.8 $Y2=1.245
r111 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.725 $Y=1.32
+ $X2=2.385 $Y2=1.32
r112 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.31 $Y=2.275
+ $X2=2.31 $Y2=1.685
r113 2 26 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r114 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%A_627_153# 1 2 8 11 15 16 18 20 22 24 25 26
+ 27 30 34 37 39 42 46 50 51
c107 8 0 2.78233e-20 $X=3.21 $Y=1.535
r108 46 48 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0.58
+ $X2=4.005 $Y2=0.745
r109 43 56 23.3527 $w=2.58e-07 $l=1.25e-07 $layer=POLY_cond $X=4.635 $Y=1.16
+ $X2=4.635 $Y2=1.035
r110 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.16 $X2=4.635 $Y2=1.16
r111 40 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=1.16
+ $X2=4.03 $Y2=1.16
r112 40 42 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.115 $Y=1.16
+ $X2=4.635 $Y2=1.16
r113 39 50 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.03 $Y=1.535
+ $X2=4.005 $Y2=1.7
r114 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=1.325
+ $X2=4.03 $Y2=1.16
r115 38 39 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.03 $Y=1.325
+ $X2=4.03 $Y2=1.535
r116 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=1.16
r117 37 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=0.745
r118 32 50 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=1.865
+ $X2=4.005 $Y2=1.7
r119 32 34 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.005 $Y=1.865
+ $X2=4.005 $Y2=2.27
r120 30 52 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.44 $Y=1.7
+ $X2=3.21 $Y2=1.7
r121 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.7 $X2=3.44 $Y2=1.7
r122 27 50 0.463323 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.895 $Y=1.7
+ $X2=4.005 $Y2=1.7
r123 27 29 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.895 $Y=1.7
+ $X2=3.44 $Y2=1.7
r124 25 26 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=3.242 $Y=0.765
+ $X2=3.242 $Y2=0.915
r125 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.155 $Y=0.96
+ $X2=5.155 $Y2=0.56
r126 21 56 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.035
+ $X2=4.635 $Y2=1.035
r127 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.08 $Y=1.035
+ $X2=5.155 $Y2=0.96
r128 20 21 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=5.08 $Y=1.035
+ $X2=4.77 $Y2=1.035
r129 16 43 39.2009 $w=2.58e-07 $l=1.90526e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.635 $Y2=1.16
r130 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.69 $Y2=1.985
r131 15 25 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.275 $Y=0.445
+ $X2=3.275 $Y2=0.765
r132 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.865
+ $X2=3.21 $Y2=1.7
r133 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.21 $Y=1.865
+ $X2=3.21 $Y2=2.275
r134 8 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.535
+ $X2=3.21 $Y2=1.7
r135 8 26 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.21 $Y=1.535
+ $X2=3.21 $Y2=0.915
r136 2 50 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.485 $X2=3.98 $Y2=1.755
r137 2 34 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.485 $X2=3.98 $Y2=2.27
r138 1 46 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=3.88
+ $Y=0.235 $X2=4.005 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%A_477_413# 1 2 9 11 13 14 15 16 20 25 27 30
+ 33
c92 33 0 1.43275e-19 $X=2.905 $Y=0.995
c93 15 0 4.38576e-20 $X=4.202 $Y=1.16
r94 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.69
+ $Y=1.16 $X2=3.69 $Y2=1.16
r95 28 33 0.89609 $w=3.3e-07 $l=3.52987e-07 $layer=LI1_cond $X=3.185 $Y=1.16
+ $X2=2.905 $Y2=0.995
r96 28 30 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=3.185 $Y=1.16
+ $X2=3.69 $Y2=1.16
r97 27 34 15.7666 $w=2.47e-07 $l=3.19022e-07 $layer=LI1_cond $X=3.1 $Y=2.015
+ $X2=3.05 $Y2=2.31
r98 26 33 8.61065 $w=1.7e-07 $l=4.16233e-07 $layer=LI1_cond $X=3.1 $Y=1.325
+ $X2=2.905 $Y2=0.995
r99 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.1 $Y=1.325 $X2=3.1
+ $Y2=2.015
r100 25 33 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=0.995
+ $X2=2.905 $Y2=0.995
r101 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.99 $Y=0.535
+ $X2=2.99 $Y2=0.995
r102 20 34 1.1476 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.915 $Y=2.31
+ $X2=3.05 $Y2=2.31
r103 20 22 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=2.31
+ $X2=2.64 $Y2=2.31
r104 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=0.45
+ $X2=2.99 $Y2=0.535
r105 16 18 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.905 $Y=0.45
+ $X2=2.58 $Y2=0.45
r106 14 31 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=4.115 $Y=1.16
+ $X2=3.69 $Y2=1.16
r107 14 15 5.03009 $w=3.3e-07 $l=8.7e-08 $layer=POLY_cond $X=4.115 $Y=1.16
+ $X2=4.202 $Y2=1.16
r108 11 15 37.0704 $w=1.5e-07 $l=1.71377e-07 $layer=POLY_cond $X=4.215 $Y=0.995
+ $X2=4.202 $Y2=1.16
r109 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.215 $Y=0.995
+ $X2=4.215 $Y2=0.56
r110 7 15 37.0704 $w=1.5e-07 $l=1.70895e-07 $layer=POLY_cond $X=4.19 $Y=1.325
+ $X2=4.202 $Y2=1.16
r111 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.19 $Y=1.325
+ $X2=4.19 $Y2=1.985
r112 2 22 600 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=2.065 $X2=2.64 $Y2=2.28
r113 1 18 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.235 $X2=2.58 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%A_953_297# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 36 37 40 44 48 51 52 54 57 59 62 65 67 68
c153 59 0 3.72061e-19 $X=6.025 $Y=1.495
c154 51 0 2.01098e-19 $X=4.975 $Y=1.495
c155 40 0 1.95136e-19 $X=7.345 $Y=1.16
r156 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.415
+ $Y=1.16 $X2=6.415 $Y2=1.16
r157 60 68 1.10616 $w=2.35e-07 $l=1.15e-07 $layer=LI1_cond $X=6.14 $Y=1.172
+ $X2=6.025 $Y2=1.172
r158 60 62 13.486 $w=2.33e-07 $l=2.75e-07 $layer=LI1_cond $X=6.14 $Y=1.172
+ $X2=6.415 $Y2=1.172
r159 58 68 5.4556 $w=2.2e-07 $l=1.18e-07 $layer=LI1_cond $X=6.025 $Y=1.29
+ $X2=6.025 $Y2=1.172
r160 58 59 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.025 $Y=1.29
+ $X2=6.025 $Y2=1.495
r161 57 68 5.4556 $w=2.2e-07 $l=1.21897e-07 $layer=LI1_cond $X=6.015 $Y=1.055
+ $X2=6.025 $Y2=1.172
r162 56 57 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=6.015 $Y=0.885
+ $X2=6.015 $Y2=1.055
r163 55 67 2.40986 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.06 $Y=1.58
+ $X2=4.905 $Y2=1.58
r164 54 59 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.91 $Y=1.58
+ $X2=6.025 $Y2=1.495
r165 54 55 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=5.91 $Y=1.58
+ $X2=5.06 $Y2=1.58
r166 53 65 2.60907 $w=1.7e-07 $l=3.49929e-07 $layer=LI1_cond $X=5.06 $Y=0.8
+ $X2=4.75 $Y2=0.715
r167 52 56 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.91 $Y=0.8
+ $X2=6.015 $Y2=0.885
r168 52 53 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=5.91 $Y=0.8
+ $X2=5.06 $Y2=0.8
r169 51 67 4.02809 $w=2.27e-07 $l=1.14782e-07 $layer=LI1_cond $X=4.975 $Y=1.495
+ $X2=4.905 $Y2=1.58
r170 50 65 3.84343 $w=2.4e-07 $l=2.98119e-07 $layer=LI1_cond $X=4.975 $Y=0.885
+ $X2=4.75 $Y2=0.715
r171 50 51 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.975 $Y=0.885
+ $X2=4.975 $Y2=1.495
r172 46 67 4.02809 $w=2.27e-07 $l=9.12688e-08 $layer=LI1_cond $X=4.892 $Y=1.665
+ $X2=4.905 $Y2=1.58
r173 46 48 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=4.892 $Y=1.665
+ $X2=4.892 $Y2=2.3
r174 42 65 3.84343 $w=2.4e-07 $l=1.55e-07 $layer=LI1_cond $X=4.905 $Y=0.715
+ $X2=4.75 $Y2=0.715
r175 42 44 9.66565 $w=3.08e-07 $l=2.6e-07 $layer=LI1_cond $X=4.905 $Y=0.715
+ $X2=4.905 $Y2=0.455
r176 39 40 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.925 $Y=1.16
+ $X2=7.345 $Y2=1.16
r177 38 39 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.505 $Y=1.16
+ $X2=6.925 $Y2=1.16
r178 37 63 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.43 $Y=1.16
+ $X2=6.415 $Y2=1.16
r179 37 38 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.43 $Y=1.16
+ $X2=6.505 $Y2=1.16
r180 35 63 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=6.07 $Y=1.16
+ $X2=6.415 $Y2=1.16
r181 35 36 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.07 $Y=1.16
+ $X2=5.995 $Y2=1.16
r182 31 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=1.325
+ $X2=7.345 $Y2=1.16
r183 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.345 $Y=1.325
+ $X2=7.345 $Y2=1.985
r184 28 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=0.995
+ $X2=7.345 $Y2=1.16
r185 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.345 $Y=0.995
+ $X2=7.345 $Y2=0.56
r186 24 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=1.16
r187 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=1.985
r188 21 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=0.995
+ $X2=6.925 $Y2=1.16
r189 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.925 $Y=0.995
+ $X2=6.925 $Y2=0.56
r190 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=1.325
+ $X2=6.505 $Y2=1.16
r191 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.505 $Y=1.325
+ $X2=6.505 $Y2=1.985
r192 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=0.995
+ $X2=6.505 $Y2=1.16
r193 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.505 $Y=0.995
+ $X2=6.505 $Y2=0.56
r194 10 36 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.16
r195 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.985
r196 7 36 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=1.16
r197 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=0.56
r198 2 67 400 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.485 $X2=4.95 $Y2=1.62
r199 2 48 400 $w=1.7e-07 $l=9.02773e-07 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.485 $X2=4.95 $Y2=2.3
r200 1 44 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.235 $X2=4.945 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%VPWR 1 2 3 4 5 6 7 24 28 32 34 38 42 46 48
+ 50 54 56 61 66 74 79 84 90 93 96 99 102 105 109
c129 109 0 1.2348e-19 $X=7.59 $Y=2.72
c130 1 0 3.29888e-20 $X=0.545 $Y=1.815
r131 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r132 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r133 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r134 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r135 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r136 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r137 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r138 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r139 88 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r140 88 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r141 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r142 85 105 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.8 $Y=2.72
+ $X2=6.67 $Y2=2.72
r143 85 87 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.8 $Y=2.72
+ $X2=7.13 $Y2=2.72
r144 84 108 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.47 $Y=2.72
+ $X2=7.645 $Y2=2.72
r145 84 87 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.47 $Y=2.72
+ $X2=7.13 $Y2=2.72
r146 83 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r147 83 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r148 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r149 80 102 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.84 $Y=2.72
+ $X2=5.707 $Y2=2.72
r150 80 82 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.84 $Y=2.72
+ $X2=6.21 $Y2=2.72
r151 79 105 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.54 $Y=2.72
+ $X2=6.67 $Y2=2.72
r152 79 82 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.54 $Y=2.72
+ $X2=6.21 $Y2=2.72
r153 78 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 78 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r155 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r156 75 99 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.58 $Y=2.72
+ $X2=4.437 $Y2=2.72
r157 75 77 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.58 $Y=2.72
+ $X2=5.29 $Y2=2.72
r158 74 102 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=5.575 $Y=2.72
+ $X2=5.707 $Y2=2.72
r159 74 77 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.575 $Y=2.72
+ $X2=5.29 $Y2=2.72
r160 73 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r161 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r162 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r163 70 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r164 69 72 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r165 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r166 67 93 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.632 $Y2=2.72
r167 67 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=2.07 $Y2=2.72
r168 66 96 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=3.515 $Y2=2.72
r169 66 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.335 $Y=2.72
+ $X2=2.99 $Y2=2.72
r170 65 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r171 65 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r172 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r173 62 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r174 62 64 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r175 61 93 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=1.632 $Y2=2.72
r176 61 64 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.45 $Y=2.72 $X2=1.15
+ $Y2=2.72
r177 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r178 56 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r179 54 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r180 54 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r181 50 53 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=7.602 $Y=1.66
+ $X2=7.602 $Y2=2.34
r182 48 108 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=7.602 $Y=2.635
+ $X2=7.645 $Y2=2.72
r183 48 53 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=7.602 $Y=2.635
+ $X2=7.602 $Y2=2.34
r184 44 105 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.67 $Y=2.635
+ $X2=6.67 $Y2=2.72
r185 44 46 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.67 $Y=2.635
+ $X2=6.67 $Y2=2.34
r186 40 102 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.707 $Y=2.635
+ $X2=5.707 $Y2=2.72
r187 40 42 27.6151 $w=2.63e-07 $l=6.35e-07 $layer=LI1_cond $X=5.707 $Y=2.635
+ $X2=5.707 $Y2=2
r188 36 99 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.437 $Y=2.635
+ $X2=4.437 $Y2=2.72
r189 36 38 14.7594 $w=2.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.437 $Y=2.635
+ $X2=4.437 $Y2=2.27
r190 35 96 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.515 $Y2=2.72
r191 34 99 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=4.437 $Y2=2.72
r192 34 35 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=3.695 $Y2=2.72
r193 30 96 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.635
+ $X2=3.515 $Y2=2.72
r194 30 32 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.515 $Y=2.635
+ $X2=3.515 $Y2=2.34
r195 26 93 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.632 $Y=2.635
+ $X2=1.632 $Y2=2.72
r196 26 28 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.632 $Y=2.635
+ $X2=1.632 $Y2=2.34
r197 22 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r198 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r199 7 53 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.42
+ $Y=1.485 $X2=7.555 $Y2=2.34
r200 7 50 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.42
+ $Y=1.485 $X2=7.555 $Y2=1.66
r201 6 46 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.58
+ $Y=1.485 $X2=6.715 $Y2=2.34
r202 5 42 300 $w=1.7e-07 $l=5.91777e-07 $layer=licon1_PDIFF $count=2 $X=5.59
+ $Y=1.485 $X2=5.755 $Y2=2
r203 4 38 600 $w=1.7e-07 $l=8.56723e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.485 $X2=4.415 $Y2=2.27
r204 3 32 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=2.065 $X2=3.42 $Y2=2.34
r205 2 28 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=2.34
r206 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%GCLK 1 2 3 4 14 15 16 19 24 26 28 29 30 31
+ 32 34
c77 3 0 1.37048e-19 $X=6.07 $Y=1.485
r78 34 64 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.135 $Y=2.21
+ $X2=7.135 $Y2=2.34
r79 34 73 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=7.135 $Y=2.21
+ $X2=7.135 $Y2=2.005
r80 32 58 2.82709 $w=5.48e-07 $l=1.3e-07 $layer=LI1_cond $X=7.025 $Y=1.53
+ $X2=7.025 $Y2=1.66
r81 31 32 7.39394 $w=5.48e-07 $l=3.4e-07 $layer=LI1_cond $X=7.025 $Y=1.19
+ $X2=7.025 $Y2=1.53
r82 30 50 2.21278 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=0.8
+ $X2=7.025 $Y2=0.885
r83 30 31 6.08913 $w=5.48e-07 $l=2.8e-07 $layer=LI1_cond $X=7.025 $Y=0.91
+ $X2=7.025 $Y2=1.19
r84 30 50 0.543672 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=7.025 $Y=0.91
+ $X2=7.025 $Y2=0.885
r85 29 73 4.92088 $w=7.13e-07 $l=8.5e-08 $layer=LI1_cond $X=6.942 $Y=1.92
+ $X2=6.942 $Y2=2.005
r86 29 58 2.78771 $w=7.23e-07 $l=1.25e-07 $layer=LI1_cond $X=7.025 $Y=1.785
+ $X2=7.025 $Y2=1.66
r87 27 28 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.205 $Y=2.005
+ $X2=6.205 $Y2=2.21
r88 26 29 9.77989 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=6.37 $Y=1.92
+ $X2=6.585 $Y2=1.92
r89 26 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.37 $Y=1.92
+ $X2=6.205 $Y2=2.005
r90 22 24 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.205 $Y=0.4
+ $X2=6.375 $Y2=0.4
r91 17 30 2.21278 $w=4.4e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.135 $Y=0.715
+ $X2=7.025 $Y2=0.8
r92 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.135 $Y=0.715
+ $X2=7.135 $Y2=0.38
r93 15 30 4.90852 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=6.75 $Y=0.8
+ $X2=7.025 $Y2=0.8
r94 15 16 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.75 $Y=0.8 $X2=6.46
+ $Y2=0.8
r95 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=0.715
+ $X2=6.46 $Y2=0.8
r96 13 24 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.375 $Y=0.545
+ $X2=6.375 $Y2=0.4
r97 13 14 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.375 $Y=0.545
+ $X2=6.375 $Y2=0.715
r98 4 64 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7
+ $Y=1.485 $X2=7.135 $Y2=2.34
r99 4 58 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7
+ $Y=1.485 $X2=7.135 $Y2=1.66
r100 3 28 600 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.485 $X2=6.205 $Y2=2.29
r101 2 19 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7
+ $Y=0.235 $X2=7.135 $Y2=0.38
r102 1 22 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.07
+ $Y=0.235 $X2=6.205 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_4%VGND 1 2 3 4 5 6 7 24 28 32 34 38 42 44 48
+ 50 52 54 56 61 66 74 79 85 88 91 94 97 100 104
c131 104 0 2.71124e-20 $X=7.59 $Y=0
c132 48 0 1.95136e-19 $X=6.715 $Y=0.38
r133 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r134 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r135 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r136 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r137 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r138 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r139 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r140 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r141 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r142 83 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r143 83 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.67 $Y2=0
r144 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r145 80 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=0 $X2=6.715
+ $Y2=0
r146 80 82 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.8 $Y=0 $X2=7.13
+ $Y2=0
r147 79 103 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.47 $Y=0
+ $X2=7.645 $Y2=0
r148 79 82 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=7.13
+ $Y2=0
r149 78 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r150 78 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r151 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r152 75 94 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.58 $Y=0 $X2=4.437
+ $Y2=0
r153 75 77 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.58 $Y=0 $X2=5.29
+ $Y2=0
r154 74 97 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.73
+ $Y2=0
r155 74 77 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.29
+ $Y2=0
r156 73 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r157 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r158 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r159 70 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r160 69 72 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r161 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r162 67 88 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.617 $Y2=0
r163 67 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r164 66 91 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=3.482 $Y2=0
r165 66 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=2.99 $Y2=0
r166 65 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r167 65 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r168 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r169 62 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r170 62 64 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r171 61 88 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.617
+ $Y2=0
r172 61 64 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.15
+ $Y2=0
r173 56 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r174 56 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r175 54 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r176 54 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r177 50 103 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=7.602 $Y=0.085
+ $X2=7.645 $Y2=0
r178 50 52 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=7.602 $Y=0.085
+ $X2=7.602 $Y2=0.38
r179 46 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=0.085
+ $X2=6.715 $Y2=0
r180 46 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.715 $Y=0.085
+ $X2=6.715 $Y2=0.38
r181 45 97 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.87 $Y=0 $X2=5.73
+ $Y2=0
r182 44 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.63 $Y=0 $X2=6.715
+ $Y2=0
r183 44 45 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.63 $Y=0 $X2=5.87
+ $Y2=0
r184 40 97 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.73 $Y=0.085
+ $X2=5.73 $Y2=0
r185 40 42 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.73 $Y=0.085
+ $X2=5.73 $Y2=0.38
r186 36 94 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.437 $Y=0.085
+ $X2=4.437 $Y2=0
r187 36 38 14.7594 $w=2.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.437 $Y=0.085
+ $X2=4.437 $Y2=0.45
r188 35 91 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.482
+ $Y2=0
r189 34 94 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.437 $Y2=0
r190 34 35 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=3.65 $Y2=0
r191 30 91 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.482 $Y=0.085
+ $X2=3.482 $Y2=0
r192 30 32 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=3.482 $Y=0.085
+ $X2=3.482 $Y2=0.445
r193 26 88 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.617 $Y=0.085
+ $X2=1.617 $Y2=0
r194 26 28 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=1.617 $Y=0.085
+ $X2=1.617 $Y2=0.38
r195 22 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r196 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r197 7 52 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.42
+ $Y=0.235 $X2=7.555 $Y2=0.38
r198 6 48 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.235 $X2=6.715 $Y2=0.38
r199 5 42 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.65
+ $Y=0.235 $X2=5.785 $Y2=0.38
r200 4 38 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=4.29
+ $Y=0.235 $X2=4.425 $Y2=0.45
r201 3 32 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.235 $X2=3.485 $Y2=0.445
r202 2 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r203 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


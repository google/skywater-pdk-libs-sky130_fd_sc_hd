* File: sky130_fd_sc_hd__fa_2.pex.spice
* Created: Thu Aug 27 14:21:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__FA_2%A_80_21# 1 2 7 9 12 14 16 19 23 27 29 35 37 38
+ 39 40 43 44 45 46 48 50 54 55 58 61 67 70 71
c226 70 0 5.62553e-20 $X=5.415 $Y=1.04
c227 61 0 1.85285e-19 $X=5.77 $Y=0.85
c228 55 0 3.3579e-19 $X=2.215 $Y=0.85
c229 46 0 1.95515e-19 $X=2.072 $Y=2.08
c230 43 0 1.83284e-19 $X=1.39 $Y=1.91
c231 40 0 7.98542e-20 $X=1.305 $Y=1.58
r232 70 73 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=1.04
+ $X2=5.415 $Y2=1.205
r233 70 72 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=1.04
+ $X2=5.415 $Y2=0.875
r234 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.415
+ $Y=1.04 $X2=5.415 $Y2=1.04
r235 62 71 13.8814 $w=3.12e-07 $l=3.99687e-07 $layer=LI1_cond $X=5.77 $Y=0.945
+ $X2=5.415 $Y2=1.04
r236 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.77 $Y=0.85
+ $X2=5.77 $Y2=0.85
r237 58 76 0.199673 $w=6.11e-07 $l=1e-08 $layer=LI1_cond $X=2.07 $Y=0.595
+ $X2=2.08 $Y2=0.595
r238 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0.85
+ $X2=2.07 $Y2=0.85
r239 55 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.215 $Y=0.85
+ $X2=2.07 $Y2=0.85
r240 54 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.625 $Y=0.85
+ $X2=5.77 $Y2=0.85
r241 54 55 4.22029 $w=1.4e-07 $l=3.41e-06 $layer=MET1_cond $X=5.625 $Y=0.85
+ $X2=2.215 $Y2=0.85
r242 46 53 2.61083 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.072 $Y=2.08
+ $X2=2.072 $Y2=1.995
r243 46 48 8.51806 $w=3.43e-07 $l=2.55e-07 $layer=LI1_cond $X=2.072 $Y=2.08
+ $X2=2.072 $Y2=2.335
r244 44 53 5.28309 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.9 $Y=1.995
+ $X2=2.072 $Y2=1.995
r245 44 45 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.9 $Y=1.995
+ $X2=1.475 $Y2=1.995
r246 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.39 $Y=1.91
+ $X2=1.475 $Y2=1.995
r247 42 43 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.39 $Y=1.665
+ $X2=1.39 $Y2=1.91
r248 41 51 1.54022 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.11 $Y=1.58
+ $X2=1.007 $Y2=1.58
r249 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.305 $Y=1.58
+ $X2=1.39 $Y2=1.665
r250 40 41 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.305 $Y=1.58
+ $X2=1.11 $Y2=1.58
r251 38 58 17.8202 $w=6.11e-07 $l=6.03158e-07 $layer=LI1_cond $X=1.535 $Y=0.74
+ $X2=2.07 $Y2=0.595
r252 38 39 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.535 $Y=0.74
+ $X2=1.075 $Y2=0.74
r253 37 51 9.61743 $w=1.95e-07 $l=1.58272e-07 $layer=LI1_cond $X=0.99 $Y=1.43
+ $X2=1.007 $Y2=1.58
r254 36 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=1.245
+ $X2=0.99 $Y2=1.16
r255 36 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.99 $Y=1.245
+ $X2=0.99 $Y2=1.43
r256 35 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=1.075
+ $X2=0.99 $Y2=1.16
r257 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.99 $Y=0.825
+ $X2=1.075 $Y2=0.74
r258 34 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.99 $Y=0.825
+ $X2=0.99 $Y2=1.075
r259 32 67 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.705 $Y=1.16
+ $X2=0.895 $Y2=1.16
r260 32 64 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.705 $Y=1.16
+ $X2=0.475 $Y2=1.16
r261 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.705
+ $Y=1.16 $X2=0.705 $Y2=1.16
r262 29 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=1.16
+ $X2=0.99 $Y2=1.16
r263 29 31 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.905 $Y=1.16
+ $X2=0.705 $Y2=1.16
r264 27 73 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=5.355 $Y=2.165
+ $X2=5.355 $Y2=1.205
r265 23 72 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.355 $Y=0.445
+ $X2=5.355 $Y2=0.875
r266 17 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.325
+ $X2=0.895 $Y2=1.16
r267 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.895 $Y=1.325
+ $X2=0.895 $Y2=1.985
r268 14 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=0.995
+ $X2=0.895 $Y2=1.16
r269 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.895 $Y=0.995
+ $X2=0.895 $Y2=0.56
r270 10 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.16
r271 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.985
r272 7 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r273 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r274 2 53 600 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.855 $X2=2.08 $Y2=1.995
r275 2 48 600 $w=1.7e-07 $l=5.67098e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.855 $X2=2.08 $Y2=2.335
r276 1 76 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.235 $X2=2.08 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%A 1 3 7 11 15 19 23 27 31 33 35 36 37 38 39 40
+ 47 52 59 64 65 69 70
c266 65 0 3.76974e-20 $X=4.915 $Y=1.04
c267 47 0 1.2547e-19 $X=2.99 $Y=1.19
c268 38 0 3.10095e-19 $X=3.135 $Y=1.19
c269 37 0 1.21386e-19 $X=4.705 $Y=1.19
c270 36 0 7.98542e-20 $X=1.755 $Y=1.19
c271 23 0 7.10647e-20 $X=4.91 $Y=2.165
c272 15 0 1.95515e-19 $X=2.71 $Y=2.17
c273 11 0 1.9888e-19 $X=2.71 $Y=0.445
c274 7 0 1.3691e-19 $X=1.395 $Y=0.445
c275 3 0 1.22604e-19 $X=1.37 $Y=2.17
r276 69 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.16
+ $X2=6.795 $Y2=0.995
r277 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.795
+ $Y=1.16 $X2=6.795 $Y2=1.16
r278 64 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.915 $Y=1.04
+ $X2=4.915 $Y2=1.205
r279 64 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.915 $Y=1.04
+ $X2=4.915 $Y2=0.875
r280 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.915
+ $Y=1.04 $X2=4.915 $Y2=1.04
r281 59 62 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.195
+ $X2=2.77 $Y2=1.36
r282 59 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.195
+ $X2=2.77 $Y2=1.03
r283 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.195 $X2=2.77 $Y2=1.195
r284 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.33
+ $Y=1.16 $X2=1.33 $Y2=1.16
r285 53 70 23.2547 $w=2.78e-07 $l=5.65e-07 $layer=LI1_cond $X=6.23 $Y=1.135
+ $X2=6.795 $Y2=1.135
r286 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.23 $Y=1.19
+ $X2=6.23 $Y2=1.19
r287 49 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.85 $Y=1.19
+ $X2=4.85 $Y2=1.19
r288 47 60 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.99 $Y=1.195
+ $X2=2.77 $Y2=1.195
r289 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.19
+ $X2=2.99 $Y2=1.19
r290 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.995 $Y=1.19
+ $X2=4.85 $Y2=1.19
r291 39 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.085 $Y=1.19
+ $X2=6.23 $Y2=1.19
r292 39 40 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=6.085 $Y=1.19
+ $X2=4.995 $Y2=1.19
r293 38 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.19
+ $X2=2.99 $Y2=1.19
r294 37 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=1.19
+ $X2=4.85 $Y2=1.19
r295 37 38 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=4.705 $Y=1.19
+ $X2=3.135 $Y2=1.19
r296 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.19
+ $X2=1.61 $Y2=1.19
r297 35 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=1.19
+ $X2=2.99 $Y2=1.19
r298 35 36 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=2.845 $Y=1.19
+ $X2=1.755 $Y2=1.19
r299 33 57 11.2 $w=3.05e-07 $l=2.8e-07 $layer=LI1_cond $X=1.61 $Y=1.16 $X2=1.33
+ $Y2=1.16
r300 33 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.19
+ $X2=1.61 $Y2=1.19
r301 29 69 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.325
+ $X2=6.795 $Y2=1.16
r302 29 31 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=6.795 $Y=1.325
+ $X2=6.795 $Y2=2.17
r303 27 71 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.735 $Y=0.445
+ $X2=6.735 $Y2=0.995
r304 23 67 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=4.91 $Y=2.165
+ $X2=4.91 $Y2=1.205
r305 19 66 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.91 $Y=0.445
+ $X2=4.91 $Y2=0.875
r306 15 62 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.71 $Y=2.17
+ $X2=2.71 $Y2=1.36
r307 11 61 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=2.71 $Y=0.445
+ $X2=2.71 $Y2=1.03
r308 5 56 38.8629 $w=2.72e-07 $l=1.93959e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.332 $Y2=1.16
r309 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.395 $Y=0.995
+ $X2=1.395 $Y2=0.445
r310 1 56 38.8629 $w=2.72e-07 $l=1.83016e-07 $layer=POLY_cond $X=1.37 $Y=1.325
+ $X2=1.332 $Y2=1.16
r311 1 3 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=1.37 $Y=1.325
+ $X2=1.37 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%B 3 7 9 11 12 14 15 16 17 18 19 21 26 29 33 35
+ 36 38 39 40 41 50 51 54 59 60 61 63 65
c233 54 0 4.51526e-19 $X=1.81 $Y=1.53
c234 51 0 2.28809e-19 $X=6.69 $Y=1.53
c235 50 0 3.77214e-20 $X=6.69 $Y=1.53
c236 41 0 5.10808e-21 $X=4.075 $Y=1.53
c237 40 0 1.7744e-19 $X=6.545 $Y=1.53
c238 39 0 1.22604e-19 $X=2.215 $Y=1.53
c239 29 0 1.47587e-19 $X=6.255 $Y=0.445
c240 18 0 1.2547e-19 $X=3.205 $Y=1.695
r241 65 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.53
+ $X2=6.315 $Y2=1.695
r242 65 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.53
+ $X2=6.315 $Y2=1.365
r243 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.315
+ $Y=1.53 $X2=6.315 $Y2=1.53
r244 59 61 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.957 $Y=1.52
+ $X2=3.957 $Y2=1.355
r245 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.905
+ $Y=1.52 $X2=3.905 $Y2=1.52
r246 54 57 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.53
+ $X2=1.81 $Y2=1.695
r247 54 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.53
+ $X2=1.81 $Y2=1.365
r248 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.53 $X2=1.81 $Y2=1.53
r249 51 66 14.9023 $w=2.88e-07 $l=3.75e-07 $layer=LI1_cond $X=6.69 $Y=1.59
+ $X2=6.315 $Y2=1.59
r250 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.69 $Y=1.53
+ $X2=6.69 $Y2=1.53
r251 47 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.93 $Y=1.53
+ $X2=3.93 $Y2=1.53
r252 41 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.075 $Y=1.53
+ $X2=3.93 $Y2=1.53
r253 40 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.545 $Y=1.53
+ $X2=6.69 $Y2=1.53
r254 40 41 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=6.545 $Y=1.53
+ $X2=4.075 $Y2=1.53
r255 39 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.215 $Y=1.53
+ $X2=2.07 $Y2=1.53
r256 38 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.785 $Y=1.53
+ $X2=3.93 $Y2=1.53
r257 38 39 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=3.785 $Y=1.53
+ $X2=2.215 $Y2=1.53
r258 36 55 12.23 $w=2.43e-07 $l=2.6e-07 $layer=LI1_cond $X=2.07 $Y=1.567
+ $X2=1.81 $Y2=1.567
r259 36 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=1.53
+ $X2=2.07 $Y2=1.53
r260 33 68 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=6.255 $Y=2.17
+ $X2=6.255 $Y2=1.695
r261 29 67 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=6.255 $Y=0.445
+ $X2=6.255 $Y2=1.365
r262 26 63 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.07 $Y=2.165
+ $X2=4.07 $Y2=1.77
r263 22 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.07 $Y=0.88
+ $X2=4.07 $Y2=0.805
r264 22 61 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.07 $Y=0.88
+ $X2=4.07 $Y2=1.355
r265 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.07 $Y=0.73
+ $X2=4.07 $Y2=0.805
r266 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.07 $Y=0.73
+ $X2=4.07 $Y2=0.445
r267 17 63 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=3.957 $Y=1.695
+ $X2=3.957 $Y2=1.77
r268 17 59 25.9538 $w=3.75e-07 $l=1.75e-07 $layer=POLY_cond $X=3.957 $Y=1.695
+ $X2=3.957 $Y2=1.52
r269 17 18 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.77 $Y=1.695
+ $X2=3.205 $Y2=1.695
r270 15 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.995 $Y=0.805
+ $X2=4.07 $Y2=0.805
r271 15 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.995 $Y=0.805
+ $X2=3.205 $Y2=0.805
r272 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.13 $Y=1.77
+ $X2=3.205 $Y2=1.695
r273 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.13 $Y=1.77 $X2=3.13
+ $Y2=2.17
r274 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.13 $Y=0.73
+ $X2=3.205 $Y2=0.805
r275 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.13 $Y=0.73 $X2=3.13
+ $Y2=0.445
r276 7 56 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.87 $Y=0.445
+ $X2=1.87 $Y2=1.365
r277 3 57 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.815 $Y=2.17
+ $X2=1.815 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%CIN 3 7 11 14 20 24 26 27 29 30 31 33 34 35 37
+ 38 42 44 50 51 52 56 58 59
c228 50 0 2.2917e-19 $X=4.49 $Y=1.52
c229 44 0 1.55247e-19 $X=2.41 $Y=1.19
c230 42 0 2.45299e-20 $X=2.29 $Y=1.19
c231 34 0 7.10647e-20 $X=4.295 $Y=1.107
c232 31 0 1.35567e-19 $X=2.495 $Y=1.655
c233 29 0 2.87523e-19 $X=2.41 $Y=1.57
c234 20 0 1.8774e-19 $X=5.78 $Y=2.165
r235 59 64 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.795 $Y=1.52
+ $X2=5.795 $Y2=1.6
r236 58 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.835 $Y=1.52
+ $X2=5.835 $Y2=1.685
r237 58 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.835 $Y=1.52
+ $X2=5.835 $Y2=1.355
r238 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.835
+ $Y=1.52 $X2=5.835 $Y2=1.52
r239 52 64 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=5.795 $Y=1.87
+ $X2=5.795 $Y2=1.6
r240 50 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.49 $Y=1.52
+ $X2=4.49 $Y2=1.355
r241 49 51 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.49 $Y=1.56
+ $X2=4.655 $Y2=1.56
r242 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.49
+ $Y=1.52 $X2=4.49 $Y2=1.52
r243 46 49 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=4.38 $Y=1.56
+ $X2=4.49 $Y2=1.56
r244 41 44 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.29 $Y=1.19
+ $X2=2.41 $Y2=1.19
r245 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.19 $X2=2.29 $Y2=1.19
r246 38 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.67 $Y=1.6
+ $X2=5.795 $Y2=1.6
r247 38 51 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=5.67 $Y=1.6
+ $X2=4.655 $Y2=1.6
r248 37 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.38 $Y=1.435
+ $X2=4.38 $Y2=1.56
r249 36 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.38 $Y=1.25
+ $X2=4.38 $Y2=1.435
r250 34 36 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=4.295 $Y=1.107
+ $X2=4.38 $Y2=1.25
r251 34 35 35.5842 $w=2.83e-07 $l=8.8e-07 $layer=LI1_cond $X=4.295 $Y=1.107
+ $X2=3.415 $Y2=1.107
r252 32 35 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.33 $Y=1.25
+ $X2=3.415 $Y2=1.107
r253 32 33 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.33 $Y=1.25
+ $X2=3.33 $Y2=1.57
r254 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=1.655
+ $X2=3.33 $Y2=1.57
r255 30 31 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.245 $Y=1.655
+ $X2=2.495 $Y2=1.655
r256 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=1.57
+ $X2=2.495 $Y2=1.655
r257 28 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=1.275
+ $X2=2.41 $Y2=1.19
r258 28 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.41 $Y=1.275
+ $X2=2.41 $Y2=1.57
r259 27 56 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.495 $Y=0.88
+ $X2=4.495 $Y2=1.355
r260 26 27 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=4.492 $Y=0.73
+ $X2=4.492 $Y2=0.88
r261 24 60 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=5.895 $Y=0.445
+ $X2=5.895 $Y2=1.355
r262 20 61 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.78 $Y=2.165
+ $X2=5.78 $Y2=1.685
r263 12 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.49 $Y=1.685
+ $X2=4.49 $Y2=1.52
r264 12 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.49 $Y=1.685
+ $X2=4.49 $Y2=2.165
r265 11 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.49 $Y=0.445
+ $X2=4.49 $Y2=0.73
r266 5 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.355
+ $X2=2.29 $Y2=1.19
r267 5 7 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.29 $Y=1.355
+ $X2=2.29 $Y2=2.17
r268 1 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.025
+ $X2=2.29 $Y2=1.19
r269 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.29 $Y=1.025
+ $X2=2.29 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%A_1086_47# 1 2 7 9 12 16 18 20 21 25 28 29 30
+ 31 34 36 38 41 47 48 54 56 62
c144 48 0 1.7744e-19 $X=6.6 $Y=2.02
c145 47 0 5.62553e-20 $X=5.71 $Y=0.425
c146 34 0 3.77214e-20 $X=7.095 $Y=1.935
r147 61 62 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=7.69 $Y=1.16 $X2=7.77
+ $Y2=1.16
r148 57 59 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=7.23 $Y=1.16 $X2=7.27
+ $Y2=1.16
r149 52 54 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.095 $Y=1.555
+ $X2=7.215 $Y2=1.555
r150 45 47 3.71115 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=0.425
+ $X2=5.71 $Y2=0.425
r151 42 61 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=7.635 $Y=1.16
+ $X2=7.69 $Y2=1.16
r152 42 59 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=7.635 $Y=1.16
+ $X2=7.27 $Y2=1.16
r153 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.635
+ $Y=1.16 $X2=7.635 $Y2=1.16
r154 39 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=1.16
+ $X2=7.215 $Y2=1.16
r155 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.3 $Y=1.16
+ $X2=7.635 $Y2=1.16
r156 38 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=1.47
+ $X2=7.215 $Y2=1.555
r157 37 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=1.245
+ $X2=7.215 $Y2=1.16
r158 37 38 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.215 $Y=1.245
+ $X2=7.215 $Y2=1.47
r159 36 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=1.075
+ $X2=7.215 $Y2=1.16
r160 35 36 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.215 $Y=0.825
+ $X2=7.215 $Y2=1.075
r161 33 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=1.64
+ $X2=7.095 $Y2=1.555
r162 33 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.095 $Y=1.64
+ $X2=7.095 $Y2=1.935
r163 32 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.685 $Y=2.02
+ $X2=6.6 $Y2=2.02
r164 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.01 $Y=2.02
+ $X2=7.095 $Y2=1.935
r165 31 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.01 $Y=2.02
+ $X2=6.685 $Y2=2.02
r166 29 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.13 $Y=0.74
+ $X2=7.215 $Y2=0.825
r167 29 30 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.13 $Y=0.74
+ $X2=6.55 $Y2=0.74
r168 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.465 $Y=0.655
+ $X2=6.55 $Y2=0.74
r169 27 28 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.465 $Y=0.505
+ $X2=6.465 $Y2=0.655
r170 25 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.38 $Y=0.38
+ $X2=6.465 $Y2=0.505
r171 25 47 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=6.38 $Y=0.38
+ $X2=5.71 $Y2=0.38
r172 21 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.6 $Y2=2.02
r173 21 23 32.0311 $w=3.38e-07 $l=9.45e-07 $layer=LI1_cond $X=6.515 $Y=2.295
+ $X2=5.57 $Y2=2.295
r174 18 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.77 $Y=0.995
+ $X2=7.77 $Y2=1.16
r175 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.77 $Y=0.995
+ $X2=7.77 $Y2=0.56
r176 14 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.69 $Y=1.325
+ $X2=7.69 $Y2=1.16
r177 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.69 $Y=1.325
+ $X2=7.69 $Y2=1.985
r178 10 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.325
+ $X2=7.27 $Y2=1.16
r179 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.27 $Y=1.325
+ $X2=7.27 $Y2=1.985
r180 7 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.23 $Y=0.995
+ $X2=7.23 $Y2=1.16
r181 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.23 $Y=0.995
+ $X2=7.23 $Y2=0.56
r182 2 23 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.845 $X2=5.57 $Y2=2.3
r183 1 45 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=5.43
+ $Y=0.235 $X2=5.625 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 47 48 49
+ 52 54 59 67 72 77 87 88 96 99 102 105 108 111
r137 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r138 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r139 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r140 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r141 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r142 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r143 85 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r144 85 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r145 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r146 82 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.22 $Y=2.72
+ $X2=7.055 $Y2=2.72
r147 82 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.22 $Y=2.72
+ $X2=7.59 $Y2=2.72
r148 81 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r149 81 106 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=4.83 $Y2=2.72
r150 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r151 78 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=2.72
+ $X2=4.7 $Y2=2.72
r152 78 80 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=4.865 $Y=2.72
+ $X2=6.67 $Y2=2.72
r153 77 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.89 $Y=2.72
+ $X2=7.055 $Y2=2.72
r154 77 80 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.89 $Y=2.72
+ $X2=6.67 $Y2=2.72
r155 76 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r156 76 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r157 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r158 73 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=2.72
+ $X2=3.86 $Y2=2.72
r159 73 75 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.025 $Y=2.72
+ $X2=4.37 $Y2=2.72
r160 72 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=2.72
+ $X2=4.7 $Y2=2.72
r161 72 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=2.72
+ $X2=4.37 $Y2=2.72
r162 71 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r163 71 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r164 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r165 68 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=2.72
+ $X2=2.92 $Y2=2.72
r166 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=2.72
+ $X2=3.45 $Y2=2.72
r167 67 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.86 $Y2=2.72
r168 67 70 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.695 $Y=2.72
+ $X2=3.45 $Y2=2.72
r169 66 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r170 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r171 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r172 63 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r173 62 65 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r174 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r175 60 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=2.72
+ $X2=1.145 $Y2=2.72
r176 60 62 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.31 $Y=2.72 $X2=1.61
+ $Y2=2.72
r177 59 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.92 $Y2=2.72
r178 59 65 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.53 $Y2=2.72
r179 58 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r180 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r181 55 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.35 $Y=2.72
+ $X2=0.69 $Y2=2.72
r182 54 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=2.72
+ $X2=1.145 $Y2=2.72
r183 54 57 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.98 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 52 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r185 49 111 27.7449 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=1.96
r186 49 55 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.175 $Y=2.72
+ $X2=0.35 $Y2=2.72
r187 49 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r188 47 84 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.815 $Y=2.72
+ $X2=7.59 $Y2=2.72
r189 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=2.72
+ $X2=7.9 $Y2=2.72
r190 46 87 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.985 $Y=2.72
+ $X2=8.05 $Y2=2.72
r191 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=2.72
+ $X2=7.9 $Y2=2.72
r192 42 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=2.635 $X2=7.9
+ $Y2=2.72
r193 42 44 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.9 $Y=2.635
+ $X2=7.9 $Y2=1.96
r194 38 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=2.635
+ $X2=7.055 $Y2=2.72
r195 38 40 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.055 $Y=2.635
+ $X2=7.055 $Y2=2.36
r196 34 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=2.635
+ $X2=4.7 $Y2=2.72
r197 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.7 $Y=2.635
+ $X2=4.7 $Y2=2.36
r198 30 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=2.635
+ $X2=3.86 $Y2=2.72
r199 30 32 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.86 $Y=2.635
+ $X2=3.86 $Y2=2
r200 26 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=2.635
+ $X2=2.92 $Y2=2.72
r201 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.92 $Y=2.635
+ $X2=2.92 $Y2=2.36
r202 22 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.72
r203 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.36
r204 7 44 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.765
+ $Y=1.485 $X2=7.9 $Y2=1.96
r205 6 40 600 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_PDIFF $count=1 $X=6.87
+ $Y=1.855 $X2=7.055 $Y2=2.36
r206 5 36 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.845 $X2=4.7 $Y2=2.36
r207 4 32 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=3.735
+ $Y=1.845 $X2=3.86 $Y2=2
r208 3 28 600 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.855 $X2=2.92 $Y2=2.36
r209 2 24 600 $w=1.7e-07 $l=9.58514e-07 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.485 $X2=1.145 $Y2=2.36
r210 1 111 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%COUT 1 2 8 9 10 12 17 21 23 24 35 37
r44 37 38 4.03065 $w=2.43e-07 $l=8e-08 $layer=LI1_cond $X=0.687 $Y=1.87
+ $X2=0.687 $Y2=1.95
r45 23 37 0.141115 $w=2.43e-07 $l=3e-09 $layer=LI1_cond $X=0.687 $Y=1.867
+ $X2=0.687 $Y2=1.87
r46 23 35 5.18354 $w=2.43e-07 $l=8.7e-08 $layer=LI1_cond $X=0.687 $Y=1.867
+ $X2=0.687 $Y2=1.78
r47 23 24 13.626 $w=2.08e-07 $l=2.58e-07 $layer=LI1_cond $X=0.705 $Y=1.952
+ $X2=0.705 $Y2=2.21
r48 23 38 0.105628 $w=2.08e-07 $l=2e-09 $layer=LI1_cond $X=0.705 $Y=1.952
+ $X2=0.705 $Y2=1.95
r49 13 35 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.65 $Y=1.585
+ $X2=0.65 $Y2=1.78
r50 12 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.735
+ $X2=0.605 $Y2=0.82
r51 11 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0.485
+ $X2=0.605 $Y2=0.4
r52 11 12 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.605 $Y=0.485
+ $X2=0.605 $Y2=0.735
r53 9 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.565 $Y=1.5
+ $X2=0.65 $Y2=1.585
r54 9 10 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.565 $Y=1.5
+ $X2=0.37 $Y2=1.5
r55 8 10 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.227 $Y=1.415
+ $X2=0.37 $Y2=1.5
r56 7 17 24.661 $w=1.68e-07 $l=3.78e-07 $layer=LI1_cond $X=0.227 $Y=0.82
+ $X2=0.605 $Y2=0.82
r57 7 8 20.6227 $w=2.83e-07 $l=5.1e-07 $layer=LI1_cond $X=0.227 $Y=0.905
+ $X2=0.227 $Y2=1.415
r58 2 23 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.685 $Y2=1.96
r59 1 21 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.685 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%A_473_371# 1 2 7 10 11 12
c23 11 0 2.45299e-20 $X=2.585 $Y=2.02
r24 12 14 4.67234 $w=2.35e-07 $l=9e-08 $layer=LI1_cond $X=3.372 $Y=2.105
+ $X2=3.372 $Y2=2.195
r25 10 12 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=3.255 $Y=2.02
+ $X2=3.372 $Y2=2.105
r26 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.255 $Y=2.02
+ $X2=2.585 $Y2=2.02
r27 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.5 $Y=2.105
+ $X2=2.585 $Y2=2.02
r28 7 9 6.45882 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.5 $Y=2.105 $X2=2.5
+ $Y2=2.195
r29 2 14 600 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.855 $X2=3.34 $Y2=2.195
r30 1 9 600 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=1.855 $X2=2.5 $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%A_829_369# 1 2 9 11 12 15
c20 12 0 1.96224e-19 $X=4.365 $Y=2.02
r21 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.12 $Y=2.105
+ $X2=5.12 $Y2=2.275
r22 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=2.02
+ $X2=5.12 $Y2=2.105
r23 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.035 $Y=2.02
+ $X2=4.365 $Y2=2.02
r24 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.28 $Y=2.105
+ $X2=4.365 $Y2=2.02
r25 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.28 $Y=2.105 $X2=4.28
+ $Y2=2.275
r26 2 15 600 $w=1.7e-07 $l=4.929e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=1.845 $X2=5.12 $Y2=2.275
r27 1 9 600 $w=1.7e-07 $l=4.929e-07 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=1.845 $X2=4.28 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%SUM 1 2 10 13 14 15 18 22 23 29
c51 23 0 1.80183e-20 $X=7.52 $Y=1.795
c52 14 0 2.30507e-20 $X=7.645 $Y=1.5
r53 28 29 11.5244 $w=2.23e-07 $l=2.25e-07 $layer=LI1_cond $X=8.082 $Y=1.415
+ $X2=8.082 $Y2=1.19
r54 27 29 14.5976 $w=2.23e-07 $l=2.85e-07 $layer=LI1_cond $X=8.082 $Y=0.905
+ $X2=8.082 $Y2=1.19
r55 22 23 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.52 $Y=1.96
+ $X2=7.52 $Y2=1.795
r56 18 20 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=0.4 $X2=7.56
+ $Y2=0.485
r57 16 26 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.725 $Y=0.82
+ $X2=7.6 $Y2=0.82
r58 15 27 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=7.97 $Y=0.82
+ $X2=8.082 $Y2=0.905
r59 15 16 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.97 $Y=0.82
+ $X2=7.725 $Y2=0.82
r60 13 28 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=7.97 $Y=1.5
+ $X2=8.082 $Y2=1.415
r61 13 14 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.97 $Y=1.5
+ $X2=7.645 $Y2=1.5
r62 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.56 $Y=1.585
+ $X2=7.645 $Y2=1.5
r63 11 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.56 $Y=1.585
+ $X2=7.56 $Y2=1.795
r64 10 26 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=0.735 $X2=7.6
+ $Y2=0.82
r65 10 20 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=7.6 $Y=0.735 $X2=7.6
+ $Y2=0.485
r66 2 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.345
+ $Y=1.485 $X2=7.48 $Y2=1.96
r67 1 26 182 $w=1.7e-07 $l=6.19516e-07 $layer=licon1_NDIFF $count=1 $X=7.305
+ $Y=0.235 $X2=7.56 $Y2=0.74
r68 1 18 182 $w=1.7e-07 $l=3.27261e-07 $layer=licon1_NDIFF $count=1 $X=7.305
+ $Y=0.235 $X2=7.56 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 47 48
+ 49 52 54 59 67 72 81 91 94 97 100 104 106
r148 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r149 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r150 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r151 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r152 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r153 84 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r154 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r155 81 103 3.40825 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=7.895 $Y=0
+ $X2=8.087 $Y2=0
r156 81 83 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.895 $Y=0
+ $X2=7.59 $Y2=0
r157 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r158 80 101 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=4.83 $Y2=0
r159 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r160 77 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=0 $X2=4.7
+ $Y2=0
r161 77 79 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=4.865 $Y=0
+ $X2=6.67 $Y2=0
r162 76 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r163 76 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r164 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r165 73 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=3.86
+ $Y2=0
r166 73 75 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=4.37
+ $Y2=0
r167 72 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=0 $X2=4.7
+ $Y2=0
r168 72 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=0
+ $X2=4.37 $Y2=0
r169 71 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r170 71 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r171 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r172 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=2.92
+ $Y2=0
r173 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0
+ $X2=3.45 $Y2=0
r174 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.86
+ $Y2=0
r175 67 70 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.45
+ $Y2=0
r176 66 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r177 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r178 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r179 63 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r180 62 65 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r181 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r182 60 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.185
+ $Y2=0
r183 60 62 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.61
+ $Y2=0
r184 59 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.92
+ $Y2=0
r185 59 65 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.755 $Y=0
+ $X2=2.53 $Y2=0
r186 58 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r187 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r188 55 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.69
+ $Y2=0
r189 54 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.185
+ $Y2=0
r190 54 57 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.69
+ $Y2=0
r191 52 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r192 49 106 14.1423 $w=3.03e-07 $l=3.15e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.4
r193 49 55 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.175 $Y=0 $X2=0.35
+ $Y2=0
r194 49 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r195 47 79 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.78 $Y=0 $X2=6.67
+ $Y2=0
r196 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=0 $X2=6.945
+ $Y2=0
r197 46 83 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=7.59
+ $Y2=0
r198 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=6.945
+ $Y2=0
r199 42 103 3.40825 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=8.087 $Y2=0
r200 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0.4
r201 38 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.945 $Y=0.085
+ $X2=6.945 $Y2=0
r202 38 40 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.945 $Y=0.085
+ $X2=6.945 $Y2=0.36
r203 34 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=0.085
+ $X2=4.7 $Y2=0
r204 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.7 $Y=0.085
+ $X2=4.7 $Y2=0.36
r205 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0
r206 30 32 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.86 $Y=0.085
+ $X2=3.86 $Y2=0.405
r207 26 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0
r208 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0.36
r209 22 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r210 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.38
r211 7 44 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.845
+ $Y=0.235 $X2=7.98 $Y2=0.4
r212 6 40 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.235 $X2=6.945 $Y2=0.36
r213 5 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.565
+ $Y=0.235 $X2=4.7 $Y2=0.36
r214 4 32 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=0.235 $X2=3.86 $Y2=0.405
r215 3 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.235 $X2=2.92 $Y2=0.36
r216 2 24 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.235 $X2=1.185 $Y2=0.38
r217 1 106 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%A_473_47# 1 2 9 11 12 15
r35 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.34 $Y=0.615
+ $X2=3.34 $Y2=0.445
r36 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.255 $Y=0.7
+ $X2=3.34 $Y2=0.615
r37 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.255 $Y=0.7
+ $X2=2.585 $Y2=0.7
r38 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.5 $Y=0.615
+ $X2=2.585 $Y2=0.7
r39 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.5 $Y=0.615 $X2=2.5
+ $Y2=0.445
r40 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.34 $Y2=0.445
r41 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.235 $X2=2.5 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_2%A_829_47# 1 2 9 11 12 15
c32 12 0 1.49223e-19 $X=4.365 $Y=0.7
r33 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.12 $Y=0.615
+ $X2=5.12 $Y2=0.445
r34 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=0.7
+ $X2=5.12 $Y2=0.615
r35 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.035 $Y=0.7
+ $X2=4.365 $Y2=0.7
r36 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.28 $Y=0.615
+ $X2=4.365 $Y2=0.7
r37 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.28 $Y=0.615 $X2=4.28
+ $Y2=0.445
r38 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.985
+ $Y=0.235 $X2=5.12 $Y2=0.445
r39 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.145
+ $Y=0.235 $X2=4.28 $Y2=0.445
.ends


* File: sky130_fd_sc_hd__and4_4.pxi.spice
* Created: Tue Sep  1 18:58:13 2020
* 
x_PM_SKY130_FD_SC_HD__AND4_4%A N_A_c_72_n N_A_M1014_g N_A_M1012_g A A N_A_c_74_n
+ PM_SKY130_FD_SC_HD__AND4_4%A
x_PM_SKY130_FD_SC_HD__AND4_4%B N_B_M1007_g N_B_M1005_g B B B N_B_c_104_n
+ N_B_c_105_n N_B_c_106_n PM_SKY130_FD_SC_HD__AND4_4%B
x_PM_SKY130_FD_SC_HD__AND4_4%C N_C_M1002_g N_C_M1008_g C C C N_C_c_141_n
+ N_C_c_142_n PM_SKY130_FD_SC_HD__AND4_4%C
x_PM_SKY130_FD_SC_HD__AND4_4%D N_D_M1013_g N_D_M1009_g D N_D_c_177_n N_D_c_178_n
+ N_D_c_179_n PM_SKY130_FD_SC_HD__AND4_4%D
x_PM_SKY130_FD_SC_HD__AND4_4%A_27_47# N_A_27_47#_M1014_s N_A_27_47#_M1012_d
+ N_A_27_47#_M1008_d N_A_27_47#_c_219_n N_A_27_47#_M1001_g N_A_27_47#_M1000_g
+ N_A_27_47#_c_220_n N_A_27_47#_M1004_g N_A_27_47#_M1003_g N_A_27_47#_c_221_n
+ N_A_27_47#_M1010_g N_A_27_47#_M1006_g N_A_27_47#_c_222_n N_A_27_47#_M1015_g
+ N_A_27_47#_M1011_g N_A_27_47#_c_223_n N_A_27_47#_c_286_p N_A_27_47#_c_247_n
+ N_A_27_47#_c_262_n N_A_27_47#_c_254_n N_A_27_47#_c_231_n N_A_27_47#_c_224_n
+ N_A_27_47#_c_303_p N_A_27_47#_c_238_n N_A_27_47#_c_241_n N_A_27_47#_c_255_n
+ N_A_27_47#_c_225_n PM_SKY130_FD_SC_HD__AND4_4%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4_4%VPWR N_VPWR_M1012_s N_VPWR_M1005_d N_VPWR_M1013_d
+ N_VPWR_M1003_d N_VPWR_M1011_d N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n
+ N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n
+ N_VPWR_c_360_n VPWR N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_351_n PM_SKY130_FD_SC_HD__AND4_4%VPWR
x_PM_SKY130_FD_SC_HD__AND4_4%X N_X_M1001_d N_X_M1010_d N_X_M1000_s N_X_M1006_s
+ N_X_c_475_p N_X_c_425_n N_X_c_428_n N_X_c_429_n N_X_c_433_n N_X_c_422_n
+ N_X_c_478_p N_X_c_462_n N_X_c_443_n N_X_c_444_n N_X_c_448_n X X X N_X_c_420_n
+ X N_X_c_452_n N_X_c_424_n PM_SKY130_FD_SC_HD__AND4_4%X
x_PM_SKY130_FD_SC_HD__AND4_4%VGND N_VGND_M1009_d N_VGND_M1004_s N_VGND_M1015_s
+ N_VGND_c_494_n N_VGND_c_495_n N_VGND_c_496_n N_VGND_c_497_n VGND
+ N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n
+ N_VGND_c_503_n PM_SKY130_FD_SC_HD__AND4_4%VGND
cc_1 VNB N_A_c_72_n 0.0185096f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A 0.00891436f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_A_c_74_n 0.0427607f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB B 6.3097e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_5 VNB N_B_c_104_n 0.0210042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_B_c_105_n 0.00181441f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_7 VNB N_B_c_106_n 0.0161651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB C 0.00268159f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_9 VNB N_C_c_141_n 0.0267065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_C_c_142_n 0.0177266f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB D 0.00139692f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_12 VNB N_D_c_177_n 0.0245841f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_13 VNB N_D_c_178_n 2.98518e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_14 VNB N_D_c_179_n 0.0159796f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_15 VNB N_A_27_47#_c_219_n 0.0165762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_220_n 0.0157767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_221_n 0.0157735f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_222_n 0.0182736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_223_n 0.00252767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_224_n 0.00259677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_225_n 0.0646106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_351_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_420_n 0.00760238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB X 0.0245272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_494_n 0.00481578f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_26 VNB N_VGND_c_495_n 3.07214e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_27 VNB N_VGND_c_496_n 0.0102812f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=0.85
cc_28 VNB N_VGND_c_497_n 0.012064f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.16
cc_29 VNB N_VGND_c_498_n 0.0570348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_499_n 0.0137367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_500_n 0.010979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_501_n 0.00593471f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_502_n 0.00436184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_503_n 0.219538f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_A_M1012_g 0.0212723f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB A 0.0126677f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_37 VPB N_A_c_74_n 0.0107611f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_38 VPB N_B_M1005_g 0.0194119f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB N_B_c_104_n 0.0045041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_B_c_105_n 0.00273701f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_41 VPB N_C_M1008_g 0.0210672f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_42 VPB C 0.00269711f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_43 VPB N_C_c_141_n 0.00744369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_D_M1013_g 0.0213948f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_45 VPB N_D_c_177_n 0.00445545f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_46 VPB N_D_c_178_n 6.46466e-19 $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_47 VPB N_A_27_47#_M1000_g 0.0183432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_M1003_g 0.0184407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_M1006_g 0.0182226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_M1011_g 0.0209316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_223_n 0.00162909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_231_n 0.00173129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_225_n 0.0104094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_352_n 0.0109102f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_55 VPB N_VPWR_c_353_n 0.029337f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=0.85
cc_56 VPB N_VPWR_c_354_n 4.06069e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_355_n 0.0206692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_356_n 0.00278104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_357_n 0.0155238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_358_n 0.00161748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_359_n 0.0102077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_360_n 0.0250342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_361_n 0.0150713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_362_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_363_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_364_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_365_n 0.00353672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_351_n 0.0436365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_X_c_422_n 6.25997e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB X 0.0091442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_X_c_424_n 0.0116007f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 N_A_M1012_g N_B_M1005_g 0.0256632f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A_c_72_n B 5.15026e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A_c_74_n N_B_c_104_n 0.0303958f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_c_74_n N_B_c_105_n 3.05518e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_c_72_n N_B_c_106_n 0.0303958f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_77 A N_A_27_47#_M1014_s 0.00410489f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_78 N_A_c_72_n N_A_27_47#_c_223_n 0.0130195f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_M1012_g N_A_27_47#_c_223_n 0.0031298f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_80 A N_A_27_47#_c_223_n 0.0514557f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_c_74_n N_A_27_47#_c_223_n 0.00783512f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_c_72_n N_A_27_47#_c_238_n 0.0129857f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_83 A N_A_27_47#_c_238_n 0.0120742f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_84 N_A_c_74_n N_A_27_47#_c_238_n 0.00185364f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_M1012_g N_A_27_47#_c_241_n 0.00663833f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_86 A N_A_27_47#_c_241_n 0.0127418f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_87 A N_VPWR_M1012_s 0.00511762f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_88 N_A_M1012_g N_VPWR_c_353_n 0.00336877f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_89 A N_VPWR_c_353_n 0.0175645f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_c_74_n N_VPWR_c_353_n 0.00223275f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_M1012_g N_VPWR_c_354_n 6.13039e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_M1012_g N_VPWR_c_361_n 0.00585385f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_M1012_g N_VPWR_c_351_n 0.0114182f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_c_72_n N_VGND_c_498_n 0.00357877f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_c_72_n N_VGND_c_503_n 0.00614193f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 A N_VGND_c_503_n 0.00238628f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_97 N_B_M1005_g N_C_M1008_g 0.0249677f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_98 B C 0.0516879f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_99 N_B_c_104_n C 2.37819e-19 $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B_c_106_n C 3.88615e-19 $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B_c_104_n N_C_c_141_n 0.0204718f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B_c_105_n N_C_c_141_n 0.0025946f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_103 B N_C_c_142_n 0.00334798f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_104 N_B_c_106_n N_C_c_142_n 0.0305802f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B_M1005_g N_A_27_47#_c_223_n 0.0035847f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_106 B N_A_27_47#_c_223_n 0.0250859f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_107 N_B_c_105_n N_A_27_47#_c_223_n 0.0251942f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_108 N_B_c_106_n N_A_27_47#_c_223_n 0.00463205f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B_M1005_g N_A_27_47#_c_247_n 0.0156401f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_110 N_B_c_104_n N_A_27_47#_c_247_n 5.45329e-19 $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_111 N_B_c_105_n N_A_27_47#_c_247_n 0.0289659f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_112 B N_A_27_47#_c_238_n 0.0108787f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_113 N_B_c_106_n N_A_27_47#_c_238_n 0.00556374f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B_M1005_g N_VPWR_c_354_n 0.00895008f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B_M1005_g N_VPWR_c_361_n 0.00544582f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B_M1005_g N_VPWR_c_351_n 0.00914755f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_117 B A_188_47# 0.00511697f $X=1.07 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_118 B N_VGND_c_498_n 0.0105283f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_119 N_B_c_106_n N_VGND_c_498_n 0.0052149f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_120 B N_VGND_c_503_n 0.012118f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_121 N_B_c_106_n N_VGND_c_503_n 0.00919877f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_122 N_C_M1008_g N_D_M1013_g 0.0230105f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_123 C D 0.0386614f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_124 N_C_c_142_n D 2.20254e-19 $X=1.452 $Y=0.995 $X2=0 $Y2=0
cc_125 C N_D_c_177_n 0.00230308f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_126 N_C_c_141_n N_D_c_177_n 0.01913f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_127 N_C_c_142_n N_D_c_177_n 6.69542e-19 $X=1.452 $Y=0.995 $X2=0 $Y2=0
cc_128 N_C_c_141_n N_D_c_178_n 3.43759e-19 $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_129 C N_D_c_179_n 0.00751095f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_130 N_C_c_142_n N_D_c_179_n 0.021064f $X=1.452 $Y=0.995 $X2=0 $Y2=0
cc_131 N_C_M1008_g N_A_27_47#_c_247_n 0.0199527f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_132 C N_A_27_47#_c_247_n 0.0019493f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_133 C N_A_27_47#_c_254_n 0.0044525f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_134 C N_A_27_47#_c_255_n 0.015435f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_135 N_C_c_141_n N_A_27_47#_c_255_n 0.00134283f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_136 N_C_M1008_g N_VPWR_c_354_n 0.00991765f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_137 N_C_M1008_g N_VPWR_c_355_n 0.00544582f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_138 N_C_M1008_g N_VPWR_c_351_n 0.00949094f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_139 C A_285_47# 0.00997671f $X=1.53 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_140 C N_VGND_c_498_n 0.00850155f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_141 N_C_c_142_n N_VGND_c_498_n 0.00573703f $X=1.452 $Y=0.995 $X2=0 $Y2=0
cc_142 C N_VGND_c_503_n 0.00983203f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_143 N_C_c_142_n N_VGND_c_503_n 0.0110688f $X=1.452 $Y=0.995 $X2=0 $Y2=0
cc_144 D N_A_27_47#_c_219_n 0.00349482f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_145 N_D_c_177_n N_A_27_47#_c_219_n 0.0230918f $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_146 N_D_c_178_n N_A_27_47#_c_219_n 0.00140868f $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_147 N_D_c_179_n N_A_27_47#_c_219_n 0.0187559f $X=1.99 $Y=0.965 $X2=0 $Y2=0
cc_148 N_D_M1013_g N_A_27_47#_M1000_g 0.0226397f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_149 N_D_M1013_g N_A_27_47#_c_262_n 0.00942752f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_150 N_D_M1013_g N_A_27_47#_c_254_n 0.0175363f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_151 D N_A_27_47#_c_254_n 0.00250919f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_152 N_D_c_177_n N_A_27_47#_c_254_n 0.00173976f $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_153 N_D_c_178_n N_A_27_47#_c_254_n 0.0107433f $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_154 N_D_M1013_g N_A_27_47#_c_231_n 0.0032894f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_155 N_D_c_178_n N_A_27_47#_c_231_n 0.00139276f $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_156 N_D_c_177_n N_A_27_47#_c_224_n 0.001398f $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_157 N_D_c_178_n N_A_27_47#_c_224_n 0.0170805f $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_158 N_D_c_178_n N_A_27_47#_c_225_n 2.13568e-19 $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_159 N_D_M1013_g N_VPWR_c_354_n 9.90489e-19 $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_160 N_D_M1013_g N_VPWR_c_355_n 0.00585385f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_161 N_D_M1013_g N_VPWR_c_356_n 0.00314448f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_162 N_D_M1013_g N_VPWR_c_351_n 0.0110904f $X=1.93 $Y=1.985 $X2=0 $Y2=0
cc_163 D N_VGND_M1009_d 0.00277396f $X=1.98 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_164 D N_VGND_c_494_n 0.00664987f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_165 N_D_c_177_n N_VGND_c_494_n 2.5741e-19 $X=1.99 $Y=1.16 $X2=0 $Y2=0
cc_166 N_D_c_179_n N_VGND_c_494_n 0.00314761f $X=1.99 $Y=0.965 $X2=0 $Y2=0
cc_167 D N_VGND_c_498_n 0.00161159f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_168 N_D_c_179_n N_VGND_c_498_n 0.00483472f $X=1.99 $Y=0.965 $X2=0 $Y2=0
cc_169 D N_VGND_c_503_n 0.00326954f $X=1.98 $Y=0.765 $X2=0 $Y2=0
cc_170 N_D_c_179_n N_VGND_c_503_n 0.00784665f $X=1.99 $Y=0.965 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_247_n N_VPWR_M1005_d 0.00456664f $X=1.455 $Y=1.58 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_254_n N_VPWR_M1013_d 0.00717557f $X=2.245 $Y=1.58 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_247_n N_VPWR_c_354_n 0.0122127f $X=1.455 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_262_n N_VPWR_c_355_n 0.0123145f $X=1.56 $Y=1.96 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1000_g N_VPWR_c_356_n 0.0103414f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_27_47#_M1003_g N_VPWR_c_356_n 4.71995e-19 $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_254_n N_VPWR_c_356_n 0.0177361f $X=2.245 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A_27_47#_M1000_g N_VPWR_c_357_n 0.00505556f $X=2.41 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1003_g N_VPWR_c_357_n 0.00541359f $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_M1003_g N_VPWR_c_358_n 0.00143109f $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1006_g N_VPWR_c_358_n 0.0106721f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1011_g N_VPWR_c_358_n 6.27883e-19 $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_M1006_g N_VPWR_c_360_n 6.0901e-19 $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1011_g N_VPWR_c_360_n 0.0112954f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_286_p N_VPWR_c_361_n 0.012815f $X=0.68 $Y=1.96 $X2=0 $Y2=0
cc_186 N_A_27_47#_M1006_g N_VPWR_c_362_n 0.0046653f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_27_47#_M1011_g N_VPWR_c_362_n 0.0046653f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_27_47#_M1012_d N_VPWR_c_351_n 0.00423495f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_M1008_d N_VPWR_c_351_n 0.0118231f $X=1.425 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1000_g N_VPWR_c_351_n 0.00850607f $X=2.41 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1003_g N_VPWR_c_351_n 0.00950154f $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1006_g N_VPWR_c_351_n 0.00789179f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1011_g N_VPWR_c_351_n 0.00789179f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_286_p N_VPWR_c_351_n 0.00801045f $X=0.68 $Y=1.96 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_262_n N_VPWR_c_351_n 0.00724021f $X=1.56 $Y=1.96 $X2=0 $Y2=0
cc_196 N_A_27_47#_M1003_g N_X_c_425_n 0.00163365f $X=2.83 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_224_n N_X_c_425_n 0.00266928f $X=2.69 $Y=1.19 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_225_n N_X_c_425_n 7.69814e-19 $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_47#_M1003_g N_X_c_428_n 0.00591341f $X=2.83 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_220_n N_X_c_429_n 0.0115451f $X=2.83 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_221_n N_X_c_429_n 0.0119773f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_303_p N_X_c_429_n 0.0279003f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_225_n N_X_c_429_n 0.00207823f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_224_n N_X_c_433_n 0.00835992f $X=2.69 $Y=1.19 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_303_p N_X_c_433_n 6.00526e-19 $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_225_n N_X_c_433_n 0.0021683f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_27_47#_M1000_g N_X_c_422_n 0.0012453f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1003_g N_X_c_422_n 0.00210743f $X=2.83 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_254_n N_X_c_422_n 0.0123221f $X=2.245 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_231_n N_X_c_422_n 6.66456e-19 $X=2.33 $Y=1.495 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_224_n N_X_c_422_n 0.00580825f $X=2.69 $Y=1.19 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_303_p N_X_c_422_n 0.00475276f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_225_n N_X_c_422_n 0.00118648f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_222_n N_X_c_443_n 0.0151481f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_27_47#_M1000_g N_X_c_444_n 0.00274552f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_27_47#_M1003_g N_X_c_444_n 0.00332394f $X=2.83 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_27_47#_M1006_g N_X_c_444_n 4.84566e-19 $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_254_n N_X_c_444_n 6.60394e-19 $X=2.245 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_303_p N_X_c_448_n 0.009137f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_225_n N_X_c_448_n 0.00216957f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_222_n X 0.0244128f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_303_p X 0.0156897f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_27_47#_M1003_g N_X_c_452_n 0.0107675f $X=2.83 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_27_47#_M1006_g N_X_c_452_n 0.014091f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_303_p N_X_c_452_n 0.0470531f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_225_n N_X_c_452_n 0.00205251f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1011_g N_X_c_424_n 0.0218965f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_225_n N_X_c_424_n 0.00207434f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_223_n A_109_47# 0.00292611f $X=0.585 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_230 N_A_27_47#_c_238_n A_109_47# 0.00449329f $X=0.585 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_231 N_A_27_47#_c_219_n N_VGND_c_494_n 0.00165501f $X=2.41 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_224_n N_VGND_c_494_n 0.0023793f $X=2.69 $Y=1.19 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_219_n N_VGND_c_495_n 5.22831e-19 $X=2.41 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_220_n N_VGND_c_495_n 0.00676788f $X=2.83 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_221_n N_VGND_c_495_n 0.00669652f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_222_n N_VGND_c_495_n 5.10275e-19 $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_221_n N_VGND_c_497_n 5.10275e-19 $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_222_n N_VGND_c_497_n 0.00779801f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_238_n N_VGND_c_498_n 0.0289623f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_219_n N_VGND_c_499_n 0.00583607f $X=2.41 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_220_n N_VGND_c_499_n 0.00339951f $X=2.83 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_221_n N_VGND_c_500_n 0.00339951f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_222_n N_VGND_c_500_n 0.00339951f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_M1014_s N_VGND_c_503_n 0.00231556f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_219_n N_VGND_c_503_n 0.0105612f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_220_n N_VGND_c_503_n 0.00395374f $X=2.83 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_221_n N_VGND_c_503_n 0.00395374f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_222_n N_VGND_c_503_n 0.00395374f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_238_n N_VGND_c_503_n 0.0179555f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_250 N_VPWR_c_351_n N_X_M1000_s 0.0038878f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_251 N_VPWR_c_351_n N_X_M1006_s 0.00562358f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_252 N_VPWR_c_357_n N_X_c_428_n 0.0151443f $X=2.955 $Y=2.72 $X2=0 $Y2=0
cc_253 N_VPWR_c_351_n N_X_c_428_n 0.00934466f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_254 N_VPWR_c_362_n N_X_c_462_n 0.0114421f $X=3.715 $Y=2.72 $X2=0 $Y2=0
cc_255 N_VPWR_c_351_n N_X_c_462_n 0.00647979f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_256 N_VPWR_M1011_d X 6.00252e-19 $X=3.745 $Y=1.485 $X2=0 $Y2=0
cc_257 N_VPWR_M1003_d N_X_c_452_n 0.003186f $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_258 N_VPWR_c_358_n N_X_c_452_n 0.01423f $X=3.04 $Y=2 $X2=0 $Y2=0
cc_259 N_VPWR_M1011_d N_X_c_424_n 0.00392904f $X=3.745 $Y=1.485 $X2=0 $Y2=0
cc_260 N_VPWR_c_360_n N_X_c_424_n 0.022628f $X=3.88 $Y=2 $X2=0 $Y2=0
cc_261 N_X_c_429_n N_VGND_M1004_s 0.00336061f $X=3.375 $Y=0.725 $X2=0 $Y2=0
cc_262 N_X_c_420_n N_VGND_M1015_s 0.00291581f $X=3.925 $Y=0.81 $X2=0 $Y2=0
cc_263 X N_VGND_M1015_s 3.27674e-19 $X=3.905 $Y=0.85 $X2=0 $Y2=0
cc_264 N_X_c_429_n N_VGND_c_495_n 0.0159876f $X=3.375 $Y=0.725 $X2=0 $Y2=0
cc_265 N_X_c_443_n N_VGND_c_497_n 0.00203332f $X=3.8 $Y=0.725 $X2=0 $Y2=0
cc_266 N_X_c_420_n N_VGND_c_497_n 0.0205549f $X=3.925 $Y=0.81 $X2=0 $Y2=0
cc_267 N_X_c_475_p N_VGND_c_499_n 0.0112345f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_268 N_X_c_429_n N_VGND_c_499_n 0.0024142f $X=3.375 $Y=0.725 $X2=0 $Y2=0
cc_269 N_X_c_429_n N_VGND_c_500_n 0.0024142f $X=3.375 $Y=0.725 $X2=0 $Y2=0
cc_270 N_X_c_478_p N_VGND_c_500_n 0.0112345f $X=3.46 $Y=0.42 $X2=0 $Y2=0
cc_271 N_X_c_443_n N_VGND_c_500_n 0.0024142f $X=3.8 $Y=0.725 $X2=0 $Y2=0
cc_272 N_X_M1001_d N_VGND_c_503_n 0.00406206f $X=2.485 $Y=0.235 $X2=0 $Y2=0
cc_273 N_X_M1010_d N_VGND_c_503_n 0.00250055f $X=3.325 $Y=0.235 $X2=0 $Y2=0
cc_274 N_X_c_475_p N_VGND_c_503_n 0.00643596f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_275 N_X_c_429_n N_VGND_c_503_n 0.00979235f $X=3.375 $Y=0.725 $X2=0 $Y2=0
cc_276 N_X_c_478_p N_VGND_c_503_n 0.00643596f $X=3.46 $Y=0.42 $X2=0 $Y2=0
cc_277 N_X_c_443_n N_VGND_c_503_n 0.0045422f $X=3.8 $Y=0.725 $X2=0 $Y2=0
cc_278 N_X_c_420_n N_VGND_c_503_n 0.00141083f $X=3.925 $Y=0.81 $X2=0 $Y2=0
cc_279 A_109_47# N_VGND_c_503_n 0.0061253f $X=0.545 $Y=0.235 $X2=1.55 $Y2=1.96
cc_280 A_188_47# N_VGND_c_503_n 0.00404868f $X=0.94 $Y=0.235 $X2=0 $Y2=0
cc_281 A_285_47# N_VGND_c_503_n 0.00936282f $X=1.425 $Y=0.235 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__xor3_2.spice
* Created: Thu Aug 27 14:50:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__xor3_2.pex.spice"
.subckt sky130_fd_sc_hd__xor3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1010 N_X_M1010_d N_A_120_21#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1010_d N_A_120_21#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.175105 PD=0.92 PS=1.36075 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75000.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1019 N_A_358_93#_M1019_d N_C_M1019_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1764 AS=0.113145 PD=1.68 PS=0.879252 NRD=38.568 NRS=61.248 M=1 R=2.8
+ SA=75001.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_120_21#_M1005_d N_C_M1005_g N_A_496_49#_M1005_s VNB NSHORT L=0.15
+ W=0.64 AD=0.128 AS=0.1728 PD=1.04 PS=1.82 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1021 N_A_478_325#_M1021_d N_A_358_93#_M1021_g N_A_120_21#_M1005_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3168 AS=0.128 PD=2.27 PS=1.04 NRD=38.436 NRS=23.436 M=1
+ R=4.26667 SA=75000.7 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_919_297#_M1001_d N_B_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1653 AS=0.195 PD=1.82 PS=1.9 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_496_49#_M1008_d N_B_M1008_g N_A_1023_365#_M1008_s VNB NSHORT L=0.15
+ W=0.64 AD=0.221766 AS=0.1628 PD=1.50943 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1004 N_A_1290_49#_M1004_d N_A_919_297#_M1004_g N_A_496_49#_M1008_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.152666 AS=0.145534 PD=1.0183 PS=0.990566 NRD=88.14
+ NRS=95.712 M=1 R=2.8 SA=75000.9 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1013 N_A_478_325#_M1013_d N_B_M1013_g N_A_1290_49#_M1004_d VNB NSHORT L=0.15
+ W=0.64 AD=0.145368 AS=0.232634 PD=1.13548 PS=1.5517 NRD=0.936 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_1023_365#_M1023_d N_A_919_297#_M1023_g N_A_478_325#_M1013_d VNB
+ NSHORT L=0.15 W=0.6 AD=0.106452 AS=0.136282 PD=0.958065 PS=1.06452 NRD=15
+ NRS=32.988 M=1 R=4 SA=75001.9 SB=75001.1 A=0.09 P=1.5 MULT=1
MM1022 N_VGND_M1022_d N_A_M1022_g N_A_1023_365#_M1023_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.113548 PD=0.91 PS=1.02194 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_1290_49#_M1020_d N_A_1023_365#_M1020_g N_VGND_M1022_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_120_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_120_21#_M1006_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.257927 AS=0.135 PD=1.76829 PS=1.27 NRD=15.7403 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1007 N_A_358_93#_M1007_d N_C_M1007_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1792 AS=0.165073 PD=1.84 PS=1.13171 NRD=0 NRS=62.449 M=1 R=4.26667
+ SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_120_21#_M1009_d N_C_M1009_g N_A_478_325#_M1009_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1596 AS=0.2688 PD=1.22 PS=2.32 NRD=9.3772 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1000 N_A_496_49#_M1000_d N_A_358_93#_M1000_g N_A_120_21#_M1009_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.441 AS=0.1596 PD=2.73 PS=1.22 NRD=57.4452 NRS=14.0658 M=1
+ R=5.6 SA=75000.8 SB=75000.4 A=0.126 P=1.98 MULT=1
MM1002 N_A_919_297#_M1002_d N_B_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2526 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1018 N_A_478_325#_M1018_d N_B_M1018_g N_A_1023_365#_M1018_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.278335 AS=0.3536 PD=1.64595 PS=2.53 NRD=46.886 NRS=37.5088 M=1
+ R=5.6 SA=75000.3 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1016 N_A_1290_49#_M1016_d N_A_919_297#_M1016_g N_A_478_325#_M1018_d VPB
+ PHIGHVT L=0.15 W=0.64 AD=0.246 AS=0.212065 PD=1.525 PS=1.25405 NRD=138.511
+ NRS=40.0107 M=1 R=4.26667 SA=75001.1 SB=75002 A=0.096 P=1.58 MULT=1
MM1014 N_A_496_49#_M1014_d N_B_M1014_g N_A_1290_49#_M1016_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.126097 AS=0.246 PD=1.04216 PS=1.525 NRD=43.7143 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_1023_365#_M1011_d N_A_919_297#_M1011_g N_A_496_49#_M1014_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.156587 AS=0.165503 PD=1.23717 PS=1.36784
+ NRD=30.8108 NRS=0 M=1 R=5.6 SA=75001.6 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g N_A_1023_365#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.186413 PD=1.27 PS=1.47283 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_A_1290_49#_M1012_d N_A_1023_365#_M1012_g N_VPWR_M1017_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.265 AS=0.135 PD=2.53 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.3759 P=22.37
*
.include "sky130_fd_sc_hd__xor3_2.pxi.spice"
*
.ends
*
*

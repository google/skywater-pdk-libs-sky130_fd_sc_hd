* File: sky130_fd_sc_hd__sedfxtp_4.pex.spice
* Created: Thu Aug 27 14:48:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%CLK 1 2 3 5 6 8 11 13
c40 1 0 2.71124e-20 $X=0.31 $Y=1.325
r41 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r42 9 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.47 $Y2=1.665
r43 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r44 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r45 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r46 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r47 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r48 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r49 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_27_47# 1 2 9 13 17 21 25 27 31 35 39 40
+ 41 44 46 48 51 54 56 57 58 59 60 67 69 74 82 85 89
c275 89 0 1.92554e-19 $X=10.175 $Y=1.41
c276 51 0 1.74912e-19 $X=7.28 $Y=0.87
c277 48 0 1.43548e-19 $X=7.45 $Y=0.845
c278 44 0 1.8506e-19 $X=0.73 $Y=1.795
c279 41 0 5.65522e-20 $X=0.615 $Y=1.88
r280 88 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.175 $Y=1.41
+ $X2=10.175 $Y2=1.575
r281 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.175
+ $Y=1.41 $X2=10.175 $Y2=1.41
r282 85 88 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=10.175 $Y=1.32
+ $X2=10.175 $Y2=1.41
r283 79 82 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=7.61 $Y=1.74
+ $X2=7.705 $Y2=1.74
r284 70 89 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=10.185 $Y=1.87
+ $X2=10.185 $Y2=1.41
r285 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.185 $Y=1.87
+ $X2=10.185 $Y2=1.87
r286 67 96 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=7.595 $Y=1.83
+ $X2=7.535 $Y2=1.83
r287 67 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.705
+ $Y=1.74 $X2=7.705 $Y2=1.74
r288 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=1.87
+ $X2=7.595 $Y2=1.87
r289 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=1.87
+ $X2=0.72 $Y2=1.87
r290 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.74 $Y=1.87
+ $X2=7.595 $Y2=1.87
r291 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.04 $Y=1.87
+ $X2=10.185 $Y2=1.87
r292 59 60 2.84653 $w=1.4e-07 $l=2.3e-06 $layer=MET1_cond $X=10.04 $Y=1.87
+ $X2=7.74 $Y2=1.87
r293 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.865 $Y=1.87
+ $X2=0.72 $Y2=1.87
r294 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=1.87
+ $X2=7.595 $Y2=1.87
r295 57 58 8.14974 $w=1.4e-07 $l=6.585e-06 $layer=MET1_cond $X=7.45 $Y=1.87
+ $X2=0.865 $Y2=1.87
r296 54 96 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.535 $Y=1.655
+ $X2=7.535 $Y2=1.83
r297 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.535 $Y=0.955
+ $X2=7.535 $Y2=1.655
r298 51 77 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.28 $Y=0.87
+ $X2=7.28 $Y2=0.735
r299 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.28
+ $Y=0.87 $X2=7.28 $Y2=0.87
r300 48 53 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.45 $Y=0.845
+ $X2=7.535 $Y2=0.955
r301 48 50 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=7.45 $Y=0.845
+ $X2=7.28 $Y2=0.845
r302 47 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r303 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r304 44 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r305 44 46 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r306 43 46 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.73 $Y=0.805
+ $X2=0.73 $Y2=1.235
r307 42 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r308 41 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r309 41 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.345 $Y2=1.88
r310 39 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.73 $Y2=0.805
r311 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r312 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r313 33 35 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r314 29 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=10.81 $Y=1.245
+ $X2=10.81 $Y2=0.415
r315 28 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.31 $Y=1.32
+ $X2=10.175 $Y2=1.32
r316 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.735 $Y=1.32
+ $X2=10.81 $Y2=1.245
r317 27 28 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=10.735 $Y=1.32
+ $X2=10.31 $Y2=1.32
r318 25 90 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=10.18 $Y=2.275
+ $X2=10.18 $Y2=1.575
r319 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.61 $Y=1.905
+ $X2=7.61 $Y2=1.74
r320 19 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.61 $Y=1.905
+ $X2=7.61 $Y2=2.275
r321 17 77 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.29 $Y=0.415
+ $X2=7.29 $Y2=0.735
r322 11 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r323 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r324 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r325 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r326 2 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r327 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%D 3 7 9 12 13 16
c51 7 0 5.26342e-20 $X=1.83 $Y=2.165
r52 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.78
+ $Y=1.145 $X2=1.78 $Y2=1.145
r53 11 16 70.9845 $w=3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.765 $Y=1.5
+ $X2=1.765 $Y2=1.145
r54 11 12 43.217 $w=3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.765 $Y=1.5 $X2=1.765
+ $Y2=1.65
r55 9 16 2.99935 $w=3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.765 $Y=1.13 $X2=1.765
+ $Y2=1.145
r56 9 10 43.217 $w=3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.765 $Y=1.13 $X2=1.765
+ $Y2=0.98
r57 7 12 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.83 $Y=2.165
+ $X2=1.83 $Y2=1.65
r58 3 10 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.83 $Y=0.445
+ $X2=1.83 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_423_343# 1 2 7 9 12 16 20 23 26 27 36
c88 27 0 1.67735e-19 $X=3.55 $Y=1.01
c89 23 0 5.26342e-20 $X=2.932 $Y=1.355
c90 20 0 1.1082e-19 $X=2.92 $Y=0.51
r91 30 33 10.7351 $w=3.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.58 $Y=1.537
+ $X2=2.92 $Y2=1.537
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.52 $X2=2.58 $Y2=1.52
r93 27 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.01
+ $X2=3.55 $Y2=0.845
r94 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.01 $X2=3.55 $Y2=1.01
r95 24 36 0.565906 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=3.085 $Y=1.01
+ $X2=2.932 $Y2=1.01
r96 24 26 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.085 $Y=1.01
+ $X2=3.55 $Y2=1.01
r97 23 33 0.378885 $w=3.63e-07 $l=1.2e-08 $layer=LI1_cond $X=2.932 $Y=1.537
+ $X2=2.92 $Y2=1.537
r98 22 36 6.17543 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=2.932 $Y=1.175
+ $X2=2.932 $Y2=1.01
r99 22 23 6.8013 $w=3.03e-07 $l=1.8e-07 $layer=LI1_cond $X=2.932 $Y=1.175
+ $X2=2.932 $Y2=1.355
r100 18 36 6.17543 $w=2.65e-07 $l=1.83916e-07 $layer=LI1_cond $X=2.892 $Y=0.845
+ $X2=2.932 $Y2=1.01
r101 18 20 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=2.892 $Y=0.845
+ $X2=2.892 $Y2=0.51
r102 14 33 1.32393 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=2.92 $Y=1.72
+ $X2=2.92 $Y2=1.537
r103 14 16 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.92 $Y=1.72
+ $X2=2.92 $Y2=1.99
r104 12 40 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.57 $Y=0.445
+ $X2=3.57 $Y2=0.845
r105 7 31 69.3653 $w=2.71e-07 $l=4.76833e-07 $layer=POLY_cond $X=2.19 $Y=1.77
+ $X2=2.58 $Y2=1.577
r106 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.19 $Y=1.77
+ $X2=2.19 $Y2=2.165
r107 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.795
+ $Y=1.845 $X2=2.92 $Y2=1.99
r108 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.92 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%DE 3 5 6 9 12 15 17 21 23 24 25
c85 6 0 1.1082e-19 $X=2.455 $Y=0.925
r86 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.01 $X2=2.29 $Y2=1.01
r87 27 29 13.5393 $w=3.56e-07 $l=1e-07 $layer=POLY_cond $X=2.19 $Y=0.992
+ $X2=2.29 $Y2=0.992
r88 25 30 5.12336 $w=3.81e-07 $l=1.6e-07 $layer=LI1_cond $X=2.337 $Y=0.85
+ $X2=2.337 $Y2=1.01
r89 19 21 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.57 $Y=1.61
+ $X2=3.57 $Y2=2.165
r90 18 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.205 $Y=1.535
+ $X2=3.13 $Y2=1.535
r91 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.495 $Y=1.535
+ $X2=3.57 $Y2=1.61
r92 17 18 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.495 $Y=1.535
+ $X2=3.205 $Y2=1.535
r93 13 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.61
+ $X2=3.13 $Y2=1.535
r94 13 15 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.13 $Y=1.61
+ $X2=3.13 $Y2=2.165
r95 12 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.46
+ $X2=3.13 $Y2=1.535
r96 11 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1 $X2=3.13
+ $Y2=0.925
r97 11 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.13 $Y=1 $X2=3.13
+ $Y2=1.46
r98 7 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=0.85 $X2=3.13
+ $Y2=0.925
r99 7 9 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.13 $Y=0.85 $X2=3.13
+ $Y2=0.445
r100 6 29 38.8573 $w=3.56e-07 $l=1.95653e-07 $layer=POLY_cond $X=2.455 $Y=0.925
+ $X2=2.29 $Y2=0.992
r101 5 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=0.925
+ $X2=3.13 $Y2=0.925
r102 5 6 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.055 $Y=0.925 $X2=2.455
+ $Y2=0.925
r103 1 27 23.0368 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.19 $Y=0.81
+ $X2=2.19 $Y2=0.992
r104 1 3 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.19 $Y=0.81 $X2=2.19
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_791_264# 1 2 9 13 17 21 23 26 30 34 40
+ 41 44 46 47 48 51 54 55
c190 47 0 6.12178e-20 $X=11.94 $Y=0.85
c191 21 0 2.06462e-20 $X=11.285 $Y=0.445
c192 9 0 5.58337e-20 $X=4.08 $Y=0.445
r193 60 62 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=11.17 $Y=1.74
+ $X2=11.285 $Y2=1.74
r194 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.085 $Y=0.85
+ $X2=12.085 $Y2=0.85
r195 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.89 $Y=0.85
+ $X2=3.89 $Y2=0.85
r196 48 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.035 $Y=0.85
+ $X2=3.89 $Y2=0.85
r197 47 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.94 $Y=0.85
+ $X2=12.085 $Y2=0.85
r198 47 48 9.7834 $w=1.4e-07 $l=7.905e-06 $layer=MET1_cond $X=11.94 $Y=0.85
+ $X2=4.035 $Y2=0.85
r199 46 55 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=12.085 $Y=0.825
+ $X2=12.085 $Y2=0.85
r200 43 55 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=12.085 $Y=1.53
+ $X2=12.085 $Y2=0.85
r201 43 44 6.82437 $w=2.65e-07 $l=2.21346e-07 $layer=LI1_cond $X=12.085 $Y=1.53
+ $X2=12.01 $Y2=1.717
r202 41 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=1.485
+ $X2=4.09 $Y2=1.65
r203 41 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=1.485
+ $X2=4.09 $Y2=1.32
r204 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.485 $X2=4.09 $Y2=1.485
r205 37 51 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.89 $Y=1.32
+ $X2=3.89 $Y2=0.85
r206 36 40 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.89 $Y=1.485 $X2=4.09
+ $Y2=1.485
r207 36 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=1.485
+ $X2=3.89 $Y2=1.32
r208 32 46 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.015 $Y=0.66
+ $X2=12.015 $Y2=0.825
r209 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.015 $Y=0.66
+ $X2=12.015 $Y2=0.385
r210 28 44 6.82437 $w=2.65e-07 $l=1.88e-07 $layer=LI1_cond $X=12.01 $Y=1.905
+ $X2=12.01 $Y2=1.717
r211 28 30 2.88111 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=12.01 $Y=1.905
+ $X2=12.01 $Y2=1.99
r212 26 62 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=11.365 $Y=1.74
+ $X2=11.285 $Y2=1.74
r213 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.365
+ $Y=1.74 $X2=11.365 $Y2=1.74
r214 23 44 0.127723 $w=3.75e-07 $l=1.7e-07 $layer=LI1_cond $X=11.84 $Y=1.717
+ $X2=12.01 $Y2=1.717
r215 23 25 14.5976 $w=3.73e-07 $l=4.75e-07 $layer=LI1_cond $X=11.84 $Y=1.717
+ $X2=11.365 $Y2=1.717
r216 19 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.285 $Y=1.575
+ $X2=11.285 $Y2=1.74
r217 19 21 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=11.285 $Y=1.575
+ $X2=11.285 $Y2=0.445
r218 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.17 $Y=1.905
+ $X2=11.17 $Y2=1.74
r219 15 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=11.17 $Y=1.905
+ $X2=11.17 $Y2=2.275
r220 13 59 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.08 $Y=2.165
+ $X2=4.08 $Y2=1.65
r221 9 58 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.08 $Y=0.445
+ $X2=4.08 $Y2=1.32
r222 2 30 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.88
+ $Y=1.845 $X2=12.005 $Y2=1.99
r223 1 34 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=11.89
+ $Y=0.235 $X2=12.015 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_885_21# 1 2 7 9 10 11 13 16 18 21 28 30
+ 31 35 36 39 40
c129 36 0 4.70699e-20 $X=6.5 $Y=1.52
c130 21 0 1.41479e-20 $X=5.13 $Y=0.34
c131 18 0 5.87547e-20 $X=5.26 $Y=0.385
r132 36 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.5 $Y=1.52
+ $X2=6.5 $Y2=1.685
r133 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.5
+ $Y=1.52 $X2=6.5 $Y2=1.52
r134 33 35 17.4682 $w=1.98e-07 $l=3.15e-07 $layer=LI1_cond $X=6.485 $Y=1.835
+ $X2=6.485 $Y2=1.52
r135 32 39 2.83584 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=5.59 $Y=1.92
+ $X2=5.372 $Y2=1.92
r136 31 33 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.385 $Y=1.92
+ $X2=6.485 $Y2=1.835
r137 31 32 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.385 $Y=1.92
+ $X2=5.59 $Y2=1.92
r138 30 39 3.64284 $w=2.55e-07 $l=1.70276e-07 $layer=LI1_cond $X=5.505 $Y=1.835
+ $X2=5.372 $Y2=1.92
r139 30 40 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.505 $Y=1.835
+ $X2=5.505 $Y2=0.935
r140 26 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.425 $Y=0.77
+ $X2=5.425 $Y2=0.935
r141 26 28 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=5.425 $Y=0.77
+ $X2=5.425 $Y2=0.75
r142 25 28 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.425 $Y=0.515
+ $X2=5.425 $Y2=0.75
r143 21 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=0.34
+ $X2=5.13 $Y2=0.505
r144 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=0.34 $X2=5.13 $Y2=0.34
r145 18 25 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=5.26 $Y=0.385
+ $X2=5.425 $Y2=0.515
r146 18 20 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.26 $Y=0.385
+ $X2=5.13 $Y2=0.385
r147 16 46 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.56 $Y=2.165
+ $X2=6.56 $Y2=1.685
r148 13 43 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.07 $Y=0.765
+ $X2=5.07 $Y2=0.505
r149 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.995 $Y=0.84
+ $X2=5.07 $Y2=0.765
r150 10 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.995 $Y=0.84
+ $X2=4.575 $Y2=0.84
r151 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.5 $Y=0.765
+ $X2=4.575 $Y2=0.84
r152 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.5 $Y=0.765 $X2=4.5
+ $Y2=0.445
r153 2 39 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=5.195
+ $Y=1.845 $X2=5.32 $Y2=2
r154 1 28 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.3
+ $Y=0.595 $X2=5.425 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%SCD 3 7 9 12
c48 3 0 1.76561e-19 $X=6.055 $Y=0.805
r49 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.02 $Y=1.52
+ $X2=6.02 $Y2=1.685
r50 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.02 $Y=1.52
+ $X2=6.02 $Y2=1.355
r51 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.02
+ $Y=1.52 $X2=6.02 $Y2=1.52
r52 9 13 8.67485 $w=4.53e-07 $l=3.3e-07 $layer=LI1_cond $X=5.987 $Y=1.19
+ $X2=5.987 $Y2=1.52
r53 7 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.08 $Y=2.165
+ $X2=6.08 $Y2=1.685
r54 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.055 $Y=0.805
+ $X2=6.055 $Y2=1.355
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%SCE 3 5 6 9 14 15 16 19 21 25 26
r94 24 26 67.5777 $w=2.96e-07 $l=4.15e-07 $layer=POLY_cond $X=5.12 $Y=1.332
+ $X2=5.535 $Y2=1.332
r95 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.44 $X2=5.12 $Y2=1.44
r96 21 25 4.60977 $w=2.23e-07 $l=9e-08 $layer=LI1_cond $X=5.137 $Y=1.53
+ $X2=5.137 $Y2=1.44
r97 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.415 $Y=0.255
+ $X2=6.415 $Y2=0.805
r98 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.34 $Y=0.18
+ $X2=6.415 $Y2=0.255
r99 15 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=6.34 $Y=0.18
+ $X2=5.71 $Y2=0.18
r100 12 26 16.2838 $w=2.96e-07 $l=2.87687e-07 $layer=POLY_cond $X=5.635 $Y=1.09
+ $X2=5.535 $Y2=1.332
r101 12 14 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.635 $Y=1.09
+ $X2=5.635 $Y2=0.805
r102 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.635 $Y=0.255
+ $X2=5.71 $Y2=0.18
r103 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.635 $Y=0.255
+ $X2=5.635 $Y2=0.805
r104 7 26 18.6531 $w=1.5e-07 $l=2.43e-07 $layer=POLY_cond $X=5.535 $Y=1.575
+ $X2=5.535 $Y2=1.332
r105 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.535 $Y=1.575
+ $X2=5.535 $Y2=2.165
r106 5 24 38.5718 $w=2.96e-07 $l=2.36525e-07 $layer=POLY_cond $X=4.955 $Y=1.5
+ $X2=5.12 $Y2=1.332
r107 5 6 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.955 $Y=1.5 $X2=4.615
+ $Y2=1.5
r108 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.54 $Y=1.575
+ $X2=4.615 $Y2=1.5
r109 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.54 $Y=1.575
+ $X2=4.54 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_193_47# 1 2 9 11 15 17 19 22 26 27 30 31
+ 32 33 42 43 45 49 58 62
c216 43 0 2.06462e-20 $X=10.605 $Y=1.53
c217 33 0 1.37287e-19 $X=7.33 $Y=1.53
c218 32 0 3.76247e-20 $X=10.46 $Y=1.53
c219 22 0 1.92554e-19 $X=10.6 $Y=2.275
c220 11 0 1.43548e-19 $X=7.655 $Y=1.29
r221 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.685
+ $Y=1.74 $X2=10.685 $Y2=1.74
r222 55 58 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=10.6 $Y=1.74
+ $X2=10.685 $Y2=1.74
r223 48 50 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.18 $Y=1.35
+ $X2=7.18 $Y2=1.485
r224 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.18
+ $Y=1.35 $X2=7.18 $Y2=1.35
r225 45 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=7.18 $Y=1.29 $X2=7.18
+ $Y2=1.35
r226 43 59 7.56291 $w=3.18e-07 $l=2.1e-07 $layer=LI1_cond $X=10.61 $Y=1.53
+ $X2=10.61 $Y2=1.74
r227 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.605 $Y=1.53
+ $X2=10.605 $Y2=1.53
r228 40 49 10.7912 $w=1.83e-07 $l=1.8e-07 $layer=LI1_cond $X=7.187 $Y=1.53
+ $X2=7.187 $Y2=1.35
r229 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.185 $Y=1.53
+ $X2=7.185 $Y2=1.53
r230 36 66 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.1 $Y=1.53 $X2=1.1
+ $Y2=1.96
r231 36 62 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.1 $Y=1.53
+ $X2=1.1 $Y2=0.51
r232 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=1.53 $X2=1.1
+ $Y2=1.53
r233 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.33 $Y=1.53
+ $X2=7.185 $Y2=1.53
r234 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.46 $Y=1.53
+ $X2=10.605 $Y2=1.53
r235 32 33 3.87375 $w=1.4e-07 $l=3.13e-06 $layer=MET1_cond $X=10.46 $Y=1.53
+ $X2=7.33 $Y2=1.53
r236 31 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=1.53
+ $X2=1.1 $Y2=1.53
r237 30 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.04 $Y=1.53
+ $X2=7.185 $Y2=1.53
r238 30 31 7.17202 $w=1.4e-07 $l=5.795e-06 $layer=MET1_cond $X=7.04 $Y=1.53
+ $X2=1.245 $Y2=1.53
r239 29 43 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=10.61 $Y=1.035
+ $X2=10.61 $Y2=1.53
r240 27 51 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=10.39 $Y=0.87
+ $X2=10.28 $Y2=0.87
r241 26 29 5.41706 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=10.537 $Y=0.87
+ $X2=10.537 $Y2=1.035
r242 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.39
+ $Y=0.87 $X2=10.39 $Y2=0.87
r243 20 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.6 $Y=1.875
+ $X2=10.6 $Y2=1.74
r244 20 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.6 $Y=1.875
+ $X2=10.6 $Y2=2.275
r245 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.28 $Y=0.705
+ $X2=10.28 $Y2=0.87
r246 17 19 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.28 $Y=0.705
+ $X2=10.28 $Y2=0.415
r247 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=7.73 $Y=1.215
+ $X2=7.73 $Y2=0.415
r248 12 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=1.29
+ $X2=7.18 $Y2=1.29
r249 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.655 $Y=1.29
+ $X2=7.73 $Y2=1.215
r250 11 12 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.655 $Y=1.29
+ $X2=7.345 $Y2=1.29
r251 9 50 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.155 $Y=2.275
+ $X2=7.155 $Y2=1.485
r252 2 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r253 1 62 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_1610_159# 1 2 9 13 17 21 25 27 28 32 36
+ 40 41 47 55
c118 40 0 6.28645e-20 $X=9.66 $Y=1.21
r119 49 50 5.12431 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=9.032 $Y=1.21
+ $X2=9.032 $Y2=1.375
r120 45 55 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=8.255 $Y=0.93
+ $X2=8.26 $Y2=0.93
r121 45 52 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=8.255 $Y=0.93
+ $X2=8.125 $Y2=0.93
r122 44 47 4.13427 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.255 $Y=0.93
+ $X2=8.37 $Y2=0.93
r123 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.255
+ $Y=0.93 $X2=8.255 $Y2=0.93
r124 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.66
+ $Y=1.21 $X2=9.66 $Y2=1.21
r125 38 49 1.93884 $w=3.3e-07 $l=2.03e-07 $layer=LI1_cond $X=9.235 $Y=1.21
+ $X2=9.032 $Y2=1.21
r126 38 40 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=9.235 $Y=1.21
+ $X2=9.66 $Y2=1.21
r127 36 50 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=8.995 $Y=1.88
+ $X2=8.995 $Y2=1.375
r128 30 32 10.6708 $w=4.03e-07 $l=3.75e-07 $layer=LI1_cond $X=9.032 $Y=0.765
+ $X2=9.032 $Y2=0.39
r129 28 49 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=9.032 $Y=0.915
+ $X2=9.032 $Y2=1.21
r130 28 30 4.26831 $w=4.03e-07 $l=1.5e-07 $layer=LI1_cond $X=9.032 $Y=0.915
+ $X2=9.032 $Y2=0.765
r131 28 47 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=8.83 $Y=0.915
+ $X2=8.37 $Y2=0.915
r132 26 41 6.10776 $w=2.75e-07 $l=2.8e-08 $layer=POLY_cond $X=9.662 $Y=1.238
+ $X2=9.662 $Y2=1.21
r133 26 27 42.1909 $w=2.75e-07 $l=1.37e-07 $layer=POLY_cond $X=9.662 $Y=1.238
+ $X2=9.662 $Y2=1.375
r134 25 41 35.9921 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.662 $Y=1.045
+ $X2=9.662 $Y2=1.21
r135 24 25 45.0266 $w=2.75e-07 $l=1.5e-07 $layer=POLY_cond $X=9.697 $Y=0.895
+ $X2=9.697 $Y2=1.045
r136 21 24 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=9.795 $Y=0.445
+ $X2=9.795 $Y2=0.895
r137 17 27 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=9.725 $Y=2.275
+ $X2=9.725 $Y2=1.375
r138 11 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.26 $Y=0.795
+ $X2=8.26 $Y2=0.93
r139 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=8.26 $Y=0.795
+ $X2=8.26 $Y2=0.445
r140 7 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.125 $Y=1.065
+ $X2=8.125 $Y2=0.93
r141 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=8.125 $Y=1.065
+ $X2=8.125 $Y2=2.275
r142 2 36 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.86
+ $Y=1.735 $X2=8.995 $Y2=1.88
r143 1 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.93
+ $Y=0.235 $X2=9.065 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_1446_413# 1 2 8 11 15 16 17 18 19 20 24
+ 29 31 33
c106 29 0 1.40584e-19 $X=7.895 $Y=1.315
c107 17 0 6.28645e-20 $X=8.82 $Y=1.1
r108 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.575
+ $Y=1.41 $X2=8.575 $Y2=1.41
r109 33 35 20.25 $w=2.44e-07 $l=4.05e-07 $layer=LI1_cond $X=8.17 $Y=1.41
+ $X2=8.575 $Y2=1.41
r110 30 33 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.17 $Y=1.575
+ $X2=8.17 $Y2=1.41
r111 30 31 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.17 $Y=1.575
+ $X2=8.17 $Y2=2.175
r112 29 33 13.75 $w=2.44e-07 $l=2.75e-07 $layer=LI1_cond $X=7.895 $Y=1.41
+ $X2=8.17 $Y2=1.41
r113 28 29 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.895 $Y=0.565
+ $X2=7.895 $Y2=1.315
r114 24 28 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=7.81 $Y=0.41
+ $X2=7.895 $Y2=0.565
r115 24 26 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=7.81 $Y=0.41
+ $X2=7.5 $Y2=0.41
r116 20 31 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=8.085 $Y=2.275
+ $X2=8.17 $Y2=2.175
r117 20 22 39.0955 $w=1.98e-07 $l=7.05e-07 $layer=LI1_cond $X=8.085 $Y=2.275
+ $X2=7.38 $Y2=2.275
r118 18 36 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=8.71 $Y=1.41
+ $X2=8.575 $Y2=1.41
r119 18 19 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=8.71 $Y=1.41
+ $X2=8.785 $Y2=1.41
r120 16 17 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=8.82 $Y=0.95
+ $X2=8.82 $Y2=1.1
r121 15 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.855 $Y=0.555
+ $X2=8.855 $Y2=0.95
r122 9 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.785 $Y=1.545
+ $X2=8.785 $Y2=1.41
r123 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=8.785 $Y=1.545
+ $X2=8.785 $Y2=2.11
r124 8 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.785 $Y=1.275
+ $X2=8.785 $Y2=1.41
r125 8 17 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=8.785 $Y=1.275
+ $X2=8.785 $Y2=1.1
r126 2 22 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=2.065 $X2=7.38 $Y2=2.275
r127 1 26 182 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.5 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_2051_413# 1 2 9 13 15 17 19 22 24 26 29
+ 31 33 36 38 40 43 45 46 50 52 56 61 63 66 69
c152 69 0 1.78258e-19 $X=11.025 $Y=1.16
r153 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.725
+ $Y=1.16 $X2=11.725 $Y2=1.16
r154 64 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.11 $Y=1.16
+ $X2=11.025 $Y2=1.16
r155 64 66 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=11.11 $Y=1.16
+ $X2=11.725 $Y2=1.16
r156 62 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.025 $Y=1.325
+ $X2=11.025 $Y2=1.16
r157 62 63 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=11.025 $Y=1.325
+ $X2=11.025 $Y2=2.165
r158 61 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.025 $Y=0.995
+ $X2=11.025 $Y2=1.16
r159 60 61 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=11.025 $Y=0.535
+ $X2=11.025 $Y2=0.995
r160 56 60 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=10.94 $Y=0.432
+ $X2=11.025 $Y2=0.535
r161 56 58 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=10.94 $Y=0.432
+ $X2=10.505 $Y2=0.432
r162 52 63 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=10.94 $Y=2.26
+ $X2=11.025 $Y2=2.165
r163 52 54 32.1053 $w=1.88e-07 $l=5.5e-07 $layer=LI1_cond $X=10.94 $Y=2.26
+ $X2=10.39 $Y2=2.26
r164 49 50 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=13.55 $Y=1.16
+ $X2=13.97 $Y2=1.16
r165 48 49 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=13.13 $Y=1.16
+ $X2=13.55 $Y2=1.16
r166 47 48 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.71 $Y=1.16
+ $X2=13.13 $Y2=1.16
r167 45 67 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=12.15 $Y=1.16
+ $X2=11.725 $Y2=1.16
r168 45 46 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.15 $Y=1.16
+ $X2=12.225 $Y2=1.16
r169 41 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.97 $Y=1.325
+ $X2=13.97 $Y2=1.16
r170 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.97 $Y=1.325
+ $X2=13.97 $Y2=1.985
r171 38 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.97 $Y=0.995
+ $X2=13.97 $Y2=1.16
r172 38 40 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.97 $Y=0.995
+ $X2=13.97 $Y2=0.56
r173 34 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.55 $Y=1.325
+ $X2=13.55 $Y2=1.16
r174 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.55 $Y=1.325
+ $X2=13.55 $Y2=1.985
r175 31 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.55 $Y=0.995
+ $X2=13.55 $Y2=1.16
r176 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.55 $Y=0.995
+ $X2=13.55 $Y2=0.56
r177 27 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.13 $Y=1.325
+ $X2=13.13 $Y2=1.16
r178 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.13 $Y=1.325
+ $X2=13.13 $Y2=1.985
r179 24 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.13 $Y=0.995
+ $X2=13.13 $Y2=1.16
r180 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.13 $Y=0.995
+ $X2=13.13 $Y2=0.56
r181 20 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.71 $Y=1.325
+ $X2=12.71 $Y2=1.16
r182 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.71 $Y=1.325
+ $X2=12.71 $Y2=1.985
r183 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.71 $Y=0.995
+ $X2=12.71 $Y2=1.16
r184 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.71 $Y=0.995
+ $X2=12.71 $Y2=0.56
r185 16 46 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.3 $Y=1.16
+ $X2=12.225 $Y2=1.16
r186 15 47 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.635 $Y=1.16
+ $X2=12.71 $Y2=1.16
r187 15 16 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=12.635 $Y=1.16
+ $X2=12.3 $Y2=1.16
r188 11 46 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.225 $Y=1.325
+ $X2=12.225 $Y2=1.16
r189 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=12.225 $Y=1.325
+ $X2=12.225 $Y2=2.165
r190 7 46 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.225 $Y=0.995
+ $X2=12.225 $Y2=1.16
r191 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=12.225 $Y=0.995
+ $X2=12.225 $Y2=0.445
r192 2 54 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=10.255
+ $Y=2.065 $X2=10.39 $Y2=2.26
r193 1 58 182 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_NDIFF $count=1 $X=10.355
+ $Y=0.235 $X2=10.505 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49
+ 51 55 59 63 69 75 80 81 83 84 86 87 89 90 92 93 94 96 108 112 117 142 143 146
+ 149 152 155 158
c210 143 0 1.8506e-19 $X=14.49 $Y=2.72
c211 41 0 1.67735e-19 $X=3.35 $Y=1.99
c212 1 0 5.65522e-20 $X=0.545 $Y=1.815
r213 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r214 156 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r215 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r216 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r217 149 150 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r218 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r219 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r220 140 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=14.49 $Y2=2.72
r221 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r222 137 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=14.03 $Y2=2.72
r223 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r224 134 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=13.11 $Y2=2.72
r225 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r226 131 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r227 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r228 128 131 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=11.27 $Y2=2.72
r229 128 159 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r230 127 130 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=9.89 $Y=2.72
+ $X2=11.27 $Y2=2.72
r231 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r232 125 158 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.66 $Y=2.72
+ $X2=9.515 $Y2=2.72
r233 125 127 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.66 $Y=2.72
+ $X2=9.89 $Y2=2.72
r234 124 156 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r235 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r236 121 124 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=8.05 $Y2=2.72
r237 121 153 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r238 120 123 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=8.05 $Y2=2.72
r239 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r240 118 152 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=6.01 $Y=2.72
+ $X2=5.837 $Y2=2.72
r241 118 120 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.01 $Y=2.72
+ $X2=6.21 $Y2=2.72
r242 117 155 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=8.425 $Y=2.72
+ $X2=8.542 $Y2=2.72
r243 117 123 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.425 $Y=2.72
+ $X2=8.05 $Y2=2.72
r244 116 153 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r245 116 150 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=3.45 $Y2=2.72
r246 115 116 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r247 113 149 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.46 $Y=2.72
+ $X2=3.362 $Y2=2.72
r248 113 115 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=3.46 $Y=2.72
+ $X2=5.29 $Y2=2.72
r249 112 152 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=5.665 $Y=2.72
+ $X2=5.837 $Y2=2.72
r250 112 115 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.665 $Y=2.72
+ $X2=5.29 $Y2=2.72
r251 111 150 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r252 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r253 108 149 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.362 $Y2=2.72
r254 108 110 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=2.99 $Y2=2.72
r255 107 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r256 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r257 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r258 104 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r259 103 106 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r260 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r261 101 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r262 101 103 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r263 96 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r264 96 98 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r265 94 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r266 94 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r267 92 139 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.095 $Y=2.72
+ $X2=14.03 $Y2=2.72
r268 92 93 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=14.095 $Y=2.72
+ $X2=14.225 $Y2=2.72
r269 91 142 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=14.355 $Y=2.72
+ $X2=14.49 $Y2=2.72
r270 91 93 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=14.355 $Y=2.72
+ $X2=14.225 $Y2=2.72
r271 89 136 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=13.255 $Y=2.72
+ $X2=13.11 $Y2=2.72
r272 89 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.255 $Y=2.72
+ $X2=13.34 $Y2=2.72
r273 88 139 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=13.425 $Y=2.72
+ $X2=14.03 $Y2=2.72
r274 88 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.425 $Y=2.72
+ $X2=13.34 $Y2=2.72
r275 86 133 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.35 $Y=2.72
+ $X2=12.19 $Y2=2.72
r276 86 87 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=12.35 $Y=2.72
+ $X2=12.467 $Y2=2.72
r277 85 136 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=12.585 $Y=2.72
+ $X2=13.11 $Y2=2.72
r278 85 87 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=12.585 $Y=2.72
+ $X2=12.467 $Y2=2.72
r279 83 130 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=11.28 $Y=2.72
+ $X2=11.27 $Y2=2.72
r280 83 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.28 $Y=2.72
+ $X2=11.41 $Y2=2.72
r281 82 133 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.54 $Y=2.72
+ $X2=12.19 $Y2=2.72
r282 82 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.54 $Y=2.72
+ $X2=11.41 $Y2=2.72
r283 80 106 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r284 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.4 $Y2=2.72
r285 79 110 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.99 $Y2=2.72
r286 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.4 $Y2=2.72
r287 75 78 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=14.225 $Y=1.63
+ $X2=14.225 $Y2=2.31
r288 73 93 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=14.225 $Y=2.635
+ $X2=14.225 $Y2=2.72
r289 73 78 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=14.225 $Y=2.635
+ $X2=14.225 $Y2=2.31
r290 69 72 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=13.34 $Y=1.63
+ $X2=13.34 $Y2=2.31
r291 67 90 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.34 $Y=2.635
+ $X2=13.34 $Y2=2.72
r292 67 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.34 $Y=2.635
+ $X2=13.34 $Y2=2.31
r293 63 66 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=12.467 $Y=1.63
+ $X2=12.467 $Y2=1.97
r294 61 87 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=12.467 $Y=2.635
+ $X2=12.467 $Y2=2.72
r295 61 66 32.6117 $w=2.33e-07 $l=6.65e-07 $layer=LI1_cond $X=12.467 $Y=2.635
+ $X2=12.467 $Y2=1.97
r296 57 84 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.41 $Y=2.635
+ $X2=11.41 $Y2=2.72
r297 57 59 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=11.41 $Y=2.635
+ $X2=11.41 $Y2=2.3
r298 53 158 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=2.635
+ $X2=9.515 $Y2=2.72
r299 53 55 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=9.515 $Y=2.635
+ $X2=9.515 $Y2=2.275
r300 52 155 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=8.66 $Y=2.72
+ $X2=8.542 $Y2=2.72
r301 51 158 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.37 $Y=2.72
+ $X2=9.515 $Y2=2.72
r302 51 52 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=9.37 $Y=2.72
+ $X2=8.66 $Y2=2.72
r303 47 155 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.542 $Y=2.635
+ $X2=8.542 $Y2=2.72
r304 47 49 31.1405 $w=2.33e-07 $l=6.35e-07 $layer=LI1_cond $X=8.542 $Y=2.635
+ $X2=8.542 $Y2=2
r305 43 152 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.837 $Y=2.635
+ $X2=5.837 $Y2=2.72
r306 43 45 9.85422 $w=3.43e-07 $l=2.95e-07 $layer=LI1_cond $X=5.837 $Y=2.635
+ $X2=5.837 $Y2=2.34
r307 39 149 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.362 $Y=2.635
+ $X2=3.362 $Y2=2.72
r308 39 41 36.6853 $w=1.93e-07 $l=6.45e-07 $layer=LI1_cond $X=3.362 $Y=2.635
+ $X2=3.362 $Y2=1.99
r309 35 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.635 $X2=2.4
+ $Y2=2.72
r310 35 37 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.4 $Y=2.635
+ $X2=2.4 $Y2=2
r311 31 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r312 31 33 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r313 10 78 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=14.045
+ $Y=1.485 $X2=14.19 $Y2=2.31
r314 10 75 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=14.045
+ $Y=1.485 $X2=14.19 $Y2=1.63
r315 9 72 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=13.205
+ $Y=1.485 $X2=13.34 $Y2=2.31
r316 9 69 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.205
+ $Y=1.485 $X2=13.34 $Y2=1.63
r317 8 66 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=12.3
+ $Y=1.845 $X2=12.5 $Y2=1.97
r318 8 63 600 $w=1.7e-07 $l=2.98706e-07 $layer=licon1_PDIFF $count=1 $X=12.3
+ $Y=1.845 $X2=12.5 $Y2=1.63
r319 7 59 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=11.245
+ $Y=2.065 $X2=11.385 $Y2=2.3
r320 6 55 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=9.39
+ $Y=2.065 $X2=9.515 $Y2=2.275
r321 5 49 300 $w=1.7e-07 $l=3.76098e-07 $layer=licon1_PDIFF $count=2 $X=8.2
+ $Y=2.065 $X2=8.545 $Y2=2
r322 4 45 600 $w=1.7e-07 $l=5.84423e-07 $layer=licon1_PDIFF $count=1 $X=5.61
+ $Y=1.845 $X2=5.805 $Y2=2.34
r323 3 41 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.205
+ $Y=1.845 $X2=3.35 $Y2=1.99
r324 2 37 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.845 $X2=2.4 $Y2=2
r325 1 33 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_299_47# 1 2 3 4 20 21 24 25 29 36 38 40
+ 43 48
c117 38 0 1.82232e-19 $X=4.27 $Y=0.51
r118 38 40 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.27 $Y=0.51
+ $X2=4.125 $Y2=0.51
r119 38 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.27 $Y=0.51
+ $X2=4.27 $Y2=0.51
r120 36 40 2.17465 $w=1.85e-07 $l=2.54e-06 $layer=MET1_cond $X=1.585 $Y=0.487
+ $X2=4.125 $Y2=0.487
r121 34 48 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.44 $Y=0.385
+ $X2=1.62 $Y2=0.385
r122 33 36 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.44 $Y=0.51
+ $X2=1.585 $Y2=0.51
r123 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.44 $Y=0.51
+ $X2=1.44 $Y2=0.51
r124 28 43 22.8354 $w=2.68e-07 $l=5.35e-07 $layer=LI1_cond $X=4.28 $Y=0.98
+ $X2=4.28 $Y2=0.445
r125 28 29 8.82932 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.33 $Y=0.98
+ $X2=4.33 $Y2=1.15
r126 25 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.43 $Y=1.82
+ $X2=4.43 $Y2=1.15
r127 24 25 9.05087 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=4.32 $Y=2 $X2=4.32
+ $Y2=1.82
r128 20 21 7.04283 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=1.57 $Y=1.99 $X2=1.57
+ $Y2=1.89
r129 13 34 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.44 $Y=0.515
+ $X2=1.44 $Y2=0.385
r130 13 21 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=1.44 $Y=0.515
+ $X2=1.44 $Y2=1.89
r131 4 24 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=4.155
+ $Y=1.845 $X2=4.29 $Y2=2
r132 3 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r133 2 43 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.235 $X2=4.29 $Y2=0.445
r134 1 48 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%A_915_47# 1 2 3 4 15 18 20 23 29 31 34 35
+ 37 40 47 49 51 54 60
c131 49 0 2.68486e-19 $X=6.615 $Y=0.51
c132 29 0 5.58337e-20 $X=4.725 $Y=0.825
r133 49 51 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.615 $Y=0.51
+ $X2=6.47 $Y2=0.51
r134 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.615 $Y=0.51
+ $X2=6.615 $Y2=0.51
r135 47 51 1.39126 $w=1.85e-07 $l=1.625e-06 $layer=MET1_cond $X=4.845 $Y=0.487
+ $X2=6.47 $Y2=0.487
r136 44 47 0.0991101 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.7 $Y=0.51
+ $X2=4.845 $Y2=0.51
r137 44 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.7 $Y=0.51 $X2=4.7
+ $Y2=0.51
r138 37 38 7.33994 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.84 $Y=2.34
+ $X2=6.84 $Y2=2.15
r139 35 40 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.84 $Y=1.185
+ $X2=6.84 $Y2=1.865
r140 31 32 4.83766 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.8 $Y=2.34 $X2=4.8
+ $Y2=2.21
r141 29 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.77 $Y=0.825
+ $X2=4.77 $Y2=1.785
r142 28 54 11.0909 $w=1.98e-07 $l=2e-07 $layer=LI1_cond $X=4.695 $Y=0.645
+ $X2=4.695 $Y2=0.445
r143 28 29 10.2632 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=4.725 $Y=0.645
+ $X2=4.725 $Y2=0.825
r144 26 38 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=6.88 $Y=2 $X2=6.88
+ $Y2=2.15
r145 23 40 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.88 $Y=1.99
+ $X2=6.88 $Y2=1.865
r146 23 26 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=6.88 $Y=1.99
+ $X2=6.88 $Y2=2
r147 20 35 9.81506 $w=4.08e-07 $l=2.05e-07 $layer=LI1_cond $X=6.72 $Y=0.98
+ $X2=6.72 $Y2=1.185
r148 19 60 9.29389 $w=3.08e-07 $l=2.5e-07 $layer=LI1_cond $X=6.72 $Y=0.41
+ $X2=6.97 $Y2=0.41
r149 19 50 3.90344 $w=3.08e-07 $l=1.05e-07 $layer=LI1_cond $X=6.72 $Y=0.41
+ $X2=6.615 $Y2=0.41
r150 19 20 11.665 $w=4.08e-07 $l=4.15e-07 $layer=LI1_cond $X=6.72 $Y=0.565
+ $X2=6.72 $Y2=0.98
r151 18 32 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.825 $Y=2
+ $X2=4.825 $Y2=2.21
r152 15 34 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=4.825 $Y=1.925
+ $X2=4.825 $Y2=1.785
r153 15 18 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=4.825 $Y=1.925
+ $X2=4.825 $Y2=2
r154 4 37 600 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_PDIFF $count=1 $X=6.635
+ $Y=1.845 $X2=6.84 $Y2=2.34
r155 4 26 600 $w=1.7e-07 $l=2.71662e-07 $layer=licon1_PDIFF $count=1 $X=6.635
+ $Y=1.845 $X2=6.84 $Y2=2
r156 3 31 600 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.845 $X2=4.8 $Y2=2.34
r157 3 18 600 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.845 $X2=4.8 $Y2=2
r158 2 60 91 $w=1.7e-07 $l=5.64978e-07 $layer=licon1_NDIFF $count=2 $X=6.49
+ $Y=0.595 $X2=6.97 $Y2=0.41
r159 1 54 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.575
+ $Y=0.235 $X2=4.71 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%Q 1 2 3 4 15 19 23 27 31 35 36
r48 31 33 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.76 $Y=1.63
+ $X2=13.76 $Y2=2.31
r49 29 35 3.71613 $w=3.3e-07 $l=1.13e-07 $layer=LI1_cond $X=13.76 $Y=1.295
+ $X2=13.76 $Y2=1.182
r50 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.76 $Y=1.295
+ $X2=13.76 $Y2=1.63
r51 25 35 3.71613 $w=3.3e-07 $l=1.12e-07 $layer=LI1_cond $X=13.76 $Y=1.07
+ $X2=13.76 $Y2=1.182
r52 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=13.76 $Y=1.07
+ $X2=13.76 $Y2=0.395
r53 24 36 2.75166 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=13.085 $Y=1.182
+ $X2=12.92 $Y2=1.182
r54 23 35 2.75166 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=13.595 $Y=1.182
+ $X2=13.76 $Y2=1.182
r55 23 24 26.122 $w=2.23e-07 $l=5.1e-07 $layer=LI1_cond $X=13.595 $Y=1.182
+ $X2=13.085 $Y2=1.182
r56 19 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=12.92 $Y=1.63
+ $X2=12.92 $Y2=2.31
r57 17 36 3.71613 $w=3.3e-07 $l=1.13e-07 $layer=LI1_cond $X=12.92 $Y=1.295
+ $X2=12.92 $Y2=1.182
r58 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.92 $Y=1.295
+ $X2=12.92 $Y2=1.63
r59 13 36 3.71613 $w=3.3e-07 $l=1.12e-07 $layer=LI1_cond $X=12.92 $Y=1.07
+ $X2=12.92 $Y2=1.182
r60 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.92 $Y=1.07
+ $X2=12.92 $Y2=0.395
r61 4 33 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=13.625
+ $Y=1.485 $X2=13.76 $Y2=2.31
r62 4 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.625
+ $Y=1.485 $X2=13.76 $Y2=1.63
r63 3 21 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=12.785
+ $Y=1.485 $X2=12.92 $Y2=2.31
r64 3 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.785
+ $Y=1.485 $X2=12.92 $Y2=1.63
r65 2 27 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=13.625
+ $Y=0.235 $X2=13.76 $Y2=0.395
r66 1 15 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=12.785
+ $Y=0.235 $X2=12.92 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__SEDFXTP_4%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49
+ 53 57 61 67 71 74 75 77 78 80 81 83 84 86 87 89 90 92 93 94 96 108 116 143 144
+ 147 150 153
c236 144 0 1.44919e-19 $X=14.49 $Y=0
c237 116 0 1.67078e-19 $X=8.245 $Y=0
c238 77 0 1.82232e-19 $X=5.76 $Y=0
r239 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r240 150 151 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r241 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r242 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r243 141 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=14.49 $Y2=0
r244 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r245 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=14.03 $Y2=0
r246 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r247 135 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=13.11 $Y2=0
r248 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r249 132 135 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=12.19 $Y2=0
r250 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r251 129 132 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=11.27 $Y2=0
r252 128 131 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=11.27 $Y2=0
r253 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r254 126 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r255 126 154 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.51 $Y2=0
r256 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r257 123 153 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=8.64 $Y=0
+ $X2=8.442 $Y2=0
r258 123 125 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.64 $Y=0
+ $X2=9.43 $Y2=0
r259 122 154 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r260 121 122 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r261 119 122 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=8.05 $Y2=0
r262 118 121 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=8.05 $Y2=0
r263 118 119 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r264 116 153 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=8.245 $Y=0
+ $X2=8.442 $Y2=0
r265 116 121 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.245 $Y=0
+ $X2=8.05 $Y2=0
r266 115 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r267 115 151 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=3.45 $Y2=0
r268 114 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r269 112 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=3.35 $Y2=0
r270 112 114 145.813 $w=1.68e-07 $l=2.235e-06 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=5.75 $Y2=0
r271 111 151 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.45 $Y2=0
r272 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r273 108 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.35 $Y2=0
r274 108 110 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=2.99 $Y2=0
r275 107 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r276 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r277 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r278 104 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r279 103 106 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r280 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r281 101 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r282 101 103 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r283 96 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r284 96 98 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r285 94 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r286 94 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r287 92 140 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.095 $Y=0
+ $X2=14.03 $Y2=0
r288 92 93 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=14.095 $Y=0
+ $X2=14.225 $Y2=0
r289 91 143 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=14.355 $Y=0
+ $X2=14.49 $Y2=0
r290 91 93 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=14.355 $Y=0
+ $X2=14.225 $Y2=0
r291 89 137 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=13.255 $Y=0
+ $X2=13.11 $Y2=0
r292 89 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.255 $Y=0
+ $X2=13.34 $Y2=0
r293 88 140 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=13.425 $Y=0
+ $X2=14.03 $Y2=0
r294 88 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.425 $Y=0
+ $X2=13.34 $Y2=0
r295 86 134 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.35 $Y=0
+ $X2=12.19 $Y2=0
r296 86 87 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=12.35 $Y=0
+ $X2=12.467 $Y2=0
r297 85 137 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=12.585 $Y=0
+ $X2=13.11 $Y2=0
r298 85 87 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=12.585 $Y=0
+ $X2=12.467 $Y2=0
r299 83 131 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=11.35 $Y=0 $X2=11.27
+ $Y2=0
r300 83 84 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=11.35 $Y=0
+ $X2=11.507 $Y2=0
r301 82 134 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=11.665 $Y=0
+ $X2=12.19 $Y2=0
r302 82 84 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=11.665 $Y=0
+ $X2=11.507 $Y2=0
r303 80 125 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=9.465 $Y=0
+ $X2=9.43 $Y2=0
r304 80 81 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=9.465 $Y=0
+ $X2=9.602 $Y2=0
r305 79 128 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.74 $Y=0 $X2=9.89
+ $Y2=0
r306 79 81 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=9.74 $Y=0 $X2=9.602
+ $Y2=0
r307 77 114 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.76 $Y=0 $X2=5.75
+ $Y2=0
r308 77 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.76 $Y=0 $X2=5.885
+ $Y2=0
r309 76 118 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.01 $Y=0 $X2=6.21
+ $Y2=0
r310 76 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.01 $Y=0 $X2=5.885
+ $Y2=0
r311 74 106 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0
+ $X2=2.07 $Y2=0
r312 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.4
+ $Y2=0
r313 73 110 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=0
+ $X2=2.99 $Y2=0
r314 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.4
+ $Y2=0
r315 69 93 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=14.225 $Y=0.085
+ $X2=14.225 $Y2=0
r316 69 71 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=14.225 $Y=0.085
+ $X2=14.225 $Y2=0.395
r317 65 90 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.34 $Y=0.085
+ $X2=13.34 $Y2=0
r318 65 67 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=13.34 $Y=0.085
+ $X2=13.34 $Y2=0.395
r319 61 63 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=12.467 $Y=0.395
+ $X2=12.467 $Y2=0.735
r320 59 87 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=12.467 $Y=0.085
+ $X2=12.467 $Y2=0
r321 59 61 15.2024 $w=2.33e-07 $l=3.1e-07 $layer=LI1_cond $X=12.467 $Y=0.085
+ $X2=12.467 $Y2=0.395
r322 55 84 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=11.507 $Y=0.085
+ $X2=11.507 $Y2=0
r323 55 57 13.3537 $w=3.13e-07 $l=3.65e-07 $layer=LI1_cond $X=11.507 $Y=0.085
+ $X2=11.507 $Y2=0.45
r324 51 81 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.602 $Y=0.085
+ $X2=9.602 $Y2=0
r325 51 53 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=9.602 $Y=0.085
+ $X2=9.602 $Y2=0.45
r326 47 153 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=8.442 $Y=0.085
+ $X2=8.442 $Y2=0
r327 47 49 9.77388 $w=3.93e-07 $l=3.35e-07 $layer=LI1_cond $X=8.442 $Y=0.085
+ $X2=8.442 $Y2=0.42
r328 43 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=0.085
+ $X2=5.885 $Y2=0
r329 43 45 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=5.885 $Y=0.085
+ $X2=5.885 $Y2=0.74
r330 39 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r331 39 41 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.445
r332 35 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=0.085 $X2=2.4
+ $Y2=0
r333 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.4 $Y=0.085
+ $X2=2.4 $Y2=0.38
r334 31 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r335 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r336 10 71 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=14.045
+ $Y=0.235 $X2=14.19 $Y2=0.395
r337 9 67 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=13.205
+ $Y=0.235 $X2=13.34 $Y2=0.395
r338 8 63 182 $w=1.7e-07 $l=5.91608e-07 $layer=licon1_NDIFF $count=1 $X=12.3
+ $Y=0.235 $X2=12.5 $Y2=0.735
r339 8 61 182 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_NDIFF $count=1 $X=12.3
+ $Y=0.235 $X2=12.5 $Y2=0.395
r340 7 57 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=11.36
+ $Y=0.235 $X2=11.495 $Y2=0.45
r341 6 53 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=9.46
+ $Y=0.235 $X2=9.585 $Y2=0.45
r342 5 49 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=8.335
+ $Y=0.235 $X2=8.475 $Y2=0.42
r343 4 45 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.71
+ $Y=0.595 $X2=5.845 $Y2=0.74
r344 3 41 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.235 $X2=3.35 $Y2=0.445
r345 2 37 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.4 $Y2=0.38
r346 1 33 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


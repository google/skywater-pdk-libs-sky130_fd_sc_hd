* File: sky130_fd_sc_hd__a211o_1.pxi.spice
* Created: Thu Aug 27 13:59:19 2020
* 
x_PM_SKY130_FD_SC_HD__A211O_1%A_80_21# N_A_80_21#_M1008_d N_A_80_21#_M1007_d
+ N_A_80_21#_M1002_d N_A_80_21#_c_57_n N_A_80_21#_M1004_g N_A_80_21#_M1006_g
+ N_A_80_21#_c_58_n N_A_80_21#_c_59_n N_A_80_21#_c_67_p N_A_80_21#_c_128_p
+ N_A_80_21#_c_64_n N_A_80_21#_c_107_p N_A_80_21#_c_68_p N_A_80_21#_c_60_n
+ N_A_80_21#_c_65_n N_A_80_21#_c_135_p N_A_80_21#_c_84_p
+ PM_SKY130_FD_SC_HD__A211O_1%A_80_21#
x_PM_SKY130_FD_SC_HD__A211O_1%A2 N_A2_c_151_n N_A2_M1003_g N_A2_M1009_g A2
+ N_A2_c_153_n PM_SKY130_FD_SC_HD__A211O_1%A2
x_PM_SKY130_FD_SC_HD__A211O_1%A1 N_A1_M1008_g N_A1_M1005_g A1 N_A1_c_184_n
+ N_A1_c_185_n N_A1_c_186_n PM_SKY130_FD_SC_HD__A211O_1%A1
x_PM_SKY130_FD_SC_HD__A211O_1%B1 N_B1_M1001_g N_B1_M1000_g B1 N_B1_c_220_n
+ N_B1_c_221_n PM_SKY130_FD_SC_HD__A211O_1%B1
x_PM_SKY130_FD_SC_HD__A211O_1%C1 N_C1_c_252_n N_C1_M1007_g N_C1_M1002_g C1
+ N_C1_c_254_n PM_SKY130_FD_SC_HD__A211O_1%C1
x_PM_SKY130_FD_SC_HD__A211O_1%X N_X_M1004_s N_X_M1006_s X X X X X X N_X_c_278_n
+ X PM_SKY130_FD_SC_HD__A211O_1%X
x_PM_SKY130_FD_SC_HD__A211O_1%VPWR N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_c_294_n
+ N_VPWR_c_295_n VPWR N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n
+ N_VPWR_c_293_n N_VPWR_c_300_n N_VPWR_c_301_n VPWR
+ PM_SKY130_FD_SC_HD__A211O_1%VPWR
x_PM_SKY130_FD_SC_HD__A211O_1%A_217_297# N_A_217_297#_M1009_s
+ N_A_217_297#_M1005_d N_A_217_297#_c_342_n N_A_217_297#_c_343_n
+ N_A_217_297#_c_347_n N_A_217_297#_c_348_n N_A_217_297#_c_350_n
+ PM_SKY130_FD_SC_HD__A211O_1%A_217_297#
x_PM_SKY130_FD_SC_HD__A211O_1%VGND N_VGND_M1004_d N_VGND_M1001_d N_VGND_c_372_n
+ VGND N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ N_VGND_c_377_n N_VGND_c_378_n VGND PM_SKY130_FD_SC_HD__A211O_1%VGND
cc_1 VNB N_A_80_21#_c_57_n 0.0230993f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_58_n 0.00417714f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_3 VNB N_A_80_21#_c_59_n 0.0352812f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_4 VNB N_A_80_21#_c_60_n 0.00773822f $X=-0.19 $Y=-0.24 $X2=2.86 $Y2=0.72
cc_5 VNB N_A2_c_151_n 0.0196207f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.235
cc_6 VNB A2 0.00251915f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A2_c_153_n 0.0273788f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_8 VNB N_A1_c_184_n 0.018091f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_9 VNB N_A1_c_185_n 0.00463632f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_10 VNB N_A1_c_186_n 0.0166822f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.325
cc_11 VNB B1 0.00198956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_220_n 0.0200322f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_13 VNB N_B1_c_221_n 0.0167989f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.325
cc_14 VNB N_C1_c_252_n 0.0224365f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.235
cc_15 VNB C1 0.0125508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_C1_c_254_n 0.0324824f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.325
cc_17 VNB N_X_c_278_n 0.0421698f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.72
cc_18 VNB N_VPWR_c_293_n 0.136896f $X=-0.19 $Y=-0.24 $X2=2.95 $Y2=1.85
cc_19 VNB N_VGND_c_372_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_373_n 0.0249845f $X=-0.19 $Y=-0.24 $X2=0.712 $Y2=1.505
cc_21 VNB N_VGND_c_374_n 0.015399f $X=-0.19 $Y=-0.24 $X2=0.825 $Y2=1.595
cc_22 VNB N_VGND_c_375_n 0.182222f $X=-0.19 $Y=-0.24 $X2=2.042 $Y2=0.625
cc_23 VNB N_VGND_c_376_n 0.0182722f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.72
cc_24 VNB N_VGND_c_377_n 0.0206035f $X=-0.19 $Y=-0.24 $X2=2.972 $Y2=0.53
cc_25 VNB N_VGND_c_378_n 0.00436092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A_80_21#_M1006_g 0.0255235f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_27 VPB N_A_80_21#_c_58_n 0.00348844f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_28 VPB N_A_80_21#_c_59_n 0.00961799f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_29 VPB N_A_80_21#_c_64_n 0.0238817f $X=-0.19 $Y=1.305 $X2=2.805 $Y2=1.595
cc_30 VPB N_A_80_21#_c_65_n 0.0285321f $X=-0.19 $Y=1.305 $X2=2.96 $Y2=1.85
cc_31 VPB N_A2_M1009_g 0.023267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB A2 6.43935e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A2_c_153_n 0.00788481f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_34 VPB N_A1_M1005_g 0.0191523f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A1_c_184_n 0.00387688f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_36 VPB N_A1_c_185_n 0.00286372f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_37 VPB N_B1_M1000_g 0.0197252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB B1 0.00198956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_B1_c_220_n 0.0039962f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_40 VPB N_C1_M1002_g 0.0267587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB C1 0.00185686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_C1_c_254_n 0.00818673f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_43 VPB X 0.0294769f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_44 VPB N_X_c_278_n 0.00882641f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.72
cc_45 VPB X 0.0065071f $X=-0.19 $Y=1.305 $X2=2.96 $Y2=0.53
cc_46 VPB N_VPWR_c_294_n 0.00776473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_295_n 4.14e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_48 VPB N_VPWR_c_296_n 0.0153767f $X=-0.19 $Y=1.305 $X2=0.712 $Y2=0.815
cc_49 VPB N_VPWR_c_297_n 0.0154602f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.72
cc_50 VPB N_VPWR_c_298_n 0.0403087f $X=-0.19 $Y=1.305 $X2=2.95 $Y2=1.685
cc_51 VPB N_VPWR_c_293_n 0.0532622f $X=-0.19 $Y=1.305 $X2=2.95 $Y2=1.85
cc_52 VPB N_VPWR_c_300_n 0.00510842f $X=-0.19 $Y=1.305 $X2=2.972 $Y2=0.625
cc_53 VPB N_VPWR_c_301_n 0.00436092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_217_297#_c_342_n 0.00282128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_217_297#_c_343_n 0.00348313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 N_A_80_21#_c_58_n N_A2_c_151_n 0.00437041f $X=0.685 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_57 N_A_80_21#_c_67_p N_A2_c_151_n 0.0190268f $X=1.915 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_58 N_A_80_21#_c_68_p N_A2_c_151_n 0.0013729f $X=2.07 $Y=0.53 $X2=-0.19
+ $Y2=-0.24
cc_59 N_A_80_21#_c_58_n N_A2_M1009_g 0.00437041f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_80_21#_c_64_n N_A2_M1009_g 0.0172214f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_58_n A2 0.0234667f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_59_n A2 0.0011295f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_67_p A2 0.0197483f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_64_n A2 0.0197541f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_58_n N_A2_c_153_n 9.64614e-19 $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_59_n N_A2_c_153_n 0.016491f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_67_p N_A2_c_153_n 0.005898f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_64_n N_A2_c_153_n 0.00589186f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_64_n N_A1_M1005_g 0.0109073f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_67_p N_A1_c_184_n 0.0014309f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_64_n N_A1_c_184_n 0.00143053f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_67_p N_A1_c_185_n 0.0270648f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_64_n N_A1_c_185_n 0.0355909f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_84_p N_A1_c_185_n 0.00917945f $X=2.042 $Y=0.72 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_67_p N_A1_c_186_n 0.00949049f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_68_p N_A1_c_186_n 0.00695673f $X=2.07 $Y=0.53 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_84_p N_A1_c_186_n 0.00151611f $X=2.042 $Y=0.72 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_64_n N_B1_M1000_g 0.0157981f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_65_n N_B1_M1000_g 0.00259861f $X=2.96 $Y=1.85 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_64_n B1 0.0274253f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_60_n B1 0.0275154f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_64_n N_B1_c_220_n 0.00209973f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_60_n N_B1_c_220_n 0.00210097f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_60_n N_B1_c_221_n 0.0123748f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_60_n N_C1_c_252_n 0.0164214f $X=2.86 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_80_21#_c_64_n N_C1_M1002_g 0.0202735f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_65_n N_C1_M1002_g 0.0144531f $X=2.96 $Y=1.85 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_64_n C1 0.0180533f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_60_n C1 0.0167689f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_64_n N_C1_c_254_n 0.00607929f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_60_n N_C1_c_254_n 0.00512329f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_57_n N_X_c_278_n 0.0158608f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_80_21#_M1006_g N_X_c_278_n 0.00527573f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_58_n N_X_c_278_n 0.0469962f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_59_n N_X_c_278_n 0.0120011f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_80_21#_M1006_g X 0.00299028f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_107_p N_VPWR_M1006_d 0.0047055f $X=0.825 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_80_21#_c_64_n N_VPWR_M1009_d 0.00359948f $X=2.805 $Y=1.595 $X2=0 $Y2=0
cc_99 N_A_80_21#_M1006_g N_VPWR_c_294_n 0.013979f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_59_n N_VPWR_c_294_n 8.30886e-19 $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_64_n N_VPWR_c_294_n 0.00195776f $X=2.805 $Y=1.595 $X2=0
+ $Y2=0
cc_102 N_A_80_21#_c_107_p N_VPWR_c_294_n 0.0156852f $X=0.825 $Y=1.595 $X2=0
+ $Y2=0
cc_103 N_A_80_21#_M1006_g N_VPWR_c_296_n 0.00486043f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_A_80_21#_c_65_n N_VPWR_c_298_n 0.0171566f $X=2.96 $Y=1.85 $X2=0 $Y2=0
cc_105 N_A_80_21#_M1002_d N_VPWR_c_293_n 0.00214551f $X=2.82 $Y=1.485 $X2=0
+ $Y2=0
cc_106 N_A_80_21#_M1006_g N_VPWR_c_293_n 0.00915791f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_107 N_A_80_21#_c_65_n N_VPWR_c_293_n 0.0109745f $X=2.96 $Y=1.85 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_64_n N_A_217_297#_M1009_s 0.00489425f $X=2.805 $Y=1.595
+ $X2=-0.19 $Y2=-0.24
cc_109 N_A_80_21#_c_64_n N_A_217_297#_M1005_d 0.00618192f $X=2.805 $Y=1.595
+ $X2=0 $Y2=0
cc_110 N_A_80_21#_c_64_n N_A_217_297#_c_342_n 0.0193105f $X=2.805 $Y=1.595 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_c_64_n N_A_217_297#_c_347_n 0.0317761f $X=2.805 $Y=1.595 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_c_64_n N_A_217_297#_c_348_n 0.0146073f $X=2.805 $Y=1.595 $X2=0
+ $Y2=0
cc_113 N_A_80_21#_c_65_n N_A_217_297#_c_348_n 0.00669316f $X=2.96 $Y=1.85 $X2=0
+ $Y2=0
cc_114 N_A_80_21#_c_65_n N_A_217_297#_c_350_n 0.00968233f $X=2.96 $Y=1.85 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_c_64_n A_472_297# 0.00957289f $X=2.805 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_80_21#_c_58_n N_VGND_M1004_d 0.00112378f $X=0.685 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_117 N_A_80_21#_c_67_p N_VGND_M1004_d 0.0185063f $X=1.915 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_80_21#_c_128_p N_VGND_M1004_d 0.00461432f $X=0.825 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_80_21#_c_60_n N_VGND_M1001_d 0.00405337f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_60_n N_VGND_c_372_n 0.0162239f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_67_p N_VGND_c_373_n 0.00892803f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_68_p N_VGND_c_373_n 0.0141293f $X=2.07 $Y=0.53 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_60_n N_VGND_c_373_n 0.00274625f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_60_n N_VGND_c_374_n 0.00274625f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_135_p N_VGND_c_374_n 0.0140055f $X=2.96 $Y=0.53 $X2=0 $Y2=0
cc_126 N_A_80_21#_M1008_d N_VGND_c_375_n 0.0023835f $X=1.93 $Y=0.235 $X2=0 $Y2=0
cc_127 N_A_80_21#_M1007_d N_VGND_c_375_n 0.00226911f $X=2.82 $Y=0.235 $X2=0
+ $Y2=0
cc_128 N_A_80_21#_c_57_n N_VGND_c_375_n 0.0121086f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_67_p N_VGND_c_375_n 0.0171709f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_128_p N_VGND_c_375_n 0.00126116f $X=0.825 $Y=0.72 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_c_68_p N_VGND_c_375_n 0.00957785f $X=2.07 $Y=0.53 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_60_n N_VGND_c_375_n 0.0104498f $X=2.86 $Y=0.72 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_135_p N_VGND_c_375_n 0.00849891f $X=2.96 $Y=0.53 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_57_n N_VGND_c_376_n 0.00549284f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_135 N_A_80_21#_c_57_n N_VGND_c_377_n 0.00897449f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_136 N_A_80_21#_c_59_n N_VGND_c_377_n 7.65257e-19 $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_67_p N_VGND_c_377_n 0.0356257f $X=1.915 $Y=0.72 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_128_p N_VGND_c_377_n 0.0182131f $X=0.825 $Y=0.72 $X2=0 $Y2=0
cc_139 N_A_80_21#_c_68_p N_VGND_c_377_n 0.00549328f $X=2.07 $Y=0.53 $X2=0 $Y2=0
cc_140 N_A_80_21#_c_67_p A_300_47# 0.00466022f $X=1.915 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A2_M1009_g N_A1_M1005_g 0.0454923f $X=1.425 $Y=1.985 $X2=0 $Y2=0
cc_142 A2 N_A1_c_184_n 2.10318e-19 $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A2_c_153_n N_A1_c_184_n 0.0214364f $X=1.425 $Y=1.16 $X2=0 $Y2=0
cc_144 A2 N_A1_c_185_n 0.0244989f $X=1.075 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A2_c_153_n N_A1_c_185_n 0.00860595f $X=1.425 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A2_c_151_n N_A1_c_186_n 0.0411168f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A2_M1009_g N_VPWR_c_294_n 0.00200931f $X=1.425 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A2_M1009_g N_VPWR_c_295_n 0.00677631f $X=1.425 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A2_M1009_g N_VPWR_c_297_n 0.0035231f $X=1.425 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A2_M1009_g N_VPWR_c_293_n 0.00539272f $X=1.425 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A2_M1009_g N_A_217_297#_c_347_n 0.0111161f $X=1.425 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A2_c_151_n N_VGND_c_373_n 0.00422911f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A2_c_151_n N_VGND_c_375_n 0.00485693f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A2_c_151_n N_VGND_c_377_n 0.0130985f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A1_M1005_g N_B1_M1000_g 0.0273063f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A1_c_184_n B1 3.23374e-19 $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_c_185_n B1 0.0267586f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A1_c_184_n N_B1_c_220_n 0.0202199f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A1_c_185_n N_B1_c_220_n 0.00212673f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A1_c_186_n N_B1_c_221_n 0.0238819f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A1_M1005_g N_VPWR_c_295_n 0.00755649f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A1_M1005_g N_VPWR_c_298_n 0.0035231f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A1_M1005_g N_VPWR_c_293_n 0.00411837f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A1_M1005_g N_A_217_297#_c_347_n 0.0111161f $X=1.855 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A1_c_186_n N_VGND_c_372_n 0.001215f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_186_n N_VGND_c_373_n 0.00418729f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A1_c_186_n N_VGND_c_375_n 0.00589251f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A1_c_186_n N_VGND_c_377_n 0.00170554f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B1_c_221_n N_C1_c_252_n 0.0235362f $X=2.325 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_170 N_B1_M1000_g N_C1_M1002_g 0.0512625f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_171 B1 C1 0.023898f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_172 N_B1_c_220_n C1 2.16206e-19 $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_173 B1 N_C1_c_254_n 0.00807514f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_174 N_B1_c_220_n N_C1_c_254_n 0.0214364f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_175 N_B1_M1000_g N_VPWR_c_295_n 0.00110171f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B1_M1000_g N_VPWR_c_298_n 0.00549284f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B1_M1000_g N_VPWR_c_293_n 0.0100645f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_178 N_B1_M1000_g N_A_217_297#_c_348_n 0.00455091f $X=2.285 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_B1_M1000_g N_A_217_297#_c_350_n 0.00675953f $X=2.285 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_B1_c_221_n N_VGND_c_372_n 0.00686288f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B1_c_221_n N_VGND_c_373_n 0.00394671f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B1_c_221_n N_VGND_c_375_n 0.00458871f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_183 N_C1_M1002_g N_VPWR_c_298_n 0.00564326f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_184 N_C1_M1002_g N_VPWR_c_293_n 0.0114172f $X=2.745 $Y=1.985 $X2=0 $Y2=0
cc_185 N_C1_M1002_g N_A_217_297#_c_348_n 6.92141e-19 $X=2.745 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_C1_M1002_g N_A_217_297#_c_350_n 0.00108796f $X=2.745 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_C1_c_252_n N_VGND_c_372_n 0.00748124f $X=2.745 $Y=0.995 $X2=0 $Y2=0
cc_188 N_C1_c_252_n N_VGND_c_374_n 0.00394671f $X=2.745 $Y=0.995 $X2=0 $Y2=0
cc_189 N_C1_c_252_n N_VGND_c_375_n 0.00553087f $X=2.745 $Y=0.995 $X2=0 $Y2=0
cc_190 X N_VPWR_c_296_n 0.0170803f $X=0.135 $Y=1.785 $X2=0 $Y2=0
cc_191 N_X_M1006_s N_VPWR_c_293_n 0.00369911f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_192 X N_VPWR_c_293_n 0.0100807f $X=0.135 $Y=1.785 $X2=0 $Y2=0
cc_193 N_X_M1004_s N_VGND_c_375_n 0.00213747f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_194 N_X_c_278_n N_VGND_c_375_n 0.0125813f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_195 N_X_c_278_n N_VGND_c_376_n 0.0201263f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_196 N_VPWR_c_293_n N_A_217_297#_M1009_s 0.00228308f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_197 N_VPWR_c_293_n N_A_217_297#_M1005_d 0.00238138f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_294_n N_A_217_297#_c_342_n 0.0147176f $X=0.69 $Y=2 $X2=0 $Y2=0
cc_199 N_VPWR_c_294_n N_A_217_297#_c_343_n 0.0271924f $X=0.69 $Y=2 $X2=0 $Y2=0
cc_200 N_VPWR_c_297_n N_A_217_297#_c_343_n 0.0165739f $X=1.475 $Y=2.72 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_293_n N_A_217_297#_c_343_n 0.00985117f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_202 N_VPWR_M1009_d N_A_217_297#_c_347_n 0.00352445f $X=1.5 $Y=1.485 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_295_n N_A_217_297#_c_347_n 0.0162814f $X=1.64 $Y=2.36 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_297_n N_A_217_297#_c_347_n 0.00256868f $X=1.475 $Y=2.72 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_298_n N_A_217_297#_c_347_n 0.00256868f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_293_n N_A_217_297#_c_347_n 0.0100249f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_298_n N_A_217_297#_c_350_n 0.0146245f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_293_n N_A_217_297#_c_350_n 0.00966897f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_293_n A_472_297# 0.0132511f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_210 N_VGND_c_375_n A_300_47# 0.00322965f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

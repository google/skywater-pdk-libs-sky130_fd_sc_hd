* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=1.879e+12p ps=1.667e+07u
M1001 VPWR a_1429_21# a_1341_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.848e+11p ps=1.72e+06u
M1002 VGND a_648_21# a_582_47# VNB nshort w=420000u l=150000u
+  ad=1.0626e+12p pd=1.148e+07u as=1.341e+11p ps=1.5e+06u
M1003 a_1160_47# a_648_21# VGND VNB nshort w=640000u l=150000u
+  ad=1.87e+11p pd=1.93e+06u as=0p ps=0u
M1004 a_1663_329# a_1255_47# a_1429_21# VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=2.457e+11p ps=2.34e+06u
M1005 a_648_21# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.94e+11p pd=2.46e+06u as=0p ps=0u
M1006 a_381_47# D VGND VNB nshort w=420000u l=150000u
+  ad=1.32e+11p pd=1.49e+06u as=0p ps=0u
M1007 VPWR a_942_21# a_1663_329# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_1429_21# a_2136_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1009 VGND a_1429_21# a_1364_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1010 a_1429_21# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_1429_21# a_2136_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1012 a_558_413# a_27_47# a_474_413# VPB phighvt w=420000u l=150000u
+  ad=1.89e+11p pd=1.74e+06u as=1.134e+11p ps=1.38e+06u
M1013 VPWR CLK a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1014 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1015 VPWR a_942_21# a_892_329# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1016 a_474_413# a_193_47# a_381_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.323e+11p ps=1.47e+06u
M1017 VGND RESET_B a_942_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1018 a_1341_413# a_193_47# a_1255_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1019 a_788_47# a_942_21# a_648_21# VNB nshort w=640000u l=150000u
+  ad=3.684e+11p pd=3.78e+06u as=1.728e+11p ps=1.82e+06u
M1020 a_381_47# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_648_21# a_558_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_892_329# a_474_413# a_648_21# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_648_21# a_474_413# a_788_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1364_47# a_27_47# a_1255_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.422e+11p ps=1.51e+06u
M1025 a_1545_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=4.062e+11p pd=3.96e+06u as=0p ps=0u
M1026 a_582_47# a_193_47# a_474_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.368e+11p ps=1.48e+06u
M1027 a_1255_47# a_193_47# a_1160_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1429_21# a_1255_47# a_1545_47# VNB nshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1029 a_788_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1113_329# a_648_21# VPWR VPB phighvt w=840000u l=150000u
+  ad=3.486e+11p pd=2.82e+06u as=0p ps=0u
M1031 a_1255_47# a_27_47# a_1113_329# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_474_413# a_27_47# a_381_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q a_2136_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1034 VPWR RESET_B a_942_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1035 Q_N a_1429_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1036 a_1545_47# a_942_21# a_1429_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1038 Q a_2136_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1039 Q_N a_1429_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__nand2b_4.pxi.spice
* Created: Tue Sep  1 19:15:56 2020
* 
x_PM_SKY130_FD_SC_HD__NAND2B_4%A_N N_A_N_M1017_g N_A_N_M1014_g A_N N_A_N_c_93_n
+ PM_SKY130_FD_SC_HD__NAND2B_4%A_N
x_PM_SKY130_FD_SC_HD__NAND2B_4%A_27_47# N_A_27_47#_M1017_s N_A_27_47#_M1014_s
+ N_A_27_47#_M1002_g N_A_27_47#_M1000_g N_A_27_47#_M1003_g N_A_27_47#_M1012_g
+ N_A_27_47#_M1007_g N_A_27_47#_M1015_g N_A_27_47#_M1010_g N_A_27_47#_M1016_g
+ N_A_27_47#_c_125_n N_A_27_47#_c_137_n N_A_27_47#_c_126_n N_A_27_47#_c_127_n
+ N_A_27_47#_c_128_n N_A_27_47#_c_129_n N_A_27_47#_c_139_n N_A_27_47#_c_130_n
+ N_A_27_47#_c_131_n N_A_27_47#_c_132_n PM_SKY130_FD_SC_HD__NAND2B_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND2B_4%B N_B_M1004_g N_B_M1001_g N_B_M1008_g N_B_M1005_g
+ N_B_M1011_g N_B_M1006_g N_B_M1013_g N_B_M1009_g B B B B N_B_c_247_n
+ N_B_c_248_n PM_SKY130_FD_SC_HD__NAND2B_4%B
x_PM_SKY130_FD_SC_HD__NAND2B_4%VPWR N_VPWR_M1014_d N_VPWR_M1000_s N_VPWR_M1012_s
+ N_VPWR_M1016_s N_VPWR_M1005_s N_VPWR_M1009_s N_VPWR_c_327_n N_VPWR_c_328_n
+ N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n
+ N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n
+ N_VPWR_c_339_n N_VPWR_c_340_n VPWR N_VPWR_c_341_n N_VPWR_c_342_n
+ N_VPWR_c_343_n N_VPWR_c_326_n PM_SKY130_FD_SC_HD__NAND2B_4%VPWR
x_PM_SKY130_FD_SC_HD__NAND2B_4%Y N_Y_M1002_s N_Y_M1007_s N_Y_M1000_d N_Y_M1015_d
+ N_Y_M1001_d N_Y_M1006_d N_Y_c_407_n N_Y_c_409_n N_Y_c_426_n N_Y_c_410_n
+ N_Y_c_433_n N_Y_c_436_n N_Y_c_411_n N_Y_c_412_n N_Y_c_459_n N_Y_c_413_n
+ N_Y_c_414_n Y Y Y N_Y_c_446_n PM_SKY130_FD_SC_HD__NAND2B_4%Y
x_PM_SKY130_FD_SC_HD__NAND2B_4%VGND N_VGND_M1017_d N_VGND_M1004_s N_VGND_M1011_s
+ N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n
+ N_VGND_c_507_n N_VGND_c_508_n VGND N_VGND_c_509_n N_VGND_c_510_n
+ N_VGND_c_511_n N_VGND_c_512_n PM_SKY130_FD_SC_HD__NAND2B_4%VGND
x_PM_SKY130_FD_SC_HD__NAND2B_4%A_215_47# N_A_215_47#_M1002_d N_A_215_47#_M1003_d
+ N_A_215_47#_M1010_d N_A_215_47#_M1008_d N_A_215_47#_M1013_d
+ N_A_215_47#_c_575_n N_A_215_47#_c_576_n N_A_215_47#_c_588_n
+ N_A_215_47#_c_595_n N_A_215_47#_c_577_n N_A_215_47#_c_578_n
+ N_A_215_47#_c_602_n N_A_215_47#_c_579_n N_A_215_47#_c_580_n
+ N_A_215_47#_c_581_n PM_SKY130_FD_SC_HD__NAND2B_4%A_215_47#
cc_1 VNB N_A_N_M1017_g 0.0265299f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB A_N 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_93_n 0.0377473f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_47#_M1002_g 0.0216349f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_47#_M1000_g 5.60601e-19 $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_6 VNB N_A_27_47#_M1003_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1012_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1007_g 0.0172529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1015_g 4.47552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1010_g 0.0173402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1016_g 4.3327e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_125_n 0.0183479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_126_n 0.00446253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_127_n 6.46682e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_128_n 0.0112315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_129_n 0.0116177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_130_n 0.00228535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_131_n 0.0328703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_132_n 0.0593722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_M1004_g 0.0177114f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_B_M1001_g 4.70147e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_22 VNB N_B_M1008_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_23 VNB N_B_M1005_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_24 VNB N_B_M1011_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_B_M1006_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B_M1013_g 0.0237242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_B_M1009_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB B 0.0159396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_B_c_247_n 0.0583981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_B_c_248_n 0.0366487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_326_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_407_n 0.00505016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB Y 0.00123574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_502_n 0.00482655f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_35 VNB N_VGND_c_503_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_504_n 0.00179046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_505_n 0.057292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_506_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_507_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_508_n 0.00340168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_509_n 0.017162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_510_n 0.0210728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_511_n 0.271667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_512_n 0.00372004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_215_47#_c_575_n 0.00232453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_215_47#_c_576_n 0.00646531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_215_47#_c_577_n 0.00354457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_215_47#_c_578_n 0.00218776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_215_47#_c_579_n 0.0128501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_215_47#_c_580_n 0.0175671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_215_47#_c_581_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VPB N_A_N_M1014_g 0.0305238f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_53 VPB N_A_N_c_93_n 0.00668925f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_54 VPB N_A_27_47#_M1000_g 0.0239395f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_55 VPB N_A_27_47#_M1012_g 0.0191612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_M1015_g 0.019143f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_M1016_g 0.0190705f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_137_n 0.0315997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_127_n 0.00391998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_139_n 0.013161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_B_M1001_g 0.0196376f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_62 VPB N_B_M1005_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_63 VPB N_B_M1006_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_B_M1009_g 0.0274817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_327_n 0.0100313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_328_n 0.00732817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_329_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_330_n 0.00412115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_331_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_332_n 0.0152212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_333_n 0.043309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_334_n 0.00605347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_335_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_336_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_337_n 0.0182802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_338_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_339_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_340_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_341_n 0.0178188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_342_n 0.0189004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_343_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_326_n 0.0484366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_Y_c_409_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_Y_c_410_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_Y_c_411_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_Y_c_412_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_Y_c_413_n 0.005634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_Y_c_414_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB Y 0.00133154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB Y 6.61229e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 N_A_N_M1017_g N_A_27_47#_c_125_n 0.00717364f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_92 N_A_N_M1014_g N_A_27_47#_c_137_n 0.0106812f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_N_M1017_g N_A_27_47#_c_126_n 0.00599295f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_94 N_A_N_c_93_n N_A_27_47#_c_127_n 0.0063209f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_N_M1017_g N_A_27_47#_c_129_n 0.0130359f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_96 A_N N_A_27_47#_c_129_n 0.0239253f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_97 N_A_N_c_93_n N_A_27_47#_c_129_n 0.00669833f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_N_M1014_g N_A_27_47#_c_139_n 0.0168408f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_99 A_N N_A_27_47#_c_139_n 0.024207f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A_N_c_93_n N_A_27_47#_c_139_n 0.00648679f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_101 A_N N_A_27_47#_c_130_n 0.0167772f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A_N_c_93_n N_A_27_47#_c_130_n 0.00240443f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_N_c_93_n N_A_27_47#_c_131_n 0.00567041f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_N_M1014_g N_VPWR_c_327_n 0.0048073f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_N_M1014_g N_VPWR_c_328_n 0.00354484f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_N_M1014_g N_VPWR_c_341_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_N_M1014_g N_VPWR_c_326_n 0.0117818f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_N_M1017_g N_VGND_c_502_n 0.00442456f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_N_M1017_g N_VGND_c_509_n 0.00421248f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A_N_M1017_g N_VGND_c_511_n 0.00799131f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_111 N_A_N_M1017_g N_A_215_47#_c_576_n 0.00337712f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A_27_47#_M1010_g N_B_M1004_g 0.0182436f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_27_47#_M1016_g N_B_M1001_g 0.0182436f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_132_n B 7.64104e-19 $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_132_n N_B_c_247_n 0.0182436f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_139_n N_VPWR_M1014_d 0.00432882f $X=0.695 $Y=1.555 $X2=-0.19
+ $Y2=-0.24
cc_117 N_A_27_47#_M1000_g N_VPWR_c_328_n 0.00424918f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_c_137_n N_VPWR_c_328_n 0.00556717f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_128_n N_VPWR_c_328_n 0.0256544f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_139_n N_VPWR_c_328_n 0.0174601f $X=0.695 $Y=1.555 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_131_n N_VPWR_c_328_n 0.0063996f $X=1.335 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1012_g N_VPWR_c_329_n 0.00146448f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_M1015_g N_VPWR_c_329_n 0.00268723f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_M1016_g N_VPWR_c_330_n 0.00468711f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_128_n N_VPWR_c_334_n 0.00701209f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_139_n N_VPWR_c_334_n 0.0147376f $X=0.695 $Y=1.555 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_M1000_g N_VPWR_c_335_n 0.00541359f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_M1012_g N_VPWR_c_335_n 0.00541359f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_M1015_g N_VPWR_c_337_n 0.00541359f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_27_47#_M1016_g N_VPWR_c_337_n 0.00518588f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_c_137_n N_VPWR_c_341_n 0.0213966f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_132 N_A_27_47#_M1014_s N_VPWR_c_326_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_M1000_g N_VPWR_c_326_n 0.0108276f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_27_47#_M1012_g N_VPWR_c_326_n 0.00950154f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_27_47#_M1015_g N_VPWR_c_326_n 0.00950154f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_M1016_g N_VPWR_c_326_n 0.0090482f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_137_n N_VPWR_c_326_n 0.0126193f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1002_g N_Y_c_407_n 0.00398755f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A_27_47#_M1003_g N_Y_c_407_n 0.0112239f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1007_g N_Y_c_407_n 0.0125587f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_128_n N_Y_c_407_n 0.0555084f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_132_n N_Y_c_407_n 0.00415773f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_27_47#_M1000_g N_Y_c_409_n 0.0033016f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_27_47#_M1012_g N_Y_c_409_n 0.00149073f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_128_n N_Y_c_409_n 0.026643f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_132_n N_Y_c_409_n 0.00206439f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_27_47#_M1000_g N_Y_c_426_n 0.00902485f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_27_47#_M1012_g N_Y_c_426_n 0.00975139f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_27_47#_M1015_g N_Y_c_426_n 6.1949e-19 $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_27_47#_M1012_g N_Y_c_410_n 0.0120357f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_27_47#_M1015_g N_Y_c_410_n 0.0130373f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_128_n N_Y_c_410_n 0.0304181f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_132_n N_Y_c_410_n 0.0019951f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_27_47#_M1012_g N_Y_c_433_n 6.19133e-19 $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_27_47#_M1015_g N_Y_c_433_n 0.00975139f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_27_47#_M1016_g N_Y_c_433_n 0.0107205f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_27_47#_M1016_g N_Y_c_436_n 6.13802e-19 $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_27_47#_M1016_g N_Y_c_413_n 0.014195f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_27_47#_M1007_g Y 0.00309532f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A_27_47#_M1015_g Y 0.00387565f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_27_47#_M1010_g Y 0.00333298f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_27_47#_M1016_g Y 0.00418035f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_128_n Y 0.0155586f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_132_n Y 0.0208995f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_27_47#_M1015_g Y 0.00180793f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_27_47#_M1016_g Y 0.0013666f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_27_47#_M1010_g N_Y_c_446_n 0.00395781f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_129_n N_VGND_M1017_d 0.0043755f $X=0.695 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_27_47#_M1002_g N_VGND_c_502_n 0.00205426f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_128_n N_VGND_c_502_n 3.11831e-19 $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_129_n N_VGND_c_502_n 0.0139975f $X=0.695 $Y=0.81 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1002_g N_VGND_c_505_n 0.00357877f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A_27_47#_M1003_g N_VGND_c_505_n 0.00357877f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1007_g N_VGND_c_505_n 0.00357877f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1010_g N_VGND_c_505_n 0.00357877f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_125_n N_VGND_c_509_n 0.0208545f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_129_n N_VGND_c_509_n 0.00207273f $X=0.695 $Y=0.81 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_M1017_s N_VGND_c_511_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1002_g N_VGND_c_511_n 0.00655123f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1003_g N_VGND_c_511_n 0.00522516f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_27_47#_M1007_g N_VGND_c_511_n 0.00522516f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1010_g N_VGND_c_511_n 0.00528897f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_125_n N_VGND_c_511_n 0.0124928f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_129_n N_VGND_c_511_n 0.00467649f $X=0.695 $Y=0.81 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_M1002_g N_A_215_47#_c_576_n 4.61765e-19 $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_125_n N_A_215_47#_c_576_n 0.00500305f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_128_n N_A_215_47#_c_576_n 0.0201437f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_129_n N_A_215_47#_c_576_n 0.0119729f $X=0.695 $Y=0.81 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_131_n N_A_215_47#_c_576_n 0.00588114f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1002_g N_A_215_47#_c_588_n 0.0103313f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1003_g N_A_215_47#_c_588_n 0.00866705f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1007_g N_A_215_47#_c_588_n 0.00866705f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1010_g N_A_215_47#_c_588_n 0.0119423f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_128_n N_A_215_47#_c_588_n 0.00348394f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_132_n N_A_215_47#_c_588_n 2.87379e-19 $X=2.67 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_M1010_g N_A_215_47#_c_577_n 7.98062e-19 $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_197 N_B_M1001_g N_VPWR_c_330_n 0.00148704f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B_M1005_g N_VPWR_c_331_n 0.00146448f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B_M1006_g N_VPWR_c_331_n 0.00268723f $X=3.945 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B_M1009_g N_VPWR_c_333_n 0.0266148f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_201 B N_VPWR_c_333_n 0.0218086f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_202 N_B_c_248_n N_VPWR_c_333_n 0.00557f $X=4.605 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B_M1001_g N_VPWR_c_339_n 0.00541359f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_204 N_B_M1005_g N_VPWR_c_339_n 0.00541359f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B_M1006_g N_VPWR_c_342_n 0.00541359f $X=3.945 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B_M1009_g N_VPWR_c_342_n 0.00541359f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B_M1001_g N_VPWR_c_326_n 0.00956534f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B_M1005_g N_VPWR_c_326_n 0.00950154f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B_M1006_g N_VPWR_c_326_n 0.00950154f $X=3.945 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B_M1009_g N_VPWR_c_326_n 0.0108063f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B_M1001_g N_Y_c_433_n 6.34334e-19 $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B_M1001_g N_Y_c_436_n 0.00978018f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B_M1005_g N_Y_c_436_n 0.00975139f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B_M1006_g N_Y_c_436_n 6.1949e-19 $X=3.945 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B_M1005_g N_Y_c_411_n 0.0120357f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B_M1006_g N_Y_c_411_n 0.0120357f $X=3.945 $Y=1.985 $X2=0 $Y2=0
cc_217 B N_Y_c_411_n 0.0366837f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_218 N_B_c_247_n N_Y_c_411_n 0.0019951f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_219 N_B_M1006_g N_Y_c_412_n 0.00149073f $X=3.945 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B_M1009_g N_Y_c_412_n 0.00527256f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_221 B N_Y_c_412_n 0.026643f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_222 N_B_c_247_n N_Y_c_412_n 0.00206439f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B_M1005_g N_Y_c_459_n 6.1949e-19 $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_224 N_B_M1006_g N_Y_c_459_n 0.00975139f $X=3.945 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B_M1009_g N_Y_c_459_n 0.00964729f $X=4.365 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B_M1001_g N_Y_c_413_n 0.0135551f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B_M1001_g N_Y_c_414_n 0.00155569f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_228 N_B_M1005_g N_Y_c_414_n 0.00149073f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_229 B N_Y_c_414_n 0.0262578f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_230 N_B_c_247_n N_Y_c_414_n 0.00206439f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B_M1004_g Y 0.00258377f $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_232 B Y 0.00626938f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_233 N_B_M1004_g N_VGND_c_503_n 0.00268723f $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_234 N_B_M1008_g N_VGND_c_503_n 0.00146448f $X=3.525 $Y=0.56 $X2=0 $Y2=0
cc_235 N_B_M1011_g N_VGND_c_504_n 0.00150833f $X=3.945 $Y=0.56 $X2=0 $Y2=0
cc_236 N_B_M1013_g N_VGND_c_504_n 0.00849805f $X=4.365 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B_M1004_g N_VGND_c_505_n 0.00420723f $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B_M1008_g N_VGND_c_507_n 0.00422241f $X=3.525 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B_M1011_g N_VGND_c_507_n 0.00422241f $X=3.945 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B_M1013_g N_VGND_c_510_n 0.00377504f $X=4.365 $Y=0.56 $X2=0 $Y2=0
cc_241 N_B_M1004_g N_VGND_c_511_n 0.00576944f $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B_M1008_g N_VGND_c_511_n 0.00569656f $X=3.525 $Y=0.56 $X2=0 $Y2=0
cc_243 N_B_M1011_g N_VGND_c_511_n 0.00569656f $X=3.945 $Y=0.56 $X2=0 $Y2=0
cc_244 N_B_M1013_g N_VGND_c_511_n 0.00559784f $X=4.365 $Y=0.56 $X2=0 $Y2=0
cc_245 N_B_M1004_g N_A_215_47#_c_595_n 0.00244813f $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_246 N_B_M1004_g N_A_215_47#_c_577_n 0.00528137f $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_247 N_B_M1008_g N_A_215_47#_c_577_n 4.58193e-19 $X=3.525 $Y=0.56 $X2=0 $Y2=0
cc_248 N_B_M1004_g N_A_215_47#_c_578_n 0.0100507f $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_249 N_B_M1008_g N_A_215_47#_c_578_n 0.0088553f $X=3.525 $Y=0.56 $X2=0 $Y2=0
cc_250 B N_A_215_47#_c_578_n 0.029722f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_251 N_B_c_247_n N_A_215_47#_c_578_n 0.00205999f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B_M1004_g N_A_215_47#_c_602_n 5.19281e-19 $X=3.105 $Y=0.56 $X2=0 $Y2=0
cc_253 N_B_M1008_g N_A_215_47#_c_602_n 0.00620543f $X=3.525 $Y=0.56 $X2=0 $Y2=0
cc_254 N_B_M1011_g N_A_215_47#_c_602_n 0.00649586f $X=3.945 $Y=0.56 $X2=0 $Y2=0
cc_255 N_B_M1013_g N_A_215_47#_c_602_n 4.57134e-19 $X=4.365 $Y=0.56 $X2=0 $Y2=0
cc_256 N_B_M1011_g N_A_215_47#_c_579_n 0.00890471f $X=3.945 $Y=0.56 $X2=0 $Y2=0
cc_257 N_B_M1013_g N_A_215_47#_c_579_n 0.0144772f $X=4.365 $Y=0.56 $X2=0 $Y2=0
cc_258 B N_A_215_47#_c_579_n 0.0712575f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_259 N_B_c_247_n N_A_215_47#_c_579_n 0.00205999f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B_c_248_n N_A_215_47#_c_579_n 0.00773686f $X=4.605 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B_M1013_g N_A_215_47#_c_580_n 0.011215f $X=4.365 $Y=0.56 $X2=0 $Y2=0
cc_262 N_B_M1008_g N_A_215_47#_c_581_n 0.00116017f $X=3.525 $Y=0.56 $X2=0 $Y2=0
cc_263 N_B_M1011_g N_A_215_47#_c_581_n 0.00116017f $X=3.945 $Y=0.56 $X2=0 $Y2=0
cc_264 B N_A_215_47#_c_581_n 0.0265408f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_265 N_B_c_247_n N_A_215_47#_c_581_n 0.00213429f $X=4.44 $Y=1.16 $X2=0 $Y2=0
cc_266 N_VPWR_c_326_n N_Y_M1000_d 0.00215201f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_267 N_VPWR_c_326_n N_Y_M1015_d 0.00215201f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_268 N_VPWR_c_326_n N_Y_M1001_d 0.00215201f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_c_326_n N_Y_M1006_d 0.00215201f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_328_n N_Y_c_409_n 0.0108853f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_271 N_VPWR_c_335_n N_Y_c_426_n 0.0189039f $X=1.955 $Y=2.72 $X2=0 $Y2=0
cc_272 N_VPWR_c_326_n N_Y_c_426_n 0.0122217f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_273 N_VPWR_M1012_s N_Y_c_410_n 0.00167154f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_274 N_VPWR_c_329_n N_Y_c_410_n 0.0129161f $X=2.04 $Y=2 $X2=0 $Y2=0
cc_275 N_VPWR_c_330_n N_Y_c_433_n 0.0466782f $X=2.895 $Y=2 $X2=0 $Y2=0
cc_276 N_VPWR_c_337_n N_Y_c_433_n 0.0199266f $X=2.81 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_326_n N_Y_c_433_n 0.0127308f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_339_n N_Y_c_436_n 0.0189039f $X=3.65 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_326_n N_Y_c_436_n 0.0122217f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_M1005_s N_Y_c_411_n 0.00167154f $X=3.6 $Y=1.485 $X2=0 $Y2=0
cc_281 N_VPWR_c_331_n N_Y_c_411_n 0.0129161f $X=3.735 $Y=2 $X2=0 $Y2=0
cc_282 N_VPWR_c_333_n N_Y_c_412_n 0.0123489f $X=4.685 $Y=1.66 $X2=0 $Y2=0
cc_283 N_VPWR_c_333_n N_Y_c_459_n 0.0547633f $X=4.685 $Y=1.66 $X2=0 $Y2=0
cc_284 N_VPWR_c_342_n N_Y_c_459_n 0.0189039f $X=4.52 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_326_n N_Y_c_459_n 0.0122217f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_M1016_s N_Y_c_413_n 0.00209012f $X=2.745 $Y=1.485 $X2=0 $Y2=0
cc_287 N_VPWR_c_330_n N_Y_c_413_n 0.0134129f $X=2.895 $Y=2 $X2=0 $Y2=0
cc_288 N_Y_M1002_s N_VGND_c_511_n 0.00216833f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_289 N_Y_M1007_s N_VGND_c_511_n 0.00216833f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_290 N_Y_c_407_n N_A_215_47#_M1003_d 0.00162207f $X=2.375 $Y=0.77 $X2=0 $Y2=0
cc_291 N_Y_c_407_n N_A_215_47#_c_576_n 0.0120104f $X=2.375 $Y=0.77 $X2=0 $Y2=0
cc_292 N_Y_M1002_s N_A_215_47#_c_588_n 0.00305599f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_293 N_Y_M1007_s N_A_215_47#_c_588_n 0.00305226f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_294 N_Y_c_407_n N_A_215_47#_c_588_n 0.0447682f $X=2.375 $Y=0.77 $X2=0 $Y2=0
cc_295 N_Y_c_446_n N_A_215_47#_c_588_n 0.0154172f $X=2.507 $Y=0.905 $X2=0 $Y2=0
cc_296 N_Y_c_413_n N_A_215_47#_c_577_n 0.00933129f $X=3.15 $Y=1.555 $X2=0 $Y2=0
cc_297 N_Y_c_446_n N_A_215_47#_c_577_n 0.0230641f $X=2.507 $Y=0.905 $X2=0 $Y2=0
cc_298 N_Y_c_413_n N_A_215_47#_c_578_n 0.00240615f $X=3.15 $Y=1.555 $X2=0 $Y2=0
cc_299 N_VGND_c_511_n N_A_215_47#_M1002_d 0.00209324f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_300 N_VGND_c_511_n N_A_215_47#_M1003_d 0.00215227f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_c_511_n N_A_215_47#_M1010_d 0.00227252f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_511_n N_A_215_47#_M1008_d 0.00215201f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_303 N_VGND_c_511_n N_A_215_47#_M1013_d 0.00354473f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_502_n N_A_215_47#_c_575_n 0.0135471f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_305 N_VGND_c_505_n N_A_215_47#_c_575_n 0.0173346f $X=3.23 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_511_n N_A_215_47#_c_575_n 0.00961661f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_502_n N_A_215_47#_c_576_n 0.00470956f $X=0.68 $Y=0.38 $X2=0
+ $Y2=0
cc_308 N_VGND_c_505_n N_A_215_47#_c_588_n 0.0837338f $X=3.23 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_511_n N_A_215_47#_c_588_n 0.0540361f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_505_n N_A_215_47#_c_595_n 0.015453f $X=3.23 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_511_n N_A_215_47#_c_595_n 0.00940698f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_M1004_s N_A_215_47#_c_578_n 0.00162148f $X=3.18 $Y=0.235 $X2=0
+ $Y2=0
cc_313 N_VGND_c_503_n N_A_215_47#_c_578_n 0.0122675f $X=3.315 $Y=0.38 $X2=0
+ $Y2=0
cc_314 N_VGND_c_505_n N_A_215_47#_c_578_n 0.00203746f $X=3.23 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_507_n N_A_215_47#_c_578_n 0.00203746f $X=4.07 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_511_n N_A_215_47#_c_578_n 0.00845923f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_507_n N_A_215_47#_c_602_n 0.0188551f $X=4.07 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_c_511_n N_A_215_47#_c_602_n 0.0122069f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_M1011_s N_A_215_47#_c_579_n 0.00162148f $X=4.02 $Y=0.235 $X2=0
+ $Y2=0
cc_320 N_VGND_c_504_n N_A_215_47#_c_579_n 0.0136249f $X=4.155 $Y=0.38 $X2=0
+ $Y2=0
cc_321 N_VGND_c_507_n N_A_215_47#_c_579_n 0.00203746f $X=4.07 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_510_n N_A_215_47#_c_579_n 0.00257231f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_511_n N_A_215_47#_c_579_n 0.00981815f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_324 N_VGND_c_504_n N_A_215_47#_c_580_n 0.0186968f $X=4.155 $Y=0.38 $X2=0
+ $Y2=0
cc_325 N_VGND_c_510_n N_A_215_47#_c_580_n 0.0230148f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_511_n N_A_215_47#_c_580_n 0.0126169f $X=4.83 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a311o_1.spice.SKY130_FD_SC_HD__A311O_1.pxi
* Created: Thu Aug 27 14:03:54 2020
* 
x_PM_SKY130_FD_SC_HD__A311O_1%A_75_199# N_A_75_199#_M1008_d N_A_75_199#_M1010_d
+ N_A_75_199#_M1000_d N_A_75_199#_M1011_g N_A_75_199#_M1004_g N_A_75_199#_c_64_n
+ N_A_75_199#_c_69_p N_A_75_199#_c_139_p N_A_75_199#_c_68_p N_A_75_199#_c_115_p
+ N_A_75_199#_c_82_p N_A_75_199#_c_83_p N_A_75_199#_c_149_p N_A_75_199#_c_150_p
+ N_A_75_199#_c_98_p N_A_75_199#_c_102_p N_A_75_199#_c_87_p N_A_75_199#_c_153_p
+ N_A_75_199#_c_128_p N_A_75_199#_c_59_n N_A_75_199#_c_60_n N_A_75_199#_c_61_n
+ N_A_75_199#_c_62_n PM_SKY130_FD_SC_HD__A311O_1%A_75_199#
x_PM_SKY130_FD_SC_HD__A311O_1%A3 N_A3_M1006_g N_A3_M1009_g A3 N_A3_c_170_n
+ N_A3_c_171_n PM_SKY130_FD_SC_HD__A311O_1%A3
x_PM_SKY130_FD_SC_HD__A311O_1%A2 N_A2_M1002_g N_A2_c_204_n N_A2_M1005_g A2 A2
+ N_A2_c_206_n PM_SKY130_FD_SC_HD__A311O_1%A2
x_PM_SKY130_FD_SC_HD__A311O_1%A1 N_A1_M1008_g N_A1_M1007_g A1 A1 N_A1_c_244_n
+ N_A1_c_245_n PM_SKY130_FD_SC_HD__A311O_1%A1
x_PM_SKY130_FD_SC_HD__A311O_1%B1 N_B1_M1001_g N_B1_M1003_g B1 N_B1_c_282_n
+ N_B1_c_283_n PM_SKY130_FD_SC_HD__A311O_1%B1
x_PM_SKY130_FD_SC_HD__A311O_1%C1 N_C1_c_315_n N_C1_M1010_g N_C1_M1000_g C1
+ N_C1_c_317_n PM_SKY130_FD_SC_HD__A311O_1%C1
x_PM_SKY130_FD_SC_HD__A311O_1%X N_X_M1011_s N_X_M1004_s N_X_c_340_n X X
+ N_X_c_343_n PM_SKY130_FD_SC_HD__A311O_1%X
x_PM_SKY130_FD_SC_HD__A311O_1%VPWR N_VPWR_M1004_d N_VPWR_M1002_d N_VPWR_c_360_n
+ VPWR N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_359_n N_VPWR_c_364_n
+ N_VPWR_c_365_n N_VPWR_c_366_n PM_SKY130_FD_SC_HD__A311O_1%VPWR
x_PM_SKY130_FD_SC_HD__A311O_1%A_201_297# N_A_201_297#_M1006_d
+ N_A_201_297#_M1007_d N_A_201_297#_c_412_n N_A_201_297#_c_423_n
+ N_A_201_297#_c_413_n N_A_201_297#_c_414_n N_A_201_297#_c_418_n
+ PM_SKY130_FD_SC_HD__A311O_1%A_201_297#
x_PM_SKY130_FD_SC_HD__A311O_1%VGND N_VGND_M1011_d N_VGND_M1001_d N_VGND_c_436_n
+ N_VGND_c_437_n VGND N_VGND_c_438_n N_VGND_c_439_n N_VGND_c_440_n
+ N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n PM_SKY130_FD_SC_HD__A311O_1%VGND
cc_1 VNB N_A_75_199#_c_59_n 0.00258127f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_2 VNB N_A_75_199#_c_60_n 0.0224102f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_3 VNB N_A_75_199#_c_61_n 0.00179679f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_4 VNB N_A_75_199#_c_62_n 0.0200973f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_5 VNB A3 0.00318933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A3_c_170_n 0.0201001f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_7 VNB N_A3_c_171_n 0.0178305f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_8 VNB N_A2_c_204_n 0.0187111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB A2 8.57749e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A2_c_206_n 0.0340812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A1 0.00408269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A1_c_244_n 0.0221071f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_13 VNB N_A1_c_245_n 0.0182188f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_14 VNB B1 0.00526451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_282_n 0.021217f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_B1_c_283_n 0.0182079f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_17 VNB N_C1_c_315_n 0.0234517f $X=-0.19 $Y=-0.24 $X2=2.245 $Y2=0.235
cc_18 VNB C1 0.00250714f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_C1_c_317_n 0.0454144f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_20 VNB N_X_c_340_n 0.0164574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB X 0.0275837f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_22 VNB N_VPWR_c_359_n 0.155873f $X=-0.19 $Y=-0.24 $X2=1.175 $Y2=0.655
cc_23 VNB N_VGND_c_436_n 0.00280508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_437_n 0.00561682f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_25 VNB N_VGND_c_438_n 0.0179052f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.825
cc_26 VNB N_VGND_c_439_n 0.0422313f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=0.74
cc_27 VNB N_VGND_c_440_n 0.0181454f $X=-0.19 $Y=-0.24 $X2=2.495 $Y2=0.74
cc_28 VNB N_VGND_c_441_n 0.201321f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=0.655
cc_29 VNB N_VGND_c_442_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_443_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=3.42 $Y2=1.96
cc_31 VPB N_A_75_199#_M1004_g 0.0215974f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_32 VPB N_A_75_199#_c_64_n 0.00148103f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.495
cc_33 VPB N_A_75_199#_c_60_n 0.00477141f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_34 VPB N_A3_M1006_g 0.0199422f $X=-0.19 $Y=1.305 $X2=3.285 $Y2=1.485
cc_35 VPB A3 0.00119915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A3_c_170_n 0.00406586f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_37 VPB N_A2_M1002_g 0.022489f $X=-0.19 $Y=1.305 $X2=3.285 $Y2=1.485
cc_38 VPB A2 0.00180717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A2_c_206_n 0.0090653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A1_M1007_g 0.022442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB A1 0.00196188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A1_c_244_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_43 VPB N_B1_M1003_g 0.0212531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB B1 0.0025273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B1_c_282_n 0.00406871f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_46 VPB N_C1_M1000_g 0.0277972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB C1 0.00250714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_C1_c_317_n 0.0110162f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_49 VPB X 0.0263273f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_50 VPB N_X_c_343_n 0.0187759f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.495
cc_51 VPB N_VPWR_c_360_n 0.00451452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_361_n 0.0181203f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_53 VPB N_VPWR_c_362_n 0.0457592f $X=-0.19 $Y=1.305 $X2=1.175 $Y2=0.425
cc_54 VPB N_VPWR_c_359_n 0.0453291f $X=-0.19 $Y=1.305 $X2=1.175 $Y2=0.655
cc_55 VPB N_VPWR_c_364_n 0.00468472f $X=-0.19 $Y=1.305 $X2=2.41 $Y2=0.425
cc_56 VPB N_VPWR_c_365_n 0.0153924f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=0.42
cc_57 VPB N_VPWR_c_366_n 0.0121855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 N_A_75_199#_M1004_g N_A3_M1006_g 0.0409774f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_59 N_A_75_199#_c_64_n N_A3_M1006_g 0.00286631f $X=0.65 $Y=1.495 $X2=0 $Y2=0
cc_60 N_A_75_199#_c_68_p N_A3_M1006_g 0.0159367f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_61 N_A_75_199#_c_69_p A3 0.0238966f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_62 N_A_75_199#_c_68_p A3 0.0228962f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_63 N_A_75_199#_c_59_n A3 0.0259822f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_75_199#_c_60_n A3 3.17302e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_75_199#_c_69_p N_A3_c_170_n 7.8959e-19 $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A_75_199#_c_68_p N_A3_c_170_n 0.00270331f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_67 N_A_75_199#_c_59_n N_A3_c_170_n 0.00286631f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_75_199#_c_60_n N_A3_c_170_n 0.0201765f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_75_199#_c_69_p N_A3_c_171_n 0.0118097f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A_75_199#_c_61_n N_A3_c_171_n 0.00365933f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_75_199#_c_62_n N_A3_c_171_n 0.0216921f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_75_199#_c_68_p N_A2_M1002_g 0.0163476f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_73 N_A_75_199#_c_69_p N_A2_c_204_n 0.00337726f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_75_199#_c_82_p N_A2_c_204_n 0.00499994f $X=1.175 $Y=0.655 $X2=0 $Y2=0
cc_75 N_A_75_199#_c_83_p N_A2_c_204_n 0.0139399f $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_76 N_A_75_199#_c_69_p A2 0.00445101f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_75_199#_c_68_p A2 0.0138341f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_75_199#_c_83_p A2 0.00558195f $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_79 N_A_75_199#_c_87_p A2 4.63021e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A_75_199#_c_68_p N_A2_c_206_n 0.00320276f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_75_199#_c_83_p N_A2_c_206_n 0.00347432f $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_82 N_A_75_199#_c_68_p N_A1_M1007_g 0.0119552f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A_75_199#_c_68_p A1 0.0222334f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_75_199#_c_83_p A1 0.00863216f $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_85 N_A_75_199#_c_87_p A1 0.0047963f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_75_199#_c_68_p N_A1_c_244_n 0.00185413f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A_75_199#_c_83_p N_A1_c_244_n 5.16916e-19 $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_88 N_A_75_199#_c_87_p N_A1_c_244_n 0.00103814f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A_75_199#_c_83_p N_A1_c_245_n 0.0102159f $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_90 N_A_75_199#_c_98_p N_A1_c_245_n 0.00454252f $X=2.41 $Y=0.655 $X2=0 $Y2=0
cc_91 N_A_75_199#_c_87_p N_A1_c_245_n 0.0036954f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_75_199#_c_68_p N_B1_M1003_g 0.0164907f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_93 N_A_75_199#_c_68_p B1 0.0331921f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_75_199#_c_102_p B1 0.0331921f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_75_199#_c_68_p N_B1_c_282_n 0.00256542f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_75_199#_c_102_p N_B1_c_282_n 0.00256542f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_75_199#_c_98_p N_B1_c_283_n 0.00367216f $X=2.41 $Y=0.655 $X2=0 $Y2=0
cc_98 N_A_75_199#_c_102_p N_B1_c_283_n 0.0130752f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_75_199#_c_102_p N_C1_c_315_n 0.015943f $X=3.335 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_75_199#_c_68_p N_C1_M1000_g 0.0190583f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A_75_199#_c_68_p C1 0.0127812f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A_75_199#_c_102_p C1 0.012603f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_75_199#_c_68_p N_C1_c_317_n 0.00163209f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_104 N_A_75_199#_c_102_p N_C1_c_317_n 0.0016034f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_75_199#_M1004_g X 0.0127682f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_75_199#_c_64_n X 0.00771894f $X=0.65 $Y=1.495 $X2=0 $Y2=0
cc_107 N_A_75_199#_c_115_p X 0.00839607f $X=0.735 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_75_199#_c_59_n X 0.0246821f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_75_199#_c_60_n X 0.00753248f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_75_199#_c_61_n X 0.00679878f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_75_199#_c_62_n X 0.00588184f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_75_199#_M1004_g N_X_c_343_n 0.00591964f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_75_199#_c_68_p N_VPWR_M1004_d 0.00237295f $X=3.335 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_75_199#_c_115_p N_VPWR_M1004_d 0.00204415f $X=0.735 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_75_199#_c_68_p N_VPWR_M1002_d 0.0182316f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_75_199#_M1004_g N_VPWR_c_360_n 0.00295236f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_75_199#_c_68_p N_VPWR_c_360_n 0.00223369f $X=3.335 $Y=1.58 $X2=0
+ $Y2=0
cc_118 N_A_75_199#_c_115_p N_VPWR_c_360_n 0.00424438f $X=0.735 $Y=1.58 $X2=0
+ $Y2=0
cc_119 N_A_75_199#_M1004_g N_VPWR_c_361_n 0.00579532f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_75_199#_c_128_p N_VPWR_c_362_n 0.0116048f $X=3.42 $Y=1.96 $X2=0 $Y2=0
cc_121 N_A_75_199#_M1000_d N_VPWR_c_359_n 0.00525232f $X=3.285 $Y=1.485 $X2=0
+ $Y2=0
cc_122 N_A_75_199#_M1004_g N_VPWR_c_359_n 0.0113774f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_75_199#_c_128_p N_VPWR_c_359_n 0.00646998f $X=3.42 $Y=1.96 $X2=0
+ $Y2=0
cc_124 N_A_75_199#_c_68_p N_A_201_297#_M1006_d 0.00513636f $X=3.335 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_125 N_A_75_199#_c_68_p N_A_201_297#_M1007_d 0.00603821f $X=3.335 $Y=1.58
+ $X2=0 $Y2=0
cc_126 N_A_75_199#_c_68_p N_A_201_297#_c_412_n 0.0164137f $X=3.335 $Y=1.58 $X2=0
+ $Y2=0
cc_127 N_A_75_199#_c_68_p N_A_201_297#_c_413_n 0.0588346f $X=3.335 $Y=1.58 $X2=0
+ $Y2=0
cc_128 N_A_75_199#_c_68_p N_A_201_297#_c_414_n 0.0155382f $X=3.335 $Y=1.58 $X2=0
+ $Y2=0
cc_129 N_A_75_199#_c_68_p A_544_297# 0.0150353f $X=3.335 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_75_199#_c_69_p N_VGND_M1011_d 0.00298535f $X=1.09 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_75_199#_c_139_p N_VGND_M1011_d 0.00244383f $X=0.735 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_132 N_A_75_199#_c_61_n N_VGND_M1011_d 6.77745e-19 $X=0.58 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_75_199#_c_102_p N_VGND_M1001_d 0.00663989f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_134 N_A_75_199#_c_69_p N_VGND_c_436_n 0.00862459f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_75_199#_c_139_p N_VGND_c_436_n 0.0102004f $X=0.735 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_75_199#_c_62_n N_VGND_c_436_n 0.00419788f $X=0.51 $Y=0.995 $X2=0
+ $Y2=0
cc_137 N_A_75_199#_c_102_p N_VGND_c_437_n 0.023107f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_75_199#_c_62_n N_VGND_c_438_n 0.00585385f $X=0.51 $Y=0.995 $X2=0
+ $Y2=0
cc_139 N_A_75_199#_c_69_p N_VGND_c_439_n 0.0023303f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_75_199#_c_83_p N_VGND_c_439_n 0.0604556f $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_141 N_A_75_199#_c_149_p N_VGND_c_439_n 0.0115639f $X=1.26 $Y=0.34 $X2=0 $Y2=0
cc_142 N_A_75_199#_c_150_p N_VGND_c_439_n 0.0118015f $X=2.41 $Y=0.425 $X2=0
+ $Y2=0
cc_143 N_A_75_199#_c_102_p N_VGND_c_439_n 0.00357612f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_75_199#_c_102_p N_VGND_c_440_n 0.00317056f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_75_199#_c_153_p N_VGND_c_440_n 0.011459f $X=3.42 $Y=0.42 $X2=0 $Y2=0
cc_146 N_A_75_199#_M1008_d N_VGND_c_441_n 0.00288515f $X=2.245 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_75_199#_M1010_d N_VGND_c_441_n 0.00370147f $X=3.285 $Y=0.235 $X2=0
+ $Y2=0
cc_148 N_A_75_199#_c_69_p N_VGND_c_441_n 0.0049831f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_75_199#_c_139_p N_VGND_c_441_n 0.00148234f $X=0.735 $Y=0.74 $X2=0
+ $Y2=0
cc_150 N_A_75_199#_c_83_p N_VGND_c_441_n 0.0382243f $X=2.325 $Y=0.34 $X2=0 $Y2=0
cc_151 N_A_75_199#_c_149_p N_VGND_c_441_n 0.00651702f $X=1.26 $Y=0.34 $X2=0
+ $Y2=0
cc_152 N_A_75_199#_c_150_p N_VGND_c_441_n 0.00651702f $X=2.41 $Y=0.425 $X2=0
+ $Y2=0
cc_153 N_A_75_199#_c_102_p N_VGND_c_441_n 0.0140331f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_75_199#_c_153_p N_VGND_c_441_n 0.00644035f $X=3.42 $Y=0.42 $X2=0
+ $Y2=0
cc_155 N_A_75_199#_c_62_n N_VGND_c_441_n 0.0117628f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_75_199#_c_69_p A_208_47# 0.00433146f $X=1.09 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_157 N_A_75_199#_c_82_p A_208_47# 0.00332487f $X=1.175 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_75_199#_c_83_p A_208_47# 0.00436823f $X=2.325 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_75_199#_c_149_p A_208_47# 0.00295929f $X=1.26 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_75_199#_c_83_p A_315_47# 0.0161421f $X=2.325 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A3_M1006_g N_A2_M1002_g 0.0209845f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A3_c_171_n N_A2_c_204_n 0.0239268f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_163 A3 A2 0.0178071f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A3_c_170_n A2 2.7047e-19 $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A3_c_171_n A2 9.12855e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_166 A3 N_A2_c_206_n 0.00273103f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A3_c_170_n N_A2_c_206_n 0.0207913f $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A3_M1006_g X 0.0012238f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A3_M1006_g N_VPWR_c_360_n 0.00161095f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A3_M1006_g N_VPWR_c_359_n 0.0106809f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A3_M1006_g N_VPWR_c_365_n 0.00585385f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A3_M1006_g N_VPWR_c_366_n 5.29988e-19 $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A3_c_171_n N_VGND_c_436_n 0.00794968f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A3_c_171_n N_VGND_c_439_n 0.00341689f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A3_c_171_n N_VGND_c_441_n 0.004321f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A2_M1002_g N_A1_M1007_g 0.0180875f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_c_204_n A1 6.93106e-19 $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_178 A2 A1 0.0312956f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_179 N_A2_c_206_n A1 0.00267575f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_180 A2 N_A1_c_244_n 3.30734e-19 $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_181 N_A2_c_206_n N_A1_c_244_n 0.0113969f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A2_c_204_n N_A1_c_245_n 0.0204534f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_183 A2 N_A1_c_245_n 8.21275e-19 $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A2_M1002_g N_VPWR_c_359_n 0.00425215f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A2_M1002_g N_VPWR_c_365_n 0.00348405f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A2_M1002_g N_VPWR_c_366_n 0.00816283f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A2_M1002_g N_A_201_297#_c_413_n 0.0111521f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A2_c_204_n N_VGND_c_436_n 0.00111186f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A2_c_204_n N_VGND_c_439_n 0.00357877f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A2_c_204_n N_VGND_c_441_n 0.00610311f $X=1.5 $Y=0.995 $X2=0 $Y2=0
cc_191 A2 A_315_47# 0.00258742f $X=1.525 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_192 N_A1_M1007_g N_B1_M1003_g 0.0220328f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_193 A1 B1 0.0158025f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_194 N_A1_c_244_n B1 0.0010569f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_195 A1 N_B1_c_282_n 0.00107131f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_196 N_A1_c_244_n N_B1_c_282_n 0.019867f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_197 A1 N_B1_c_283_n 9.17638e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_198 N_A1_c_245_n N_B1_c_283_n 0.0187941f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A1_M1007_g N_VPWR_c_362_n 0.00348405f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A1_M1007_g N_VPWR_c_359_n 0.00424101f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A1_M1007_g N_VPWR_c_366_n 0.00920925f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A1_M1007_g N_A_201_297#_c_413_n 0.0111521f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A1_c_245_n N_VGND_c_439_n 0.00357877f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A1_c_245_n N_VGND_c_441_n 0.00592608f $X=2.225 $Y=0.995 $X2=0 $Y2=0
cc_205 A1 A_315_47# 0.00238581f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_206 N_B1_c_283_n N_C1_c_315_n 0.0240541f $X=2.705 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_207 N_B1_M1003_g N_C1_M1000_g 0.0370246f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_208 B1 C1 0.0190675f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_209 N_B1_c_282_n C1 2.22562e-19 $X=2.705 $Y=1.16 $X2=0 $Y2=0
cc_210 B1 N_C1_c_317_n 0.00361954f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_211 N_B1_c_282_n N_C1_c_317_n 0.0132908f $X=2.705 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B1_M1003_g N_VPWR_c_362_n 0.00579312f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1003_g N_VPWR_c_359_n 0.0111099f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1003_g N_VPWR_c_366_n 0.00107507f $X=2.645 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_M1003_g N_A_201_297#_c_414_n 0.00348987f $X=2.645 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_B1_M1003_g N_A_201_297#_c_418_n 0.0083653f $X=2.645 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_B1_c_283_n N_VGND_c_437_n 0.00461366f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_283_n N_VGND_c_439_n 0.00428022f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_283_n N_VGND_c_441_n 0.00625899f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_220 N_C1_M1000_g N_VPWR_c_362_n 0.00585385f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_221 N_C1_M1000_g N_VPWR_c_359_n 0.0120456f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_222 N_C1_M1000_g N_A_201_297#_c_414_n 7.46923e-19 $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_C1_M1000_g N_A_201_297#_c_418_n 0.0020408f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_224 N_C1_c_315_n N_VGND_c_437_n 0.0046597f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_225 N_C1_c_315_n N_VGND_c_440_n 0.00428022f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_226 N_C1_c_315_n N_VGND_c_441_n 0.00704399f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_227 N_X_c_343_n N_VPWR_c_361_n 0.0173518f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_228 N_X_M1004_s N_VPWR_c_359_n 0.00232276f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_229 N_X_c_343_n N_VPWR_c_359_n 0.0126588f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_230 N_X_c_340_n N_VGND_c_438_n 0.0195709f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_231 N_X_M1011_s N_VGND_c_441_n 0.00209319f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_232 N_X_c_340_n N_VGND_c_441_n 0.0117951f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_233 N_VPWR_c_359_n N_A_201_297#_M1006_d 0.00330569f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_234 N_VPWR_c_359_n N_A_201_297#_M1007_d 0.0029666f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_359_n N_A_201_297#_c_423_n 0.0095318f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_365_n N_A_201_297#_c_423_n 0.0157576f $X=1.455 $Y=2.53 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_366_n N_A_201_297#_c_423_n 0.0154636f $X=2.125 $Y=2.53 $X2=0
+ $Y2=0
cc_238 N_VPWR_M1002_d N_A_201_297#_c_413_n 0.0134402f $X=1.485 $Y=1.485 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_362_n N_A_201_297#_c_413_n 0.00241441f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_359_n N_A_201_297#_c_413_n 0.0121417f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_365_n N_A_201_297#_c_413_n 0.00226665f $X=1.455 $Y=2.53 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_366_n N_A_201_297#_c_413_n 0.0303091f $X=2.125 $Y=2.53 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_362_n N_A_201_297#_c_418_n 0.0153379f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_359_n N_A_201_297#_c_418_n 0.00944122f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_366_n N_A_201_297#_c_418_n 0.0148615f $X=2.125 $Y=2.53 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_359_n A_544_297# 0.0177487f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_247 N_VGND_c_441_n A_208_47# 0.00328857f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_248 N_VGND_c_441_n A_315_47# 0.00420294f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__dlrtn_1.spice.SKY130_FD_SC_HD__DLRTN_1.pxi
* Created: Thu Aug 27 14:17:07 2020
* 
x_PM_SKY130_FD_SC_HD__DLRTN_1%GATE_N N_GATE_N_c_136_n N_GATE_N_c_131_n
+ N_GATE_N_M1019_g N_GATE_N_c_137_n N_GATE_N_M1011_g N_GATE_N_c_132_n
+ N_GATE_N_c_138_n GATE_N GATE_N N_GATE_N_c_134_n N_GATE_N_c_135_n
+ PM_SKY130_FD_SC_HD__DLRTN_1%GATE_N
x_PM_SKY130_FD_SC_HD__DLRTN_1%A_27_47# N_A_27_47#_M1019_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1012_g N_A_27_47#_M1000_g N_A_27_47#_M1016_g N_A_27_47#_M1003_g
+ N_A_27_47#_c_328_p N_A_27_47#_c_175_n N_A_27_47#_c_176_n N_A_27_47#_c_186_n
+ N_A_27_47#_c_187_n N_A_27_47#_c_188_n N_A_27_47#_c_177_n N_A_27_47#_c_178_n
+ N_A_27_47#_c_179_n N_A_27_47#_c_180_n N_A_27_47#_c_190_n N_A_27_47#_c_191_n
+ N_A_27_47#_c_192_n N_A_27_47#_c_193_n N_A_27_47#_c_194_n N_A_27_47#_c_181_n
+ N_A_27_47#_c_182_n N_A_27_47#_c_196_n N_A_27_47#_c_183_n
+ PM_SKY130_FD_SC_HD__DLRTN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRTN_1%D N_D_M1004_g N_D_M1018_g D N_D_c_343_n
+ N_D_c_344_n PM_SKY130_FD_SC_HD__DLRTN_1%D
x_PM_SKY130_FD_SC_HD__DLRTN_1%A_299_47# N_A_299_47#_M1004_s N_A_299_47#_M1018_s
+ N_A_299_47#_M1009_g N_A_299_47#_M1014_g N_A_299_47#_c_389_n
+ N_A_299_47#_c_382_n N_A_299_47#_c_390_n N_A_299_47#_c_391_n
+ N_A_299_47#_c_383_n N_A_299_47#_c_384_n N_A_299_47#_c_385_n
+ N_A_299_47#_c_386_n N_A_299_47#_c_387_n PM_SKY130_FD_SC_HD__DLRTN_1%A_299_47#
x_PM_SKY130_FD_SC_HD__DLRTN_1%A_193_47# N_A_193_47#_M1012_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1001_g N_A_193_47#_c_464_n N_A_193_47#_c_465_n
+ N_A_193_47#_M1007_g N_A_193_47#_c_471_n N_A_193_47#_c_467_n
+ N_A_193_47#_c_473_n N_A_193_47#_c_474_n N_A_193_47#_c_475_n
+ N_A_193_47#_c_476_n N_A_193_47#_c_477_n N_A_193_47#_c_478_n
+ N_A_193_47#_c_479_n PM_SKY130_FD_SC_HD__DLRTN_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRTN_1%A_724_21# N_A_724_21#_M1008_s N_A_724_21#_M1002_d
+ N_A_724_21#_M1017_g N_A_724_21#_M1006_g N_A_724_21#_M1010_g
+ N_A_724_21#_M1015_g N_A_724_21#_c_586_n N_A_724_21#_c_587_n
+ N_A_724_21#_c_578_n N_A_724_21#_c_597_p N_A_724_21#_c_579_n
+ N_A_724_21#_c_647_p N_A_724_21#_c_617_p N_A_724_21#_c_580_n
+ N_A_724_21#_c_581_n N_A_724_21#_c_625_p N_A_724_21#_c_582_n
+ PM_SKY130_FD_SC_HD__DLRTN_1%A_724_21#
x_PM_SKY130_FD_SC_HD__DLRTN_1%A_561_413# N_A_561_413#_M1016_d
+ N_A_561_413#_M1001_d N_A_561_413#_M1008_g N_A_561_413#_M1002_g
+ N_A_561_413#_c_674_n N_A_561_413#_c_675_n N_A_561_413#_c_682_n
+ N_A_561_413#_c_685_n N_A_561_413#_c_676_n N_A_561_413#_c_680_n
+ N_A_561_413#_c_677_n N_A_561_413#_c_678_n
+ PM_SKY130_FD_SC_HD__DLRTN_1%A_561_413#
x_PM_SKY130_FD_SC_HD__DLRTN_1%RESET_B N_RESET_B_M1005_g N_RESET_B_M1013_g
+ RESET_B RESET_B N_RESET_B_c_759_n N_RESET_B_c_760_n RESET_B
+ PM_SKY130_FD_SC_HD__DLRTN_1%RESET_B
x_PM_SKY130_FD_SC_HD__DLRTN_1%VPWR N_VPWR_M1011_d N_VPWR_M1018_d N_VPWR_M1006_d
+ N_VPWR_M1002_s N_VPWR_M1013_d N_VPWR_c_796_n N_VPWR_c_797_n N_VPWR_c_798_n
+ N_VPWR_c_799_n N_VPWR_c_800_n VPWR N_VPWR_c_801_n N_VPWR_c_802_n
+ N_VPWR_c_803_n N_VPWR_c_804_n N_VPWR_c_795_n N_VPWR_c_806_n N_VPWR_c_807_n
+ N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n
+ PM_SKY130_FD_SC_HD__DLRTN_1%VPWR
x_PM_SKY130_FD_SC_HD__DLRTN_1%Q N_Q_M1010_d N_Q_M1015_d Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HD__DLRTN_1%Q
x_PM_SKY130_FD_SC_HD__DLRTN_1%VGND N_VGND_M1019_d N_VGND_M1004_d N_VGND_M1017_d
+ N_VGND_M1005_d N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n VGND
+ N_VGND_c_912_n N_VGND_c_913_n N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n
+ N_VGND_c_917_n N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_920_n N_VGND_c_921_n
+ PM_SKY130_FD_SC_HD__DLRTN_1%VGND
cc_1 VNB N_GATE_N_c_131_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_N_c_132_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_134_n 0.0212744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_135_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1012_g 0.0397896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_175_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_8 VNB N_A_27_47#_c_176_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_177_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_178_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_179_n 0.0271287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_180_n 0.00378537f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_181_n 0.0230671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_182_n 0.0176114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_183_n 0.00459588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1004_g 0.025905f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_17 VNB N_D_M1018_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_343_n 0.00407935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_19 VNB N_D_c_344_n 0.0421785f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_20 VNB N_A_299_47#_M1014_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_299_47#_c_382_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_383_n 0.00496114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_47#_c_384_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_24 VNB N_A_299_47#_c_385_n 0.00265154f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_25 VNB N_A_299_47#_c_386_n 0.0274388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_299_47#_c_387_n 0.01709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_464_n 0.0133385f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_28 VNB N_A_193_47#_c_465_n 0.00520223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_M1007_g 0.0463933f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_30 VNB N_A_193_47#_c_467_n 0.0140955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_724_21#_M1017_g 0.0519341f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_32 VNB N_A_724_21#_c_578_n 0.00495607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_724_21#_c_579_n 0.00327629f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_724_21#_c_580_n 0.00361772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_724_21#_c_581_n 0.0300539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_724_21#_c_582_n 0.0222331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_561_413#_M1008_g 0.0239171f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_38 VNB N_A_561_413#_M1002_g 4.97209e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_39 VNB N_A_561_413#_c_674_n 0.0530275f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_40 VNB N_A_561_413#_c_675_n 0.00717034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_561_413#_c_676_n 0.00804154f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_42 VNB N_A_561_413#_c_677_n 0.0116303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_561_413#_c_678_n 0.00312597f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_44 VNB RESET_B 0.00868437f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_45 VNB N_RESET_B_c_759_n 0.0213453f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_46 VNB N_RESET_B_c_760_n 0.0192228f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_47 VNB N_VPWR_c_795_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB Q 0.0398558f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_49 VNB N_VGND_c_909_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_50 VNB N_VGND_c_910_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_51 VNB N_VGND_c_911_n 0.00592465f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_52 VNB N_VGND_c_912_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_53 VNB N_VGND_c_913_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_914_n 0.0412073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_915_n 0.0157049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_916_n 0.334293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_917_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_918_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_919_n 0.00507544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_920_n 0.0259335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_921_n 0.0161685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VPB N_GATE_N_c_136_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_63 VPB N_GATE_N_c_137_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_64 VPB N_GATE_N_c_138_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_65 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_66 VPB N_GATE_N_c_134_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_67 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_68 VPB N_A_27_47#_M1003_g 0.0212472f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_69 VPB N_A_27_47#_c_186_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_187_n 0.00556025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_188_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_177_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_190_n 0.0280095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_191_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_192_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_193_n 0.0035222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_194_n 0.0037442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_181_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_196_n 0.0328957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_183_n 2.971e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_D_M1018_g 0.0462846f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_82 VPB N_D_c_343_n 0.00235013f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_83 VPB N_A_299_47#_M1014_g 0.0366887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_299_47#_c_389_n 0.00712099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_299_47#_c_390_n 0.00415091f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_86 VPB N_A_299_47#_c_391_n 0.00290124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_299_47#_c_384_n 0.00361895f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_88 VPB N_A_193_47#_M1001_g 0.0316829f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_89 VPB N_A_193_47#_c_464_n 0.0172364f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_90 VPB N_A_193_47#_c_465_n 0.00687211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_193_47#_c_471_n 0.0117991f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_92 VPB N_A_193_47#_c_467_n 0.00804665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_193_47#_c_473_n 0.00293933f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_94 VPB N_A_193_47#_c_474_n 0.00515533f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_95 VPB N_A_193_47#_c_475_n 0.00238602f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_96 VPB N_A_193_47#_c_476_n 0.00711634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_193_47#_c_477_n 0.00114133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_193_47#_c_478_n 0.0104341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_193_47#_c_479_n 0.0126899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_724_21#_M1017_g 0.019403f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_101 VPB N_A_724_21#_M1006_g 0.0275278f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_102 VPB N_A_724_21#_M1015_g 0.0255236f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_103 VPB N_A_724_21#_c_586_n 0.00648694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_724_21#_c_587_n 0.0414704f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_105 VPB N_A_724_21#_c_580_n 0.00229942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_724_21#_c_581_n 0.0070014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_561_413#_M1002_g 0.026671f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_108 VPB N_A_561_413#_c_680_n 0.00517422f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_109 VPB N_A_561_413#_c_678_n 0.00493415f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_110 VPB N_RESET_B_M1013_g 0.0224286f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_111 VPB RESET_B 0.00549261f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_112 VPB N_RESET_B_c_759_n 0.00413333f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_113 VPB N_VPWR_c_796_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_797_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_798_n 0.00761302f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_116 VPB N_VPWR_c_799_n 0.00598254f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_117 VPB N_VPWR_c_800_n 0.00111355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_801_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_802_n 0.0295132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_803_n 0.0406078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_804_n 0.0150987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_795_n 0.0582089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_806_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_807_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_808_n 0.00555175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_809_n 0.00417584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_810_n 0.0129339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_811_n 0.0158867f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB Q 0.0464482f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_130 N_GATE_N_c_131_n N_A_27_47#_M1012_g 0.0187834f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_131 N_GATE_N_c_135_n N_A_27_47#_M1012_g 0.0041981f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_132 N_GATE_N_c_138_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_133 N_GATE_N_c_134_n N_A_27_47#_M1000_g 0.00527228f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_134 N_GATE_N_c_131_n N_A_27_47#_c_175_n 0.00663556f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_135 N_GATE_N_c_132_n N_A_27_47#_c_175_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_136 N_GATE_N_c_132_n N_A_27_47#_c_176_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_137 GATE_N N_A_27_47#_c_176_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_138 N_GATE_N_c_134_n N_A_27_47#_c_176_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_139 N_GATE_N_c_137_n N_A_27_47#_c_186_n 0.0135489f $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_140 N_GATE_N_c_138_n N_A_27_47#_c_186_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_141 N_GATE_N_c_137_n N_A_27_47#_c_188_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_142 N_GATE_N_c_138_n N_A_27_47#_c_188_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_143 GATE_N N_A_27_47#_c_188_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_144 N_GATE_N_c_134_n N_A_27_47#_c_188_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_145 N_GATE_N_c_134_n N_A_27_47#_c_177_n 0.00319708f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_146 N_GATE_N_c_132_n N_A_27_47#_c_178_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_147 GATE_N N_A_27_47#_c_178_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_148 N_GATE_N_c_135_n N_A_27_47#_c_178_n 0.0015185f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_149 N_GATE_N_c_136_n N_A_27_47#_c_191_n 0.0033897f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_150 N_GATE_N_c_138_n N_A_27_47#_c_191_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_151 GATE_N N_A_27_47#_c_191_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_152 N_GATE_N_c_136_n N_A_27_47#_c_192_n 7.60515e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_153 N_GATE_N_c_138_n N_A_27_47#_c_192_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_154 GATE_N N_A_27_47#_c_181_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_155 N_GATE_N_c_134_n N_A_27_47#_c_181_n 0.0165992f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_156 N_GATE_N_c_137_n N_VPWR_c_796_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_157 N_GATE_N_c_137_n N_VPWR_c_801_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_158 N_GATE_N_c_137_n N_VPWR_c_795_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_159 N_GATE_N_c_131_n N_VGND_c_909_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_160 N_GATE_N_c_131_n N_VGND_c_912_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_161 N_GATE_N_c_132_n N_VGND_c_912_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_162 N_GATE_N_c_131_n N_VGND_c_916_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_190_n N_D_M1018_g 0.00583826f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_190_n N_D_c_343_n 0.0087134f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_165 N_A_27_47#_M1012_g N_D_c_344_n 0.00520956f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_190_n N_A_299_47#_M1014_g 0.00493352f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_183_n N_A_299_47#_M1014_g 0.00369716f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_168 N_A_27_47#_c_190_n N_A_299_47#_c_390_n 0.0116478f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_190_n N_A_299_47#_c_391_n 0.0115067f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_179_n N_A_299_47#_c_383_n 9.56555e-19 $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_180_n N_A_299_47#_c_383_n 0.0129081f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_190_n N_A_299_47#_c_383_n 0.00675641f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_183_n N_A_299_47#_c_383_n 0.00178567f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_174 N_A_27_47#_c_190_n N_A_299_47#_c_384_n 0.0108506f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_179_n N_A_299_47#_c_386_n 0.0117556f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_180_n N_A_299_47#_c_386_n 9.50608e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_190_n N_A_299_47#_c_386_n 0.00107604f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_183_n N_A_299_47#_c_386_n 9.9633e-19 $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_179_n N_A_299_47#_c_387_n 0.00200147f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_180_n N_A_299_47#_c_387_n 2.04855e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_182_n N_A_299_47#_c_387_n 0.0197936f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_M1003_g N_A_193_47#_M1001_g 0.014011f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_187_n N_A_193_47#_M1001_g 0.00220245f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_180_n N_A_193_47#_c_464_n 7.03475e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_190_n N_A_193_47#_c_464_n 0.00144279f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_193_n N_A_193_47#_c_464_n 0.00140497f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_194_n N_A_193_47#_c_464_n 0.0049391f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_196_n N_A_193_47#_c_464_n 0.0184089f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_183_n N_A_193_47#_c_464_n 0.01293f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_179_n N_A_193_47#_c_465_n 0.0186665f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_180_n N_A_193_47#_c_465_n 0.00136525f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_179_n N_A_193_47#_M1007_g 0.0192792f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_180_n N_A_193_47#_M1007_g 0.00256423f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_182_n N_A_193_47#_M1007_g 0.0126141f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_183_n N_A_193_47#_M1007_g 0.0048126f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_190_n N_A_193_47#_c_471_n 0.00274258f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_193_n N_A_193_47#_c_471_n 7.88621e-19 $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_194_n N_A_193_47#_c_471_n 0.00220245f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_196_n N_A_193_47#_c_471_n 0.0160512f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_M1012_g N_A_193_47#_c_467_n 0.00779983f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_175_n N_A_193_47#_c_467_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_177_n N_A_193_47#_c_467_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_178_n N_A_193_47#_c_467_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_190_n N_A_193_47#_c_467_n 0.0184539f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_191_n N_A_193_47#_c_467_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_192_n N_A_193_47#_c_467_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_186_n N_A_193_47#_c_473_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_190_n N_A_193_47#_c_473_n 0.00195186f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_181_n N_A_193_47#_c_473_n 0.00779983f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_190_n N_A_193_47#_c_474_n 0.0871075f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_M1000_g N_A_193_47#_c_475_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_186_n N_A_193_47#_c_475_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_190_n N_A_193_47#_c_475_n 0.0259095f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_192_n N_A_193_47#_c_475_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_M1000_g N_A_193_47#_c_476_n 0.00779983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_187_n N_A_193_47#_c_477_n 0.00155445f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_190_n N_A_193_47#_c_477_n 0.0255946f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_190_n N_A_193_47#_c_478_n 0.00169866f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_193_n N_A_193_47#_c_478_n 0.00124306f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_183_n N_A_193_47#_c_478_n 0.00220245f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_221 N_A_27_47#_c_179_n N_A_193_47#_c_479_n 4.0812e-19 $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_180_n N_A_193_47#_c_479_n 0.00161882f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_190_n N_A_193_47#_c_479_n 0.0240266f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_193_n N_A_193_47#_c_479_n 0.00272314f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_196_n N_A_193_47#_c_479_n 2.5966e-19 $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_183_n N_A_193_47#_c_479_n 0.0454941f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_194_n N_A_724_21#_M1017_g 4.9921e-19 $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_183_n N_A_724_21#_M1017_g 2.17095e-19 $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_229 N_A_27_47#_M1003_g N_A_724_21#_M1006_g 0.0313447f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_187_n N_A_724_21#_c_587_n 8.09252e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_196_n N_A_724_21#_c_587_n 0.0313447f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_179_n N_A_561_413#_c_682_n 0.00144439f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_180_n N_A_561_413#_c_682_n 0.0162478f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_182_n N_A_561_413#_c_682_n 0.00412044f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_M1003_g N_A_561_413#_c_685_n 0.0116262f $X=3.335 $Y=2.275
+ $X2=0 $Y2=0
cc_236 N_A_27_47#_c_187_n N_A_561_413#_c_685_n 0.016081f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_193_n N_A_561_413#_c_685_n 0.00173361f $X=3.015 $Y=1.53
+ $X2=0 $Y2=0
cc_238 N_A_27_47#_c_196_n N_A_561_413#_c_685_n 0.00111122f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_239 N_A_27_47#_c_180_n N_A_561_413#_c_676_n 0.0204123f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_193_n N_A_561_413#_c_680_n 0.00130345f $X=3.015 $Y=1.53
+ $X2=0 $Y2=0
cc_241 N_A_27_47#_c_194_n N_A_561_413#_c_680_n 0.0359174f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_196_n N_A_561_413#_c_680_n 0.00856317f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_243 N_A_27_47#_c_183_n N_A_561_413#_c_680_n 0.00353544f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_244 N_A_27_47#_c_180_n N_A_561_413#_c_677_n 6.41977e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_196_n N_A_561_413#_c_677_n 0.00316305f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_246 N_A_27_47#_c_183_n N_A_561_413#_c_677_n 0.0176273f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_247 N_A_27_47#_c_186_n N_VPWR_M1011_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_248 N_A_27_47#_M1000_g N_VPWR_c_796_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_186_n N_VPWR_c_796_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_188_n N_VPWR_c_796_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_191_n N_VPWR_c_796_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_190_n N_VPWR_c_797_n 0.0019389f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_186_n N_VPWR_c_801_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_188_n N_VPWR_c_801_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_255 N_A_27_47#_M1000_g N_VPWR_c_802_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1003_g N_VPWR_c_803_n 0.00366111f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1000_g N_VPWR_c_795_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1003_g N_VPWR_c_795_n 0.00549379f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_186_n N_VPWR_c_795_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_188_n N_VPWR_c_795_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_175_n N_VGND_M1019_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_262 N_A_27_47#_M1012_g N_VGND_c_909_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_175_n N_VGND_c_909_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_177_n N_VGND_c_909_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_181_n N_VGND_c_909_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_182_n N_VGND_c_910_n 0.00174223f $X=2.8 $Y=0.705 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_328_p N_VGND_c_912_n 0.00713694f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_175_n N_VGND_c_912_n 0.00243651f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1012_g N_VGND_c_913_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_179_n N_VGND_c_914_n 9.43262e-19 $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_180_n N_VGND_c_914_n 0.00182549f $X=3.01 $Y=0.87 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_182_n N_VGND_c_914_n 0.00425892f $X=2.8 $Y=0.705 $X2=0 $Y2=0
cc_273 N_A_27_47#_M1019_s N_VGND_c_916_n 0.003754f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_274 N_A_27_47#_M1012_g N_VGND_c_916_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_328_p N_VGND_c_916_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_175_n N_VGND_c_916_n 0.00549708f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_179_n N_VGND_c_916_n 0.00121904f $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_180_n N_VGND_c_916_n 0.00328555f $X=3.01 $Y=0.87 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_182_n N_VGND_c_916_n 0.00628992f $X=2.8 $Y=0.705 $X2=0 $Y2=0
cc_280 N_D_c_344_n N_A_299_47#_M1014_g 0.0382098f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_281 N_D_M1018_g N_A_299_47#_c_389_n 0.012851f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_282 N_D_M1004_g N_A_299_47#_c_382_n 0.0144498f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_283 N_D_c_343_n N_A_299_47#_c_382_n 0.00627239f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_284 N_D_c_344_n N_A_299_47#_c_382_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_285 N_D_M1018_g N_A_299_47#_c_390_n 0.00794545f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_286 N_D_M1018_g N_A_299_47#_c_391_n 0.00412429f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_287 N_D_c_343_n N_A_299_47#_c_391_n 0.0229667f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_288 N_D_c_344_n N_A_299_47#_c_391_n 0.00131849f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_289 N_D_M1004_g N_A_299_47#_c_383_n 0.00563568f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_290 N_D_c_343_n N_A_299_47#_c_383_n 0.0107593f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_291 N_D_c_343_n N_A_299_47#_c_384_n 0.0164827f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_292 N_D_c_344_n N_A_299_47#_c_384_n 0.00552652f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_293 N_D_M1004_g N_A_299_47#_c_385_n 0.00120855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_294 N_D_c_343_n N_A_299_47#_c_385_n 0.0138491f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_295 N_D_c_344_n N_A_299_47#_c_385_n 0.0042466f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_296 N_D_M1004_g N_A_299_47#_c_386_n 0.0197208f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_297 N_D_M1004_g N_A_299_47#_c_387_n 0.015283f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_298 N_D_M1004_g N_A_193_47#_c_467_n 0.00203374f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_299 N_D_M1018_g N_A_193_47#_c_467_n 0.00459933f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_300 N_D_c_343_n N_A_193_47#_c_467_n 0.0209974f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_301 N_D_c_344_n N_A_193_47#_c_467_n 0.00256393f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_302 N_D_M1018_g N_A_193_47#_c_473_n 0.00134564f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_303 N_D_M1018_g N_A_193_47#_c_474_n 0.00294239f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_304 N_D_M1018_g N_VPWR_c_797_n 0.00304701f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_305 N_D_M1018_g N_VPWR_c_802_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_306 N_D_M1018_g N_VPWR_c_795_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_307 N_D_M1004_g N_VGND_c_910_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_308 N_D_M1004_g N_VGND_c_913_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_309 N_D_M1004_g N_VGND_c_916_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_310 N_D_c_344_n N_VGND_c_916_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_311 N_A_299_47#_M1014_g N_A_193_47#_M1001_g 0.0342299f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_312 N_A_299_47#_M1014_g N_A_193_47#_c_465_n 0.0248238f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_313 N_A_299_47#_c_389_n N_A_193_47#_c_467_n 0.0010921f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_314 N_A_299_47#_c_391_n N_A_193_47#_c_467_n 0.00859001f $X=1.785 $Y=1.58
+ $X2=0 $Y2=0
cc_315 N_A_299_47#_c_385_n N_A_193_47#_c_467_n 0.0191833f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_316 N_A_299_47#_c_389_n N_A_193_47#_c_473_n 0.0471072f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_317 N_A_299_47#_M1014_g N_A_193_47#_c_474_n 0.00365242f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_318 N_A_299_47#_c_389_n N_A_193_47#_c_474_n 0.022748f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_319 N_A_299_47#_c_390_n N_A_193_47#_c_474_n 0.00551435f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_320 N_A_299_47#_c_389_n N_A_193_47#_c_475_n 0.00273055f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_321 N_A_299_47#_M1014_g N_A_193_47#_c_477_n 0.00149195f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_322 N_A_299_47#_M1014_g N_A_193_47#_c_479_n 0.00673436f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_323 N_A_299_47#_c_390_n N_A_193_47#_c_479_n 0.00754519f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_324 N_A_299_47#_c_384_n N_A_193_47#_c_479_n 0.00645446f $X=2.055 $Y=1.495
+ $X2=0 $Y2=0
cc_325 N_A_299_47#_c_387_n N_A_561_413#_c_682_n 6.54613e-19 $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_326 N_A_299_47#_M1014_g N_VPWR_c_797_n 0.0223997f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_327 N_A_299_47#_c_389_n N_VPWR_c_797_n 0.0232987f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_328 N_A_299_47#_c_390_n N_VPWR_c_797_n 0.013562f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_329 N_A_299_47#_c_389_n N_VPWR_c_802_n 0.0159418f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_330 N_A_299_47#_M1014_g N_VPWR_c_803_n 0.00212864f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_331 N_A_299_47#_M1018_s N_VPWR_c_795_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_332 N_A_299_47#_M1014_g N_VPWR_c_795_n 0.00262666f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_333 N_A_299_47#_c_389_n N_VPWR_c_795_n 0.00576627f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_334 N_A_299_47#_c_383_n N_VGND_M1004_d 0.00156939f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_382_n N_VGND_c_910_n 0.00259081f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_336 N_A_299_47#_c_383_n N_VGND_c_910_n 0.0141976f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_337 N_A_299_47#_c_387_n N_VGND_c_910_n 0.00964732f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_382_n N_VGND_c_913_n 0.00255672f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_339 N_A_299_47#_c_385_n N_VGND_c_913_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_340 N_A_299_47#_c_386_n N_VGND_c_914_n 9.84895e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_341 N_A_299_47#_c_387_n N_VGND_c_914_n 0.0046653f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_342 N_A_299_47#_M1004_s N_VGND_c_916_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_343 N_A_299_47#_c_382_n N_VGND_c_916_n 0.00473142f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_344 N_A_299_47#_c_383_n N_VGND_c_916_n 0.00552372f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_345 N_A_299_47#_c_385_n N_VGND_c_916_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_c_386_n N_VGND_c_916_n 0.00117722f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_347 N_A_299_47#_c_387_n N_VGND_c_916_n 0.00454932f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_348 N_A_193_47#_M1007_g N_A_724_21#_M1017_g 0.0428016f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_349 N_A_193_47#_M1007_g N_A_561_413#_c_682_n 0.0125275f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_350 N_A_193_47#_M1001_g N_A_561_413#_c_685_n 0.00281839f $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_351 N_A_193_47#_M1007_g N_A_561_413#_c_676_n 0.0058879f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_352 N_A_193_47#_M1001_g N_A_561_413#_c_680_n 8.05921e-19 $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_353 N_A_193_47#_c_464_n N_A_561_413#_c_680_n 6.71539e-19 $X=3.145 $Y=1.32
+ $X2=0 $Y2=0
cc_354 N_A_193_47#_c_464_n N_A_561_413#_c_677_n 9.06019e-19 $X=3.145 $Y=1.32
+ $X2=0 $Y2=0
cc_355 N_A_193_47#_M1007_g N_A_561_413#_c_677_n 0.00230714f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_356 N_A_193_47#_c_474_n N_VPWR_M1018_d 6.81311e-19 $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_357 N_A_193_47#_c_476_n N_VPWR_c_796_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_358 N_A_193_47#_M1001_g N_VPWR_c_797_n 0.00357414f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_359 N_A_193_47#_c_474_n N_VPWR_c_797_n 0.0171797f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_360 N_A_193_47#_c_477_n N_VPWR_c_797_n 0.0013481f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_361 N_A_193_47#_c_479_n N_VPWR_c_797_n 0.00972665f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_362 N_A_193_47#_c_476_n N_VPWR_c_802_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_363 N_A_193_47#_M1001_g N_VPWR_c_803_n 0.00487021f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_364 N_A_193_47#_c_479_n N_VPWR_c_803_n 0.00456724f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_365 N_A_193_47#_M1001_g N_VPWR_c_795_n 0.00815857f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_366 N_A_193_47#_c_474_n N_VPWR_c_795_n 0.0516753f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_367 N_A_193_47#_c_475_n N_VPWR_c_795_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_368 N_A_193_47#_c_476_n N_VPWR_c_795_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_369 N_A_193_47#_c_477_n N_VPWR_c_795_n 0.0151013f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_479_n N_VPWR_c_795_n 0.00403974f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_c_474_n A_465_369# 0.00119229f $X=2.41 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_372 N_A_193_47#_c_477_n A_465_369# 0.00120144f $X=2.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_373 N_A_193_47#_c_479_n A_465_369# 0.0030615f $X=2.67 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_374 N_A_193_47#_M1007_g N_VGND_c_911_n 0.0017297f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_375 N_A_193_47#_c_467_n N_VGND_c_913_n 0.00732874f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_376 N_A_193_47#_M1007_g N_VGND_c_914_n 0.0037981f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_M1012_d N_VGND_c_916_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_378 N_A_193_47#_M1007_g N_VGND_c_916_n 0.00555936f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_467_n N_VGND_c_916_n 0.00616598f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_380 N_A_724_21#_c_578_n N_A_561_413#_M1008_g 0.0073654f $X=4.425 $Y=0.4 $X2=0
+ $Y2=0
cc_381 N_A_724_21#_c_597_p N_A_561_413#_M1008_g 0.00820318f $X=5.605 $Y=0.74
+ $X2=0 $Y2=0
cc_382 N_A_724_21#_c_579_n N_A_561_413#_M1008_g 8.67038e-19 $X=4.59 $Y=0.74
+ $X2=0 $Y2=0
cc_383 N_A_724_21#_c_586_n N_A_561_413#_M1002_g 0.0167742f $X=4.75 $Y=1.7 $X2=0
+ $Y2=0
cc_384 N_A_724_21#_c_587_n N_A_561_413#_M1002_g 0.00640354f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_385 N_A_724_21#_M1017_g N_A_561_413#_c_674_n 0.017529f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_386 N_A_724_21#_c_586_n N_A_561_413#_c_674_n 0.00837083f $X=4.75 $Y=1.7 $X2=0
+ $Y2=0
cc_387 N_A_724_21#_c_587_n N_A_561_413#_c_674_n 0.00424117f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_388 N_A_724_21#_c_579_n N_A_561_413#_c_674_n 0.00920019f $X=4.59 $Y=0.74
+ $X2=0 $Y2=0
cc_389 N_A_724_21#_M1017_g N_A_561_413#_c_682_n 0.00158904f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_390 N_A_724_21#_M1006_g N_A_561_413#_c_685_n 0.00369776f $X=3.695 $Y=2.275
+ $X2=0 $Y2=0
cc_391 N_A_724_21#_M1017_g N_A_561_413#_c_676_n 0.0109933f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_392 N_A_724_21#_M1017_g N_A_561_413#_c_680_n 0.0114233f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_393 N_A_724_21#_M1006_g N_A_561_413#_c_680_n 0.0143765f $X=3.695 $Y=2.275
+ $X2=0 $Y2=0
cc_394 N_A_724_21#_c_586_n N_A_561_413#_c_680_n 0.0249855f $X=4.75 $Y=1.7 $X2=0
+ $Y2=0
cc_395 N_A_724_21#_c_587_n N_A_561_413#_c_680_n 0.00797618f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_396 N_A_724_21#_M1017_g N_A_561_413#_c_677_n 0.00552416f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_397 N_A_724_21#_M1017_g N_A_561_413#_c_678_n 0.0170195f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_398 N_A_724_21#_c_586_n N_A_561_413#_c_678_n 0.0352918f $X=4.75 $Y=1.7 $X2=0
+ $Y2=0
cc_399 N_A_724_21#_c_587_n N_A_561_413#_c_678_n 0.00594586f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_400 N_A_724_21#_c_579_n N_A_561_413#_c_678_n 0.00652597f $X=4.59 $Y=0.74
+ $X2=0 $Y2=0
cc_401 N_A_724_21#_c_617_p N_RESET_B_M1013_g 0.0189052f $X=5.605 $Y=1.7 $X2=0
+ $Y2=0
cc_402 N_A_724_21#_c_580_n N_RESET_B_M1013_g 0.00560495f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_403 N_A_724_21#_c_586_n RESET_B 0.0131995f $X=4.75 $Y=1.7 $X2=0 $Y2=0
cc_404 N_A_724_21#_c_597_p RESET_B 0.057366f $X=5.605 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A_724_21#_c_579_n RESET_B 0.00496106f $X=4.59 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A_724_21#_c_617_p RESET_B 0.0299357f $X=5.605 $Y=1.7 $X2=0 $Y2=0
cc_407 N_A_724_21#_c_580_n RESET_B 0.028948f $X=5.84 $Y=1.16 $X2=0 $Y2=0
cc_408 N_A_724_21#_c_581_n RESET_B 0.00118675f $X=5.84 $Y=1.16 $X2=0 $Y2=0
cc_409 N_A_724_21#_c_625_p RESET_B 0.0127852f $X=4.845 $Y=1.755 $X2=0 $Y2=0
cc_410 N_A_724_21#_c_597_p N_RESET_B_c_759_n 0.00144439f $X=5.605 $Y=0.74 $X2=0
+ $Y2=0
cc_411 N_A_724_21#_c_617_p N_RESET_B_c_759_n 0.00139346f $X=5.605 $Y=1.7 $X2=0
+ $Y2=0
cc_412 N_A_724_21#_c_580_n N_RESET_B_c_759_n 7.78563e-19 $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_413 N_A_724_21#_c_581_n N_RESET_B_c_759_n 0.00628892f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_414 N_A_724_21#_c_578_n N_RESET_B_c_760_n 0.00151191f $X=4.425 $Y=0.4 $X2=0
+ $Y2=0
cc_415 N_A_724_21#_c_597_p N_RESET_B_c_760_n 0.0135455f $X=5.605 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A_724_21#_c_580_n N_RESET_B_c_760_n 0.00453224f $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_417 N_A_724_21#_c_586_n N_VPWR_M1002_s 0.00664759f $X=4.75 $Y=1.7 $X2=0 $Y2=0
cc_418 N_A_724_21#_c_617_p N_VPWR_M1013_d 0.0258799f $X=5.605 $Y=1.7 $X2=0 $Y2=0
cc_419 N_A_724_21#_c_580_n N_VPWR_M1013_d 9.71909e-19 $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_420 N_A_724_21#_M1006_g N_VPWR_c_798_n 0.0045387f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_421 N_A_724_21#_c_586_n N_VPWR_c_798_n 0.0157229f $X=4.75 $Y=1.7 $X2=0 $Y2=0
cc_422 N_A_724_21#_c_587_n N_VPWR_c_798_n 0.00522755f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_423 N_A_724_21#_c_586_n N_VPWR_c_800_n 0.0123588f $X=4.75 $Y=1.7 $X2=0 $Y2=0
cc_424 N_A_724_21#_M1006_g N_VPWR_c_803_n 0.00541489f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_425 N_A_724_21#_M1015_g N_VPWR_c_804_n 0.0046653f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_A_724_21#_M1002_d N_VPWR_c_795_n 0.00270514f $X=4.71 $Y=1.485 $X2=0
+ $Y2=0
cc_427 N_A_724_21#_M1006_g N_VPWR_c_795_n 0.0106979f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_428 N_A_724_21#_M1015_g N_VPWR_c_795_n 0.00879747f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_429 N_A_724_21#_c_586_n N_VPWR_c_795_n 0.0142526f $X=4.75 $Y=1.7 $X2=0 $Y2=0
cc_430 N_A_724_21#_c_587_n N_VPWR_c_795_n 0.00110429f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_431 N_A_724_21#_c_647_p N_VPWR_c_795_n 0.00724021f $X=4.845 $Y=2.27 $X2=0
+ $Y2=0
cc_432 N_A_724_21#_c_617_p N_VPWR_c_795_n 0.00858141f $X=5.605 $Y=1.7 $X2=0
+ $Y2=0
cc_433 N_A_724_21#_c_647_p N_VPWR_c_810_n 0.0121054f $X=4.845 $Y=2.27 $X2=0
+ $Y2=0
cc_434 N_A_724_21#_M1015_g N_VPWR_c_811_n 0.0120904f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_435 N_A_724_21#_c_617_p N_VPWR_c_811_n 0.039787f $X=5.605 $Y=1.7 $X2=0 $Y2=0
cc_436 N_A_724_21#_c_580_n Q 0.0503644f $X=5.84 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_724_21#_c_582_n Q 0.0210305f $X=5.875 $Y=0.995 $X2=0 $Y2=0
cc_438 N_A_724_21#_c_597_p N_VGND_M1005_d 0.0194842f $X=5.605 $Y=0.74 $X2=0
+ $Y2=0
cc_439 N_A_724_21#_c_580_n N_VGND_M1005_d 9.59589e-19 $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_440 N_A_724_21#_M1017_g N_VGND_c_911_n 0.0115393f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_441 N_A_724_21#_c_578_n N_VGND_c_911_n 0.0230011f $X=4.425 $Y=0.4 $X2=0 $Y2=0
cc_442 N_A_724_21#_M1017_g N_VGND_c_914_n 0.0046653f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_443 N_A_724_21#_c_582_n N_VGND_c_915_n 0.0046653f $X=5.875 $Y=0.995 $X2=0
+ $Y2=0
cc_444 N_A_724_21#_M1008_s N_VGND_c_916_n 0.00209319f $X=4.3 $Y=0.235 $X2=0
+ $Y2=0
cc_445 N_A_724_21#_M1017_g N_VGND_c_916_n 0.00813035f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_446 N_A_724_21#_c_578_n N_VGND_c_916_n 0.0131361f $X=4.425 $Y=0.4 $X2=0 $Y2=0
cc_447 N_A_724_21#_c_597_p N_VGND_c_916_n 0.0166334f $X=5.605 $Y=0.74 $X2=0
+ $Y2=0
cc_448 N_A_724_21#_c_582_n N_VGND_c_916_n 0.00891004f $X=5.875 $Y=0.995 $X2=0
+ $Y2=0
cc_449 N_A_724_21#_c_578_n N_VGND_c_920_n 0.0222092f $X=4.425 $Y=0.4 $X2=0 $Y2=0
cc_450 N_A_724_21#_c_597_p N_VGND_c_920_n 0.00732922f $X=5.605 $Y=0.74 $X2=0
+ $Y2=0
cc_451 N_A_724_21#_c_578_n N_VGND_c_921_n 0.0075261f $X=4.425 $Y=0.4 $X2=0 $Y2=0
cc_452 N_A_724_21#_c_597_p N_VGND_c_921_n 0.056372f $X=5.605 $Y=0.74 $X2=0 $Y2=0
cc_453 N_A_724_21#_c_581_n N_VGND_c_921_n 6.30284e-19 $X=5.84 $Y=1.16 $X2=0
+ $Y2=0
cc_454 N_A_724_21#_c_582_n N_VGND_c_921_n 0.0161125f $X=5.875 $Y=0.995 $X2=0
+ $Y2=0
cc_455 N_A_724_21#_c_597_p A_942_47# 0.00444569f $X=5.605 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_456 N_A_561_413#_M1002_g N_RESET_B_M1013_g 0.0244797f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_457 N_A_561_413#_M1008_g RESET_B 0.0031979f $X=4.635 $Y=0.56 $X2=0 $Y2=0
cc_458 N_A_561_413#_M1002_g RESET_B 0.00344736f $X=4.635 $Y=1.985 $X2=0 $Y2=0
cc_459 N_A_561_413#_c_674_n RESET_B 0.00709738f $X=4.56 $Y=1.16 $X2=0 $Y2=0
cc_460 N_A_561_413#_c_675_n RESET_B 0.00640764f $X=4.635 $Y=1.16 $X2=0 $Y2=0
cc_461 N_A_561_413#_c_678_n RESET_B 0.0254879f $X=4.145 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_561_413#_M1008_g N_RESET_B_c_759_n 0.020192f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_463 N_A_561_413#_M1008_g N_RESET_B_c_760_n 0.0424171f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_464 N_A_561_413#_c_685_n N_VPWR_c_797_n 0.00489615f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_465 N_A_561_413#_M1002_g N_VPWR_c_798_n 0.00105344f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_466 N_A_561_413#_M1002_g N_VPWR_c_800_n 0.00858459f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_467 N_A_561_413#_c_685_n N_VPWR_c_803_n 0.0343719f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_468 N_A_561_413#_M1001_d N_VPWR_c_795_n 0.00699187f $X=2.805 $Y=2.065 $X2=0
+ $Y2=0
cc_469 N_A_561_413#_M1002_g N_VPWR_c_795_n 0.00477699f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_470 N_A_561_413#_c_685_n N_VPWR_c_795_n 0.0265731f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_471 N_A_561_413#_M1002_g N_VPWR_c_810_n 0.00505556f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_472 N_A_561_413#_M1002_g N_VPWR_c_811_n 5.94208e-19 $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_A_561_413#_c_685_n A_682_413# 0.00145479f $X=3.48 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_474 N_A_561_413#_c_680_n A_682_413# 0.00208506f $X=3.565 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_475 N_A_561_413#_c_682_n N_VGND_c_910_n 0.00209539f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_476 N_A_561_413#_M1008_g N_VGND_c_911_n 0.00234993f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_477 N_A_561_413#_c_674_n N_VGND_c_911_n 0.00160278f $X=4.56 $Y=1.16 $X2=0
+ $Y2=0
cc_478 N_A_561_413#_c_682_n N_VGND_c_911_n 0.010424f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_479 N_A_561_413#_c_678_n N_VGND_c_911_n 0.0113448f $X=4.145 $Y=1.16 $X2=0
+ $Y2=0
cc_480 N_A_561_413#_c_682_n N_VGND_c_914_n 0.0221606f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_481 N_A_561_413#_M1016_d N_VGND_c_916_n 0.00237979f $X=2.865 $Y=0.235 $X2=0
+ $Y2=0
cc_482 N_A_561_413#_M1008_g N_VGND_c_916_n 0.00709954f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_483 N_A_561_413#_c_682_n N_VGND_c_916_n 0.0222941f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_484 N_A_561_413#_M1008_g N_VGND_c_920_n 0.00415469f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_485 N_A_561_413#_M1008_g N_VGND_c_921_n 0.00189265f $X=4.635 $Y=0.56 $X2=0
+ $Y2=0
cc_486 N_A_561_413#_c_682_n A_659_47# 0.00365607f $X=3.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_487 N_A_561_413#_c_676_n A_659_47# 0.00149829f $X=3.415 $Y=1.025 $X2=-0.19
+ $Y2=-0.24
cc_488 N_RESET_B_M1013_g N_VPWR_c_800_n 5.73883e-19 $X=5.055 $Y=1.985 $X2=0
+ $Y2=0
cc_489 N_RESET_B_M1013_g N_VPWR_c_795_n 0.00475773f $X=5.055 $Y=1.985 $X2=0
+ $Y2=0
cc_490 N_RESET_B_M1013_g N_VPWR_c_810_n 0.00505556f $X=5.055 $Y=1.985 $X2=0
+ $Y2=0
cc_491 N_RESET_B_M1013_g N_VPWR_c_811_n 0.0175119f $X=5.055 $Y=1.985 $X2=0 $Y2=0
cc_492 N_RESET_B_c_760_n N_VGND_c_916_n 0.00389423f $X=5.065 $Y=0.995 $X2=0
+ $Y2=0
cc_493 N_RESET_B_c_760_n N_VGND_c_920_n 0.00327422f $X=5.065 $Y=0.995 $X2=0
+ $Y2=0
cc_494 N_RESET_B_c_760_n N_VGND_c_921_n 0.0176784f $X=5.065 $Y=0.995 $X2=0 $Y2=0
cc_495 N_VPWR_c_795_n A_465_369# 0.00373974f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_496 N_VPWR_c_795_n A_682_413# 0.00170472f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_497 N_VPWR_c_795_n N_Q_M1015_d 0.00383158f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_498 N_VPWR_c_804_n Q 0.0169196f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_499 N_VPWR_c_795_n Q 0.00988906f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_500 Q N_VGND_c_915_n 0.00880728f $X=6.15 $Y=0.425 $X2=0 $Y2=0
cc_501 N_Q_M1010_d N_VGND_c_916_n 0.00405593f $X=6.045 $Y=0.235 $X2=0 $Y2=0
cc_502 Q N_VGND_c_916_n 0.00906349f $X=6.15 $Y=0.425 $X2=0 $Y2=0
cc_503 N_VGND_c_916_n A_465_47# 0.0139156f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_504 N_VGND_c_916_n A_659_47# 0.00687059f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_505 N_VGND_c_916_n A_942_47# 0.00323135f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__or2_2.pxi.spice
* Created: Thu Aug 27 14:42:41 2020
* 
x_PM_SKY130_FD_SC_HD__OR2_2%B N_B_M1007_g N_B_M1004_g B B N_B_c_46_n
+ PM_SKY130_FD_SC_HD__OR2_2%B
x_PM_SKY130_FD_SC_HD__OR2_2%A N_A_M1006_g N_A_M1001_g A A N_A_c_73_n
+ PM_SKY130_FD_SC_HD__OR2_2%A
x_PM_SKY130_FD_SC_HD__OR2_2%A_39_297# N_A_39_297#_M1007_d N_A_39_297#_M1004_s
+ N_A_39_297#_c_106_n N_A_39_297#_M1000_g N_A_39_297#_M1002_g
+ N_A_39_297#_c_107_n N_A_39_297#_M1003_g N_A_39_297#_M1005_g
+ N_A_39_297#_c_108_n N_A_39_297#_c_130_n N_A_39_297#_c_114_n
+ N_A_39_297#_c_109_n N_A_39_297#_c_124_n N_A_39_297#_c_110_n
+ PM_SKY130_FD_SC_HD__OR2_2%A_39_297#
x_PM_SKY130_FD_SC_HD__OR2_2%VPWR N_VPWR_M1001_d N_VPWR_M1005_d N_VPWR_c_176_n
+ N_VPWR_c_177_n N_VPWR_c_178_n VPWR N_VPWR_c_179_n N_VPWR_c_180_n
+ N_VPWR_c_181_n N_VPWR_c_175_n PM_SKY130_FD_SC_HD__OR2_2%VPWR
x_PM_SKY130_FD_SC_HD__OR2_2%X N_X_M1000_d N_X_M1002_s N_X_c_204_n X N_X_c_219_n
+ PM_SKY130_FD_SC_HD__OR2_2%X
x_PM_SKY130_FD_SC_HD__OR2_2%VGND N_VGND_M1007_s N_VGND_M1006_d N_VGND_M1003_s
+ N_VGND_c_236_n N_VGND_c_237_n N_VGND_c_238_n N_VGND_c_239_n N_VGND_c_240_n
+ VGND N_VGND_c_241_n N_VGND_c_242_n N_VGND_c_243_n N_VGND_c_244_n
+ PM_SKY130_FD_SC_HD__OR2_2%VGND
cc_1 VNB N_B_M1007_g 0.0331249f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB B 0.0113985f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_B_c_46_n 0.0459535f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_4 VNB N_A_M1006_g 0.0288484f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB A 0.00409615f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_6 VNB N_A_c_73_n 0.0209416f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_7 VNB N_A_39_297#_c_106_n 0.0166586f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.695
cc_8 VNB N_A_39_297#_c_107_n 0.0190315f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_9 VNB N_A_39_297#_c_108_n 0.00421483f $X=-0.19 $Y=-0.24 $X2=0.247 $Y2=1.16
cc_10 VNB N_A_39_297#_c_109_n 5.05956e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_39_297#_c_110_n 0.0355374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_175_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_X_c_204_n 0.00802153f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_14 VNB X 0.020816f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_15 VNB N_VGND_c_236_n 0.0101374f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_16 VNB N_VGND_c_237_n 0.0191673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_238_n 0.00264128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_239_n 0.0106755f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_19 VNB N_VGND_c_240_n 0.0126448f $X=-0.19 $Y=-0.24 $X2=0.247 $Y2=0.85
cc_20 VNB N_VGND_c_241_n 0.0190583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_242_n 0.0121091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_243_n 0.00479031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_244_n 0.142076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VPB N_B_M1004_g 0.0272501f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.695
cc_25 VPB B 0.00176543f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_26 VPB N_B_c_46_n 0.0118142f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_27 VPB N_A_M1001_g 0.0208486f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.695
cc_28 VPB A 0.00300939f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_29 VPB N_A_c_73_n 0.00456039f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_30 VPB N_A_39_297#_M1002_g 0.0212926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_39_297#_M1005_g 0.0229705f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_39_297#_c_108_n 0.00161876f $X=-0.19 $Y=1.305 $X2=0.247 $Y2=1.16
cc_33 VPB N_A_39_297#_c_114_n 0.0157579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_39_297#_c_109_n 9.43842e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_39_297#_c_110_n 0.0047903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_176_n 0.00416524f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_37 VPB N_VPWR_c_177_n 0.0110934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_178_n 0.00416524f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_39 VPB N_VPWR_c_179_n 0.0371475f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_40 VPB N_VPWR_c_180_n 0.0172154f $X=-0.19 $Y=1.305 $X2=0.247 $Y2=1.16
cc_41 VPB N_VPWR_c_181_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_175_n 0.0755826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB X 0.0307062f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_44 N_B_M1007_g N_A_M1006_g 0.0223994f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_45 N_B_M1004_g N_A_M1001_g 0.0319815f $X=0.53 $Y=1.695 $X2=0 $Y2=0
cc_46 N_B_M1007_g A 2.10173e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_47 N_B_c_46_n A 3.15735e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_48 N_B_c_46_n N_A_c_73_n 0.0319815f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_49 N_B_M1007_g N_A_39_297#_c_108_n 0.0121126f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_50 N_B_M1004_g N_A_39_297#_c_108_n 0.00838774f $X=0.53 $Y=1.695 $X2=0 $Y2=0
cc_51 B N_A_39_297#_c_108_n 0.0393703f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_52 N_B_c_46_n N_A_39_297#_c_108_n 0.010132f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_53 N_B_M1004_g N_A_39_297#_c_114_n 0.0170135f $X=0.53 $Y=1.695 $X2=0 $Y2=0
cc_54 B N_A_39_297#_c_114_n 0.0155318f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_55 N_B_c_46_n N_A_39_297#_c_114_n 0.0049962f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_56 N_B_M1007_g N_A_39_297#_c_124_n 0.00397816f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_57 N_B_M1004_g N_VPWR_c_179_n 0.00327927f $X=0.53 $Y=1.695 $X2=0 $Y2=0
cc_58 N_B_M1004_g N_VPWR_c_175_n 0.00417489f $X=0.53 $Y=1.695 $X2=0 $Y2=0
cc_59 N_B_M1007_g N_VGND_c_237_n 0.00448362f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_60 B N_VGND_c_237_n 0.0166603f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_61 N_B_c_46_n N_VGND_c_237_n 0.00179184f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B_M1007_g N_VGND_c_241_n 0.00541359f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_63 N_B_M1007_g N_VGND_c_244_n 0.0104829f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_64 B N_VGND_c_244_n 7.6743e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_A_39_297#_c_106_n 0.0206998f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_66 A N_A_39_297#_c_106_n 0.00497619f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_A_39_297#_M1002_g 0.0200395f $X=0.89 $Y=1.695 $X2=0 $Y2=0
cc_68 N_A_M1006_g N_A_39_297#_c_108_n 0.0105175f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_69 A N_A_39_297#_c_108_n 0.0429397f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_70 N_A_M1001_g N_A_39_297#_c_130_n 0.0159541f $X=0.89 $Y=1.695 $X2=0 $Y2=0
cc_71 A N_A_39_297#_c_130_n 0.0296821f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_72 N_A_c_73_n N_A_39_297#_c_130_n 7.21566e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1001_g N_A_39_297#_c_114_n 9.34042e-19 $X=0.89 $Y=1.695 $X2=0 $Y2=0
cc_74 N_A_M1001_g N_A_39_297#_c_109_n 8.0108e-19 $X=0.89 $Y=1.695 $X2=0 $Y2=0
cc_75 A N_A_39_297#_c_109_n 0.0253715f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_c_73_n N_A_39_297#_c_109_n 2.49936e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_73_n N_A_39_297#_c_110_n 0.0183045f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_VPWR_c_176_n 0.00442731f $X=0.89 $Y=1.695 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_VPWR_c_179_n 0.00327927f $X=0.89 $Y=1.695 $X2=0 $Y2=0
cc_80 N_A_M1001_g N_VPWR_c_175_n 0.00417489f $X=0.89 $Y=1.695 $X2=0 $Y2=0
cc_81 A X 0.0048433f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_82 A N_VGND_M1006_d 0.00266597f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_VGND_c_238_n 0.00644978f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_84 A N_VGND_c_238_n 0.0195582f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_85 N_A_c_73_n N_VGND_c_238_n 2.29546e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_M1006_g N_VGND_c_241_n 0.00585385f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_M1006_g N_VGND_c_244_n 0.00787418f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_88 A N_VGND_c_244_n 0.00716308f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_89 N_A_39_297#_c_130_n A_121_297# 0.00473129f $X=1.445 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_90 N_A_39_297#_c_114_n A_121_297# 0.00144354f $X=0.695 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_39_297#_c_130_n N_VPWR_M1001_d 0.00715465f $X=1.445 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_39_297#_M1002_g N_VPWR_c_176_n 0.00316354f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_93 N_A_39_297#_c_130_n N_VPWR_c_176_n 0.0131801f $X=1.445 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_39_297#_M1005_g N_VPWR_c_178_n 0.00316354f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_95 N_A_39_297#_M1002_g N_VPWR_c_180_n 0.00540367f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_96 N_A_39_297#_M1005_g N_VPWR_c_180_n 0.00421248f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_97 N_A_39_297#_M1002_g N_VPWR_c_175_n 0.0107815f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_98 N_A_39_297#_M1005_g N_VPWR_c_175_n 0.00667935f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_99 N_A_39_297#_c_130_n N_X_M1002_s 0.00242555f $X=1.445 $Y=1.58 $X2=0 $Y2=0
cc_100 N_A_39_297#_c_107_n N_X_c_204_n 0.0116408f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_39_297#_c_109_n N_X_c_204_n 0.00764635f $X=1.53 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_39_297#_c_110_n N_X_c_204_n 0.00191734f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_39_297#_c_106_n X 5.77812e-19 $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_39_297#_M1002_g X 0.00354274f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_39_297#_c_107_n X 0.00721277f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_39_297#_M1005_g X 0.0315154f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_39_297#_c_130_n X 0.0235405f $X=1.445 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_39_297#_c_109_n X 0.0370288f $X=1.53 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_39_297#_c_110_n X 0.0158158f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_39_297#_M1002_g N_X_c_219_n 0.00535723f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_39_297#_M1005_g N_X_c_219_n 0.0109535f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_39_297#_c_106_n N_VGND_c_238_n 0.00997997f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_113 N_A_39_297#_c_107_n N_VGND_c_238_n 8.96527e-19 $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_114 N_A_39_297#_c_106_n N_VGND_c_240_n 8.65114e-19 $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_A_39_297#_c_107_n N_VGND_c_240_n 0.00885796f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_116 N_A_39_297#_c_124_n N_VGND_c_241_n 0.0163547f $X=0.68 $Y=0.43 $X2=0 $Y2=0
cc_117 N_A_39_297#_c_106_n N_VGND_c_242_n 0.0046653f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_118 N_A_39_297#_c_107_n N_VGND_c_242_n 0.00341574f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_119 N_A_39_297#_M1007_d N_VGND_c_244_n 0.00249917f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_120 N_A_39_297#_c_106_n N_VGND_c_244_n 0.00796766f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_121 N_A_39_297#_c_107_n N_VGND_c_244_n 0.00402423f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_A_39_297#_c_124_n N_VGND_c_244_n 0.0108145f $X=0.68 $Y=0.43 $X2=0 $Y2=0
cc_123 N_VPWR_c_175_n N_X_M1002_s 0.00215201f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_124 N_VPWR_M1005_d X 0.00593212f $X=1.89 $Y=1.485 $X2=0 $Y2=0
cc_125 N_VPWR_c_177_n X 0.00159763f $X=2.025 $Y=2.635 $X2=0 $Y2=0
cc_126 N_VPWR_c_178_n X 0.0126475f $X=2.025 $Y=2.34 $X2=0 $Y2=0
cc_127 N_VPWR_c_180_n X 0.00205878f $X=1.94 $Y=2.72 $X2=0 $Y2=0
cc_128 N_VPWR_c_175_n X 0.00741106f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_129 N_VPWR_c_180_n N_X_c_219_n 0.0184921f $X=1.94 $Y=2.72 $X2=0 $Y2=0
cc_130 N_VPWR_c_175_n N_X_c_219_n 0.012098f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_131 N_X_c_204_n N_VGND_M1003_s 0.00292162f $X=1.605 $Y=0.565 $X2=0 $Y2=0
cc_132 X N_VGND_M1003_s 2.61253e-19 $X=1.99 $Y=1.785 $X2=0 $Y2=0
cc_133 N_X_c_204_n N_VGND_c_239_n 4.88604e-19 $X=1.605 $Y=0.565 $X2=0 $Y2=0
cc_134 N_X_c_204_n N_VGND_c_240_n 0.0229176f $X=1.605 $Y=0.565 $X2=0 $Y2=0
cc_135 N_X_c_204_n N_VGND_c_242_n 0.00848422f $X=1.605 $Y=0.565 $X2=0 $Y2=0
cc_136 N_X_M1000_d N_VGND_c_244_n 0.0042048f $X=1.47 $Y=0.235 $X2=0 $Y2=0
cc_137 N_X_c_204_n N_VGND_c_244_n 0.0126564f $X=1.605 $Y=0.565 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__clkinv_2.spice.pex
* Created: Thu Aug 27 14:12:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKINV_2%A 3 7 11 13 15 19 21 22 23
r49 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1
+ $Y=1.16 $X2=1 $Y2=1.16
r50 32 34 10.3656 $w=2.79e-07 $l=6e-08 $layer=POLY_cond $X=0.94 $Y=1.16 $X2=1
+ $Y2=1.16
r51 28 30 30.233 $w=2.79e-07 $l=1.75e-07 $layer=POLY_cond $X=0.32 $Y=1.16
+ $X2=0.495 $Y2=1.16
r52 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.16 $X2=0.32 $Y2=1.16
r53 23 35 7.68295 $w=2.23e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=1.177 $X2=1
+ $Y2=1.177
r54 22 35 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=0.69 $Y=1.177 $X2=1
+ $Y2=1.177
r55 22 29 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.69 $Y=1.177
+ $X2=0.32 $Y2=1.177
r56 21 29 4.60977 $w=2.23e-07 $l=9e-08 $layer=LI1_cond $X=0.23 $Y=1.177 $X2=0.32
+ $Y2=1.177
r57 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.37 $Y=1.025
+ $X2=1.37 $Y2=0.445
r58 13 17 2.5914 $w=2.79e-07 $l=1.5e-08 $layer=POLY_cond $X=1.355 $Y=1.16
+ $X2=1.37 $Y2=1.16
r59 13 34 61.3298 $w=2.79e-07 $l=3.55e-07 $layer=POLY_cond $X=1.355 $Y=1.16
+ $X2=1 $Y2=1.16
r60 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.355 $Y=1.295
+ $X2=1.355 $Y2=1.985
r61 9 32 17.2686 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.94 $Y=1.015
+ $X2=0.94 $Y2=1.16
r62 9 11 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.94 $Y=1.015
+ $X2=0.94 $Y2=0.445
r63 5 32 2.5914 $w=2.79e-07 $l=1.5e-08 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.94 $Y2=1.16
r64 5 30 74.2867 $w=2.79e-07 $l=4.3e-07 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.495 $Y2=1.16
r65 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.925 $Y=1.295
+ $X2=0.925 $Y2=1.985
r66 1 30 17.2686 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.495 $Y=1.305
+ $X2=0.495 $Y2=1.16
r67 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.495 $Y=1.305
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_2%Y 1 2 3 12 14 15 18 22 24 25 26 28 29 30 31
+ 37 38
c50 37 0 8.53357e-20 $X=1.615 $Y=0.895
r51 31 38 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=1.545
+ $X2=1.615 $Y2=1.46
r52 31 38 0.329269 $w=2.78e-07 $l=8e-09 $layer=LI1_cond $X=1.615 $Y=1.452
+ $X2=1.615 $Y2=1.46
r53 30 31 10.7836 $w=2.78e-07 $l=2.62e-07 $layer=LI1_cond $X=1.615 $Y=1.19
+ $X2=1.615 $Y2=1.452
r54 29 37 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.81
+ $X2=1.615 $Y2=0.895
r55 29 30 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=0.915
+ $X2=1.615 $Y2=1.19
r56 29 37 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=1.615 $Y=0.915
+ $X2=1.615 $Y2=0.895
r57 27 28 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.27 $Y=1.545
+ $X2=1.14 $Y2=1.545
r58 26 31 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.475 $Y=1.545
+ $X2=1.615 $Y2=1.545
r59 26 27 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.475 $Y=1.545
+ $X2=1.27 $Y2=1.545
r60 24 29 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=1.615 $Y2=0.81
r61 24 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.475 $Y=0.81
+ $X2=1.25 $Y2=0.81
r62 20 25 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.137 $Y=0.725
+ $X2=1.25 $Y2=0.81
r63 20 22 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=1.137 $Y=0.725
+ $X2=1.137 $Y2=0.445
r64 16 28 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.63
+ $X2=1.14 $Y2=1.545
r65 16 18 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=1.14 $Y=1.63 $X2=1.14
+ $Y2=1.83
r66 14 28 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.01 $Y=1.545
+ $X2=1.14 $Y2=1.545
r67 14 15 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.01 $Y=1.545 $X2=0.41
+ $Y2=1.545
r68 10 15 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.282 $Y=1.63
+ $X2=0.41 $Y2=1.545
r69 10 12 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=0.282 $Y=1.63
+ $X2=0.282 $Y2=1.83
r70 3 18 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.485 $X2=1.14 $Y2=1.83
r71 2 12 300 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=1.83
r72 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.155 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_2%VPWR 1 2 9 11 13 15 17 22 28 32
r27 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r29 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r32 23 28 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.84 $Y=2.72 $X2=0.71
+ $Y2=2.72
r33 23 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.84 $Y=2.72
+ $X2=1.15 $Y2=2.72
r34 22 31 4.00962 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.44 $Y=2.72 $X2=1.64
+ $Y2=2.72
r35 22 25 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 17 28 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.58 $Y=2.72 $X2=0.71
+ $Y2=2.72
r37 17 19 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.58 $Y=2.72
+ $X2=0.23 $Y2=2.72
r38 15 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r39 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r40 11 31 3.1676 $w=2.55e-07 $l=1.15888e-07 $layer=LI1_cond $X=1.567 $Y=2.635
+ $X2=1.64 $Y2=2.72
r41 11 13 30.2799 $w=2.53e-07 $l=6.7e-07 $layer=LI1_cond $X=1.567 $Y=2.635
+ $X2=1.567 $Y2=1.965
r42 7 28 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.72
r43 7 9 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=0.71 $Y=2.635 $X2=0.71
+ $Y2=1.965
r44 2 13 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=1.43
+ $Y=1.485 $X2=1.57 $Y2=1.965
r45 1 9 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.485 $X2=0.71 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_2%VGND 1 2 9 11 13 15 17 22 28 32
c24 11 0 8.53357e-20 $X=1.585 $Y=0.085
r25 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r26 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r27 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r28 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r29 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r30 23 28 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.707
+ $Y2=0
r31 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.15
+ $Y2=0
r32 22 31 4.79676 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.63
+ $Y2=0
r33 22 25 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.15
+ $Y2=0
r34 17 28 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.707
+ $Y2=0
r35 17 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.23
+ $Y2=0
r36 15 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r37 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r38 11 31 2.96942 $w=3.3e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.63 $Y2=0
r39 11 13 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.585 $Y2=0.39
r40 7 28 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0
r41 7 9 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0.445
r42 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.39
r43 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.725 $Y2=0.445
.ends


* File: sky130_fd_sc_hd__a311oi_2.pxi.spice
* Created: Thu Aug 27 14:04:21 2020
* 
x_PM_SKY130_FD_SC_HD__A311OI_2%A3 N_A3_c_71_n N_A3_M1009_g N_A3_M1006_g
+ N_A3_c_72_n N_A3_M1019_g N_A3_M1017_g A3 A3 N_A3_c_73_n
+ PM_SKY130_FD_SC_HD__A311OI_2%A3
x_PM_SKY130_FD_SC_HD__A311OI_2%A2 N_A2_c_107_n N_A2_M1015_g N_A2_M1002_g
+ N_A2_c_108_n N_A2_M1016_g N_A2_M1018_g A2 A2 N_A2_c_109_n N_A2_c_110_n
+ PM_SKY130_FD_SC_HD__A311OI_2%A2
x_PM_SKY130_FD_SC_HD__A311OI_2%A1 N_A1_M1000_g N_A1_M1003_g N_A1_c_153_n
+ N_A1_M1010_g N_A1_c_154_n N_A1_M1012_g A1 A1 A1 N_A1_c_156_n
+ PM_SKY130_FD_SC_HD__A311OI_2%A1
x_PM_SKY130_FD_SC_HD__A311OI_2%B1 N_B1_c_201_n N_B1_M1007_g N_B1_M1001_g
+ N_B1_c_202_n N_B1_M1011_g N_B1_M1005_g B1 B1 N_B1_c_204_n
+ PM_SKY130_FD_SC_HD__A311OI_2%B1
x_PM_SKY130_FD_SC_HD__A311OI_2%C1 N_C1_c_251_n N_C1_M1008_g N_C1_M1004_g
+ N_C1_c_252_n N_C1_M1013_g N_C1_M1014_g C1 C1 C1 N_C1_c_253_n N_C1_c_278_p
+ N_C1_c_254_n PM_SKY130_FD_SC_HD__A311OI_2%C1
x_PM_SKY130_FD_SC_HD__A311OI_2%VPWR N_VPWR_M1006_d N_VPWR_M1017_d N_VPWR_M1018_s
+ N_VPWR_M1003_d N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n
+ N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n
+ VPWR N_VPWR_c_308_n N_VPWR_c_309_n N_VPWR_c_298_n N_VPWR_c_311_n
+ PM_SKY130_FD_SC_HD__A311OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A311OI_2%A_109_297# N_A_109_297#_M1006_s
+ N_A_109_297#_M1002_d N_A_109_297#_M1000_s N_A_109_297#_M1001_s
+ N_A_109_297#_c_404_n N_A_109_297#_c_376_n N_A_109_297#_c_377_n
+ N_A_109_297#_c_381_n N_A_109_297#_c_382_n N_A_109_297#_c_413_n
+ N_A_109_297#_c_375_n N_A_109_297#_c_384_n N_A_109_297#_c_391_n
+ N_A_109_297#_c_395_n PM_SKY130_FD_SC_HD__A311OI_2%A_109_297#
x_PM_SKY130_FD_SC_HD__A311OI_2%A_641_297# N_A_641_297#_M1001_d
+ N_A_641_297#_M1005_d N_A_641_297#_M1014_s N_A_641_297#_c_424_n
+ N_A_641_297#_c_427_n N_A_641_297#_c_431_n N_A_641_297#_c_433_n
+ N_A_641_297#_c_428_n PM_SKY130_FD_SC_HD__A311OI_2%A_641_297#
x_PM_SKY130_FD_SC_HD__A311OI_2%Y N_Y_M1010_d N_Y_M1012_d N_Y_M1011_s N_Y_M1013_d
+ N_Y_M1004_d N_Y_c_460_n N_Y_c_467_n N_Y_c_469_n N_Y_c_480_n N_Y_c_481_n
+ N_Y_c_486_n N_Y_c_521_p N_Y_c_473_n N_Y_c_474_n Y Y Y Y N_Y_c_476_n Y
+ N_Y_c_495_n Y PM_SKY130_FD_SC_HD__A311OI_2%Y
x_PM_SKY130_FD_SC_HD__A311OI_2%A_27_47# N_A_27_47#_M1009_d N_A_27_47#_M1019_d
+ N_A_27_47#_M1016_d N_A_27_47#_c_555_p N_A_27_47#_c_537_n N_A_27_47#_c_541_n
+ N_A_27_47#_c_553_p N_A_27_47#_c_536_n N_A_27_47#_c_547_n
+ PM_SKY130_FD_SC_HD__A311OI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__A311OI_2%VGND N_VGND_M1009_s N_VGND_M1007_d N_VGND_M1008_s
+ N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n
+ VGND N_VGND_c_572_n N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n
+ N_VGND_c_576_n N_VGND_c_577_n PM_SKY130_FD_SC_HD__A311OI_2%VGND
x_PM_SKY130_FD_SC_HD__A311OI_2%A_277_47# N_A_277_47#_M1015_s N_A_277_47#_M1010_s
+ N_A_277_47#_c_649_n PM_SKY130_FD_SC_HD__A311OI_2%A_277_47#
cc_1 VNB N_A3_c_71_n 0.0217541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A3_c_72_n 0.0160222f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A3_c_73_n 0.0620421f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_4 VNB N_A2_c_107_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_A2_c_108_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_6 VNB N_A2_c_109_n 0.00377146f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_7 VNB N_A2_c_110_n 0.0330528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_c_153_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_9 VNB N_A1_c_154_n 0.0165278f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_10 VNB A1 0.0029391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_156_n 0.0607174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_201_n 0.0162993f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_B1_c_202_n 0.0178799f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_14 VNB B1 0.00508059f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_15 VNB N_B1_c_204_n 0.0338659f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_16 VNB N_C1_c_251_n 0.0178426f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_17 VNB N_C1_c_252_n 0.0217503f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_18 VNB N_C1_c_253_n 0.0578954f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_19 VNB N_C1_c_254_n 0.00887859f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_20 VNB N_VPWR_c_298_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_460_n 0.00208149f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_22 VNB Y 0.00938422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_536_n 0.00220864f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_24 VNB N_VGND_c_567_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_25 VNB N_VGND_c_568_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_26 VNB N_VGND_c_569_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_570_n 0.0644097f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_28 VNB N_VGND_c_571_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_29 VNB N_VGND_c_572_n 0.01517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_573_n 0.0179279f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_574_n 0.01517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_575_n 0.2816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_576_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_577_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_277_47#_c_649_n 0.00653612f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_36 VPB N_A3_M1006_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A3_M1017_g 0.0185651f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_38 VPB N_A3_c_73_n 0.0138306f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_39 VPB N_A2_M1002_g 0.018686f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_40 VPB N_A2_M1018_g 0.0189137f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_41 VPB N_A2_c_109_n 0.00205765f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_42 VPB N_A2_c_110_n 0.00522588f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A1_M1000_g 0.0187928f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_44 VPB N_A1_M1003_g 0.02509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB A1 0.00124565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A1_c_156_n 0.018442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_B1_M1001_g 0.0259823f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_48 VPB N_B1_M1005_g 0.0210669f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_49 VPB B1 0.0012492f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_50 VPB N_B1_c_204_n 0.00549678f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_51 VPB N_C1_M1004_g 0.0210057f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_52 VPB N_C1_M1014_g 0.021871f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_53 VPB C1 0.0142061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_C1_c_253_n 0.0136341f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_55 VPB N_VPWR_c_299_n 0.0100141f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_56 VPB N_VPWR_c_300_n 0.0423786f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_57 VPB N_VPWR_c_301_n 3.17494e-19 $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_58 VPB N_VPWR_c_302_n 3.03604e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_303_n 0.0102455f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_60 VPB N_VPWR_c_304_n 0.0128097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_305_n 0.00463502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_306_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_307_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_308_n 0.0160841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_309_n 0.0636651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_298_n 0.0529832f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_311_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_109_297#_c_375_n 0.0119483f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_69 VPB N_A_641_297#_c_424_n 0.00292106f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_70 VPB Y 0.00432102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 N_A3_c_72_n N_A2_c_107_n 0.023564f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_72 N_A3_M1017_g N_A2_M1002_g 0.023564f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 A3 N_A2_c_109_n 0.0215092f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A3_c_73_n N_A2_c_109_n 0.00347698f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_75 A3 N_A2_c_110_n 2.50845e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A3_c_73_n N_A2_c_110_n 0.023564f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A3_M1006_g N_VPWR_c_300_n 0.00311793f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_78 A3 N_VPWR_c_300_n 0.0169901f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A3_c_73_n N_VPWR_c_300_n 0.00596154f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A3_M1006_g N_VPWR_c_301_n 6.41958e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A3_M1017_g N_VPWR_c_301_n 0.0103454f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A3_M1006_g N_VPWR_c_308_n 0.00585385f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A3_M1017_g N_VPWR_c_308_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A3_M1006_g N_VPWR_c_298_n 0.0114913f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A3_M1017_g N_VPWR_c_298_n 0.00789179f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A3_M1017_g N_A_109_297#_c_376_n 0.0181226f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_87 A3 N_A_109_297#_c_377_n 0.00996364f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_88 N_A3_c_73_n N_A_109_297#_c_377_n 0.00200701f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A3_c_71_n N_A_27_47#_c_537_n 0.0127525f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A3_c_72_n N_A_27_47#_c_537_n 0.0160373f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_91 A3 N_A_27_47#_c_537_n 0.0278215f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A3_c_73_n N_A_27_47#_c_537_n 0.00201785f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_93 A3 N_A_27_47#_c_541_n 0.0135367f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_94 N_A3_c_73_n N_A_27_47#_c_541_n 0.00391331f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A3_c_71_n N_VGND_c_567_n 0.00837154f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A3_c_72_n N_VGND_c_567_n 0.00787405f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A3_c_72_n N_VGND_c_570_n 0.00341689f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A3_c_71_n N_VGND_c_572_n 0.00341689f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A3_c_71_n N_VGND_c_575_n 0.00493711f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A3_c_72_n N_VGND_c_575_n 0.00401011f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A2_M1018_g N_A1_M1000_g 0.0275979f $X=1.74 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A2_c_109_n A1 0.0263518f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A2_c_110_n A1 0.0026202f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A2_c_109_n N_A1_c_156_n 3.20936e-19 $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A2_c_110_n N_A1_c_156_n 0.016449f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A2_M1002_g N_VPWR_c_301_n 0.0101944f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A2_M1018_g N_VPWR_c_301_n 6.04015e-19 $X=1.74 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A2_M1002_g N_VPWR_c_302_n 6.13705e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A2_M1018_g N_VPWR_c_302_n 0.0104116f $X=1.74 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A2_M1002_g N_VPWR_c_304_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A2_M1018_g N_VPWR_c_304_n 0.0046653f $X=1.74 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A2_M1002_g N_VPWR_c_298_n 0.00791817f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A2_M1018_g N_VPWR_c_298_n 0.00791817f $X=1.74 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A2_M1002_g N_A_109_297#_c_376_n 0.0145497f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A2_c_109_n N_A_109_297#_c_376_n 0.0183405f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A2_M1018_g N_A_109_297#_c_381_n 0.00498027f $X=1.74 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A2_M1018_g N_A_109_297#_c_382_n 0.0149234f $X=1.74 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A2_c_109_n N_A_109_297#_c_382_n 0.00900104f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A2_c_109_n N_A_109_297#_c_384_n 0.0101997f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A2_c_110_n N_A_109_297#_c_384_n 0.00226621f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A2_c_107_n N_A_27_47#_c_536_n 0.011504f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A2_c_108_n N_A_27_47#_c_536_n 0.00841904f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A2_c_109_n N_A_27_47#_c_536_n 0.0392679f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A2_c_110_n N_A_27_47#_c_536_n 0.00201785f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A2_c_109_n N_A_27_47#_c_547_n 0.010813f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A2_c_107_n N_VGND_c_567_n 0.00116167f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A2_c_107_n N_VGND_c_570_n 0.00416042f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A2_c_108_n N_VGND_c_570_n 0.00368123f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_107_n N_VGND_c_575_n 0.00574236f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A2_c_108_n N_VGND_c_575_n 0.00662341f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A2_c_107_n N_A_277_47#_c_649_n 0.00248308f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A2_c_108_n N_A_277_47#_c_649_n 0.0101206f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A1_c_154_n N_B1_c_201_n 0.0224159f $X=3.09 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_134 A1 B1 0.0200511f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_135 N_A1_c_156_n B1 0.00263292f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_136 A1 N_B1_c_204_n 3.70222e-19 $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A1_c_156_n N_B1_c_204_n 0.0177772f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A1_M1000_g N_VPWR_c_302_n 0.010251f $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A1_M1003_g N_VPWR_c_302_n 6.10071e-19 $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A1_M1000_g N_VPWR_c_303_n 6.0901e-19 $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A1_M1003_g N_VPWR_c_303_n 0.0112954f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_VPWR_c_306_n 0.0046653f $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A1_M1003_g N_VPWR_c_306_n 0.0046653f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A1_M1000_g N_VPWR_c_298_n 0.00789179f $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1003_g N_VPWR_c_298_n 0.00789179f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1000_g N_A_109_297#_c_382_n 0.0146058f $X=2.18 $Y=1.985 $X2=0 $Y2=0
cc_147 A1 N_A_109_297#_c_382_n 0.0139037f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A1_M1003_g N_A_109_297#_c_375_n 0.0166344f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_149 A1 N_A_109_297#_c_375_n 0.0321066f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A1_c_156_n N_A_109_297#_c_375_n 0.0123611f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_151 A1 N_A_109_297#_c_391_n 0.00996364f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A1_c_156_n N_A_109_297#_c_391_n 0.00200701f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A1_c_153_n N_Y_c_460_n 0.00841904f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_c_154_n N_Y_c_460_n 0.0130837f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_155 A1 N_Y_c_460_n 0.0537496f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_c_156_n N_Y_c_460_n 0.00944635f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_c_154_n N_Y_c_467_n 0.00513804f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_158 A1 N_A_27_47#_c_536_n 0.00823827f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A1_c_154_n N_VGND_c_568_n 0.00111602f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A1_c_153_n N_VGND_c_570_n 0.00368123f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A1_c_154_n N_VGND_c_570_n 0.00416042f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A1_c_153_n N_VGND_c_575_n 0.00662341f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_154_n N_VGND_c_575_n 0.00581458f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A1_c_153_n N_A_277_47#_c_649_n 0.0101206f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_154_n N_A_277_47#_c_649_n 0.00256936f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_166 A1 N_A_277_47#_c_649_n 0.00615361f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A1_c_156_n N_A_277_47#_c_649_n 0.004081f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B1_c_202_n N_C1_c_251_n 0.0132267f $X=3.96 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_169 N_B1_M1005_g N_C1_M1004_g 0.0132267f $X=3.96 $Y=1.985 $X2=0 $Y2=0
cc_170 N_B1_c_204_n N_C1_c_253_n 0.0132267f $X=3.96 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B1_M1001_g N_VPWR_c_303_n 0.0089414f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_172 N_B1_M1001_g N_VPWR_c_309_n 0.00366111f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B1_M1005_g N_VPWR_c_309_n 0.00366111f $X=3.96 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B1_M1001_g N_VPWR_c_298_n 0.00656615f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_175 N_B1_M1005_g N_VPWR_c_298_n 0.00582333f $X=3.96 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B1_M1001_g N_A_109_297#_c_375_n 0.0109097f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_177 B1 N_A_109_297#_c_375_n 0.00864271f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_178 N_B1_M1001_g N_A_109_297#_c_395_n 0.0124037f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_179 N_B1_M1005_g N_A_109_297#_c_395_n 0.00970367f $X=3.96 $Y=1.985 $X2=0
+ $Y2=0
cc_180 B1 N_A_109_297#_c_395_n 0.0158881f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_181 N_B1_c_204_n N_A_109_297#_c_395_n 0.0019817f $X=3.96 $Y=1.16 $X2=0 $Y2=0
cc_182 N_B1_M1001_g N_A_641_297#_c_424_n 0.00922647f $X=3.54 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_B1_M1005_g N_A_641_297#_c_424_n 0.0146424f $X=3.96 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_M1005_g N_A_641_297#_c_427_n 0.00669554f $X=3.96 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_B1_M1005_g N_A_641_297#_c_428_n 0.00117077f $X=3.96 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_B1_c_201_n N_Y_c_467_n 0.00448007f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B1_c_201_n N_Y_c_469_n 0.0116758f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_202_n N_Y_c_469_n 0.0126169f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_189 B1 N_Y_c_469_n 0.0403452f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_190 N_B1_c_204_n N_Y_c_469_n 0.00201785f $X=3.96 $Y=1.16 $X2=0 $Y2=0
cc_191 B1 N_Y_c_473_n 8.56474e-19 $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_192 N_B1_M1005_g N_Y_c_474_n 2.89812e-19 $X=3.96 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B1_M1005_g Y 7.53471e-19 $X=3.96 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B1_M1005_g N_Y_c_476_n 0.00289868f $X=3.96 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_c_202_n Y 0.00382311f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_196 B1 Y 0.024605f $X=3.87 $Y=1.105 $X2=0 $Y2=0
cc_197 N_B1_c_204_n Y 0.00537446f $X=3.96 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B1_c_201_n N_VGND_c_568_n 0.00793987f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_c_202_n N_VGND_c_568_n 0.00799974f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B1_c_202_n N_VGND_c_569_n 8.50269e-19 $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B1_c_201_n N_VGND_c_570_n 0.00341689f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_202_n N_VGND_c_573_n 0.00341689f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B1_c_201_n N_VGND_c_575_n 0.00408232f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B1_c_202_n N_VGND_c_575_n 0.004507f $X=3.96 $Y=0.995 $X2=0 $Y2=0
cc_205 N_C1_M1004_g N_VPWR_c_309_n 0.00366111f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_206 N_C1_M1014_g N_VPWR_c_309_n 0.00366111f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_207 N_C1_M1004_g N_VPWR_c_298_n 0.00582333f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_208 N_C1_M1014_g N_VPWR_c_298_n 0.00619429f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_209 N_C1_M1004_g N_A_109_297#_c_395_n 0.00113094f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_210 C1 N_A_641_297#_M1014_s 0.0051341f $X=5.2 $Y=1.445 $X2=0 $Y2=0
cc_211 N_C1_M1004_g N_A_641_297#_c_427_n 0.00637525f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_C1_M1004_g N_A_641_297#_c_431_n 0.0122673f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_213 N_C1_M1014_g N_A_641_297#_c_431_n 0.0115247f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_214 C1 N_A_641_297#_c_433_n 0.0143639f $X=5.2 $Y=1.445 $X2=0 $Y2=0
cc_215 N_C1_c_253_n N_A_641_297#_c_433_n 6.58607e-19 $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_216 N_C1_M1004_g N_A_641_297#_c_428_n 0.00111203f $X=4.63 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_C1_c_251_n N_Y_c_480_n 0.0054658f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_218 N_C1_c_251_n N_Y_c_481_n 0.017154f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_219 N_C1_c_252_n N_Y_c_481_n 0.0132219f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_220 N_C1_c_253_n N_Y_c_481_n 0.00601443f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_221 N_C1_c_278_p N_Y_c_481_n 0.0195031f $X=5.175 $Y=1.185 $X2=0 $Y2=0
cc_222 N_C1_c_254_n N_Y_c_481_n 0.010476f $X=5.292 $Y=1.295 $X2=0 $Y2=0
cc_223 N_C1_M1004_g N_Y_c_486_n 0.0114962f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_224 N_C1_M1004_g N_Y_c_474_n 0.00447346f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_225 N_C1_M1014_g N_Y_c_474_n 0.00737576f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_226 N_C1_c_253_n N_Y_c_474_n 0.00210713f $X=5.05 $Y=1.16 $X2=0 $Y2=0
cc_227 N_C1_c_278_p N_Y_c_474_n 0.014536f $X=5.175 $Y=1.185 $X2=0 $Y2=0
cc_228 N_C1_M1004_g Y 0.00391878f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_229 N_C1_M1014_g Y 0.00331573f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_230 N_C1_c_251_n Y 0.0158151f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_231 N_C1_c_278_p Y 0.0130519f $X=5.175 $Y=1.185 $X2=0 $Y2=0
cc_232 N_C1_M1004_g N_Y_c_495_n 0.00284346f $X=4.63 $Y=1.985 $X2=0 $Y2=0
cc_233 N_C1_M1014_g N_Y_c_495_n 0.00245403f $X=5.05 $Y=1.985 $X2=0 $Y2=0
cc_234 N_C1_c_251_n N_VGND_c_568_n 8.5189e-19 $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_235 N_C1_c_251_n N_VGND_c_569_n 0.00922541f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_236 N_C1_c_252_n N_VGND_c_569_n 0.00837154f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_237 N_C1_c_251_n N_VGND_c_573_n 0.00341689f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_238 N_C1_c_252_n N_VGND_c_574_n 0.00341689f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_239 N_C1_c_251_n N_VGND_c_575_n 0.00457046f $X=4.63 $Y=0.995 $X2=0 $Y2=0
cc_240 N_C1_c_252_n N_VGND_c_575_n 0.00493711f $X=5.05 $Y=0.995 $X2=0 $Y2=0
cc_241 N_VPWR_c_298_n N_A_109_297#_M1006_s 0.00562358f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_242 N_VPWR_c_298_n N_A_109_297#_M1002_d 0.00605104f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_298_n N_A_109_297#_M1000_s 0.00562358f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_298_n N_A_109_297#_M1001_s 0.00219239f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_308_n N_A_109_297#_c_404_n 0.0113958f $X=0.935 $Y=2.72 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_298_n N_A_109_297#_c_404_n 0.00646998f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_247 N_VPWR_M1017_d N_A_109_297#_c_376_n 0.00447418f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_301_n N_A_109_297#_c_376_n 0.0170259f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_249 N_VPWR_c_302_n N_A_109_297#_c_381_n 0.0390324f $X=1.95 $Y=2 $X2=0 $Y2=0
cc_250 N_VPWR_c_304_n N_A_109_297#_c_381_n 0.0116048f $X=1.785 $Y=2.72 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_298_n N_A_109_297#_c_381_n 0.00646998f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_252 N_VPWR_M1018_s N_A_109_297#_c_382_n 0.00736233f $X=1.815 $Y=1.485 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_302_n N_A_109_297#_c_382_n 0.018653f $X=1.95 $Y=2 $X2=0 $Y2=0
cc_254 N_VPWR_c_306_n N_A_109_297#_c_413_n 0.0113958f $X=2.645 $Y=2.72 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_298_n N_A_109_297#_c_413_n 0.00646998f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_256 N_VPWR_M1003_d N_A_109_297#_c_375_n 0.00494461f $X=2.675 $Y=1.485 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_303_n N_A_109_297#_c_375_n 0.0219767f $X=2.81 $Y=2 $X2=0 $Y2=0
cc_258 N_VPWR_c_303_n N_A_109_297#_c_395_n 0.00511749f $X=2.81 $Y=2 $X2=0 $Y2=0
cc_259 N_VPWR_c_298_n N_A_641_297#_M1001_d 0.00211652f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_260 N_VPWR_c_298_n N_A_641_297#_M1005_d 0.00421956f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_298_n N_A_641_297#_M1014_s 0.00348623f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_303_n N_A_641_297#_c_424_n 0.0148612f $X=2.81 $Y=2 $X2=0 $Y2=0
cc_263 N_VPWR_c_309_n N_A_641_297#_c_424_n 0.0432961f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_298_n N_A_641_297#_c_424_n 0.0336003f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_309_n N_A_641_297#_c_431_n 0.043459f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_266 N_VPWR_c_298_n N_A_641_297#_c_431_n 0.0317771f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_309_n N_A_641_297#_c_428_n 0.0228518f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_298_n N_A_641_297#_c_428_n 0.0126396f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_298_n N_Y_M1004_d 0.00219239f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_270 N_A_109_297#_c_375_n N_A_641_297#_M1001_d 0.0118636f $X=3.585 $Y=1.66
+ $X2=-0.19 $Y2=1.305
cc_271 N_A_109_297#_M1001_s N_A_641_297#_c_424_n 0.00325424f $X=3.615 $Y=1.485
+ $X2=0 $Y2=0
cc_272 N_A_109_297#_c_375_n N_A_641_297#_c_424_n 0.0119326f $X=3.585 $Y=1.66
+ $X2=0 $Y2=0
cc_273 N_A_109_297#_c_395_n N_A_641_297#_c_424_n 0.0157268f $X=3.75 $Y=1.66
+ $X2=0 $Y2=0
cc_274 N_A_109_297#_c_395_n N_A_641_297#_c_427_n 0.0118727f $X=3.75 $Y=1.66
+ $X2=0 $Y2=0
cc_275 N_A_109_297#_c_395_n N_Y_c_476_n 0.00530715f $X=3.75 $Y=1.66 $X2=0 $Y2=0
cc_276 N_A_641_297#_c_431_n N_Y_M1004_d 0.00325424f $X=5.175 $Y=2.34 $X2=0 $Y2=0
cc_277 N_A_641_297#_M1005_d N_Y_c_486_n 0.00126758f $X=4.035 $Y=1.485 $X2=0
+ $Y2=0
cc_278 N_A_641_297#_c_431_n N_Y_c_486_n 0.0032538f $X=5.175 $Y=2.34 $X2=0 $Y2=0
cc_279 N_A_641_297#_M1005_d N_Y_c_476_n 0.00623313f $X=4.035 $Y=1.485 $X2=0
+ $Y2=0
cc_280 N_A_641_297#_c_427_n N_Y_c_476_n 0.0124446f $X=4.275 $Y=2 $X2=0 $Y2=0
cc_281 N_A_641_297#_c_431_n N_Y_c_476_n 0.00111169f $X=5.175 $Y=2.34 $X2=0 $Y2=0
cc_282 N_A_641_297#_M1005_d Y 7.22859e-19 $X=4.035 $Y=1.485 $X2=0 $Y2=0
cc_283 N_A_641_297#_c_427_n N_Y_c_495_n 0.0109026f $X=4.275 $Y=2 $X2=0 $Y2=0
cc_284 N_A_641_297#_c_431_n N_Y_c_495_n 0.0169852f $X=5.175 $Y=2.34 $X2=0 $Y2=0
cc_285 N_Y_c_460_n N_A_27_47#_c_536_n 0.0145425f $X=3.235 $Y=0.74 $X2=0 $Y2=0
cc_286 N_Y_c_469_n N_VGND_M1007_d 0.00313177f $X=4.085 $Y=0.74 $X2=0 $Y2=0
cc_287 N_Y_c_481_n N_VGND_M1008_s 0.00338858f $X=5.175 $Y=0.74 $X2=0 $Y2=0
cc_288 N_Y_c_467_n N_VGND_c_568_n 0.0148352f $X=3.32 $Y=0.42 $X2=0 $Y2=0
cc_289 N_Y_c_469_n N_VGND_c_568_n 0.0145262f $X=4.085 $Y=0.74 $X2=0 $Y2=0
cc_290 N_Y_c_480_n N_VGND_c_569_n 0.00771043f $X=4.17 $Y=0.42 $X2=0 $Y2=0
cc_291 N_Y_c_481_n N_VGND_c_569_n 0.0145262f $X=5.175 $Y=0.74 $X2=0 $Y2=0
cc_292 N_Y_c_460_n N_VGND_c_570_n 0.00261494f $X=3.235 $Y=0.74 $X2=0 $Y2=0
cc_293 N_Y_c_467_n N_VGND_c_570_n 0.0116627f $X=3.32 $Y=0.42 $X2=0 $Y2=0
cc_294 N_Y_c_469_n N_VGND_c_570_n 0.00242316f $X=4.085 $Y=0.74 $X2=0 $Y2=0
cc_295 N_Y_c_469_n N_VGND_c_573_n 0.00881568f $X=4.085 $Y=0.74 $X2=0 $Y2=0
cc_296 N_Y_c_480_n N_VGND_c_573_n 0.0111777f $X=4.17 $Y=0.42 $X2=0 $Y2=0
cc_297 N_Y_c_481_n N_VGND_c_574_n 0.0023303f $X=5.175 $Y=0.74 $X2=0 $Y2=0
cc_298 N_Y_c_521_p N_VGND_c_574_n 0.011459f $X=5.26 $Y=0.42 $X2=0 $Y2=0
cc_299 N_Y_M1010_d N_VGND_c_575_n 0.00213436f $X=2.335 $Y=0.235 $X2=0 $Y2=0
cc_300 N_Y_M1012_d N_VGND_c_575_n 0.00288092f $X=3.165 $Y=0.235 $X2=0 $Y2=0
cc_301 N_Y_M1011_s N_VGND_c_575_n 0.00557668f $X=4.035 $Y=0.235 $X2=0 $Y2=0
cc_302 N_Y_M1013_d N_VGND_c_575_n 0.00370147f $X=5.125 $Y=0.235 $X2=0 $Y2=0
cc_303 N_Y_c_460_n N_VGND_c_575_n 0.00607196f $X=3.235 $Y=0.74 $X2=0 $Y2=0
cc_304 N_Y_c_467_n N_VGND_c_575_n 0.00644035f $X=3.32 $Y=0.42 $X2=0 $Y2=0
cc_305 N_Y_c_469_n N_VGND_c_575_n 0.021179f $X=4.085 $Y=0.74 $X2=0 $Y2=0
cc_306 N_Y_c_480_n N_VGND_c_575_n 0.00638388f $X=4.17 $Y=0.42 $X2=0 $Y2=0
cc_307 N_Y_c_481_n N_VGND_c_575_n 0.00557926f $X=5.175 $Y=0.74 $X2=0 $Y2=0
cc_308 N_Y_c_521_p N_VGND_c_575_n 0.00644035f $X=5.26 $Y=0.42 $X2=0 $Y2=0
cc_309 N_Y_c_460_n N_A_277_47#_M1010_s 0.00309864f $X=3.235 $Y=0.74 $X2=0 $Y2=0
cc_310 N_Y_M1010_d N_A_277_47#_c_649_n 0.00484155f $X=2.335 $Y=0.235 $X2=0 $Y2=0
cc_311 N_Y_c_460_n N_A_277_47#_c_649_n 0.0372984f $X=3.235 $Y=0.74 $X2=0 $Y2=0
cc_312 N_Y_c_467_n N_A_277_47#_c_649_n 0.0121093f $X=3.32 $Y=0.42 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_537_n N_VGND_M1009_s 0.00313177f $X=1.015 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_314 N_A_27_47#_c_537_n N_VGND_c_567_n 0.0145262f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_27_47#_c_537_n N_VGND_c_570_n 0.0023303f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_553_p N_VGND_c_570_n 0.0112554f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_536_n N_VGND_c_570_n 0.00233958f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_27_47#_c_555_p N_VGND_c_572_n 0.011459f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_319 N_A_27_47#_c_537_n N_VGND_c_572_n 0.0023303f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_27_47#_M1009_d N_VGND_c_575_n 0.00370147f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_M1019_d N_VGND_c_575_n 0.00252188f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_M1016_d N_VGND_c_575_n 0.00213436f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_555_p N_VGND_c_575_n 0.00644035f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_324 N_A_27_47#_c_537_n N_VGND_c_575_n 0.00970918f $X=1.015 $Y=0.74 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_553_p N_VGND_c_575_n 0.00644035f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_326 N_A_27_47#_c_536_n N_VGND_c_575_n 0.00551407f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A_27_47#_c_536_n N_A_277_47#_M1015_s 0.00309864f $X=1.94 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_328 N_A_27_47#_M1016_d N_A_277_47#_c_649_n 0.00507876f $X=1.805 $Y=0.235
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_536_n N_A_277_47#_c_649_n 0.0372984f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_VGND_c_575_n N_A_277_47#_M1015_s 0.00218617f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_331 N_VGND_c_575_n N_A_277_47#_M1010_s 0.00218617f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_332 N_VGND_c_570_n N_A_277_47#_c_649_n 0.073805f $X=3.585 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_575_n N_A_277_47#_c_649_n 0.0590677f $X=5.29 $Y=0 $X2=0 $Y2=0

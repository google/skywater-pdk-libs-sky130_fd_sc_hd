* File: sky130_fd_sc_hd__sdfbbn_1.pxi.spice
* Created: Thu Aug 27 14:45:18 2020
* 
x_PM_SKY130_FD_SC_HD__SDFBBN_1%CLK_N N_CLK_N_c_313_n N_CLK_N_c_308_n
+ N_CLK_N_M1045_g N_CLK_N_c_314_n N_CLK_N_M1025_g N_CLK_N_c_309_n
+ N_CLK_N_c_315_n CLK_N CLK_N N_CLK_N_c_311_n N_CLK_N_c_312_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%CLK_N
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_27_47# N_A_27_47#_M1045_s N_A_27_47#_M1025_s
+ N_A_27_47#_M1026_g N_A_27_47#_M1000_g N_A_27_47#_M1039_g N_A_27_47#_c_354_n
+ N_A_27_47#_c_355_n N_A_27_47#_M1044_g N_A_27_47#_c_357_n N_A_27_47#_c_358_n
+ N_A_27_47#_M1010_g N_A_27_47#_M1019_g N_A_27_47#_c_359_n N_A_27_47#_c_360_n
+ N_A_27_47#_c_361_n N_A_27_47#_c_381_n N_A_27_47#_c_362_n N_A_27_47#_c_363_n
+ N_A_27_47#_c_364_n N_A_27_47#_c_382_n N_A_27_47#_c_383_n N_A_27_47#_c_384_n
+ N_A_27_47#_c_365_n N_A_27_47#_c_366_n N_A_27_47#_c_367_n N_A_27_47#_c_368_n
+ N_A_27_47#_c_369_n N_A_27_47#_c_370_n N_A_27_47#_c_371_n N_A_27_47#_c_372_n
+ N_A_27_47#_c_373_n N_A_27_47#_c_374_n N_A_27_47#_c_375_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%SCD N_SCD_c_639_n N_SCD_c_640_n N_SCD_c_641_n
+ N_SCD_M1007_g N_SCD_M1033_g SCD SCD N_SCD_c_646_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%SCD
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_423_315# N_A_423_315#_M1041_s
+ N_A_423_315#_M1034_s N_A_423_315#_c_697_n N_A_423_315#_M1038_g
+ N_A_423_315#_c_698_n N_A_423_315#_c_699_n N_A_423_315#_M1042_g
+ N_A_423_315#_c_757_p N_A_423_315#_c_700_n N_A_423_315#_c_691_n
+ N_A_423_315#_c_692_n N_A_423_315#_c_701_n N_A_423_315#_c_693_n
+ N_A_423_315#_c_694_n N_A_423_315#_c_703_n N_A_423_315#_c_695_n
+ N_A_423_315#_c_704_n N_A_423_315#_c_696_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_423_315#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%SCE N_SCE_c_804_n N_SCE_M1013_g N_SCE_c_805_n
+ N_SCE_c_806_n N_SCE_M1041_g N_SCE_c_807_n N_SCE_c_814_n N_SCE_c_815_n
+ N_SCE_M1034_g N_SCE_c_816_n N_SCE_c_817_n N_SCE_M1021_g N_SCE_c_808_n
+ N_SCE_c_809_n N_SCE_c_819_n SCE SCE SCE N_SCE_c_811_n N_SCE_c_812_n SCE
+ PM_SKY130_FD_SC_HD__SDFBBN_1%SCE
x_PM_SKY130_FD_SC_HD__SDFBBN_1%D N_D_M1027_g N_D_M1017_g D D N_D_c_923_n
+ N_D_c_924_n PM_SKY130_FD_SC_HD__SDFBBN_1%D
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_193_47# N_A_193_47#_M1026_d N_A_193_47#_M1000_d
+ N_A_193_47#_c_976_n N_A_193_47#_M1014_g N_A_193_47#_M1011_g
+ N_A_193_47#_M1031_g N_A_193_47#_c_977_n N_A_193_47#_c_978_n
+ N_A_193_47#_M1024_g N_A_193_47#_c_980_n N_A_193_47#_c_981_n
+ N_A_193_47#_c_982_n N_A_193_47#_c_989_n N_A_193_47#_c_990_n
+ N_A_193_47#_c_991_n N_A_193_47#_c_992_n N_A_193_47#_c_993_n
+ N_A_193_47#_c_994_n N_A_193_47#_c_995_n N_A_193_47#_c_996_n
+ N_A_193_47#_c_997_n N_A_193_47#_c_998_n N_A_193_47#_c_983_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_1102_21# N_A_1102_21#_M1040_d
+ N_A_1102_21#_M1012_d N_A_1102_21#_M1009_g N_A_1102_21#_M1035_g
+ N_A_1102_21#_M1047_g N_A_1102_21#_c_1202_n N_A_1102_21#_M1016_g
+ N_A_1102_21#_c_1211_n N_A_1102_21#_c_1260_p N_A_1102_21#_c_1223_n
+ N_A_1102_21#_c_1203_n N_A_1102_21#_c_1204_n N_A_1102_21#_c_1205_n
+ N_A_1102_21#_c_1213_n N_A_1102_21#_c_1214_n N_A_1102_21#_c_1228_n
+ N_A_1102_21#_c_1206_n N_A_1102_21#_c_1207_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_1102_21#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%SET_B N_SET_B_M1004_g N_SET_B_c_1349_n
+ N_SET_B_M1012_g N_SET_B_M1006_g N_SET_B_M1008_g SET_B N_SET_B_c_1354_n
+ N_SET_B_c_1355_n N_SET_B_c_1356_n N_SET_B_c_1357_n N_SET_B_c_1358_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%SET_B
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_917_47# N_A_917_47#_M1014_d N_A_917_47#_M1039_d
+ N_A_917_47#_M1040_g N_A_917_47#_c_1479_n N_A_917_47#_M1036_g
+ N_A_917_47#_c_1490_n N_A_917_47#_c_1495_n N_A_917_47#_c_1485_n
+ N_A_917_47#_c_1498_n N_A_917_47#_c_1480_n N_A_917_47#_c_1481_n
+ N_A_917_47#_c_1482_n PM_SKY130_FD_SC_HD__SDFBBN_1%A_917_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_1396_21# N_A_1396_21#_M1015_s
+ N_A_1396_21#_M1005_s N_A_1396_21#_M1032_g N_A_1396_21#_M1030_g
+ N_A_1396_21#_M1028_g N_A_1396_21#_M1029_g N_A_1396_21#_c_1593_n
+ N_A_1396_21#_c_1594_n N_A_1396_21#_c_1602_n N_A_1396_21#_c_1603_n
+ N_A_1396_21#_c_1595_n N_A_1396_21#_c_1596_n N_A_1396_21#_c_1605_n
+ N_A_1396_21#_c_1606_n N_A_1396_21#_c_1607_n N_A_1396_21#_c_1608_n
+ N_A_1396_21#_c_1597_n N_A_1396_21#_c_1598_n N_A_1396_21#_c_1599_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_1396_21#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_1887_21# N_A_1887_21#_M1020_d
+ N_A_1887_21#_M1008_d N_A_1887_21#_M1003_g N_A_1887_21#_M1043_g
+ N_A_1887_21#_c_1753_n N_A_1887_21#_M1001_g N_A_1887_21#_M1037_g
+ N_A_1887_21#_c_1754_n N_A_1887_21#_c_1755_n N_A_1887_21#_c_1756_n
+ N_A_1887_21#_c_1757_n N_A_1887_21#_M1046_g N_A_1887_21#_c_1767_n
+ N_A_1887_21#_M1022_g N_A_1887_21#_c_1758_n N_A_1887_21#_c_1759_n
+ N_A_1887_21#_c_1768_n N_A_1887_21#_c_1769_n N_A_1887_21#_c_1770_n
+ N_A_1887_21#_c_1771_n N_A_1887_21#_c_1829_p N_A_1887_21#_c_1877_p
+ N_A_1887_21#_c_1800_n N_A_1887_21#_c_1760_n N_A_1887_21#_c_1773_n
+ N_A_1887_21#_c_1774_n N_A_1887_21#_c_1817_n N_A_1887_21#_c_1793_n
+ N_A_1887_21#_c_1820_n N_A_1887_21#_c_1761_n N_A_1887_21#_c_1762_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_1887_21#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_1714_47# N_A_1714_47#_M1010_d
+ N_A_1714_47#_M1031_d N_A_1714_47#_M1020_g N_A_1714_47#_M1023_g
+ N_A_1714_47#_c_1945_n N_A_1714_47#_c_1948_n N_A_1714_47#_c_1934_n
+ N_A_1714_47#_c_1940_n N_A_1714_47#_c_1935_n N_A_1714_47#_c_1936_n
+ N_A_1714_47#_c_1937_n N_A_1714_47#_c_1938_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_1714_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%RESET_B N_RESET_B_M1015_g N_RESET_B_M1005_g
+ RESET_B N_RESET_B_c_2034_n PM_SKY130_FD_SC_HD__SDFBBN_1%RESET_B
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_2596_47# N_A_2596_47#_M1046_s
+ N_A_2596_47#_M1022_s N_A_2596_47#_M1018_g N_A_2596_47#_M1002_g
+ N_A_2596_47#_c_2068_n N_A_2596_47#_c_2074_n N_A_2596_47#_c_2069_n
+ N_A_2596_47#_c_2070_n N_A_2596_47#_c_2071_n N_A_2596_47#_c_2072_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_2596_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%VPWR N_VPWR_M1025_d N_VPWR_M1033_s N_VPWR_M1034_d
+ N_VPWR_M1035_d N_VPWR_M1030_d N_VPWR_M1043_d N_VPWR_M1028_d N_VPWR_M1005_d
+ N_VPWR_M1022_d N_VPWR_c_2121_n N_VPWR_c_2122_n N_VPWR_c_2123_n N_VPWR_c_2124_n
+ N_VPWR_c_2125_n N_VPWR_c_2126_n N_VPWR_c_2127_n N_VPWR_c_2128_n
+ N_VPWR_c_2129_n N_VPWR_c_2130_n VPWR VPWR N_VPWR_c_2131_n N_VPWR_c_2132_n
+ N_VPWR_c_2133_n N_VPWR_c_2134_n N_VPWR_c_2135_n N_VPWR_c_2136_n
+ N_VPWR_c_2137_n N_VPWR_c_2138_n N_VPWR_c_2120_n N_VPWR_c_2140_n
+ N_VPWR_c_2141_n N_VPWR_c_2142_n N_VPWR_c_2143_n N_VPWR_c_2144_n
+ N_VPWR_c_2145_n N_VPWR_c_2146_n PM_SKY130_FD_SC_HD__SDFBBN_1%VPWR
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_453_47# N_A_453_47#_M1013_d N_A_453_47#_M1027_d
+ N_A_453_47#_M1038_d N_A_453_47#_M1017_d N_A_453_47#_c_2328_n
+ N_A_453_47#_c_2329_n N_A_453_47#_c_2330_n N_A_453_47#_c_2338_n
+ N_A_453_47#_c_2339_n N_A_453_47#_c_2331_n N_A_453_47#_c_2348_n
+ N_A_453_47#_c_2349_n N_A_453_47#_c_2340_n N_A_453_47#_c_2332_n
+ N_A_453_47#_c_2333_n N_A_453_47#_c_2334_n N_A_453_47#_c_2335_n
+ N_A_453_47#_c_2336_n PM_SKY130_FD_SC_HD__SDFBBN_1%A_453_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%Q_N N_Q_N_M1001_d N_Q_N_M1037_d N_Q_N_c_2490_n
+ N_Q_N_c_2487_n Q_N Q_N Q_N N_Q_N_c_2489_n Q_N PM_SKY130_FD_SC_HD__SDFBBN_1%Q_N
x_PM_SKY130_FD_SC_HD__SDFBBN_1%Q N_Q_M1018_d N_Q_M1002_d N_Q_c_2517_n
+ N_Q_c_2520_n N_Q_c_2518_n Q Q Q PM_SKY130_FD_SC_HD__SDFBBN_1%Q
x_PM_SKY130_FD_SC_HD__SDFBBN_1%VGND N_VGND_M1045_d N_VGND_M1007_s N_VGND_M1041_d
+ N_VGND_M1009_d N_VGND_M1016_s N_VGND_M1003_d N_VGND_M1015_d N_VGND_M1046_d
+ N_VGND_c_2533_n N_VGND_c_2534_n N_VGND_c_2535_n N_VGND_c_2536_n
+ N_VGND_c_2537_n N_VGND_c_2538_n N_VGND_c_2539_n N_VGND_c_2540_n
+ N_VGND_c_2541_n N_VGND_c_2542_n N_VGND_c_2543_n N_VGND_c_2544_n
+ N_VGND_c_2545_n N_VGND_c_2546_n VGND VGND N_VGND_c_2547_n N_VGND_c_2548_n
+ N_VGND_c_2549_n N_VGND_c_2550_n N_VGND_c_2551_n N_VGND_c_2552_n
+ N_VGND_c_2553_n N_VGND_c_2554_n N_VGND_c_2555_n N_VGND_c_2556_n
+ N_VGND_c_2557_n N_VGND_c_2558_n PM_SKY130_FD_SC_HD__SDFBBN_1%VGND
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_1241_47# N_A_1241_47#_M1004_d
+ N_A_1241_47#_M1032_d N_A_1241_47#_c_2756_n N_A_1241_47#_c_2759_n
+ N_A_1241_47#_c_2766_n PM_SKY130_FD_SC_HD__SDFBBN_1%A_1241_47#
x_PM_SKY130_FD_SC_HD__SDFBBN_1%A_2004_47# N_A_2004_47#_M1006_d
+ N_A_2004_47#_M1029_d N_A_2004_47#_c_2790_n N_A_2004_47#_c_2786_n
+ PM_SKY130_FD_SC_HD__SDFBBN_1%A_2004_47#
cc_1 VNB N_CLK_N_c_308_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_N_c_309_n 0.022961f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK_N 0.0164093f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_N_c_311_n 0.0195341f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_CLK_N_c_312_n 0.0141401f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1026_g 0.0381872f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_354_n 0.0129551f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_A_27_47#_c_355_n 0.00459297f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_9 VNB N_A_27_47#_M1044_g 0.0215804f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_10 VNB N_A_27_47#_c_357_n 0.00887161f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_11 VNB N_A_27_47#_c_358_n 0.018237f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_12 VNB N_A_27_47#_c_359_n 0.0110359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_360_n 7.55444e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_361_n 0.00777415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_362_n 0.00302102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_363_n 0.0314088f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_364_n 0.00454848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_365_n 0.0331664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_366_n 0.00310819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_367_n 0.00103865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_368_n 0.0218696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_369_n 0.00113053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_370_n 0.00292248f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_371_n 0.00300617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_372_n 0.00196881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_373_n 0.00147534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_374_n 0.0239438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_375_n 0.0265632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_SCD_c_639_n 0.0205861f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_30 VNB N_SCD_c_640_n 0.0270831f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.07
cc_31 VNB N_SCD_c_641_n 0.0174657f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_32 VNB SCD 0.00341923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_423_315#_c_691_n 0.00241998f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_34 VNB N_A_423_315#_c_692_n 6.63947e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_35 VNB N_A_423_315#_c_693_n 0.00853678f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_36 VNB N_A_423_315#_c_694_n 0.00305016f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_37 VNB N_A_423_315#_c_695_n 0.0277476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_423_315#_c_696_n 0.0158279f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_SCE_c_804_n 0.0168392f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_40 VNB N_SCE_c_805_n 0.0413612f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.59
cc_41 VNB N_SCE_c_806_n 0.0177358f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_42 VNB N_SCE_c_807_n 0.0243731f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_43 VNB N_SCE_c_808_n 0.00422122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_SCE_c_809_n 0.00782164f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_45 VNB SCE 0.00160574f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_46 VNB N_SCE_c_811_n 0.0357353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_SCE_c_812_n 0.00372596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB SCE 0.00326522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_D_M1027_g 0.044552f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_50 VNB N_A_193_47#_c_976_n 0.0182085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_51 VNB N_A_193_47#_c_977_n 0.0123509f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_52 VNB N_A_193_47#_c_978_n 0.00338667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_193_47#_M1024_g 0.0470486f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_54 VNB N_A_193_47#_c_980_n 0.00248736f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_55 VNB N_A_193_47#_c_981_n 0.00245151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_193_47#_c_982_n 0.0361921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_193_47#_c_983_n 0.017705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1102_21#_M1009_g 0.0391229f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_59 VNB N_A_1102_21#_c_1202_n 0.0193514f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_60 VNB N_A_1102_21#_c_1203_n 0.00172002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1102_21#_c_1204_n 0.00168282f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_62 VNB N_A_1102_21#_c_1205_n 0.0120378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1102_21#_c_1206_n 0.00605681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1102_21#_c_1207_n 0.0322423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_SET_B_M1004_g 0.020438f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_66 VNB N_SET_B_c_1349_n 0.0333483f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_67 VNB N_SET_B_M1012_g 0.00707886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_68 VNB N_SET_B_M1006_g 0.0200592f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_69 VNB N_SET_B_M1008_g 0.00796403f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_70 VNB SET_B 0.00789765f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_71 VNB N_SET_B_c_1354_n 0.0157323f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_72 VNB N_SET_B_c_1355_n 0.0019592f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_73 VNB N_SET_B_c_1356_n 0.00209085f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_74 VNB N_SET_B_c_1357_n 0.00534937f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_75 VNB N_SET_B_c_1358_n 0.0320885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_917_47#_M1040_g 0.025905f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_77 VNB N_A_917_47#_c_1479_n 0.0122117f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_78 VNB N_A_917_47#_c_1480_n 0.00794493f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_79 VNB N_A_917_47#_c_1481_n 0.00813299f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_80 VNB N_A_917_47#_c_1482_n 0.00378595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1396_21#_M1032_g 0.0290696f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_82 VNB N_A_1396_21#_M1029_g 0.0279648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1396_21#_c_1593_n 0.0112366f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_84 VNB N_A_1396_21#_c_1594_n 0.00216934f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_85 VNB N_A_1396_21#_c_1595_n 0.00260218f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_86 VNB N_A_1396_21#_c_1596_n 9.08783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1396_21#_c_1597_n 0.0242128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1396_21#_c_1598_n 0.0195979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1396_21#_c_1599_n 0.00516403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1887_21#_M1003_g 0.0443092f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_91 VNB N_A_1887_21#_c_1753_n 0.0204895f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_92 VNB N_A_1887_21#_c_1754_n 0.053914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_1887_21#_c_1755_n 0.00812918f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_94 VNB N_A_1887_21#_c_1756_n 4.83843e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_95 VNB N_A_1887_21#_c_1757_n 0.0183894f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_96 VNB N_A_1887_21#_c_1758_n 0.0180373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_1887_21#_c_1759_n 0.00820903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_1887_21#_c_1760_n 0.0032181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_1887_21#_c_1761_n 0.00274082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_1887_21#_c_1762_n 0.0150907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_1714_47#_M1020_g 0.022372f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_102 VNB N_A_1714_47#_c_1934_n 0.0117442f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_103 VNB N_A_1714_47#_c_1935_n 0.0114112f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_104 VNB N_A_1714_47#_c_1936_n 4.78869e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_A_1714_47#_c_1937_n 0.00178317f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_106 VNB N_A_1714_47#_c_1938_n 0.0176282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_RESET_B_M1015_g 0.0349589f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_108 VNB RESET_B 0.00386832f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_109 VNB N_RESET_B_c_2034_n 0.028487f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_110 VNB N_A_2596_47#_c_2068_n 0.0072656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_A_2596_47#_c_2069_n 0.00526785f $X=-0.19 $Y=-0.24 $X2=0.24
+ $Y2=1.235
cc_112 VNB N_A_2596_47#_c_2070_n 0.0253082f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_113 VNB N_A_2596_47#_c_2071_n 2.89573e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_114 VNB N_A_2596_47#_c_2072_n 0.0201038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VPWR_c_2120_n 0.592346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_A_453_47#_c_2328_n 0.00501575f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_117 VNB N_A_453_47#_c_2329_n 0.00527679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_A_453_47#_c_2330_n 0.00546227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_A_453_47#_c_2331_n 0.0044763f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_120 VNB N_A_453_47#_c_2332_n 0.00719271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_A_453_47#_c_2333_n 0.00101315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_A_453_47#_c_2334_n 0.00683943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_A_453_47#_c_2335_n 0.00268493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_A_453_47#_c_2336_n 0.00894414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_Q_N_c_2487_n 0.00377264f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_126 VNB Q_N 0.00140118f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_127 VNB N_Q_N_c_2489_n 0.00366681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_Q_c_2517_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_129 VNB N_Q_c_2518_n 0.0244322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB Q 0.0155218f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_131 VNB N_VGND_c_2533_n 4.08532e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_132 VNB N_VGND_c_2534_n 0.00948744f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_133 VNB N_VGND_c_2535_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2536_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2537_n 0.00562688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2538_n 0.00244296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2539_n 0.00555851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2540_n 0.00259569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2541_n 0.0578465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2542_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2543_n 0.0398903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2544_n 0.00540406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2545_n 0.0404697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2546_n 0.0037591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2547_n 0.0147647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2548_n 0.0157857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2549_n 0.0402043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2550_n 0.0540515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2551_n 0.0289512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2552_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2553_n 0.65913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2554_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2555_n 0.00526527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2556_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2557_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2558_n 0.00430718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_157 VPB N_CLK_N_c_313_n 0.0118979f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_158 VPB N_CLK_N_c_314_n 0.0186097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_159 VPB N_CLK_N_c_315_n 0.0238007f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_160 VPB CLK_N 0.0154846f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_161 VPB N_CLK_N_c_311_n 0.0100928f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_162 VPB N_A_27_47#_M1000_g 0.0375468f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_163 VPB N_A_27_47#_M1039_g 0.0466111f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_164 VPB N_A_27_47#_c_354_n 0.0179398f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_165 VPB N_A_27_47#_c_355_n 0.00349583f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_166 VPB N_A_27_47#_M1019_g 0.0221986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_27_47#_c_381_n 0.0018848f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_27_47#_c_382_n 0.0038403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_27_47#_c_383_n 0.0288235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_27_47#_c_384_n 0.0294336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_27_47#_c_370_n 0.00321856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_27_47#_c_373_n 2.53141e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_27_47#_c_374_n 0.0119971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_SCD_c_640_n 0.00121161f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.07
cc_175 VPB N_SCD_M1033_g 0.0216746f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_176 VPB SCD 0.00516166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_SCD_c_646_n 0.0412346f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_178 VPB N_A_423_315#_c_697_n 0.0182151f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_179 VPB N_A_423_315#_c_698_n 0.0313294f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_180 VPB N_A_423_315#_c_699_n 0.00762464f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_181 VPB N_A_423_315#_c_700_n 0.00342623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_423_315#_c_701_n 0.00510623f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_183 VPB N_A_423_315#_c_694_n 0.00541848f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_184 VPB N_A_423_315#_c_703_n 0.00313836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_423_315#_c_704_n 0.0336341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_SCE_c_814_n 0.0251528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_SCE_c_815_n 0.0173084f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_188 VPB N_SCE_c_816_n 0.02507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_SCE_c_817_n 0.0144409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_SCE_c_809_n 0.0101059f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_191 VPB N_SCE_c_819_n 0.0054195f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_192 VPB SCE 0.00817088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_D_M1027_g 0.00332407f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_194 VPB N_D_M1017_g 0.0342848f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_195 VPB D 0.00446496f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_196 VPB N_D_c_923_n 0.0380878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_D_c_924_n 0.00243882f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_198 VPB N_A_193_47#_M1011_g 0.0215674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_193_47#_M1031_g 0.020906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_193_47#_c_977_n 0.017753f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_201 VPB N_A_193_47#_c_978_n 0.00403587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_193_47#_c_980_n 0.00290906f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_203 VPB N_A_193_47#_c_989_n 0.0289063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_193_47#_c_990_n 0.00491076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_193_47#_c_991_n 0.0082441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_193_47#_c_992_n 0.00165593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_193_47#_c_993_n 0.00361706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_193_47#_c_994_n 0.026688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_193_47#_c_995_n 0.00617568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_193_47#_c_996_n 0.0282388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_A_193_47#_c_997_n 0.00514398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_193_47#_c_998_n 0.0125285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_193_47#_c_983_n 0.0180042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_1102_21#_M1009_g 0.0151853f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_215 VPB N_A_1102_21#_M1035_g 0.0210587f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_216 VPB N_A_1102_21#_M1047_g 0.0317411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_217 VPB N_A_1102_21#_c_1211_n 0.00546651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_1102_21#_c_1204_n 0.00530406f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_219 VPB N_A_1102_21#_c_1213_n 0.0059313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1102_21#_c_1214_n 0.0330038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1102_21#_c_1207_n 0.00659461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_SET_B_M1012_g 0.0510974f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_223 VPB N_SET_B_M1008_g 0.0496972f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_224 VPB N_A_917_47#_c_1479_n 0.0180645f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_225 VPB N_A_917_47#_M1036_g 0.0203673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_226 VPB N_A_917_47#_c_1485_n 0.0121294f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_227 VPB N_A_917_47#_c_1481_n 0.00821712f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_228 VPB N_A_917_47#_c_1482_n 0.00219434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_1396_21#_M1030_g 0.0205161f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_230 VPB N_A_1396_21#_M1028_g 0.0210669f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_231 VPB N_A_1396_21#_c_1602_n 0.0018943f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_232 VPB N_A_1396_21#_c_1603_n 0.0051975f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_233 VPB N_A_1396_21#_c_1596_n 0.00162652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_1396_21#_c_1605_n 0.0327539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_1396_21#_c_1606_n 0.00261931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_1396_21#_c_1607_n 0.00737873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_A_1396_21#_c_1608_n 0.00331979f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_1396_21#_c_1597_n 0.0219071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_A_1396_21#_c_1598_n 0.025869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_1396_21#_c_1599_n 0.00361429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_A_1887_21#_M1003_g 0.0159956f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_242 VPB N_A_1887_21#_M1043_g 0.021027f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_243 VPB N_A_1887_21#_M1037_g 0.0245592f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_244 VPB N_A_1887_21#_c_1756_n 0.0131751f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_245 VPB N_A_1887_21#_c_1767_n 0.0188717f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_246 VPB N_A_1887_21#_c_1768_n 0.0180742f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_A_1887_21#_c_1769_n 0.00423323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_A_1887_21#_c_1770_n 0.0329665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_A_1887_21#_c_1771_n 0.00304218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_A_1887_21#_c_1760_n 0.00331106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_A_1887_21#_c_1773_n 0.0072909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_A_1887_21#_c_1774_n 0.0016887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_A_1887_21#_c_1761_n 2.41561e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_A_1887_21#_c_1762_n 0.00402209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_A_1714_47#_M1023_g 0.021833f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_256 VPB N_A_1714_47#_c_1940_n 0.0117899f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_257 VPB N_A_1714_47#_c_1935_n 0.00583428f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_258 VPB N_A_1714_47#_c_1936_n 7.45241e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_A_1714_47#_c_1937_n 0.00126723f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_260 VPB N_A_1714_47#_c_1938_n 0.00898586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_RESET_B_M1005_g 0.0248581f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_262 VPB RESET_B 9.55576e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_263 VPB N_RESET_B_c_2034_n 0.00925958f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_264 VPB N_A_2596_47#_M1002_g 0.024323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_A_2596_47#_c_2074_n 0.0132727f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_266 VPB N_A_2596_47#_c_2069_n 0.00532263f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_267 VPB N_A_2596_47#_c_2070_n 0.00545303f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_268 VPB N_VPWR_c_2121_n 0.00105358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_2122_n 0.00871789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_2123_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_2124_n 0.00313724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_2125_n 0.00562862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_2126_n 0.00349941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_2127_n 0.0292737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_2128_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_2129_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_2130_n 0.022998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_2131_n 0.0147455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_2132_n 0.0156521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_2133_n 0.0421083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_2134_n 0.0533335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_2135_n 0.0591311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_2136_n 0.0306954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_2137_n 0.0293379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_2138_n 0.0152168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_2120_n 0.0748962f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_2140_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_2141_n 0.00579271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_2142_n 0.0043639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_2143_n 0.00609488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_2144_n 0.00928062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_2145_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_2146_n 0.00424285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_294 VPB N_A_453_47#_c_2328_n 0.00436598f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_295 VPB N_A_453_47#_c_2338_n 0.0062713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_296 VPB N_A_453_47#_c_2339_n 0.00316476f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_297 VPB N_A_453_47#_c_2340_n 0.0132288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_298 VPB N_A_453_47#_c_2334_n 0.00448045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_299 VPB N_A_453_47#_c_2335_n 0.00140728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_300 VPB N_A_453_47#_c_2336_n 3.85213e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_301 VPB N_Q_N_c_2490_n 0.00137514f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_302 VPB N_Q_N_c_2487_n 0.00384198f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_303 VPB Q_N 0.00760625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_304 VPB N_Q_c_2520_n 0.00715183f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_305 VPB N_Q_c_2518_n 0.00847384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_306 VPB Q 0.0331954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_307 N_CLK_N_c_308_n N_A_27_47#_M1026_g 0.0205277f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_308 CLK_N N_A_27_47#_M1026_g 3.07529e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_309 N_CLK_N_c_312_n N_A_27_47#_M1026_g 0.00498861f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_310 N_CLK_N_c_315_n N_A_27_47#_M1000_g 0.0275641f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_311 CLK_N N_A_27_47#_M1000_g 5.68848e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_312 N_CLK_N_c_311_n N_A_27_47#_M1000_g 0.00521293f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_313 N_CLK_N_c_308_n N_A_27_47#_c_360_n 0.00694711f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_314 N_CLK_N_c_309_n N_A_27_47#_c_360_n 0.00799602f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_315 CLK_N N_A_27_47#_c_360_n 0.00698378f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_316 N_CLK_N_c_309_n N_A_27_47#_c_361_n 0.00634383f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_317 CLK_N N_A_27_47#_c_361_n 0.021626f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_318 N_CLK_N_c_311_n N_A_27_47#_c_361_n 7.17088e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_319 N_CLK_N_c_314_n N_A_27_47#_c_381_n 0.0129659f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_320 N_CLK_N_c_315_n N_A_27_47#_c_381_n 0.0013404f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_321 CLK_N N_A_27_47#_c_381_n 0.00690269f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_322 N_CLK_N_c_314_n N_A_27_47#_c_384_n 2.2023e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_323 N_CLK_N_c_315_n N_A_27_47#_c_384_n 0.00374438f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_324 CLK_N N_A_27_47#_c_384_n 0.0227757f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_325 N_CLK_N_c_311_n N_A_27_47#_c_384_n 5.66731e-19 $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_326 N_CLK_N_c_309_n N_A_27_47#_c_366_n 0.0017166f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_327 N_CLK_N_c_312_n N_A_27_47#_c_366_n 0.00154887f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_328 N_CLK_N_c_309_n N_A_27_47#_c_370_n 0.00155723f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_329 N_CLK_N_c_315_n N_A_27_47#_c_370_n 0.0045823f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_330 CLK_N N_A_27_47#_c_370_n 0.0517134f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_331 N_CLK_N_c_311_n N_A_27_47#_c_370_n 0.00100166f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_332 N_CLK_N_c_312_n N_A_27_47#_c_370_n 0.00207651f $X=0.24 $Y=1.07 $X2=0
+ $Y2=0
cc_333 CLK_N N_A_27_47#_c_374_n 0.00162145f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_334 N_CLK_N_c_311_n N_A_27_47#_c_374_n 0.0169859f $X=0.24 $Y=1.235 $X2=0
+ $Y2=0
cc_335 N_CLK_N_c_314_n N_VPWR_c_2121_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_336 N_CLK_N_c_314_n N_VPWR_c_2131_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_337 N_CLK_N_c_314_n N_VPWR_c_2120_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_338 N_CLK_N_c_308_n N_VGND_c_2533_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_339 N_CLK_N_c_308_n N_VGND_c_2547_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_340 N_CLK_N_c_309_n N_VGND_c_2547_n 4.87495e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_341 N_CLK_N_c_308_n N_VGND_c_2553_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_342 N_A_27_47#_M1026_g N_SCD_c_639_n 0.00428787f $X=0.89 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_343 N_A_27_47#_c_365_n N_SCD_c_639_n 0.007436f $X=5.095 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_344 N_A_27_47#_c_365_n N_SCD_c_640_n 0.00364587f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_345 N_A_27_47#_c_374_n N_SCD_c_640_n 0.00428787f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_365_n SCD 0.00880959f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_347 N_A_27_47#_c_365_n N_SCD_c_646_n 0.00214559f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_348 N_A_27_47#_c_374_n N_SCD_c_646_n 0.00541562f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_349 N_A_27_47#_c_365_n N_A_423_315#_c_691_n 0.01551f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_365_n N_A_423_315#_c_692_n 0.00650835f $X=5.095 $Y=0.85
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_365_n N_A_423_315#_c_693_n 0.0219941f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_365_n N_SCE_c_805_n 0.00433321f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_353 N_A_27_47#_c_365_n N_SCE_c_807_n 0.00222485f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_365_n N_SCE_c_808_n 5.06978e-19 $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_365_n N_SCE_c_809_n 4.62069e-19 $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_356 N_A_27_47#_c_365_n SCE 0.00840674f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_365_n N_SCE_c_811_n 0.00664112f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_365_n N_SCE_c_812_n 0.0211739f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_365_n SCE 8.83519e-19 $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_360 N_A_27_47#_c_355_n N_D_M1027_g 0.00262015f $X=4.665 $Y=1.32 $X2=0 $Y2=0
cc_361 N_A_27_47#_M1039_g N_D_M1017_g 0.0168061f $X=4.59 $Y=2.275 $X2=0 $Y2=0
cc_362 N_A_27_47#_c_355_n N_D_c_923_n 0.0168061f $X=4.665 $Y=1.32 $X2=0 $Y2=0
cc_363 N_A_27_47#_M1044_g N_A_193_47#_c_976_n 0.0133222f $X=5.075 $Y=0.415 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_M1039_g N_A_193_47#_M1011_g 0.0190294f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_364_n N_A_193_47#_c_977_n 0.0110233f $X=8.937 $Y=1.305 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_382_n N_A_193_47#_c_977_n 0.00852739f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_383_n N_A_193_47#_c_977_n 0.0213022f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_373_n N_A_193_47#_c_977_n 3.23054e-19 $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_362_n N_A_193_47#_c_978_n 2.62384e-19 $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_363_n N_A_193_47#_c_978_n 0.0206253f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_364_n N_A_193_47#_c_978_n 0.00356667f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_373_n N_A_193_47#_c_978_n 9.01357e-19 $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_358_n N_A_193_47#_M1024_g 0.0131194f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_362_n N_A_193_47#_M1024_g 0.00310082f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_363_n N_A_193_47#_M1024_g 0.0213524f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_364_n N_A_193_47#_M1024_g 0.00638693f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_M1039_g N_A_193_47#_c_980_n 0.00528668f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_354_n N_A_193_47#_c_980_n 0.00831083f $X=5 $Y=1.32 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_355_n N_A_193_47#_c_980_n 0.0022386f $X=4.665 $Y=1.32 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_369_n N_A_193_47#_c_980_n 0.00410439f $X=5.385 $Y=1.19 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_375_n N_A_193_47#_c_980_n 0.00664557f $X=5.165 $Y=0.93 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_355_n N_A_193_47#_c_981_n 3.39184e-19 $X=4.665 $Y=1.32 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_M1044_g N_A_193_47#_c_981_n 0.0012712f $X=5.075 $Y=0.415 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_365_n N_A_193_47#_c_981_n 0.016789f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_367_n N_A_193_47#_c_981_n 0.00434229f $X=5.277 $Y=1.12 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_371_n N_A_193_47#_c_981_n 4.98674e-19 $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_372_n N_A_193_47#_c_981_n 0.0150146f $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_355_n N_A_193_47#_c_982_n 0.0188524f $X=4.665 $Y=1.32 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1044_g N_A_193_47#_c_982_n 0.0215913f $X=5.075 $Y=0.415 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_365_n N_A_193_47#_c_982_n 0.00704926f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_372_n N_A_193_47#_c_982_n 9.68262e-19 $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_M1039_g N_A_193_47#_c_989_n 0.00642348f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_M1000_g N_A_193_47#_c_990_n 0.00459685f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_381_n N_A_193_47#_c_990_n 0.00561563f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_370_n N_A_193_47#_c_990_n 0.00113557f $X=0.69 $Y=0.85 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_354_n N_A_193_47#_c_991_n 3.07651e-19 $X=5 $Y=1.32 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_369_n N_A_193_47#_c_991_n 0.113653f $X=5.385 $Y=1.19 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_M1039_g N_A_193_47#_c_992_n 5.24592e-19 $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_M1019_g N_A_193_47#_c_993_n 0.00133927f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_400 N_A_27_47#_c_382_n N_A_193_47#_c_993_n 0.00483121f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_383_n N_A_193_47#_c_993_n 0.00219663f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_M1039_g N_A_193_47#_c_994_n 0.0174486f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_354_n N_A_193_47#_c_994_n 0.0215712f $X=5 $Y=1.32 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_372_n N_A_193_47#_c_994_n 4.47525e-19 $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_M1039_g N_A_193_47#_c_995_n 0.00918811f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_354_n N_A_193_47#_c_995_n 0.0080751f $X=5 $Y=1.32 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_372_n N_A_193_47#_c_995_n 0.00377721f $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_M1019_g N_A_193_47#_c_996_n 0.0192968f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_382_n N_A_193_47#_c_996_n 5.88448e-19 $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_c_383_n N_A_193_47#_c_996_n 0.0169266f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_c_368_n N_A_193_47#_c_996_n 2.37019e-19 $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_M1019_g N_A_193_47#_c_997_n 6.52047e-19 $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_364_n N_A_193_47#_c_997_n 0.00682571f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_382_n N_A_193_47#_c_997_n 0.0168759f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_383_n N_A_193_47#_c_997_n 0.00153059f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_373_n N_A_193_47#_c_997_n 0.00149027f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_382_n N_A_193_47#_c_998_n 0.00347329f $X=8.955 $Y=1.74 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_M1026_g N_A_193_47#_c_983_n 0.0158807f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_360_n N_A_193_47#_c_983_n 0.011372f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_c_381_n N_A_193_47#_c_983_n 0.00862152f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_365_n N_A_193_47#_c_983_n 0.0271407f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_366_n N_A_193_47#_c_983_n 0.00145827f $X=0.835 $Y=0.85 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_370_n N_A_193_47#_c_983_n 0.0688642f $X=0.69 $Y=0.85 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_M1044_g N_A_1102_21#_M1009_g 0.0215231f $X=5.075 $Y=0.415
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_c_357_n N_A_1102_21#_M1009_g 0.0124743f $X=5.102 $Y=1.245
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_372_n N_A_1102_21#_M1009_g 7.27967e-19 $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_375_n N_A_1102_21#_M1009_g 0.0215509f $X=5.165 $Y=0.93 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_358_n N_A_1102_21#_c_1202_n 0.0328414f $X=8.495 $Y=0.705
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_362_n N_A_1102_21#_c_1202_n 0.00159059f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_368_n N_A_1102_21#_c_1211_n 0.00196084f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_368_n N_A_1102_21#_c_1223_n 0.00352482f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_368_n N_A_1102_21#_c_1203_n 0.00183112f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_368_n N_A_1102_21#_c_1204_n 0.0155502f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_c_368_n N_A_1102_21#_c_1205_n 0.00982723f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_368_n N_A_1102_21#_c_1213_n 8.24776e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_368_n N_A_1102_21#_c_1228_n 6.83984e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_437 N_A_27_47#_c_362_n N_A_1102_21#_c_1206_n 0.0111636f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_363_n N_A_1102_21#_c_1206_n 9.32912e-19 $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_364_n N_A_1102_21#_c_1206_n 0.00462764f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_368_n N_A_1102_21#_c_1206_n 0.0153364f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_373_n N_A_1102_21#_c_1206_n 0.00129536f $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_362_n N_A_1102_21#_c_1207_n 5.74798e-19 $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_363_n N_A_1102_21#_c_1207_n 0.00181008f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_364_n N_A_1102_21#_c_1207_n 0.00174717f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_368_n N_A_1102_21#_c_1207_n 0.00365485f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_373_n N_A_1102_21#_c_1207_n 6.8647e-19 $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_368_n N_SET_B_c_1349_n 0.00468202f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_368_n N_SET_B_M1012_g 0.00120025f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_368_n SET_B 0.00611649f $X=8.365 $Y=1.19 $X2=0 $Y2=0
cc_450 N_A_27_47#_c_362_n N_SET_B_c_1354_n 0.0194369f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_363_n N_SET_B_c_1354_n 0.0023248f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_364_n N_SET_B_c_1354_n 0.00534882f $X=8.937 $Y=1.305 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_c_368_n N_SET_B_c_1354_n 0.158094f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_373_n N_SET_B_c_1354_n 0.0254944f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_368_n N_SET_B_c_1355_n 0.0265126f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_368_n N_A_917_47#_M1040_g 0.00187255f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_368_n N_A_917_47#_c_1479_n 0.00397012f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_458 N_A_27_47#_M1044_g N_A_917_47#_c_1490_n 0.0126242f $X=5.075 $Y=0.415
+ $X2=0 $Y2=0
cc_459 N_A_27_47#_c_365_n N_A_917_47#_c_1490_n 0.00725231f $X=5.095 $Y=0.85
+ $X2=0 $Y2=0
cc_460 N_A_27_47#_c_371_n N_A_917_47#_c_1490_n 0.00273619f $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_372_n N_A_917_47#_c_1490_n 0.0119311f $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_375_n N_A_917_47#_c_1490_n 7.57004e-19 $X=5.165 $Y=0.93
+ $X2=0 $Y2=0
cc_463 N_A_27_47#_M1039_g N_A_917_47#_c_1495_n 0.00268255f $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_464 N_A_27_47#_M1039_g N_A_917_47#_c_1485_n 9.15899e-19 $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_465 N_A_27_47#_c_369_n N_A_917_47#_c_1485_n 3.12058e-19 $X=5.385 $Y=1.19
+ $X2=0 $Y2=0
cc_466 N_A_27_47#_c_368_n N_A_917_47#_c_1498_n 3.38709e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_467 N_A_27_47#_M1044_g N_A_917_47#_c_1480_n 0.00143591f $X=5.075 $Y=0.415
+ $X2=0 $Y2=0
cc_468 N_A_27_47#_c_357_n N_A_917_47#_c_1480_n 0.00141498f $X=5.102 $Y=1.245
+ $X2=0 $Y2=0
cc_469 N_A_27_47#_c_368_n N_A_917_47#_c_1480_n 0.015221f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_371_n N_A_917_47#_c_1480_n 0.0143356f $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_c_372_n N_A_917_47#_c_1480_n 0.0184389f $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_375_n N_A_917_47#_c_1480_n 0.00218886f $X=5.165 $Y=0.93
+ $X2=0 $Y2=0
cc_473 N_A_27_47#_c_368_n N_A_917_47#_c_1481_n 0.0396722f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_357_n N_A_917_47#_c_1482_n 0.00270419f $X=5.102 $Y=1.245
+ $X2=0 $Y2=0
cc_475 N_A_27_47#_c_368_n N_A_917_47#_c_1482_n 0.0110709f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_369_n N_A_917_47#_c_1482_n 0.00507004f $X=5.385 $Y=1.19
+ $X2=0 $Y2=0
cc_477 N_A_27_47#_c_372_n N_A_917_47#_c_1482_n 0.00228768f $X=5.24 $Y=0.85 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_368_n N_A_1396_21#_M1032_g 0.00125485f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_479 N_A_27_47#_c_368_n N_A_1396_21#_c_1596_n 0.0122882f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_480 N_A_27_47#_c_364_n N_A_1396_21#_c_1605_n 0.00715591f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_481 N_A_27_47#_c_382_n N_A_1396_21#_c_1605_n 0.0157692f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_482 N_A_27_47#_c_383_n N_A_1396_21#_c_1605_n 0.00190553f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_483 N_A_27_47#_c_368_n N_A_1396_21#_c_1605_n 0.014133f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_c_373_n N_A_1396_21#_c_1605_n 0.027417f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_368_n N_A_1396_21#_c_1606_n 0.0276968f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_486 N_A_27_47#_c_382_n N_A_1396_21#_c_1607_n 0.00264766f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_487 N_A_27_47#_c_368_n N_A_1396_21#_c_1607_n 0.00618009f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_488 N_A_27_47#_c_368_n N_A_1396_21#_c_1597_n 0.00581052f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_489 N_A_27_47#_c_382_n N_A_1887_21#_M1003_g 3.55913e-19 $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_490 N_A_27_47#_M1019_g N_A_1887_21#_M1043_g 0.0155835f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_491 N_A_27_47#_M1019_g N_A_1887_21#_c_1770_n 6.56548e-19 $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_492 N_A_27_47#_c_383_n N_A_1887_21#_c_1770_n 0.00900453f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_493 N_A_27_47#_M1019_g N_A_1714_47#_c_1945_n 0.00935459f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_494 N_A_27_47#_c_382_n N_A_1714_47#_c_1945_n 0.00669245f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_495 N_A_27_47#_c_383_n N_A_1714_47#_c_1945_n 0.0028948f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_496 N_A_27_47#_c_362_n N_A_1714_47#_c_1948_n 0.00390894f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_497 N_A_27_47#_c_363_n N_A_1714_47#_c_1948_n 0.00171906f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_498 N_A_27_47#_c_364_n N_A_1714_47#_c_1948_n 0.00314176f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_499 N_A_27_47#_c_362_n N_A_1714_47#_c_1934_n 0.011772f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_364_n N_A_1714_47#_c_1934_n 0.00837617f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_501 N_A_27_47#_c_373_n N_A_1714_47#_c_1934_n 6.65017e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_502 N_A_27_47#_M1019_g N_A_1714_47#_c_1940_n 0.00655842f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_503 N_A_27_47#_c_382_n N_A_1714_47#_c_1940_n 0.0359925f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_504 N_A_27_47#_c_383_n N_A_1714_47#_c_1940_n 0.0021011f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_505 N_A_27_47#_c_364_n N_A_1714_47#_c_1936_n 0.00588727f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_506 N_A_27_47#_c_382_n N_A_1714_47#_c_1936_n 0.00820582f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_507 N_A_27_47#_c_373_n N_A_1714_47#_c_1936_n 2.68785e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_508 N_A_27_47#_c_381_n N_VPWR_M1025_d 0.00165787f $X=0.605 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_509 N_A_27_47#_M1000_g N_VPWR_c_2121_n 0.00864163f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_c_381_n N_VPWR_c_2121_n 0.0171178f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_c_384_n N_VPWR_c_2121_n 0.0127414f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_512 N_A_27_47#_M1000_g N_VPWR_c_2122_n 0.00232641f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_c_381_n N_VPWR_c_2131_n 0.0018545f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_384_n N_VPWR_c_2131_n 0.0177604f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_515 N_A_27_47#_M1000_g N_VPWR_c_2132_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_M1039_g N_VPWR_c_2134_n 0.00541732f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_M1019_g N_VPWR_c_2135_n 0.00367119f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_518 N_A_27_47#_M1000_g N_VPWR_c_2120_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_519 N_A_27_47#_M1039_g N_VPWR_c_2120_n 0.00628048f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_520 N_A_27_47#_M1019_g N_VPWR_c_2120_n 0.00567418f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_c_381_n N_VPWR_c_2120_n 0.00505319f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_384_n N_VPWR_c_2120_n 0.00954719f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_523 N_A_27_47#_c_365_n N_A_453_47#_c_2328_n 0.00382719f $X=5.095 $Y=0.85
+ $X2=0 $Y2=0
cc_524 N_A_27_47#_c_365_n N_A_453_47#_c_2329_n 0.01951f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_525 N_A_27_47#_c_365_n N_A_453_47#_c_2330_n 0.013739f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_526 N_A_27_47#_c_365_n N_A_453_47#_c_2331_n 0.00505777f $X=5.095 $Y=0.85
+ $X2=0 $Y2=0
cc_527 N_A_27_47#_c_365_n N_A_453_47#_c_2348_n 0.00320961f $X=5.095 $Y=0.85
+ $X2=0 $Y2=0
cc_528 N_A_27_47#_M1039_g N_A_453_47#_c_2349_n 0.00733893f $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_529 N_A_27_47#_c_355_n N_A_453_47#_c_2340_n 0.00733893f $X=4.665 $Y=1.32
+ $X2=0 $Y2=0
cc_530 N_A_27_47#_c_365_n N_A_453_47#_c_2332_n 0.081679f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_531 N_A_27_47#_c_365_n N_A_453_47#_c_2333_n 0.027791f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_532 N_A_27_47#_c_365_n N_A_453_47#_c_2334_n 0.0095442f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_533 N_A_27_47#_c_355_n N_A_453_47#_c_2335_n 0.0012436f $X=4.665 $Y=1.32 $X2=0
+ $Y2=0
cc_534 N_A_27_47#_c_365_n N_A_453_47#_c_2335_n 0.0266185f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_535 N_A_27_47#_c_355_n N_A_453_47#_c_2336_n 6.16568e-19 $X=4.665 $Y=1.32
+ $X2=0 $Y2=0
cc_536 N_A_27_47#_c_365_n N_A_453_47#_c_2336_n 0.00495236f $X=5.095 $Y=0.85
+ $X2=0 $Y2=0
cc_537 N_A_27_47#_c_360_n N_VGND_M1045_d 0.00162876f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_538 N_A_27_47#_M1026_g N_VGND_c_2533_n 0.00789067f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_539 N_A_27_47#_c_360_n N_VGND_c_2533_n 0.0154833f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_540 N_A_27_47#_c_365_n N_VGND_c_2533_n 2.30481e-19 $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_541 N_A_27_47#_c_366_n N_VGND_c_2533_n 0.00116209f $X=0.835 $Y=0.85 $X2=0
+ $Y2=0
cc_542 N_A_27_47#_c_374_n N_VGND_c_2533_n 5.88506e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_543 N_A_27_47#_M1026_g N_VGND_c_2534_n 0.00327532f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_544 N_A_27_47#_c_365_n N_VGND_c_2534_n 0.00456395f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_545 N_A_27_47#_c_365_n N_VGND_c_2535_n 0.00120945f $X=5.095 $Y=0.85 $X2=0
+ $Y2=0
cc_546 N_A_27_47#_c_368_n N_VGND_c_2536_n 0.00147999f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_547 N_A_27_47#_c_358_n N_VGND_c_2537_n 0.00179515f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_548 N_A_27_47#_M1044_g N_VGND_c_2541_n 0.00359964f $X=5.075 $Y=0.415 $X2=0
+ $Y2=0
cc_549 N_A_27_47#_c_358_n N_VGND_c_2545_n 0.00435972f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_550 N_A_27_47#_c_362_n N_VGND_c_2545_n 0.00288727f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_551 N_A_27_47#_c_363_n N_VGND_c_2545_n 2.15978e-19 $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_552 N_A_27_47#_c_359_n N_VGND_c_2547_n 0.0106361f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_553 N_A_27_47#_c_360_n N_VGND_c_2547_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_554 N_A_27_47#_M1026_g N_VGND_c_2548_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_555 N_A_27_47#_M1045_s N_VGND_c_2553_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_556 N_A_27_47#_M1026_g N_VGND_c_2553_n 0.00581646f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_557 N_A_27_47#_M1044_g N_VGND_c_2553_n 0.00578342f $X=5.075 $Y=0.415 $X2=0
+ $Y2=0
cc_558 N_A_27_47#_c_358_n N_VGND_c_2553_n 0.00620849f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_559 N_A_27_47#_c_359_n N_VGND_c_2553_n 0.00898615f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_560 N_A_27_47#_c_360_n N_VGND_c_2553_n 0.00523689f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_561 N_A_27_47#_c_362_n N_VGND_c_2553_n 0.00224883f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_562 N_A_27_47#_c_365_n N_VGND_c_2553_n 0.203023f $X=5.095 $Y=0.85 $X2=0 $Y2=0
cc_563 N_A_27_47#_c_366_n N_VGND_c_2553_n 0.0131302f $X=0.835 $Y=0.85 $X2=0
+ $Y2=0
cc_564 N_A_27_47#_c_371_n N_VGND_c_2553_n 0.0153327f $X=5.24 $Y=0.85 $X2=0 $Y2=0
cc_565 N_SCD_M1033_g N_A_423_315#_c_697_n 0.0310159f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_566 N_SCD_c_646_n N_A_423_315#_c_699_n 0.0310159f $X=1.642 $Y=1.49 $X2=0
+ $Y2=0
cc_567 N_SCD_c_641_n N_SCE_c_804_n 0.0206603f $X=1.83 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_568 N_SCD_c_639_n SCE 6.2958e-19 $X=1.642 $Y=0.88 $X2=0 $Y2=0
cc_569 N_SCD_c_641_n SCE 0.00429052f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_570 N_SCD_c_639_n N_SCE_c_811_n 0.0260921f $X=1.642 $Y=0.88 $X2=0 $Y2=0
cc_571 N_SCD_c_640_n N_SCE_c_811_n 0.0081432f $X=1.642 $Y=1.325 $X2=0 $Y2=0
cc_572 N_SCD_c_639_n N_SCE_c_812_n 0.00125284f $X=1.642 $Y=0.88 $X2=0 $Y2=0
cc_573 N_SCD_c_640_n N_SCE_c_812_n 0.00414815f $X=1.642 $Y=1.325 $X2=0 $Y2=0
cc_574 SCD N_SCE_c_812_n 0.00761429f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_575 N_SCD_c_640_n SCE 0.00345389f $X=1.642 $Y=1.325 $X2=0 $Y2=0
cc_576 SCD SCE 0.0314072f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_577 N_SCD_c_646_n SCE 0.00716905f $X=1.642 $Y=1.49 $X2=0 $Y2=0
cc_578 N_SCD_M1033_g N_A_193_47#_c_989_n 0.00853668f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_579 SCD N_A_193_47#_c_989_n 0.00832905f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_580 N_SCD_c_646_n N_A_193_47#_c_989_n 0.00160021f $X=1.642 $Y=1.49 $X2=0
+ $Y2=0
cc_581 N_SCD_M1033_g N_A_193_47#_c_990_n 9.04442e-19 $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_582 N_SCD_c_639_n N_A_193_47#_c_983_n 0.00526933f $X=1.642 $Y=0.88 $X2=0
+ $Y2=0
cc_583 N_SCD_c_640_n N_A_193_47#_c_983_n 8.79848e-19 $X=1.642 $Y=1.325 $X2=0
+ $Y2=0
cc_584 N_SCD_c_641_n N_A_193_47#_c_983_n 0.00248233f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_585 N_SCD_M1033_g N_A_193_47#_c_983_n 0.00414955f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_586 SCD N_A_193_47#_c_983_n 0.0505612f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_587 N_SCD_c_646_n N_A_193_47#_c_983_n 0.00111321f $X=1.642 $Y=1.49 $X2=0
+ $Y2=0
cc_588 N_SCD_M1033_g N_VPWR_c_2122_n 0.015447f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_589 SCD N_VPWR_c_2122_n 0.0161253f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_590 N_SCD_c_646_n N_VPWR_c_2122_n 0.00306868f $X=1.642 $Y=1.49 $X2=0 $Y2=0
cc_591 N_SCD_M1033_g N_VPWR_c_2133_n 0.00442511f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_592 N_SCD_M1033_g N_VPWR_c_2120_n 0.00418686f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_593 N_SCD_M1033_g N_A_453_47#_c_2338_n 0.00153013f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_594 N_SCD_c_639_n N_VGND_c_2534_n 0.00504501f $X=1.642 $Y=0.88 $X2=0 $Y2=0
cc_595 N_SCD_c_641_n N_VGND_c_2534_n 0.00528037f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_596 SCD N_VGND_c_2534_n 0.00644652f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_597 N_SCD_c_646_n N_VGND_c_2534_n 3.43054e-19 $X=1.642 $Y=1.49 $X2=0 $Y2=0
cc_598 N_SCD_c_639_n N_VGND_c_2549_n 9.17963e-19 $X=1.642 $Y=0.88 $X2=0 $Y2=0
cc_599 N_SCD_c_641_n N_VGND_c_2549_n 0.00585144f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_600 N_SCD_c_639_n N_VGND_c_2553_n 7.68569e-19 $X=1.642 $Y=0.88 $X2=0 $Y2=0
cc_601 N_SCD_c_641_n N_VGND_c_2553_n 0.00755725f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_602 N_A_423_315#_c_698_n N_SCE_c_805_n 0.00544208f $X=2.71 $Y=1.65 $X2=0
+ $Y2=0
cc_603 N_A_423_315#_c_691_n N_SCE_c_805_n 0.0010119f $X=3.43 $Y=0.71 $X2=0 $Y2=0
cc_604 N_A_423_315#_c_692_n N_SCE_c_805_n 0.00582182f $X=3.04 $Y=0.71 $X2=0
+ $Y2=0
cc_605 N_A_423_315#_c_704_n N_SCE_c_805_n 2.44473e-19 $X=2.845 $Y=1.65 $X2=0
+ $Y2=0
cc_606 N_A_423_315#_c_691_n N_SCE_c_806_n 0.00748623f $X=3.43 $Y=0.71 $X2=0
+ $Y2=0
cc_607 N_A_423_315#_c_696_n N_SCE_c_806_n 0.0150386f $X=3.615 $Y=0.765 $X2=0
+ $Y2=0
cc_608 N_A_423_315#_c_694_n N_SCE_c_807_n 0.00144501f $X=3.517 $Y=1.575 $X2=0
+ $Y2=0
cc_609 N_A_423_315#_c_701_n N_SCE_c_814_n 0.0113843f $X=3.43 $Y=1.66 $X2=0 $Y2=0
cc_610 N_A_423_315#_c_703_n N_SCE_c_814_n 0.00376173f $X=3.14 $Y=1.74 $X2=0
+ $Y2=0
cc_611 N_A_423_315#_c_704_n N_SCE_c_814_n 0.0212597f $X=2.845 $Y=1.65 $X2=0
+ $Y2=0
cc_612 N_A_423_315#_c_701_n N_SCE_c_816_n 0.00673533f $X=3.43 $Y=1.66 $X2=0
+ $Y2=0
cc_613 N_A_423_315#_c_691_n N_SCE_c_808_n 0.00503781f $X=3.43 $Y=0.71 $X2=0
+ $Y2=0
cc_614 N_A_423_315#_c_693_n N_SCE_c_808_n 0.0058072f $X=3.517 $Y=1.095 $X2=0
+ $Y2=0
cc_615 N_A_423_315#_c_695_n N_SCE_c_808_n 0.0176611f $X=3.615 $Y=0.93 $X2=0
+ $Y2=0
cc_616 N_A_423_315#_c_691_n N_SCE_c_809_n 0.00179745f $X=3.43 $Y=0.71 $X2=0
+ $Y2=0
cc_617 N_A_423_315#_c_694_n N_SCE_c_809_n 0.0061053f $X=3.517 $Y=1.575 $X2=0
+ $Y2=0
cc_618 N_A_423_315#_c_703_n N_SCE_c_809_n 0.00427623f $X=3.14 $Y=1.74 $X2=0
+ $Y2=0
cc_619 N_A_423_315#_c_700_n N_SCE_c_819_n 0.00719381f $X=3.055 $Y=2.3 $X2=0
+ $Y2=0
cc_620 N_A_423_315#_c_699_n N_SCE_c_811_n 0.00980599f $X=2.265 $Y=1.65 $X2=0
+ $Y2=0
cc_621 N_A_423_315#_c_699_n N_SCE_c_812_n 0.00107361f $X=2.265 $Y=1.65 $X2=0
+ $Y2=0
cc_622 N_A_423_315#_c_699_n SCE 0.00452196f $X=2.265 $Y=1.65 $X2=0 $Y2=0
cc_623 N_A_423_315#_c_693_n N_D_M1027_g 0.00116781f $X=3.517 $Y=1.095 $X2=0
+ $Y2=0
cc_624 N_A_423_315#_c_694_n N_D_M1027_g 0.00156486f $X=3.517 $Y=1.575 $X2=0
+ $Y2=0
cc_625 N_A_423_315#_c_695_n N_D_M1027_g 0.0212986f $X=3.615 $Y=0.93 $X2=0 $Y2=0
cc_626 N_A_423_315#_c_696_n N_D_M1027_g 0.0279761f $X=3.615 $Y=0.765 $X2=0 $Y2=0
cc_627 N_A_423_315#_c_701_n N_D_M1017_g 3.77634e-19 $X=3.43 $Y=1.66 $X2=0 $Y2=0
cc_628 N_A_423_315#_c_701_n D 0.00500934f $X=3.43 $Y=1.66 $X2=0 $Y2=0
cc_629 N_A_423_315#_c_701_n N_D_c_923_n 2.21976e-19 $X=3.43 $Y=1.66 $X2=0 $Y2=0
cc_630 N_A_423_315#_c_694_n N_D_c_923_n 0.00127508f $X=3.517 $Y=1.575 $X2=0
+ $Y2=0
cc_631 N_A_423_315#_c_701_n N_D_c_924_n 0.00859304f $X=3.43 $Y=1.66 $X2=0 $Y2=0
cc_632 N_A_423_315#_c_694_n N_D_c_924_n 0.0128301f $X=3.517 $Y=1.575 $X2=0 $Y2=0
cc_633 N_A_423_315#_c_697_n N_A_193_47#_c_989_n 0.00680134f $X=2.19 $Y=1.725
+ $X2=0 $Y2=0
cc_634 N_A_423_315#_c_698_n N_A_193_47#_c_989_n 0.00618502f $X=2.71 $Y=1.65
+ $X2=0 $Y2=0
cc_635 N_A_423_315#_c_700_n N_A_193_47#_c_989_n 0.00727137f $X=3.055 $Y=2.3
+ $X2=0 $Y2=0
cc_636 N_A_423_315#_c_701_n N_A_193_47#_c_989_n 0.0112091f $X=3.43 $Y=1.66 $X2=0
+ $Y2=0
cc_637 N_A_423_315#_c_703_n N_A_193_47#_c_989_n 0.0189992f $X=3.14 $Y=1.74 $X2=0
+ $Y2=0
cc_638 N_A_423_315#_c_704_n N_A_193_47#_c_989_n 0.00366084f $X=2.845 $Y=1.65
+ $X2=0 $Y2=0
cc_639 N_A_423_315#_c_697_n N_VPWR_c_2122_n 0.00275879f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_640 N_A_423_315#_c_701_n N_VPWR_c_2123_n 0.00443397f $X=3.43 $Y=1.66 $X2=0
+ $Y2=0
cc_641 N_A_423_315#_c_697_n N_VPWR_c_2133_n 0.00489197f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_642 N_A_423_315#_c_700_n N_VPWR_c_2133_n 0.0114446f $X=3.055 $Y=2.3 $X2=0
+ $Y2=0
cc_643 N_A_423_315#_M1034_s N_VPWR_c_2120_n 0.00224156f $X=2.93 $Y=2.065 $X2=0
+ $Y2=0
cc_644 N_A_423_315#_c_697_n N_VPWR_c_2120_n 0.00669614f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_645 N_A_423_315#_c_700_n N_VPWR_c_2120_n 0.00304943f $X=3.055 $Y=2.3 $X2=0
+ $Y2=0
cc_646 N_A_423_315#_c_703_n N_VPWR_c_2120_n 0.00278709f $X=3.14 $Y=1.74 $X2=0
+ $Y2=0
cc_647 N_A_423_315#_c_704_n N_VPWR_c_2120_n 0.0015002f $X=2.845 $Y=1.65 $X2=0
+ $Y2=0
cc_648 N_A_423_315#_c_698_n N_A_453_47#_c_2328_n 0.00314428f $X=2.71 $Y=1.65
+ $X2=0 $Y2=0
cc_649 N_A_423_315#_c_757_p N_A_453_47#_c_2329_n 0.00184347f $X=2.955 $Y=0.47
+ $X2=0 $Y2=0
cc_650 N_A_423_315#_c_692_n N_A_453_47#_c_2329_n 0.0114152f $X=3.04 $Y=0.71
+ $X2=0 $Y2=0
cc_651 N_A_423_315#_c_693_n N_A_453_47#_c_2330_n 0.0286058f $X=3.517 $Y=1.095
+ $X2=0 $Y2=0
cc_652 N_A_423_315#_c_695_n N_A_453_47#_c_2330_n 8.18104e-19 $X=3.615 $Y=0.93
+ $X2=0 $Y2=0
cc_653 N_A_423_315#_c_696_n N_A_453_47#_c_2330_n 8.00641e-19 $X=3.615 $Y=0.765
+ $X2=0 $Y2=0
cc_654 N_A_423_315#_c_697_n N_A_453_47#_c_2338_n 0.0101367f $X=2.19 $Y=1.725
+ $X2=0 $Y2=0
cc_655 N_A_423_315#_c_698_n N_A_453_47#_c_2338_n 0.00422041f $X=2.71 $Y=1.65
+ $X2=0 $Y2=0
cc_656 N_A_423_315#_c_700_n N_A_453_47#_c_2338_n 0.0204236f $X=3.055 $Y=2.3
+ $X2=0 $Y2=0
cc_657 N_A_423_315#_c_697_n N_A_453_47#_c_2339_n 0.00286335f $X=2.19 $Y=1.725
+ $X2=0 $Y2=0
cc_658 N_A_423_315#_c_698_n N_A_453_47#_c_2339_n 0.0142188f $X=2.71 $Y=1.65
+ $X2=0 $Y2=0
cc_659 N_A_423_315#_c_703_n N_A_453_47#_c_2339_n 0.0225306f $X=3.14 $Y=1.74
+ $X2=0 $Y2=0
cc_660 N_A_423_315#_c_704_n N_A_453_47#_c_2339_n 0.0013702f $X=2.845 $Y=1.65
+ $X2=0 $Y2=0
cc_661 N_A_423_315#_c_757_p N_A_453_47#_c_2331_n 0.0191025f $X=2.955 $Y=0.47
+ $X2=0 $Y2=0
cc_662 N_A_423_315#_c_694_n N_A_453_47#_c_2340_n 0.00283705f $X=3.517 $Y=1.575
+ $X2=0 $Y2=0
cc_663 N_A_423_315#_c_691_n N_A_453_47#_c_2332_n 0.00227496f $X=3.43 $Y=0.71
+ $X2=0 $Y2=0
cc_664 N_A_423_315#_c_693_n N_A_453_47#_c_2332_n 0.0052838f $X=3.517 $Y=1.095
+ $X2=0 $Y2=0
cc_665 N_A_423_315#_c_694_n N_A_453_47#_c_2332_n 0.0152158f $X=3.517 $Y=1.575
+ $X2=0 $Y2=0
cc_666 N_A_423_315#_c_703_n N_A_453_47#_c_2332_n 0.00687783f $X=3.14 $Y=1.74
+ $X2=0 $Y2=0
cc_667 N_A_423_315#_c_691_n N_A_453_47#_c_2333_n 8.72827e-19 $X=3.43 $Y=0.71
+ $X2=0 $Y2=0
cc_668 N_A_423_315#_c_692_n N_A_453_47#_c_2333_n 7.72628e-19 $X=3.04 $Y=0.71
+ $X2=0 $Y2=0
cc_669 N_A_423_315#_c_693_n N_A_453_47#_c_2333_n 4.99861e-19 $X=3.517 $Y=1.095
+ $X2=0 $Y2=0
cc_670 N_A_423_315#_c_694_n N_A_453_47#_c_2333_n 0.00163519f $X=3.517 $Y=1.575
+ $X2=0 $Y2=0
cc_671 N_A_423_315#_c_703_n N_A_453_47#_c_2333_n 0.00260056f $X=3.14 $Y=1.74
+ $X2=0 $Y2=0
cc_672 N_A_423_315#_c_698_n N_A_453_47#_c_2334_n 0.00470255f $X=2.71 $Y=1.65
+ $X2=0 $Y2=0
cc_673 N_A_423_315#_c_691_n N_A_453_47#_c_2334_n 0.00139769f $X=3.43 $Y=0.71
+ $X2=0 $Y2=0
cc_674 N_A_423_315#_c_692_n N_A_453_47#_c_2334_n 0.00693312f $X=3.04 $Y=0.71
+ $X2=0 $Y2=0
cc_675 N_A_423_315#_c_693_n N_A_453_47#_c_2334_n 6.30058e-19 $X=3.517 $Y=1.095
+ $X2=0 $Y2=0
cc_676 N_A_423_315#_c_694_n N_A_453_47#_c_2334_n 0.0120352f $X=3.517 $Y=1.575
+ $X2=0 $Y2=0
cc_677 N_A_423_315#_c_703_n N_A_453_47#_c_2334_n 0.022707f $X=3.14 $Y=1.74 $X2=0
+ $Y2=0
cc_678 N_A_423_315#_c_694_n N_A_453_47#_c_2335_n 0.00113041f $X=3.517 $Y=1.575
+ $X2=0 $Y2=0
cc_679 N_A_423_315#_c_693_n N_A_453_47#_c_2336_n 0.00239251f $X=3.517 $Y=1.095
+ $X2=0 $Y2=0
cc_680 N_A_423_315#_c_694_n N_A_453_47#_c_2336_n 0.00632144f $X=3.517 $Y=1.575
+ $X2=0 $Y2=0
cc_681 N_A_423_315#_c_691_n N_VGND_M1041_d 0.00137857f $X=3.43 $Y=0.71 $X2=0
+ $Y2=0
cc_682 N_A_423_315#_c_693_n N_VGND_M1041_d 4.13197e-19 $X=3.517 $Y=1.095 $X2=0
+ $Y2=0
cc_683 N_A_423_315#_c_691_n N_VGND_c_2535_n 0.00965906f $X=3.43 $Y=0.71 $X2=0
+ $Y2=0
cc_684 N_A_423_315#_c_693_n N_VGND_c_2535_n 0.00479139f $X=3.517 $Y=1.095 $X2=0
+ $Y2=0
cc_685 N_A_423_315#_c_696_n N_VGND_c_2535_n 0.00923099f $X=3.615 $Y=0.765 $X2=0
+ $Y2=0
cc_686 N_A_423_315#_c_693_n N_VGND_c_2541_n 0.00162619f $X=3.517 $Y=1.095 $X2=0
+ $Y2=0
cc_687 N_A_423_315#_c_695_n N_VGND_c_2541_n 5.44271e-19 $X=3.615 $Y=0.93 $X2=0
+ $Y2=0
cc_688 N_A_423_315#_c_696_n N_VGND_c_2541_n 0.00370456f $X=3.615 $Y=0.765 $X2=0
+ $Y2=0
cc_689 N_A_423_315#_c_757_p N_VGND_c_2549_n 0.00857854f $X=2.955 $Y=0.47 $X2=0
+ $Y2=0
cc_690 N_A_423_315#_c_691_n N_VGND_c_2549_n 0.00274687f $X=3.43 $Y=0.71 $X2=0
+ $Y2=0
cc_691 N_A_423_315#_M1041_s N_VGND_c_2553_n 0.00206506f $X=2.83 $Y=0.235 $X2=0
+ $Y2=0
cc_692 N_A_423_315#_c_757_p N_VGND_c_2553_n 0.00294183f $X=2.955 $Y=0.47 $X2=0
+ $Y2=0
cc_693 N_A_423_315#_c_691_n N_VGND_c_2553_n 0.00256363f $X=3.43 $Y=0.71 $X2=0
+ $Y2=0
cc_694 N_A_423_315#_c_693_n N_VGND_c_2553_n 0.00409914f $X=3.517 $Y=1.095 $X2=0
+ $Y2=0
cc_695 N_A_423_315#_c_696_n N_VGND_c_2553_n 0.0038579f $X=3.615 $Y=0.765 $X2=0
+ $Y2=0
cc_696 N_SCE_c_807_n N_D_M1027_g 0.00182482f $X=3.165 $Y=1.255 $X2=0 $Y2=0
cc_697 N_SCE_c_809_n N_D_M1027_g 0.00117503f $X=3.265 $Y=1.33 $X2=0 $Y2=0
cc_698 N_SCE_c_814_n N_D_M1017_g 0.00220726f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_699 N_SCE_c_816_n N_D_M1017_g 0.0354143f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_700 N_SCE_c_814_n D 0.00151478f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_701 N_SCE_c_816_n D 0.0102805f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_702 N_SCE_c_809_n N_D_c_923_n 0.00587231f $X=3.265 $Y=1.33 $X2=0 $Y2=0
cc_703 N_SCE_c_814_n N_D_c_924_n 2.11412e-19 $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_704 N_SCE_c_814_n N_A_193_47#_c_989_n 0.00200713f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_705 N_SCE_c_816_n N_A_193_47#_c_989_n 0.0105806f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_706 N_SCE_c_819_n N_A_193_47#_c_989_n 0.00368443f $X=3.265 $Y=1.91 $X2=0
+ $Y2=0
cc_707 SCE N_A_193_47#_c_989_n 0.0116705f $X=2.07 $Y=1.19 $X2=0 $Y2=0
cc_708 N_SCE_c_815_n N_VPWR_c_2123_n 0.00905101f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_709 N_SCE_c_816_n N_VPWR_c_2123_n 0.00200263f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_710 N_SCE_c_817_n N_VPWR_c_2123_n 0.0091805f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_711 N_SCE_c_815_n N_VPWR_c_2133_n 0.0046653f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_712 N_SCE_c_817_n N_VPWR_c_2134_n 0.0046653f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_713 N_SCE_c_815_n N_VPWR_c_2120_n 0.00571875f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_714 N_SCE_c_817_n N_VPWR_c_2120_n 0.00446764f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_715 N_SCE_c_805_n N_A_453_47#_c_2328_n 3.82858e-19 $X=3.09 $Y=0.81 $X2=0
+ $Y2=0
cc_716 N_SCE_c_814_n N_A_453_47#_c_2328_n 0.00235072f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_717 N_SCE_c_811_n N_A_453_47#_c_2328_n 0.00100604f $X=2.242 $Y=0.81 $X2=0
+ $Y2=0
cc_718 N_SCE_c_812_n N_A_453_47#_c_2328_n 0.00608482f $X=2.23 $Y=0.985 $X2=0
+ $Y2=0
cc_719 SCE N_A_453_47#_c_2328_n 0.0211215f $X=2.07 $Y=1.19 $X2=0 $Y2=0
cc_720 N_SCE_c_804_n N_A_453_47#_c_2329_n 0.00225228f $X=2.19 $Y=0.735 $X2=0
+ $Y2=0
cc_721 N_SCE_c_805_n N_A_453_47#_c_2329_n 0.0133761f $X=3.09 $Y=0.81 $X2=0 $Y2=0
cc_722 N_SCE_c_806_n N_A_453_47#_c_2329_n 3.86943e-19 $X=3.165 $Y=0.735 $X2=0
+ $Y2=0
cc_723 N_SCE_c_807_n N_A_453_47#_c_2329_n 0.00311676f $X=3.165 $Y=1.255 $X2=0
+ $Y2=0
cc_724 SCE N_A_453_47#_c_2329_n 0.00899145f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_725 N_SCE_c_811_n N_A_453_47#_c_2329_n 0.00223737f $X=2.242 $Y=0.81 $X2=0
+ $Y2=0
cc_726 N_SCE_c_812_n N_A_453_47#_c_2329_n 0.0187098f $X=2.23 $Y=0.985 $X2=0
+ $Y2=0
cc_727 N_SCE_c_814_n N_A_453_47#_c_2338_n 0.00117937f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_728 N_SCE_c_814_n N_A_453_47#_c_2339_n 0.00155912f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_729 SCE N_A_453_47#_c_2339_n 0.0101785f $X=2.07 $Y=1.19 $X2=0 $Y2=0
cc_730 N_SCE_c_805_n N_A_453_47#_c_2331_n 9.34339e-19 $X=3.09 $Y=0.81 $X2=0
+ $Y2=0
cc_731 N_SCE_c_806_n N_A_453_47#_c_2331_n 8.53191e-19 $X=3.165 $Y=0.735 $X2=0
+ $Y2=0
cc_732 SCE N_A_453_47#_c_2331_n 0.0188601f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_733 N_SCE_c_811_n N_A_453_47#_c_2331_n 0.00554806f $X=2.242 $Y=0.81 $X2=0
+ $Y2=0
cc_734 N_SCE_c_807_n N_A_453_47#_c_2332_n 0.00270498f $X=3.165 $Y=1.255 $X2=0
+ $Y2=0
cc_735 N_SCE_c_816_n N_A_453_47#_c_2332_n 7.55221e-19 $X=3.61 $Y=1.91 $X2=0
+ $Y2=0
cc_736 N_SCE_c_809_n N_A_453_47#_c_2332_n 0.00304813f $X=3.265 $Y=1.33 $X2=0
+ $Y2=0
cc_737 N_SCE_c_805_n N_A_453_47#_c_2333_n 4.90637e-19 $X=3.09 $Y=0.81 $X2=0
+ $Y2=0
cc_738 N_SCE_c_807_n N_A_453_47#_c_2333_n 0.00243077f $X=3.165 $Y=1.255 $X2=0
+ $Y2=0
cc_739 N_SCE_c_809_n N_A_453_47#_c_2333_n 0.00129524f $X=3.265 $Y=1.33 $X2=0
+ $Y2=0
cc_740 N_SCE_c_812_n N_A_453_47#_c_2333_n 2.5364e-19 $X=2.23 $Y=0.985 $X2=0
+ $Y2=0
cc_741 N_SCE_c_805_n N_A_453_47#_c_2334_n 0.00608267f $X=3.09 $Y=0.81 $X2=0
+ $Y2=0
cc_742 N_SCE_c_807_n N_A_453_47#_c_2334_n 0.00777503f $X=3.165 $Y=1.255 $X2=0
+ $Y2=0
cc_743 N_SCE_c_806_n N_VGND_c_2535_n 0.00809491f $X=3.165 $Y=0.735 $X2=0 $Y2=0
cc_744 N_SCE_c_804_n N_VGND_c_2549_n 0.00530891f $X=2.19 $Y=0.735 $X2=0 $Y2=0
cc_745 N_SCE_c_805_n N_VGND_c_2549_n 0.00380949f $X=3.09 $Y=0.81 $X2=0 $Y2=0
cc_746 N_SCE_c_806_n N_VGND_c_2549_n 0.0038055f $X=3.165 $Y=0.735 $X2=0 $Y2=0
cc_747 SCE N_VGND_c_2549_n 0.0077098f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_748 N_SCE_c_804_n N_VGND_c_2553_n 0.00682761f $X=2.19 $Y=0.735 $X2=0 $Y2=0
cc_749 N_SCE_c_805_n N_VGND_c_2553_n 0.00266575f $X=3.09 $Y=0.81 $X2=0 $Y2=0
cc_750 N_SCE_c_806_n N_VGND_c_2553_n 0.00553323f $X=3.165 $Y=0.735 $X2=0 $Y2=0
cc_751 SCE N_VGND_c_2553_n 0.00362007f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_752 N_SCE_c_812_n N_VGND_c_2553_n 0.00202853f $X=2.23 $Y=0.985 $X2=0 $Y2=0
cc_753 SCE A_381_47# 0.00111667f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_754 N_D_M1027_g N_A_193_47#_c_976_n 0.0217263f $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_755 N_D_M1027_g N_A_193_47#_c_980_n 0.00105567f $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_756 N_D_M1027_g N_A_193_47#_c_981_n 4.84984e-19 $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_757 N_D_M1017_g N_A_193_47#_c_989_n 0.00431782f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_758 D N_A_193_47#_c_989_n 0.0220131f $X=3.825 $Y=2.125 $X2=0 $Y2=0
cc_759 N_D_c_924_n N_A_193_47#_c_989_n 0.00282913f $X=3.942 $Y=1.675 $X2=0 $Y2=0
cc_760 N_D_M1017_g N_VPWR_c_2123_n 0.00153679f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_761 D N_VPWR_c_2123_n 0.0113378f $X=3.825 $Y=2.125 $X2=0 $Y2=0
cc_762 N_D_M1017_g N_VPWR_c_2134_n 0.00544863f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_763 D N_VPWR_c_2134_n 0.00908856f $X=3.825 $Y=2.125 $X2=0 $Y2=0
cc_764 N_D_M1017_g N_VPWR_c_2120_n 0.00636867f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_765 D N_VPWR_c_2120_n 0.00400058f $X=3.825 $Y=2.125 $X2=0 $Y2=0
cc_766 N_D_M1027_g N_A_453_47#_c_2330_n 0.0103334f $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_767 N_D_M1027_g N_A_453_47#_c_2348_n 0.00528745f $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_768 N_D_M1027_g N_A_453_47#_c_2340_n 5.80007e-19 $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_769 D N_A_453_47#_c_2340_n 0.026929f $X=3.825 $Y=2.125 $X2=0 $Y2=0
cc_770 N_D_c_923_n N_A_453_47#_c_2340_n 0.00613845f $X=4.105 $Y=1.49 $X2=0 $Y2=0
cc_771 N_D_c_924_n N_A_453_47#_c_2340_n 0.0190643f $X=3.942 $Y=1.675 $X2=0 $Y2=0
cc_772 N_D_M1027_g N_A_453_47#_c_2332_n 0.001745f $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_773 N_D_c_923_n N_A_453_47#_c_2332_n 0.00455589f $X=4.105 $Y=1.49 $X2=0 $Y2=0
cc_774 N_D_c_924_n N_A_453_47#_c_2332_n 0.00746689f $X=3.942 $Y=1.675 $X2=0
+ $Y2=0
cc_775 N_D_M1027_g N_A_453_47#_c_2335_n 7.84718e-19 $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_776 N_D_c_923_n N_A_453_47#_c_2335_n 2.33386e-19 $X=4.105 $Y=1.49 $X2=0 $Y2=0
cc_777 N_D_M1027_g N_A_453_47#_c_2336_n 0.00937505f $X=4.035 $Y=0.445 $X2=0
+ $Y2=0
cc_778 N_D_c_923_n N_A_453_47#_c_2336_n 0.00309445f $X=4.105 $Y=1.49 $X2=0 $Y2=0
cc_779 N_D_c_924_n N_A_453_47#_c_2336_n 0.0101861f $X=3.942 $Y=1.675 $X2=0 $Y2=0
cc_780 D A_752_413# 0.00521948f $X=3.825 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_781 N_D_M1027_g N_VGND_c_2535_n 0.00167941f $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_782 N_D_M1027_g N_VGND_c_2541_n 0.00390689f $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_783 N_D_M1027_g N_VGND_c_2553_n 0.00551104f $X=4.035 $Y=0.445 $X2=0 $Y2=0
cc_784 N_A_193_47#_M1011_g N_A_1102_21#_M1035_g 0.0154054f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_785 N_A_193_47#_c_991_n N_A_1102_21#_M1035_g 0.00197541f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_786 N_A_193_47#_M1031_g N_A_1102_21#_M1047_g 0.0164618f $X=8.505 $Y=2.275
+ $X2=0 $Y2=0
cc_787 N_A_193_47#_c_978_n N_A_1102_21#_M1047_g 0.00557814f $X=8.58 $Y=1.32
+ $X2=0 $Y2=0
cc_788 N_A_193_47#_c_991_n N_A_1102_21#_M1047_g 0.00750594f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_789 N_A_193_47#_c_996_n N_A_1102_21#_M1047_g 0.00910409f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_790 N_A_193_47#_c_997_n N_A_1102_21#_M1047_g 0.00264318f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_791 N_A_193_47#_c_991_n N_A_1102_21#_c_1211_n 0.0240118f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_792 N_A_193_47#_c_991_n N_A_1102_21#_c_1223_n 0.0279826f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_793 N_A_193_47#_c_991_n N_A_1102_21#_c_1213_n 0.0141612f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_794 N_A_193_47#_M1011_g N_A_1102_21#_c_1214_n 8.43685e-19 $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_795 N_A_193_47#_c_991_n N_A_1102_21#_c_1214_n 0.00238493f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_796 N_A_193_47#_c_994_n N_A_1102_21#_c_1214_n 0.0103483f $X=5.04 $Y=1.74
+ $X2=0 $Y2=0
cc_797 N_A_193_47#_c_991_n N_A_1102_21#_c_1228_n 0.00959465f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_798 N_A_193_47#_c_978_n N_A_1102_21#_c_1207_n 0.0027239f $X=8.58 $Y=1.32
+ $X2=0 $Y2=0
cc_799 N_A_193_47#_M1024_g N_SET_B_c_1354_n 0.00574114f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_800 N_A_193_47#_c_976_n N_A_917_47#_c_1490_n 0.00309756f $X=4.51 $Y=0.705
+ $X2=0 $Y2=0
cc_801 N_A_193_47#_c_981_n N_A_917_47#_c_1490_n 0.00920514f $X=4.655 $Y=0.87
+ $X2=0 $Y2=0
cc_802 N_A_193_47#_c_982_n N_A_917_47#_c_1490_n 0.00120295f $X=4.655 $Y=0.87
+ $X2=0 $Y2=0
cc_803 N_A_193_47#_M1011_g N_A_917_47#_c_1495_n 0.0091014f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_804 N_A_193_47#_c_989_n N_A_917_47#_c_1495_n 2.09728e-19 $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_805 N_A_193_47#_c_991_n N_A_917_47#_c_1495_n 0.00506942f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_806 N_A_193_47#_c_992_n N_A_917_47#_c_1495_n 0.00303545f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_807 N_A_193_47#_c_994_n N_A_917_47#_c_1495_n 0.00186639f $X=5.04 $Y=1.74
+ $X2=0 $Y2=0
cc_808 N_A_193_47#_c_995_n N_A_917_47#_c_1495_n 0.0152514f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_809 N_A_193_47#_M1011_g N_A_917_47#_c_1485_n 0.0065077f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_810 N_A_193_47#_c_980_n N_A_917_47#_c_1485_n 0.0060387f $X=4.702 $Y=1.575
+ $X2=0 $Y2=0
cc_811 N_A_193_47#_c_991_n N_A_917_47#_c_1485_n 0.013911f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_812 N_A_193_47#_c_992_n N_A_917_47#_c_1485_n 0.00149623f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_813 N_A_193_47#_c_994_n N_A_917_47#_c_1485_n 0.00193983f $X=5.04 $Y=1.74
+ $X2=0 $Y2=0
cc_814 N_A_193_47#_c_995_n N_A_917_47#_c_1485_n 0.0283189f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_815 N_A_193_47#_c_991_n N_A_917_47#_c_1481_n 0.00350894f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_816 N_A_193_47#_c_980_n N_A_917_47#_c_1482_n 0.00648296f $X=4.702 $Y=1.575
+ $X2=0 $Y2=0
cc_817 N_A_193_47#_c_991_n N_A_917_47#_c_1482_n 0.00445486f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_818 N_A_193_47#_c_991_n N_A_1396_21#_M1030_g 0.00576309f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_819 N_A_193_47#_c_991_n N_A_1396_21#_c_1596_n 0.00477237f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_820 N_A_193_47#_c_977_n N_A_1396_21#_c_1605_n 0.00385681f $X=8.96 $Y=1.32
+ $X2=0 $Y2=0
cc_821 N_A_193_47#_c_991_n N_A_1396_21#_c_1605_n 0.0139809f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_822 N_A_193_47#_c_993_n N_A_1396_21#_c_1605_n 0.0255925f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_823 N_A_193_47#_c_996_n N_A_1396_21#_c_1605_n 0.00176885f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_824 N_A_193_47#_c_997_n N_A_1396_21#_c_1605_n 0.00661378f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_825 N_A_193_47#_c_998_n N_A_1396_21#_c_1605_n 0.00371524f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_826 N_A_193_47#_c_991_n N_A_1396_21#_c_1606_n 0.0264578f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_827 N_A_193_47#_c_996_n N_A_1396_21#_c_1606_n 7.96394e-19 $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_828 N_A_193_47#_c_997_n N_A_1396_21#_c_1606_n 0.00130051f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_829 N_A_193_47#_c_998_n N_A_1396_21#_c_1606_n 7.27878e-19 $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_830 N_A_193_47#_c_991_n N_A_1396_21#_c_1607_n 0.020032f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_831 N_A_193_47#_c_996_n N_A_1396_21#_c_1607_n 6.45403e-19 $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_832 N_A_193_47#_c_997_n N_A_1396_21#_c_1607_n 0.00461622f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_833 N_A_193_47#_c_998_n N_A_1396_21#_c_1607_n 0.00148716f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_834 N_A_193_47#_c_991_n N_A_1396_21#_c_1597_n 6.72943e-19 $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_835 N_A_193_47#_M1024_g N_A_1887_21#_M1003_g 0.0428093f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_836 N_A_193_47#_M1031_g N_A_1714_47#_c_1945_n 0.00496872f $X=8.505 $Y=2.275
+ $X2=0 $Y2=0
cc_837 N_A_193_47#_c_993_n N_A_1714_47#_c_1945_n 0.00187313f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_838 N_A_193_47#_c_997_n N_A_1714_47#_c_1945_n 0.00141396f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_839 N_A_193_47#_M1024_g N_A_1714_47#_c_1948_n 0.00969843f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_840 N_A_193_47#_M1024_g N_A_1714_47#_c_1934_n 0.0106063f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_841 N_A_193_47#_c_993_n N_A_1714_47#_c_1940_n 0.00214622f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_842 N_A_193_47#_c_997_n N_A_1714_47#_c_1940_n 0.0013353f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_843 N_A_193_47#_M1024_g N_A_1714_47#_c_1936_n 0.00155103f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_844 N_A_193_47#_c_991_n N_VPWR_M1030_d 0.00670518f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_845 N_A_193_47#_c_983_n N_VPWR_c_2121_n 0.0127345f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_846 N_A_193_47#_c_989_n N_VPWR_c_2122_n 0.0169174f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_847 N_A_193_47#_c_990_n N_VPWR_c_2122_n 0.00138261f $X=1.295 $Y=1.87 $X2=0
+ $Y2=0
cc_848 N_A_193_47#_c_983_n N_VPWR_c_2122_n 0.0415488f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_849 N_A_193_47#_c_989_n N_VPWR_c_2123_n 0.00464499f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_850 N_A_193_47#_c_991_n N_VPWR_c_2124_n 0.00160449f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_851 N_A_193_47#_c_991_n N_VPWR_c_2125_n 0.0137399f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_852 N_A_193_47#_c_983_n N_VPWR_c_2132_n 0.0156296f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_853 N_A_193_47#_M1011_g N_VPWR_c_2134_n 0.00367119f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_854 N_A_193_47#_M1031_g N_VPWR_c_2135_n 0.00424681f $X=8.505 $Y=2.275 $X2=0
+ $Y2=0
cc_855 N_A_193_47#_c_997_n N_VPWR_c_2135_n 0.00254851f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_856 N_A_193_47#_M1011_g N_VPWR_c_2120_n 0.00562272f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_857 N_A_193_47#_M1031_g N_VPWR_c_2120_n 0.0061745f $X=8.505 $Y=2.275 $X2=0
+ $Y2=0
cc_858 N_A_193_47#_c_989_n N_VPWR_c_2120_n 0.162881f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_859 N_A_193_47#_c_990_n N_VPWR_c_2120_n 0.0151864f $X=1.295 $Y=1.87 $X2=0
+ $Y2=0
cc_860 N_A_193_47#_c_991_n N_VPWR_c_2120_n 0.159156f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_861 N_A_193_47#_c_992_n N_VPWR_c_2120_n 0.0160117f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_862 N_A_193_47#_c_993_n N_VPWR_c_2120_n 0.0148451f $X=8.51 $Y=1.87 $X2=0
+ $Y2=0
cc_863 N_A_193_47#_c_995_n N_VPWR_c_2120_n 5.19592e-19 $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_864 N_A_193_47#_c_996_n N_VPWR_c_2120_n 3.05853e-19 $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_865 N_A_193_47#_c_997_n N_VPWR_c_2120_n 0.00131252f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_866 N_A_193_47#_c_983_n N_VPWR_c_2120_n 0.00381175f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_867 N_A_193_47#_c_989_n A_381_363# 0.00298073f $X=4.685 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_868 N_A_193_47#_c_989_n N_A_453_47#_c_2328_n 0.00420567f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_869 N_A_193_47#_c_976_n N_A_453_47#_c_2330_n 0.00289683f $X=4.51 $Y=0.705
+ $X2=0 $Y2=0
cc_870 N_A_193_47#_c_981_n N_A_453_47#_c_2330_n 0.00908369f $X=4.655 $Y=0.87
+ $X2=0 $Y2=0
cc_871 N_A_193_47#_c_989_n N_A_453_47#_c_2338_n 0.0181929f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_872 N_A_193_47#_c_989_n N_A_453_47#_c_2339_n 0.00871274f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_873 N_A_193_47#_c_989_n N_A_453_47#_c_2349_n 0.00145724f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_874 N_A_193_47#_c_980_n N_A_453_47#_c_2340_n 0.0192784f $X=4.702 $Y=1.575
+ $X2=0 $Y2=0
cc_875 N_A_193_47#_c_989_n N_A_453_47#_c_2340_n 0.0150313f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_876 N_A_193_47#_c_992_n N_A_453_47#_c_2340_n 0.00178031f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_877 N_A_193_47#_c_995_n N_A_453_47#_c_2340_n 0.0278139f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_878 N_A_193_47#_c_989_n N_A_453_47#_c_2332_n 0.0467326f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_879 N_A_193_47#_c_989_n N_A_453_47#_c_2333_n 0.0125021f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_880 N_A_193_47#_c_989_n N_A_453_47#_c_2334_n 0.00442222f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_881 N_A_193_47#_c_980_n N_A_453_47#_c_2335_n 0.00738424f $X=4.702 $Y=1.575
+ $X2=0 $Y2=0
cc_882 N_A_193_47#_c_982_n N_A_453_47#_c_2335_n 5.1224e-19 $X=4.655 $Y=0.87
+ $X2=0 $Y2=0
cc_883 N_A_193_47#_c_989_n N_A_453_47#_c_2335_n 0.0134544f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_884 N_A_193_47#_c_980_n N_A_453_47#_c_2336_n 0.0146356f $X=4.702 $Y=1.575
+ $X2=0 $Y2=0
cc_885 N_A_193_47#_c_982_n N_A_453_47#_c_2336_n 4.22252e-19 $X=4.655 $Y=0.87
+ $X2=0 $Y2=0
cc_886 N_A_193_47#_c_989_n N_A_453_47#_c_2336_n 0.00120157f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_887 N_A_193_47#_c_991_n A_1351_329# 0.00101797f $X=8.365 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_888 N_A_193_47#_c_991_n A_1572_329# 0.00532504f $X=8.365 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_889 N_A_193_47#_c_983_n N_VGND_c_2534_n 0.0209768f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_890 N_A_193_47#_M1024_g N_VGND_c_2538_n 0.00124887f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_891 N_A_193_47#_c_976_n N_VGND_c_2541_n 0.00540301f $X=4.51 $Y=0.705 $X2=0
+ $Y2=0
cc_892 N_A_193_47#_M1024_g N_VGND_c_2545_n 0.00359964f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_893 N_A_193_47#_c_983_n N_VGND_c_2548_n 0.00955835f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_894 N_A_193_47#_M1026_d N_VGND_c_2553_n 0.00217251f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_895 N_A_193_47#_c_976_n N_VGND_c_2553_n 0.00660662f $X=4.51 $Y=0.705 $X2=0
+ $Y2=0
cc_896 N_A_193_47#_M1024_g N_VGND_c_2553_n 0.00563077f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_897 N_A_193_47#_c_983_n N_VGND_c_2553_n 0.0038044f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_898 N_A_1102_21#_M1009_g N_SET_B_M1004_g 0.0153299f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_899 N_A_1102_21#_c_1203_n N_SET_B_M1004_g 6.39023e-19 $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_900 N_A_1102_21#_M1009_g N_SET_B_c_1349_n 0.0213009f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_901 N_A_1102_21#_M1009_g N_SET_B_M1012_g 0.0127011f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_902 N_A_1102_21#_M1035_g N_SET_B_M1012_g 0.0101628f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_903 N_A_1102_21#_c_1211_n N_SET_B_M1012_g 0.0159332f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_904 N_A_1102_21#_c_1260_p N_SET_B_M1012_g 0.00507112f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_905 N_A_1102_21#_c_1213_n N_SET_B_M1012_g 0.00473578f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_906 N_A_1102_21#_c_1214_n N_SET_B_M1012_g 0.0201903f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_907 N_A_1102_21#_M1009_g SET_B 6.3543e-19 $X=5.585 $Y=0.445 $X2=0 $Y2=0
cc_908 N_A_1102_21#_c_1203_n SET_B 0.00891484f $X=6.9 $Y=1.065 $X2=0 $Y2=0
cc_909 N_A_1102_21#_c_1202_n N_SET_B_c_1354_n 0.00496686f $X=7.995 $Y=0.985
+ $X2=0 $Y2=0
cc_910 N_A_1102_21#_c_1203_n N_SET_B_c_1354_n 0.0207759f $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_911 N_A_1102_21#_c_1205_n N_SET_B_c_1354_n 0.0220549f $X=7.795 $Y=0.98 $X2=0
+ $Y2=0
cc_912 N_A_1102_21#_c_1206_n N_SET_B_c_1354_n 0.0111147f $X=7.96 $Y=0.98 $X2=0
+ $Y2=0
cc_913 N_A_1102_21#_c_1203_n N_SET_B_c_1355_n 0.00235101f $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_914 N_A_1102_21#_c_1203_n N_A_917_47#_M1040_g 0.0071865f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_915 N_A_1102_21#_c_1204_n N_A_917_47#_M1040_g 0.00316772f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_916 N_A_1102_21#_c_1203_n N_A_917_47#_c_1479_n 8.58646e-19 $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_917 N_A_1102_21#_c_1204_n N_A_917_47#_c_1479_n 0.00795872f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_918 N_A_1102_21#_c_1228_n N_A_917_47#_c_1479_n 9.09922e-19 $X=6.47 $Y=1.87
+ $X2=0 $Y2=0
cc_919 N_A_1102_21#_c_1223_n N_A_917_47#_M1036_g 0.0125726f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_920 N_A_1102_21#_M1035_g N_A_917_47#_c_1495_n 0.00191115f $X=5.61 $Y=2.275
+ $X2=0 $Y2=0
cc_921 N_A_1102_21#_M1009_g N_A_917_47#_c_1485_n 0.00984954f $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_922 N_A_1102_21#_M1035_g N_A_917_47#_c_1485_n 0.00585604f $X=5.61 $Y=2.275
+ $X2=0 $Y2=0
cc_923 N_A_1102_21#_c_1213_n N_A_917_47#_c_1485_n 0.033045f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_924 N_A_1102_21#_M1009_g N_A_917_47#_c_1498_n 0.0131348f $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_925 N_A_1102_21#_M1009_g N_A_917_47#_c_1480_n 0.0106026f $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_926 N_A_1102_21#_c_1211_n N_A_917_47#_c_1481_n 0.0141289f $X=6.385 $Y=1.91
+ $X2=0 $Y2=0
cc_927 N_A_1102_21#_c_1223_n N_A_917_47#_c_1481_n 0.00218253f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_928 N_A_1102_21#_c_1204_n N_A_917_47#_c_1481_n 0.0246735f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_929 N_A_1102_21#_c_1228_n N_A_917_47#_c_1481_n 0.00650509f $X=6.47 $Y=1.87
+ $X2=0 $Y2=0
cc_930 N_A_1102_21#_M1009_g N_A_917_47#_c_1482_n 0.0106844f $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_931 N_A_1102_21#_c_1213_n N_A_917_47#_c_1482_n 0.0170209f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_932 N_A_1102_21#_c_1214_n N_A_917_47#_c_1482_n 0.0013712f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_933 N_A_1102_21#_c_1203_n N_A_1396_21#_M1032_g 0.00918226f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_934 N_A_1102_21#_c_1204_n N_A_1396_21#_M1032_g 0.00343246f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_935 N_A_1102_21#_c_1205_n N_A_1396_21#_M1032_g 0.00932512f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_936 N_A_1102_21#_c_1206_n N_A_1396_21#_M1032_g 0.00133201f $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_937 N_A_1102_21#_c_1207_n N_A_1396_21#_M1032_g 0.00183414f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_938 N_A_1102_21#_M1047_g N_A_1396_21#_M1030_g 0.0153539f $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_939 N_A_1102_21#_c_1223_n N_A_1396_21#_M1030_g 0.00219889f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_940 N_A_1102_21#_M1047_g N_A_1396_21#_c_1596_n 2.86505e-19 $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_941 N_A_1102_21#_c_1204_n N_A_1396_21#_c_1596_n 0.0307647f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_942 N_A_1102_21#_c_1205_n N_A_1396_21#_c_1596_n 0.0205705f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_943 N_A_1102_21#_c_1207_n N_A_1396_21#_c_1596_n 0.00382982f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_944 N_A_1102_21#_c_1206_n N_A_1396_21#_c_1606_n 9.59092e-19 $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_945 N_A_1102_21#_c_1207_n N_A_1396_21#_c_1606_n 0.00358318f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_946 N_A_1102_21#_M1047_g N_A_1396_21#_c_1607_n 0.0143059f $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_947 N_A_1102_21#_c_1205_n N_A_1396_21#_c_1607_n 0.00760725f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_948 N_A_1102_21#_c_1206_n N_A_1396_21#_c_1607_n 0.0207118f $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_949 N_A_1102_21#_c_1207_n N_A_1396_21#_c_1607_n 0.00632961f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_950 N_A_1102_21#_c_1204_n N_A_1396_21#_c_1597_n 0.00679802f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_951 N_A_1102_21#_c_1205_n N_A_1396_21#_c_1597_n 0.00688444f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_952 N_A_1102_21#_c_1206_n N_A_1396_21#_c_1597_n 7.55152e-19 $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_953 N_A_1102_21#_c_1207_n N_A_1396_21#_c_1597_n 0.0166785f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_954 N_A_1102_21#_M1047_g N_A_1714_47#_c_1945_n 7.04843e-19 $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_955 N_A_1102_21#_M1035_g N_VPWR_c_2124_n 0.00326498f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_956 N_A_1102_21#_c_1211_n N_VPWR_c_2124_n 0.0124698f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_957 N_A_1102_21#_c_1260_p N_VPWR_c_2124_n 0.00820313f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_958 N_A_1102_21#_c_1213_n N_VPWR_c_2124_n 0.0125544f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_959 N_A_1102_21#_c_1214_n N_VPWR_c_2124_n 7.62241e-19 $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_960 N_A_1102_21#_M1047_g N_VPWR_c_2125_n 0.0163458f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_961 N_A_1102_21#_c_1223_n N_VPWR_c_2125_n 0.0048929f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_962 N_A_1102_21#_c_1211_n N_VPWR_c_2127_n 0.00474052f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_963 N_A_1102_21#_c_1260_p N_VPWR_c_2127_n 0.00725778f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_964 N_A_1102_21#_c_1223_n N_VPWR_c_2127_n 0.00598455f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_965 N_A_1102_21#_M1035_g N_VPWR_c_2134_n 0.00535335f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_966 N_A_1102_21#_c_1213_n N_VPWR_c_2134_n 0.00111392f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_967 N_A_1102_21#_M1047_g N_VPWR_c_2135_n 0.00585385f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_968 N_A_1102_21#_M1012_d N_VPWR_c_2120_n 0.0031612f $X=6.215 $Y=2.065 $X2=0
+ $Y2=0
cc_969 N_A_1102_21#_M1035_g N_VPWR_c_2120_n 0.00664368f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_970 N_A_1102_21#_M1047_g N_VPWR_c_2120_n 0.00762825f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_971 N_A_1102_21#_c_1211_n N_VPWR_c_2120_n 0.00386836f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_972 N_A_1102_21#_c_1260_p N_VPWR_c_2120_n 0.0029026f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_973 N_A_1102_21#_c_1223_n N_VPWR_c_2120_n 0.00505387f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_974 N_A_1102_21#_c_1213_n N_VPWR_c_2120_n 0.00128163f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_975 N_A_1102_21#_c_1223_n A_1351_329# 0.00339576f $X=6.815 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_976 N_A_1102_21#_c_1204_n A_1351_329# 0.00178287f $X=6.9 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_977 N_A_1102_21#_M1009_g N_VGND_c_2536_n 0.00460185f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_978 N_A_1102_21#_c_1202_n N_VGND_c_2537_n 0.0128365f $X=7.995 $Y=0.985 $X2=0
+ $Y2=0
cc_979 N_A_1102_21#_c_1205_n N_VGND_c_2537_n 0.00451721f $X=7.795 $Y=0.98 $X2=0
+ $Y2=0
cc_980 N_A_1102_21#_c_1206_n N_VGND_c_2537_n 0.00366066f $X=7.96 $Y=0.98 $X2=0
+ $Y2=0
cc_981 N_A_1102_21#_c_1207_n N_VGND_c_2537_n 7.09376e-19 $X=7.96 $Y=1.15 $X2=0
+ $Y2=0
cc_982 N_A_1102_21#_M1009_g N_VGND_c_2541_n 0.00361677f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_983 N_A_1102_21#_c_1202_n N_VGND_c_2545_n 0.00368966f $X=7.995 $Y=0.985 $X2=0
+ $Y2=0
cc_984 N_A_1102_21#_M1040_d N_VGND_c_2553_n 0.00178362f $X=6.71 $Y=0.235 $X2=0
+ $Y2=0
cc_985 N_A_1102_21#_M1009_g N_VGND_c_2553_n 0.00583928f $X=5.585 $Y=0.445 $X2=0
+ $Y2=0
cc_986 N_A_1102_21#_c_1202_n N_VGND_c_2553_n 0.00386226f $X=7.995 $Y=0.985 $X2=0
+ $Y2=0
cc_987 N_A_1102_21#_M1040_d N_A_1241_47#_c_2756_n 0.00310223f $X=6.71 $Y=0.235
+ $X2=0 $Y2=0
cc_988 N_A_1102_21#_c_1203_n N_A_1241_47#_c_2756_n 0.0134123f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_989 N_A_1102_21#_c_1205_n N_A_1241_47#_c_2756_n 0.00259503f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_990 N_A_1102_21#_c_1202_n N_A_1241_47#_c_2759_n 0.00441801f $X=7.995 $Y=0.985
+ $X2=0 $Y2=0
cc_991 N_A_1102_21#_c_1205_n N_A_1241_47#_c_2759_n 0.0106429f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_992 N_SET_B_M1004_g N_A_917_47#_M1040_g 0.0269398f $X=6.13 $Y=0.445 $X2=0
+ $Y2=0
cc_993 N_SET_B_c_1349_n N_A_917_47#_M1040_g 0.00357471f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_994 SET_B N_A_917_47#_M1040_g 0.00241265f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_995 N_SET_B_c_1354_n N_A_917_47#_M1040_g 0.00474901f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_996 N_SET_B_c_1355_n N_A_917_47#_M1040_g 0.00138035f $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_997 N_SET_B_M1012_g N_A_917_47#_c_1479_n 0.0210777f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_998 N_SET_B_M1012_g N_A_917_47#_M1036_g 0.0228864f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_999 N_SET_B_M1004_g N_A_917_47#_c_1498_n 3.34359e-19 $X=6.13 $Y=0.445 $X2=0
+ $Y2=0
cc_1000 N_SET_B_M1004_g N_A_917_47#_c_1480_n 0.00152109f $X=6.13 $Y=0.445 $X2=0
+ $Y2=0
cc_1001 N_SET_B_c_1349_n N_A_917_47#_c_1480_n 0.00222178f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_1002 N_SET_B_M1012_g N_A_917_47#_c_1480_n 5.60873e-19 $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_1003 SET_B N_A_917_47#_c_1480_n 0.0203506f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1004 N_SET_B_c_1355_n N_A_917_47#_c_1480_n 0.00109428f $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_1005 N_SET_B_c_1349_n N_A_917_47#_c_1481_n 0.00376157f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_1006 N_SET_B_M1012_g N_A_917_47#_c_1481_n 0.0132556f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_1007 SET_B N_A_917_47#_c_1481_n 0.025593f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1008 N_SET_B_c_1354_n N_A_917_47#_c_1481_n 0.00368272f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1009 N_SET_B_c_1355_n N_A_917_47#_c_1481_n 6.67689e-19 $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_1010 N_SET_B_M1012_g N_A_917_47#_c_1482_n 4.77133e-19 $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_1011 N_SET_B_c_1354_n N_A_1396_21#_M1032_g 0.00317213f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1012 N_SET_B_c_1354_n N_A_1396_21#_c_1596_n 5.29205e-19 $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1013 N_SET_B_M1008_g N_A_1396_21#_c_1605_n 0.00584134f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_1014 N_SET_B_c_1354_n N_A_1396_21#_c_1605_n 0.0486626f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1015 N_SET_B_c_1356_n N_A_1396_21#_c_1605_n 0.0135087f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1016 N_SET_B_M1006_g N_A_1887_21#_M1003_g 0.0176601f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1017 N_SET_B_M1008_g N_A_1887_21#_M1003_g 0.0134226f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_1018 N_SET_B_c_1354_n N_A_1887_21#_M1003_g 0.0062764f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1019 N_SET_B_c_1356_n N_A_1887_21#_M1003_g 0.00136079f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1020 N_SET_B_c_1357_n N_A_1887_21#_M1003_g 0.00225723f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1021 N_SET_B_c_1358_n N_A_1887_21#_M1003_g 0.0208839f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_1022 N_SET_B_M1008_g N_A_1887_21#_M1043_g 0.0109753f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_1023 N_SET_B_M1008_g N_A_1887_21#_c_1769_n 0.00710111f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_1024 N_SET_B_M1008_g N_A_1887_21#_c_1770_n 0.0197396f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_1025 N_SET_B_M1008_g N_A_1887_21#_c_1771_n 0.0136222f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_1026 N_SET_B_c_1357_n N_A_1887_21#_c_1760_n 0.00826722f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1027 N_SET_B_M1006_g N_A_1887_21#_c_1793_n 6.76595e-19 $X=9.945 $Y=0.445
+ $X2=0 $Y2=0
cc_1028 N_SET_B_c_1356_n N_A_1887_21#_c_1793_n 2.38039e-19 $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1029 N_SET_B_c_1357_n N_A_1887_21#_c_1793_n 0.00146062f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1030 N_SET_B_M1006_g N_A_1714_47#_M1020_g 0.0178199f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1031 N_SET_B_c_1357_n N_A_1714_47#_M1020_g 0.00170615f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1032 N_SET_B_c_1358_n N_A_1714_47#_M1020_g 0.00949755f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_1033 N_SET_B_M1008_g N_A_1714_47#_M1023_g 0.0325064f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_1034 N_SET_B_c_1354_n N_A_1714_47#_c_1948_n 0.00885264f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1035 N_SET_B_c_1354_n N_A_1714_47#_c_1934_n 0.017797f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1036 N_SET_B_c_1356_n N_A_1714_47#_c_1934_n 0.0022902f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1037 N_SET_B_c_1357_n N_A_1714_47#_c_1934_n 0.0118231f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1038 N_SET_B_M1008_g N_A_1714_47#_c_1935_n 0.0117551f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_1039 N_SET_B_c_1354_n N_A_1714_47#_c_1935_n 0.00876649f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1040 N_SET_B_c_1356_n N_A_1714_47#_c_1935_n 0.00124273f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1041 N_SET_B_c_1357_n N_A_1714_47#_c_1935_n 0.0248097f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1042 N_SET_B_c_1358_n N_A_1714_47#_c_1935_n 0.00502994f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_1043 N_SET_B_c_1358_n N_A_1714_47#_c_1937_n 0.00111157f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_1044 N_SET_B_c_1358_n N_A_1714_47#_c_1938_n 0.0212871f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_1045 N_SET_B_M1012_g N_VPWR_c_2124_n 0.0094739f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_1046 N_SET_B_M1012_g N_VPWR_c_2127_n 0.00373914f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_1047 N_SET_B_M1008_g N_VPWR_c_2130_n 0.00368415f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_1048 N_SET_B_M1012_g N_VPWR_c_2120_n 0.00439789f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_1049 N_SET_B_M1008_g N_VPWR_c_2120_n 0.00444663f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_1050 N_SET_B_M1008_g N_VPWR_c_2144_n 0.00857728f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_1051 N_SET_B_c_1354_n N_VGND_M1016_s 0.00213425f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_1052 N_SET_B_M1004_g N_VGND_c_2536_n 0.0028663f $X=6.13 $Y=0.445 $X2=0 $Y2=0
cc_1053 N_SET_B_c_1349_n N_VGND_c_2536_n 8.27269e-19 $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_1054 SET_B N_VGND_c_2536_n 0.00871499f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1055 N_SET_B_c_1354_n N_VGND_c_2537_n 0.00430431f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1056 N_SET_B_M1006_g N_VGND_c_2538_n 0.00283027f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1057 N_SET_B_c_1354_n N_VGND_c_2538_n 0.00606882f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1058 N_SET_B_c_1356_n N_VGND_c_2538_n 7.41662e-19 $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1059 N_SET_B_c_1357_n N_VGND_c_2538_n 0.00350326f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1060 N_SET_B_M1004_g N_VGND_c_2543_n 0.00439071f $X=6.13 $Y=0.445 $X2=0 $Y2=0
cc_1061 SET_B N_VGND_c_2543_n 0.0034491f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1062 N_SET_B_M1006_g N_VGND_c_2550_n 0.00439071f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1063 N_SET_B_c_1357_n N_VGND_c_2550_n 0.00352663f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1064 N_SET_B_M1004_g N_VGND_c_2553_n 0.00605812f $X=6.13 $Y=0.445 $X2=0 $Y2=0
cc_1065 N_SET_B_M1006_g N_VGND_c_2553_n 0.00595439f $X=9.945 $Y=0.445 $X2=0
+ $Y2=0
cc_1066 SET_B N_VGND_c_2553_n 0.00346802f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1067 N_SET_B_c_1354_n N_VGND_c_2553_n 0.164988f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_1068 N_SET_B_c_1355_n N_VGND_c_2553_n 0.0148804f $X=6.355 $Y=0.85 $X2=0 $Y2=0
cc_1069 N_SET_B_c_1356_n N_VGND_c_2553_n 0.0141642f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1070 N_SET_B_c_1357_n N_VGND_c_2553_n 0.00284893f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1071 N_SET_B_c_1354_n N_A_1241_47#_M1004_d 0.0016435f $X=9.745 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1072 N_SET_B_c_1355_n N_A_1241_47#_M1004_d 7.95181e-19 $X=6.355 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1073 N_SET_B_c_1354_n N_A_1241_47#_M1032_d 0.00215149f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1074 N_SET_B_c_1354_n N_A_1241_47#_c_2756_n 0.00439674f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1075 N_SET_B_c_1354_n N_A_1241_47#_c_2759_n 0.00234876f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1076 SET_B N_A_1241_47#_c_2766_n 0.00141362f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1077 N_SET_B_c_1354_n N_A_1241_47#_c_2766_n 0.00613011f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1078 N_SET_B_c_1355_n N_A_1241_47#_c_2766_n 0.00187066f $X=6.355 $Y=0.85
+ $X2=0 $Y2=0
cc_1079 N_SET_B_c_1354_n A_1614_47# 0.00377207f $X=9.745 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_1080 N_SET_B_M1006_g N_A_2004_47#_c_2786_n 0.00348207f $X=9.945 $Y=0.445
+ $X2=0 $Y2=0
cc_1081 N_SET_B_c_1357_n N_A_2004_47#_c_2786_n 0.00344477f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1082 N_SET_B_c_1358_n N_A_2004_47#_c_2786_n 2.8008e-19 $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_1083 N_A_917_47#_M1040_g N_A_1396_21#_M1032_g 0.0190309f $X=6.635 $Y=0.555
+ $X2=0 $Y2=0
cc_1084 N_A_917_47#_M1036_g N_A_1396_21#_M1030_g 0.0271962f $X=6.68 $Y=2.065
+ $X2=0 $Y2=0
cc_1085 N_A_917_47#_c_1479_n N_A_1396_21#_c_1597_n 0.0489195f $X=6.68 $Y=1.485
+ $X2=0 $Y2=0
cc_1086 N_A_917_47#_M1036_g N_VPWR_c_2124_n 0.00136797f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1087 N_A_917_47#_M1036_g N_VPWR_c_2127_n 0.00432313f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1088 N_A_917_47#_c_1495_n N_VPWR_c_2134_n 0.0377433f $X=5.295 $Y=2.335 $X2=0
+ $Y2=0
cc_1089 N_A_917_47#_M1039_d N_VPWR_c_2120_n 0.00173085f $X=4.665 $Y=2.065 $X2=0
+ $Y2=0
cc_1090 N_A_917_47#_M1036_g N_VPWR_c_2120_n 0.00600471f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1091 N_A_917_47#_c_1495_n N_VPWR_c_2120_n 0.0132511f $X=5.295 $Y=2.335 $X2=0
+ $Y2=0
cc_1092 N_A_917_47#_c_1490_n N_A_453_47#_c_2348_n 0.0127229f $X=5.485 $Y=0.365
+ $X2=0 $Y2=0
cc_1093 N_A_917_47#_c_1495_n N_A_453_47#_c_2349_n 0.0123114f $X=5.295 $Y=2.335
+ $X2=0 $Y2=0
cc_1094 N_A_917_47#_c_1495_n A_1017_413# 0.00858887f $X=5.295 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1095 N_A_917_47#_c_1485_n A_1017_413# 0.00579571f $X=5.38 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1096 N_A_917_47#_c_1498_n N_VGND_c_2536_n 0.0190862f $X=5.585 $Y=0.655 $X2=0
+ $Y2=0
cc_1097 N_A_917_47#_c_1490_n N_VGND_c_2541_n 0.050218f $X=5.485 $Y=0.365 $X2=0
+ $Y2=0
cc_1098 N_A_917_47#_c_1498_n N_VGND_c_2541_n 0.0103263f $X=5.585 $Y=0.655 $X2=0
+ $Y2=0
cc_1099 N_A_917_47#_M1040_g N_VGND_c_2543_n 0.00357877f $X=6.635 $Y=0.555 $X2=0
+ $Y2=0
cc_1100 N_A_917_47#_M1014_d N_VGND_c_2553_n 0.0027411f $X=4.585 $Y=0.235 $X2=0
+ $Y2=0
cc_1101 N_A_917_47#_M1040_g N_VGND_c_2553_n 0.00542287f $X=6.635 $Y=0.555 $X2=0
+ $Y2=0
cc_1102 N_A_917_47#_c_1490_n N_VGND_c_2553_n 0.017244f $X=5.485 $Y=0.365 $X2=0
+ $Y2=0
cc_1103 N_A_917_47#_c_1498_n N_VGND_c_2553_n 0.00628076f $X=5.585 $Y=0.655 $X2=0
+ $Y2=0
cc_1104 N_A_917_47#_c_1490_n A_1030_47# 0.00710613f $X=5.485 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1105 N_A_917_47#_M1040_g N_A_1241_47#_c_2756_n 0.00692382f $X=6.635 $Y=0.555
+ $X2=0 $Y2=0
cc_1106 N_A_917_47#_M1040_g N_A_1241_47#_c_2766_n 0.00198345f $X=6.635 $Y=0.555
+ $X2=0 $Y2=0
cc_1107 N_A_917_47#_c_1479_n N_A_1241_47#_c_2766_n 0.00105819f $X=6.68 $Y=1.485
+ $X2=0 $Y2=0
cc_1108 N_A_1396_21#_c_1605_n N_A_1887_21#_M1003_g 0.00413877f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1109 N_A_1396_21#_c_1605_n N_A_1887_21#_c_1769_n 0.015309f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1110 N_A_1396_21#_c_1605_n N_A_1887_21#_c_1770_n 0.0070058f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1111 N_A_1396_21#_c_1605_n N_A_1887_21#_c_1771_n 0.010417f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1112 N_A_1396_21#_c_1605_n N_A_1887_21#_c_1800_n 0.00964432f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1113 N_A_1396_21#_M1028_g N_A_1887_21#_c_1760_n 0.012752f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1114 N_A_1396_21#_M1029_g N_A_1887_21#_c_1760_n 0.00627146f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1115 N_A_1396_21#_c_1594_n N_A_1887_21#_c_1760_n 0.0070899f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1116 N_A_1396_21#_c_1602_n N_A_1887_21#_c_1760_n 0.0127165f $X=11.355 $Y=1.66
+ $X2=0 $Y2=0
cc_1117 N_A_1396_21#_c_1605_n N_A_1887_21#_c_1760_n 0.0265111f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1118 N_A_1396_21#_c_1608_n N_A_1887_21#_c_1760_n 5.59542e-19 $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1119 N_A_1396_21#_c_1598_n N_A_1887_21#_c_1760_n 0.00913483f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1120 N_A_1396_21#_c_1599_n N_A_1887_21#_c_1760_n 0.044948f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1121 N_A_1396_21#_M1005_s N_A_1887_21#_c_1773_n 0.00479715f $X=11.555
+ $Y=1.505 $X2=0 $Y2=0
cc_1122 N_A_1396_21#_M1028_g N_A_1887_21#_c_1773_n 0.00741003f $X=10.895
+ $Y=2.065 $X2=0 $Y2=0
cc_1123 N_A_1396_21#_c_1602_n N_A_1887_21#_c_1773_n 0.0212381f $X=11.355 $Y=1.66
+ $X2=0 $Y2=0
cc_1124 N_A_1396_21#_c_1603_n N_A_1887_21#_c_1773_n 0.0321071f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1125 N_A_1396_21#_c_1605_n N_A_1887_21#_c_1773_n 0.00664652f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1126 N_A_1396_21#_c_1608_n N_A_1887_21#_c_1773_n 0.00170504f $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1127 N_A_1396_21#_c_1598_n N_A_1887_21#_c_1773_n 0.00265268f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1128 N_A_1396_21#_c_1603_n N_A_1887_21#_c_1774_n 0.00840283f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1129 N_A_1396_21#_c_1605_n N_A_1887_21#_c_1817_n 0.00453864f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1130 N_A_1396_21#_M1029_g N_A_1887_21#_c_1793_n 0.00433462f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1131 N_A_1396_21#_c_1595_n N_A_1887_21#_c_1793_n 0.00421697f $X=11.68 $Y=0.43
+ $X2=0 $Y2=0
cc_1132 N_A_1396_21#_M1028_g N_A_1887_21#_c_1820_n 0.00480312f $X=10.895
+ $Y=2.065 $X2=0 $Y2=0
cc_1133 N_A_1396_21#_M1029_g N_A_1714_47#_M1020_g 0.0269235f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1134 N_A_1396_21#_M1028_g N_A_1714_47#_M1023_g 0.039703f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1135 N_A_1396_21#_c_1605_n N_A_1714_47#_M1023_g 0.00711753f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1136 N_A_1396_21#_c_1605_n N_A_1714_47#_c_1940_n 0.0219541f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1137 N_A_1396_21#_c_1605_n N_A_1714_47#_c_1935_n 0.0228784f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1138 N_A_1396_21#_M1029_g N_A_1714_47#_c_1937_n 2.38141e-19 $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1139 N_A_1396_21#_c_1605_n N_A_1714_47#_c_1937_n 0.00714757f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1140 N_A_1396_21#_M1029_g N_A_1714_47#_c_1938_n 0.0117459f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1141 N_A_1396_21#_c_1598_n N_A_1714_47#_c_1938_n 0.039703f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1142 N_A_1396_21#_c_1593_n N_RESET_B_M1015_g 0.00688843f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1143 N_A_1396_21#_c_1595_n N_RESET_B_M1015_g 0.00291196f $X=11.68 $Y=0.43
+ $X2=0 $Y2=0
cc_1144 N_A_1396_21#_c_1599_n N_RESET_B_M1015_g 0.00237866f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1145 N_A_1396_21#_c_1603_n N_RESET_B_M1005_g 0.00360287f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1146 N_A_1396_21#_c_1608_n N_RESET_B_M1005_g 0.00264823f $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1147 N_A_1396_21#_c_1598_n N_RESET_B_M1005_g 0.0025096f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1148 N_A_1396_21#_c_1599_n N_RESET_B_M1005_g 0.00309824f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1149 N_A_1396_21#_c_1593_n RESET_B 0.0195128f $X=11.565 $Y=0.84 $X2=0 $Y2=0
cc_1150 N_A_1396_21#_c_1603_n RESET_B 0.015564f $X=11.68 $Y=1.66 $X2=0 $Y2=0
cc_1151 N_A_1396_21#_c_1598_n RESET_B 5.50348e-19 $X=10.95 $Y=1.32 $X2=0 $Y2=0
cc_1152 N_A_1396_21#_c_1599_n RESET_B 0.0185145f $X=11.165 $Y=1.32 $X2=0 $Y2=0
cc_1153 N_A_1396_21#_M1029_g N_RESET_B_c_2034_n 0.00201274f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1154 N_A_1396_21#_c_1593_n N_RESET_B_c_2034_n 0.00537728f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1155 N_A_1396_21#_c_1603_n N_RESET_B_c_2034_n 0.00527649f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1156 N_A_1396_21#_c_1598_n N_RESET_B_c_2034_n 0.0092343f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1157 N_A_1396_21#_c_1599_n N_RESET_B_c_2034_n 0.00327697f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1158 N_A_1396_21#_c_1596_n N_VPWR_M1030_d 0.00297048f $X=7.32 $Y=1.32 $X2=0
+ $Y2=0
cc_1159 N_A_1396_21#_c_1607_n N_VPWR_M1030_d 0.00221014f $X=8.05 $Y=1.53 $X2=0
+ $Y2=0
cc_1160 N_A_1396_21#_c_1602_n N_VPWR_M1028_d 0.00314302f $X=11.355 $Y=1.66 $X2=0
+ $Y2=0
cc_1161 N_A_1396_21#_M1030_g N_VPWR_c_2125_n 0.00353361f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1162 N_A_1396_21#_c_1596_n N_VPWR_c_2125_n 0.011531f $X=7.32 $Y=1.32 $X2=0
+ $Y2=0
cc_1163 N_A_1396_21#_c_1607_n N_VPWR_c_2125_n 7.83548e-19 $X=8.05 $Y=1.53 $X2=0
+ $Y2=0
cc_1164 N_A_1396_21#_c_1597_n N_VPWR_c_2125_n 0.00111411f $X=7.1 $Y=1.32 $X2=0
+ $Y2=0
cc_1165 N_A_1396_21#_M1030_g N_VPWR_c_2127_n 0.00583607f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1166 N_A_1396_21#_M1028_g N_VPWR_c_2129_n 0.0111257f $X=10.895 $Y=2.065 $X2=0
+ $Y2=0
cc_1167 N_A_1396_21#_M1028_g N_VPWR_c_2130_n 0.00339283f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1168 N_A_1396_21#_M1030_g N_VPWR_c_2120_n 0.00670824f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1169 N_A_1396_21#_M1028_g N_VPWR_c_2120_n 0.00383548f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1170 N_A_1396_21#_c_1607_n A_1572_329# 0.00272182f $X=8.05 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_1171 N_A_1396_21#_M1032_g N_VGND_c_2537_n 0.00320142f $X=7.055 $Y=0.555 $X2=0
+ $Y2=0
cc_1172 N_A_1396_21#_c_1593_n N_VGND_c_2539_n 0.00363346f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1173 N_A_1396_21#_c_1595_n N_VGND_c_2539_n 0.00651166f $X=11.68 $Y=0.43 $X2=0
+ $Y2=0
cc_1174 N_A_1396_21#_M1032_g N_VGND_c_2543_n 0.00357877f $X=7.055 $Y=0.555 $X2=0
+ $Y2=0
cc_1175 N_A_1396_21#_M1029_g N_VGND_c_2550_n 0.00357877f $X=10.95 $Y=0.555 $X2=0
+ $Y2=0
cc_1176 N_A_1396_21#_c_1593_n N_VGND_c_2550_n 0.00300947f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1177 N_A_1396_21#_c_1594_n N_VGND_c_2550_n 0.00167376f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1178 N_A_1396_21#_c_1595_n N_VGND_c_2550_n 0.0131956f $X=11.68 $Y=0.43 $X2=0
+ $Y2=0
cc_1179 N_A_1396_21#_M1015_s N_VGND_c_2553_n 0.00353057f $X=11.555 $Y=0.235
+ $X2=0 $Y2=0
cc_1180 N_A_1396_21#_M1032_g N_VGND_c_2553_n 0.00661646f $X=7.055 $Y=0.555 $X2=0
+ $Y2=0
cc_1181 N_A_1396_21#_M1029_g N_VGND_c_2553_n 0.00657041f $X=10.95 $Y=0.555 $X2=0
+ $Y2=0
cc_1182 N_A_1396_21#_c_1593_n N_VGND_c_2553_n 0.00541125f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1183 N_A_1396_21#_c_1594_n N_VGND_c_2553_n 0.00326613f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1184 N_A_1396_21#_c_1595_n N_VGND_c_2553_n 0.00796608f $X=11.68 $Y=0.43 $X2=0
+ $Y2=0
cc_1185 N_A_1396_21#_M1032_g N_A_1241_47#_c_2756_n 0.0105649f $X=7.055 $Y=0.555
+ $X2=0 $Y2=0
cc_1186 N_A_1396_21#_c_1594_n N_A_2004_47#_M1029_d 0.00388496f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1187 N_A_1396_21#_M1029_g N_A_2004_47#_c_2790_n 0.0112006f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1188 N_A_1396_21#_c_1594_n N_A_2004_47#_c_2790_n 0.0138009f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1189 N_A_1396_21#_c_1595_n N_A_2004_47#_c_2790_n 0.0150406f $X=11.68 $Y=0.43
+ $X2=0 $Y2=0
cc_1190 N_A_1396_21#_c_1598_n N_A_2004_47#_c_2790_n 5.45076e-19 $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1191 N_A_1887_21#_c_1760_n N_A_1714_47#_M1020_g 0.0029268f $X=10.817 $Y=1.915
+ $X2=0 $Y2=0
cc_1192 N_A_1887_21#_c_1793_n N_A_1714_47#_M1020_g 0.00534702f $X=10.817
+ $Y=0.687 $X2=0 $Y2=0
cc_1193 N_A_1887_21#_c_1800_n N_A_1714_47#_M1023_g 0.0118664f $X=10.73 $Y=2
+ $X2=0 $Y2=0
cc_1194 N_A_1887_21#_M1043_g N_A_1714_47#_c_1945_n 0.00204127f $X=9.515 $Y=2.275
+ $X2=0 $Y2=0
cc_1195 N_A_1887_21#_M1003_g N_A_1714_47#_c_1934_n 0.0101965f $X=9.51 $Y=0.445
+ $X2=0 $Y2=0
cc_1196 N_A_1887_21#_M1003_g N_A_1714_47#_c_1940_n 0.00912509f $X=9.51 $Y=0.445
+ $X2=0 $Y2=0
cc_1197 N_A_1887_21#_M1043_g N_A_1714_47#_c_1940_n 0.0058046f $X=9.515 $Y=2.275
+ $X2=0 $Y2=0
cc_1198 N_A_1887_21#_c_1769_n N_A_1714_47#_c_1940_n 0.0248025f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1199 N_A_1887_21#_c_1829_p N_A_1714_47#_c_1940_n 0.0135579f $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1200 N_A_1887_21#_M1003_g N_A_1714_47#_c_1935_n 0.0115262f $X=9.51 $Y=0.445
+ $X2=0 $Y2=0
cc_1201 N_A_1887_21#_c_1769_n N_A_1714_47#_c_1935_n 0.0154989f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1202 N_A_1887_21#_c_1770_n N_A_1714_47#_c_1935_n 0.00130368f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1203 N_A_1887_21#_c_1771_n N_A_1714_47#_c_1935_n 0.00635717f $X=10.24 $Y=2
+ $X2=0 $Y2=0
cc_1204 N_A_1887_21#_c_1817_n N_A_1714_47#_c_1935_n 0.00162703f $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1205 N_A_1887_21#_c_1800_n N_A_1714_47#_c_1937_n 0.00158774f $X=10.73 $Y=2
+ $X2=0 $Y2=0
cc_1206 N_A_1887_21#_c_1760_n N_A_1714_47#_c_1937_n 0.0241086f $X=10.817
+ $Y=1.915 $X2=0 $Y2=0
cc_1207 N_A_1887_21#_c_1817_n N_A_1714_47#_c_1937_n 9.97507e-19 $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1208 N_A_1887_21#_c_1760_n N_A_1714_47#_c_1938_n 0.0123488f $X=10.817
+ $Y=1.915 $X2=0 $Y2=0
cc_1209 N_A_1887_21#_c_1817_n N_A_1714_47#_c_1938_n 4.0151e-19 $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1210 N_A_1887_21#_c_1753_n N_RESET_B_M1015_g 0.0182137f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1211 N_A_1887_21#_c_1761_n N_RESET_B_M1015_g 0.00220565f $X=12.34 $Y=1.16
+ $X2=0 $Y2=0
cc_1212 N_A_1887_21#_c_1762_n N_RESET_B_M1015_g 0.0180038f $X=12.34 $Y=1.16
+ $X2=0 $Y2=0
cc_1213 N_A_1887_21#_c_1773_n N_RESET_B_M1005_g 0.0142369f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1214 N_A_1887_21#_c_1773_n RESET_B 0.00314679f $X=12.16 $Y=2 $X2=0 $Y2=0
cc_1215 N_A_1887_21#_c_1761_n RESET_B 0.0193193f $X=12.34 $Y=1.16 $X2=0 $Y2=0
cc_1216 N_A_1887_21#_c_1762_n RESET_B 7.2681e-19 $X=12.34 $Y=1.16 $X2=0 $Y2=0
cc_1217 N_A_1887_21#_M1037_g N_RESET_B_c_2034_n 0.0294485f $X=12.375 $Y=1.985
+ $X2=0 $Y2=0
cc_1218 N_A_1887_21#_c_1774_n N_RESET_B_c_2034_n 0.00991514f $X=12.245 $Y=1.915
+ $X2=0 $Y2=0
cc_1219 N_A_1887_21#_c_1761_n N_RESET_B_c_2034_n 6.95467e-19 $X=12.34 $Y=1.16
+ $X2=0 $Y2=0
cc_1220 N_A_1887_21#_c_1756_n N_A_2596_47#_M1002_g 0.0046261f $X=13.19 $Y=1.535
+ $X2=0 $Y2=0
cc_1221 N_A_1887_21#_c_1768_n N_A_2596_47#_M1002_g 0.0111659f $X=13.315 $Y=1.61
+ $X2=0 $Y2=0
cc_1222 N_A_1887_21#_c_1753_n N_A_2596_47#_c_2068_n 0.00110305f $X=12.375
+ $Y=0.995 $X2=0 $Y2=0
cc_1223 N_A_1887_21#_c_1755_n N_A_2596_47#_c_2068_n 0.00388761f $X=13.19
+ $Y=1.025 $X2=0 $Y2=0
cc_1224 N_A_1887_21#_c_1757_n N_A_2596_47#_c_2068_n 0.00984702f $X=13.315
+ $Y=0.73 $X2=0 $Y2=0
cc_1225 N_A_1887_21#_c_1758_n N_A_2596_47#_c_2068_n 0.00977969f $X=13.315
+ $Y=0.805 $X2=0 $Y2=0
cc_1226 N_A_1887_21#_M1037_g N_A_2596_47#_c_2074_n 0.00166592f $X=12.375
+ $Y=1.985 $X2=0 $Y2=0
cc_1227 N_A_1887_21#_c_1756_n N_A_2596_47#_c_2074_n 0.00715595f $X=13.19
+ $Y=1.535 $X2=0 $Y2=0
cc_1228 N_A_1887_21#_c_1767_n N_A_2596_47#_c_2074_n 0.0108344f $X=13.315
+ $Y=1.685 $X2=0 $Y2=0
cc_1229 N_A_1887_21#_c_1768_n N_A_2596_47#_c_2074_n 0.0101822f $X=13.315 $Y=1.61
+ $X2=0 $Y2=0
cc_1230 N_A_1887_21#_c_1758_n N_A_2596_47#_c_2069_n 0.00368279f $X=13.315
+ $Y=0.805 $X2=0 $Y2=0
cc_1231 N_A_1887_21#_c_1768_n N_A_2596_47#_c_2069_n 0.00324612f $X=13.315
+ $Y=1.61 $X2=0 $Y2=0
cc_1232 N_A_1887_21#_c_1755_n N_A_2596_47#_c_2070_n 0.0131356f $X=13.19 $Y=1.025
+ $X2=0 $Y2=0
cc_1233 N_A_1887_21#_c_1754_n N_A_2596_47#_c_2071_n 0.0110704f $X=13.115 $Y=1.16
+ $X2=0 $Y2=0
cc_1234 N_A_1887_21#_c_1755_n N_A_2596_47#_c_2071_n 0.00116339f $X=13.19
+ $Y=1.025 $X2=0 $Y2=0
cc_1235 N_A_1887_21#_c_1756_n N_A_2596_47#_c_2071_n 0.00116339f $X=13.19
+ $Y=1.535 $X2=0 $Y2=0
cc_1236 N_A_1887_21#_c_1759_n N_A_2596_47#_c_2071_n 0.00732445f $X=13.19 $Y=1.16
+ $X2=0 $Y2=0
cc_1237 N_A_1887_21#_c_1755_n N_A_2596_47#_c_2072_n 0.0025256f $X=13.19 $Y=1.025
+ $X2=0 $Y2=0
cc_1238 N_A_1887_21#_c_1757_n N_A_2596_47#_c_2072_n 0.0159703f $X=13.315 $Y=0.73
+ $X2=0 $Y2=0
cc_1239 N_A_1887_21#_c_1771_n N_VPWR_M1043_d 0.00124767f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1240 N_A_1887_21#_c_1829_p N_VPWR_M1043_d 0.00160397f $X=9.8 $Y=2 $X2=0 $Y2=0
cc_1241 N_A_1887_21#_c_1773_n N_VPWR_M1028_d 0.0044189f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1242 N_A_1887_21#_c_1773_n N_VPWR_M1005_d 0.00750664f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1243 N_A_1887_21#_c_1774_n N_VPWR_M1005_d 0.00487804f $X=12.245 $Y=1.915
+ $X2=0 $Y2=0
cc_1244 N_A_1887_21#_c_1767_n N_VPWR_c_2126_n 0.00444994f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1245 N_A_1887_21#_c_1773_n N_VPWR_c_2129_n 0.0844105f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1246 N_A_1887_21#_c_1771_n N_VPWR_c_2130_n 0.00359839f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1247 N_A_1887_21#_c_1877_p N_VPWR_c_2130_n 0.00713694f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1248 N_A_1887_21#_c_1800_n N_VPWR_c_2130_n 0.00458994f $X=10.73 $Y=2 $X2=0
+ $Y2=0
cc_1249 N_A_1887_21#_c_1773_n N_VPWR_c_2130_n 5.56361e-19 $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1250 N_A_1887_21#_c_1820_n N_VPWR_c_2130_n 0.00270619f $X=10.817 $Y=2 $X2=0
+ $Y2=0
cc_1251 N_A_1887_21#_M1043_g N_VPWR_c_2135_n 0.00542601f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1252 N_A_1887_21#_c_1829_p N_VPWR_c_2135_n 9.91118e-19 $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1253 N_A_1887_21#_M1037_g N_VPWR_c_2137_n 0.0046653f $X=12.375 $Y=1.985 $X2=0
+ $Y2=0
cc_1254 N_A_1887_21#_c_1767_n N_VPWR_c_2137_n 0.00464873f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1255 N_A_1887_21#_M1008_d N_VPWR_c_2120_n 0.00327257f $X=10.13 $Y=2.065 $X2=0
+ $Y2=0
cc_1256 N_A_1887_21#_M1043_g N_VPWR_c_2120_n 0.00997697f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1257 N_A_1887_21#_M1037_g N_VPWR_c_2120_n 0.00929621f $X=12.375 $Y=1.985
+ $X2=0 $Y2=0
cc_1258 N_A_1887_21#_c_1767_n N_VPWR_c_2120_n 0.00924075f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1259 N_A_1887_21#_c_1771_n N_VPWR_c_2120_n 0.00704318f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1260 N_A_1887_21#_c_1829_p N_VPWR_c_2120_n 0.00270501f $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1261 N_A_1887_21#_c_1877_p N_VPWR_c_2120_n 0.00608739f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1262 N_A_1887_21#_c_1800_n N_VPWR_c_2120_n 0.00829558f $X=10.73 $Y=2 $X2=0
+ $Y2=0
cc_1263 N_A_1887_21#_c_1773_n N_VPWR_c_2120_n 0.00701098f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1264 N_A_1887_21#_c_1820_n N_VPWR_c_2120_n 0.00481592f $X=10.817 $Y=2 $X2=0
+ $Y2=0
cc_1265 N_A_1887_21#_M1043_g N_VPWR_c_2144_n 0.00321606f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1266 N_A_1887_21#_c_1770_n N_VPWR_c_2144_n 7.01948e-19 $X=9.635 $Y=1.74 $X2=0
+ $Y2=0
cc_1267 N_A_1887_21#_c_1771_n N_VPWR_c_2144_n 0.0106677f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1268 N_A_1887_21#_c_1829_p N_VPWR_c_2144_n 0.0126362f $X=9.8 $Y=2 $X2=0 $Y2=0
cc_1269 N_A_1887_21#_c_1877_p N_VPWR_c_2144_n 0.00687131f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1270 N_A_1887_21#_M1037_g N_VPWR_c_2145_n 0.0100464f $X=12.375 $Y=1.985 $X2=0
+ $Y2=0
cc_1271 N_A_1887_21#_c_1773_n N_VPWR_c_2145_n 0.00915613f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1272 N_A_1887_21#_c_1800_n A_2122_329# 0.00202121f $X=10.73 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1273 N_A_1887_21#_c_1760_n A_2122_329# 0.0030402f $X=10.817 $Y=1.915
+ $X2=-0.19 $Y2=-0.24
cc_1274 N_A_1887_21#_c_1820_n A_2122_329# 5.84995e-19 $X=10.817 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1275 N_A_1887_21#_c_1754_n N_Q_N_c_2490_n 0.00237367f $X=13.115 $Y=1.16 $X2=0
+ $Y2=0
cc_1276 N_A_1887_21#_c_1767_n N_Q_N_c_2490_n 0.00131217f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1277 N_A_1887_21#_c_1768_n N_Q_N_c_2490_n 5.76238e-19 $X=13.315 $Y=1.61 $X2=0
+ $Y2=0
cc_1278 N_A_1887_21#_c_1753_n N_Q_N_c_2487_n 0.00547914f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1279 N_A_1887_21#_c_1754_n N_Q_N_c_2487_n 0.0206846f $X=13.115 $Y=1.16 $X2=0
+ $Y2=0
cc_1280 N_A_1887_21#_c_1756_n N_Q_N_c_2487_n 5.76238e-19 $X=13.19 $Y=1.535 $X2=0
+ $Y2=0
cc_1281 N_A_1887_21#_c_1758_n N_Q_N_c_2487_n 8.63605e-19 $X=13.315 $Y=0.805
+ $X2=0 $Y2=0
cc_1282 N_A_1887_21#_c_1774_n N_Q_N_c_2487_n 0.0126467f $X=12.245 $Y=1.915 $X2=0
+ $Y2=0
cc_1283 N_A_1887_21#_c_1761_n N_Q_N_c_2487_n 0.0224115f $X=12.34 $Y=1.16 $X2=0
+ $Y2=0
cc_1284 N_A_1887_21#_c_1762_n N_Q_N_c_2487_n 0.00302465f $X=12.34 $Y=1.16 $X2=0
+ $Y2=0
cc_1285 N_A_1887_21#_c_1754_n Q_N 0.00230535f $X=13.115 $Y=1.16 $X2=0 $Y2=0
cc_1286 N_A_1887_21#_c_1767_n Q_N 8.70693e-19 $X=13.315 $Y=1.685 $X2=0 $Y2=0
cc_1287 N_A_1887_21#_c_1757_n N_Q_N_c_2489_n 0.00104845f $X=13.315 $Y=0.73 $X2=0
+ $Y2=0
cc_1288 N_A_1887_21#_M1003_g N_VGND_c_2538_n 0.00815427f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_1289 N_A_1887_21#_c_1753_n N_VGND_c_2539_n 0.0127745f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1290 N_A_1887_21#_c_1761_n N_VGND_c_2539_n 0.0105198f $X=12.34 $Y=1.16 $X2=0
+ $Y2=0
cc_1291 N_A_1887_21#_c_1762_n N_VGND_c_2539_n 0.00200592f $X=12.34 $Y=1.16 $X2=0
+ $Y2=0
cc_1292 N_A_1887_21#_c_1757_n N_VGND_c_2540_n 0.00415965f $X=13.315 $Y=0.73
+ $X2=0 $Y2=0
cc_1293 N_A_1887_21#_M1003_g N_VGND_c_2545_n 0.00486043f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_1294 N_A_1887_21#_c_1753_n N_VGND_c_2551_n 0.0046653f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1295 N_A_1887_21#_c_1757_n N_VGND_c_2551_n 0.00533769f $X=13.315 $Y=0.73
+ $X2=0 $Y2=0
cc_1296 N_A_1887_21#_c_1758_n N_VGND_c_2551_n 2.84936e-19 $X=13.315 $Y=0.805
+ $X2=0 $Y2=0
cc_1297 N_A_1887_21#_M1020_d N_VGND_c_2553_n 0.00216833f $X=10.605 $Y=0.235
+ $X2=0 $Y2=0
cc_1298 N_A_1887_21#_M1003_g N_VGND_c_2553_n 0.00476342f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_1299 N_A_1887_21#_c_1753_n N_VGND_c_2553_n 0.00934473f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1300 N_A_1887_21#_c_1757_n N_VGND_c_2553_n 0.0109269f $X=13.315 $Y=0.73 $X2=0
+ $Y2=0
cc_1301 N_A_1887_21#_M1020_d N_A_2004_47#_c_2790_n 0.00312752f $X=10.605
+ $Y=0.235 $X2=0 $Y2=0
cc_1302 N_A_1887_21#_c_1793_n N_A_2004_47#_c_2790_n 0.0145304f $X=10.817
+ $Y=0.687 $X2=0 $Y2=0
cc_1303 N_A_1714_47#_M1023_g N_VPWR_c_2129_n 0.00209073f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1304 N_A_1714_47#_M1023_g N_VPWR_c_2130_n 0.00425094f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1305 N_A_1714_47#_c_1945_n N_VPWR_c_2135_n 0.0377433f $X=9.21 $Y=2.335 $X2=0
+ $Y2=0
cc_1306 N_A_1714_47#_M1031_d N_VPWR_c_2120_n 0.00205544f $X=8.58 $Y=2.065 $X2=0
+ $Y2=0
cc_1307 N_A_1714_47#_M1023_g N_VPWR_c_2120_n 0.00591666f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1308 N_A_1714_47#_c_1945_n N_VPWR_c_2120_n 0.0272797f $X=9.21 $Y=2.335 $X2=0
+ $Y2=0
cc_1309 N_A_1714_47#_M1023_g N_VPWR_c_2144_n 0.00144209f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1310 N_A_1714_47#_c_1945_n A_1800_413# 0.0111731f $X=9.21 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1311 N_A_1714_47#_c_1940_n A_1800_413# 0.00577347f $X=9.295 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1312 N_A_1714_47#_c_1948_n N_VGND_c_2545_n 0.0433004f $X=9.21 $Y=0.365 $X2=0
+ $Y2=0
cc_1313 N_A_1714_47#_M1020_g N_VGND_c_2550_n 0.00357877f $X=10.53 $Y=0.555 $X2=0
+ $Y2=0
cc_1314 N_A_1714_47#_M1010_d N_VGND_c_2553_n 0.00269406f $X=8.57 $Y=0.235 $X2=0
+ $Y2=0
cc_1315 N_A_1714_47#_M1020_g N_VGND_c_2553_n 0.00568671f $X=10.53 $Y=0.555 $X2=0
+ $Y2=0
cc_1316 N_A_1714_47#_c_1948_n N_VGND_c_2553_n 0.0129075f $X=9.21 $Y=0.365 $X2=0
+ $Y2=0
cc_1317 N_A_1714_47#_c_1948_n A_1822_47# 0.00370882f $X=9.21 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1318 N_A_1714_47#_c_1934_n A_1822_47# 0.00307731f $X=9.295 $Y=1.235 $X2=-0.19
+ $Y2=-0.24
cc_1319 N_A_1714_47#_M1020_g N_A_2004_47#_c_2790_n 0.0109023f $X=10.53 $Y=0.555
+ $X2=0 $Y2=0
cc_1320 N_A_1714_47#_c_1937_n N_A_2004_47#_c_2790_n 0.00298717f $X=10.475
+ $Y=1.24 $X2=0 $Y2=0
cc_1321 N_A_1714_47#_c_1937_n N_A_2004_47#_c_2786_n 0.00197757f $X=10.475
+ $Y=1.24 $X2=0 $Y2=0
cc_1322 N_A_1714_47#_c_1938_n N_A_2004_47#_c_2786_n 3.51607e-19 $X=10.475
+ $Y=1.24 $X2=0 $Y2=0
cc_1323 N_RESET_B_M1005_g N_VPWR_c_2136_n 0.00655753f $X=11.89 $Y=1.825 $X2=0
+ $Y2=0
cc_1324 N_RESET_B_M1015_g N_VGND_c_2539_n 0.00662758f $X=11.89 $Y=0.445 $X2=0
+ $Y2=0
cc_1325 N_RESET_B_M1015_g N_VGND_c_2550_n 0.00585385f $X=11.89 $Y=0.445 $X2=0
+ $Y2=0
cc_1326 N_RESET_B_M1015_g N_VGND_c_2553_n 0.0120869f $X=11.89 $Y=0.445 $X2=0
+ $Y2=0
cc_1327 N_A_2596_47#_M1002_g N_VPWR_c_2126_n 0.0142968f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1328 N_A_2596_47#_c_2074_n N_VPWR_c_2126_n 0.047587f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1329 N_A_2596_47#_c_2069_n N_VPWR_c_2126_n 0.0103596f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1330 N_A_2596_47#_c_2070_n N_VPWR_c_2126_n 0.00249491f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1331 N_A_2596_47#_c_2074_n N_VPWR_c_2137_n 0.0169293f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1332 N_A_2596_47#_M1002_g N_VPWR_c_2138_n 0.00486043f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1333 N_A_2596_47#_M1002_g N_VPWR_c_2120_n 0.0092657f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1334 N_A_2596_47#_c_2074_n N_VPWR_c_2120_n 0.0115924f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1335 N_A_2596_47#_c_2074_n N_Q_N_c_2487_n 0.0871059f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1336 N_A_2596_47#_c_2071_n N_Q_N_c_2487_n 0.0251545f $X=13.117 $Y=1.16 $X2=0
+ $Y2=0
cc_1337 N_A_2596_47#_c_2068_n N_Q_N_c_2489_n 0.0590331f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1338 N_A_2596_47#_M1002_g N_Q_c_2520_n 0.00523703f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1339 N_A_2596_47#_c_2074_n N_Q_c_2520_n 0.00411039f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1340 N_A_2596_47#_c_2069_n N_Q_c_2518_n 0.0266146f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1341 N_A_2596_47#_c_2072_n N_Q_c_2518_n 0.0212692f $X=13.72 $Y=0.995 $X2=0
+ $Y2=0
cc_1342 N_A_2596_47#_c_2068_n N_VGND_c_2540_n 0.0212529f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1343 N_A_2596_47#_c_2069_n N_VGND_c_2540_n 0.0103062f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1344 N_A_2596_47#_c_2070_n N_VGND_c_2540_n 0.00246314f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1345 N_A_2596_47#_c_2072_n N_VGND_c_2540_n 0.00939953f $X=13.72 $Y=0.995
+ $X2=0 $Y2=0
cc_1346 N_A_2596_47#_c_2068_n N_VGND_c_2551_n 0.0199778f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1347 N_A_2596_47#_c_2072_n N_VGND_c_2552_n 0.0046653f $X=13.72 $Y=0.995 $X2=0
+ $Y2=0
cc_1348 N_A_2596_47#_M1046_s N_VGND_c_2553_n 0.00210122f $X=12.98 $Y=0.235 $X2=0
+ $Y2=0
cc_1349 N_A_2596_47#_c_2068_n N_VGND_c_2553_n 0.0118987f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1350 N_A_2596_47#_c_2072_n N_VGND_c_2553_n 0.00895857f $X=13.72 $Y=0.995
+ $X2=0 $Y2=0
cc_1351 N_VPWR_c_2120_n N_A_453_47#_M1017_d 0.00314748f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1352 N_VPWR_c_2122_n N_A_453_47#_c_2338_n 0.0170763f $X=1.62 $Y=1.97 $X2=0
+ $Y2=0
cc_1353 N_VPWR_c_2133_n N_A_453_47#_c_2338_n 0.0151498f $X=3.31 $Y=2.72 $X2=0
+ $Y2=0
cc_1354 N_VPWR_c_2120_n N_A_453_47#_c_2338_n 0.00610123f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1355 N_VPWR_c_2134_n N_A_453_47#_c_2349_n 0.0146346f $X=5.705 $Y=2.72 $X2=0
+ $Y2=0
cc_1356 N_VPWR_c_2120_n N_A_453_47#_c_2349_n 0.00387733f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1357 N_VPWR_c_2120_n A_752_413# 0.00234073f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1358 N_VPWR_c_2120_n A_1017_413# 0.00350408f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1359 N_VPWR_c_2120_n A_1351_329# 0.0026811f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1360 N_VPWR_c_2120_n A_1572_329# 0.00777501f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1361 N_VPWR_c_2120_n A_1800_413# 0.00555699f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1362 N_VPWR_c_2120_n A_2122_329# 0.00245111f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1363 N_VPWR_c_2120_n N_Q_N_M1037_d 0.00387172f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1364 N_VPWR_c_2126_n Q_N 0.00154263f $X=13.575 $Y=1.94 $X2=0 $Y2=0
cc_1365 N_VPWR_c_2137_n Q_N 0.0197934f $X=13.455 $Y=2.72 $X2=0 $Y2=0
cc_1366 N_VPWR_c_2120_n Q_N 0.0108988f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1367 N_VPWR_c_2120_n N_Q_M1002_d 0.00387172f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1368 N_VPWR_c_2138_n Q 0.018001f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1369 N_VPWR_c_2120_n Q 0.00993603f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1370 N_A_453_47#_c_2331_n N_VGND_c_2535_n 0.00124227f $X=2.57 $Y=0.43 $X2=0
+ $Y2=0
cc_1371 N_A_453_47#_c_2348_n N_VGND_c_2541_n 0.0162566f $X=4.035 $Y=0.43 $X2=0
+ $Y2=0
cc_1372 N_A_453_47#_c_2331_n N_VGND_c_2549_n 0.020692f $X=2.57 $Y=0.43 $X2=0
+ $Y2=0
cc_1373 N_A_453_47#_M1013_d N_VGND_c_2553_n 0.00221188f $X=2.265 $Y=0.235 $X2=0
+ $Y2=0
cc_1374 N_A_453_47#_M1027_d N_VGND_c_2553_n 0.00297483f $X=4.11 $Y=0.235 $X2=0
+ $Y2=0
cc_1375 N_A_453_47#_c_2331_n N_VGND_c_2553_n 0.0057868f $X=2.57 $Y=0.43 $X2=0
+ $Y2=0
cc_1376 N_A_453_47#_c_2348_n N_VGND_c_2553_n 0.00600312f $X=4.035 $Y=0.43 $X2=0
+ $Y2=0
cc_1377 N_Q_N_c_2487_n N_VGND_c_2539_n 0.00205006f $X=12.642 $Y=1.63 $X2=0 $Y2=0
cc_1378 N_Q_N_c_2489_n N_VGND_c_2551_n 0.0196011f $X=12.642 $Y=0.573 $X2=0 $Y2=0
cc_1379 N_Q_N_M1001_d N_VGND_c_2553_n 0.00387172f $X=12.45 $Y=0.235 $X2=0 $Y2=0
cc_1380 N_Q_N_c_2489_n N_VGND_c_2553_n 0.010859f $X=12.642 $Y=0.573 $X2=0 $Y2=0
cc_1381 Q N_VGND_c_2552_n 0.0179467f $X=13.945 $Y=0.425 $X2=0 $Y2=0
cc_1382 N_Q_M1018_d N_VGND_c_2553_n 0.00387172f $X=13.865 $Y=0.235 $X2=0 $Y2=0
cc_1383 Q N_VGND_c_2553_n 0.00992392f $X=13.945 $Y=0.425 $X2=0 $Y2=0
cc_1384 N_VGND_c_2553_n A_381_47# 0.00165237f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1385 N_VGND_c_2553_n A_735_47# 0.00358656f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1386 N_VGND_c_2553_n A_1030_47# 0.00250526f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1387 N_VGND_c_2553_n N_A_1241_47#_M1004_d 0.00245729f $X=14.03 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1388 N_VGND_c_2553_n N_A_1241_47#_M1032_d 0.00204204f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1389 N_VGND_c_2537_n N_A_1241_47#_c_2756_n 0.0106201f $X=7.785 $Y=0.38 $X2=0
+ $Y2=0
cc_1390 N_VGND_c_2543_n N_A_1241_47#_c_2756_n 0.0113927f $X=7.62 $Y=0 $X2=0
+ $Y2=0
cc_1391 N_VGND_c_2553_n N_A_1241_47#_c_2756_n 0.00305438f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1392 N_VGND_c_2537_n N_A_1241_47#_c_2759_n 0.00222831f $X=7.785 $Y=0.38 $X2=0
+ $Y2=0
cc_1393 N_VGND_c_2543_n N_A_1241_47#_c_2766_n 0.0516775f $X=7.62 $Y=0 $X2=0
+ $Y2=0
cc_1394 N_VGND_c_2553_n N_A_1241_47#_c_2766_n 0.0150078f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1395 N_VGND_c_2553_n A_1614_47# 0.00506251f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1396 N_VGND_c_2553_n A_1822_47# 0.00257693f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1397 N_VGND_c_2553_n N_A_2004_47#_M1006_d 0.0037415f $X=14.03 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1398 N_VGND_c_2553_n N_A_2004_47#_M1029_d 0.00224765f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1399 N_VGND_c_2550_n N_A_2004_47#_c_2790_n 0.0470538f $X=12 $Y=0 $X2=0 $Y2=0
cc_1400 N_VGND_c_2553_n N_A_2004_47#_c_2790_n 0.029878f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1401 N_VGND_c_2550_n N_A_2004_47#_c_2786_n 0.0213706f $X=12 $Y=0 $X2=0 $Y2=0
cc_1402 N_VGND_c_2553_n N_A_2004_47#_c_2786_n 0.01237f $X=14.03 $Y=0 $X2=0 $Y2=0

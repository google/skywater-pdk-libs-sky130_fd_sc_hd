* NGSPICE file created from sky130_fd_sc_hd__and4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
M1000 a_27_47# C VPWR VPB phighvt w=420000u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=8.895e+11p ps=6.3e+06u
M1001 a_303_47# C a_197_47# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.596e+11p ps=1.6e+06u
M1002 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=3.9255e+11p ps=2.66e+06u
M1003 a_197_47# B a_109_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1004 VPWR B a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_47# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND D a_303_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR D a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_109_47# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1009 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__a211o_1.spice
* Created: Tue Sep  1 18:50:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a211o_1.pex.spice"
.subckt sky130_fd_sc_hd__a211o_1  VNB VPB A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_80_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.26 AS=0.17225 PD=1.45 PS=1.83 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1003 A_300_47# N_A2_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.26 PD=0.93 PS=1.45 NRD=15.684 NRS=14.76 M=1 R=4.33333 SA=75001.1
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1008 N_A_80_21#_M1008_d N_A1_M1008_g A_300_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75001.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_B1_M1001_g N_A_80_21#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.091 PD=0.96 PS=0.93 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_A_80_21#_M1007_d N_C1_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.10075 PD=1.83 PS=0.96 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75002.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_80_21#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A2_M1009_g N_A_217_297#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1005 N_A_217_297#_M1005_d N_A1_M1005_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 A_472_297# N_B1_M1000_g N_A_217_297#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.14 PD=1.31 PS=1.28 NRD=19.6803 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_80_21#_M1002_d N_C1_M1002_g A_472_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.155 PD=2.53 PS=1.31 NRD=0 NRS=19.6803 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_56 VPB 0 1.60767e-19 $X=0.135 $Y=2.635
*
.include "sky130_fd_sc_hd__a211o_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o2111ai_1.pxi.spice
* Created: Tue Sep  1 19:20:10 2020
* 
x_PM_SKY130_FD_SC_HD__O2111AI_1%D1 N_D1_M1007_g N_D1_M1002_g D1 D1 N_D1_c_55_n
+ PM_SKY130_FD_SC_HD__O2111AI_1%D1
x_PM_SKY130_FD_SC_HD__O2111AI_1%C1 N_C1_M1003_g N_C1_M1004_g C1 C1 N_C1_c_87_n
+ PM_SKY130_FD_SC_HD__O2111AI_1%C1
x_PM_SKY130_FD_SC_HD__O2111AI_1%B1 N_B1_M1005_g N_B1_M1006_g B1 B1 N_B1_c_124_n
+ N_B1_c_125_n PM_SKY130_FD_SC_HD__O2111AI_1%B1
x_PM_SKY130_FD_SC_HD__O2111AI_1%A2 N_A2_M1009_g N_A2_M1008_g A2 A2 N_A2_c_159_n
+ N_A2_c_160_n PM_SKY130_FD_SC_HD__O2111AI_1%A2
x_PM_SKY130_FD_SC_HD__O2111AI_1%A1 N_A1_M1000_g N_A1_M1001_g A1 N_A1_c_197_n
+ PM_SKY130_FD_SC_HD__O2111AI_1%A1
x_PM_SKY130_FD_SC_HD__O2111AI_1%VPWR N_VPWR_M1007_s N_VPWR_M1004_d
+ N_VPWR_M1001_d N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n
+ N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n VPWR
+ N_VPWR_c_230_n N_VPWR_c_221_n PM_SKY130_FD_SC_HD__O2111AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O2111AI_1%Y N_Y_M1002_s N_Y_M1007_d N_Y_M1006_d
+ N_Y_c_304_n N_Y_c_290_n N_Y_c_298_n N_Y_c_311_n N_Y_c_276_n N_Y_c_282_n Y Y
+ N_Y_c_275_n PM_SKY130_FD_SC_HD__O2111AI_1%Y
x_PM_SKY130_FD_SC_HD__O2111AI_1%A_343_47# N_A_343_47#_M1005_d
+ N_A_343_47#_M1000_d N_A_343_47#_c_331_n N_A_343_47#_c_344_p
+ N_A_343_47#_c_329_n N_A_343_47#_c_330_n
+ PM_SKY130_FD_SC_HD__O2111AI_1%A_343_47#
x_PM_SKY130_FD_SC_HD__O2111AI_1%VGND N_VGND_M1009_d N_VGND_c_353_n VGND
+ N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n
+ PM_SKY130_FD_SC_HD__O2111AI_1%VGND
cc_1 VNB N_D1_M1007_g 5.21268e-19 $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.985
cc_2 VNB N_D1_M1002_g 0.0209284f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=0.56
cc_3 VNB N_D1_c_55_n 0.0299139f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_4 VNB N_C1_M1003_g 0.0177335f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.985
cc_5 VNB N_C1_M1004_g 4.69323e-19 $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=0.56
cc_6 VNB C1 0.00142068f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_7 VNB N_C1_c_87_n 0.0286601f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_8 VNB N_B1_M1005_g 0.0201512f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.985
cc_9 VNB N_B1_M1006_g 4.58507e-19 $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=0.56
cc_10 VNB N_B1_c_124_n 0.0268575f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_11 VNB N_B1_c_125_n 0.00573654f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_12 VNB N_A2_M1009_g 0.0202313f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.985
cc_13 VNB N_A2_M1008_g 4.58507e-19 $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=0.56
cc_14 VNB N_A2_c_159_n 0.0254145f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.025
cc_15 VNB N_A2_c_160_n 0.00822454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_M1000_g 0.0248229f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.985
cc_17 VNB A1 0.0140665f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_18 VNB N_A1_c_197_n 0.035975f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_19 VNB N_VPWR_c_221_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB Y 0.0218527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_275_n 0.0425106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_343_47#_c_329_n 0.00868656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_343_47#_c_330_n 0.0145675f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_24 VNB N_VGND_c_353_n 0.0055721f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=0.56
cc_25 VNB N_VGND_c_354_n 0.0616997f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_26 VNB N_VGND_c_355_n 0.017407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_356_n 0.183517f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.53
cc_28 VNB N_VGND_c_357_n 0.00631048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_D1_M1007_g 0.0228639f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.985
cc_30 VPB D1 0.00286395f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_31 VPB N_C1_M1004_g 0.0206161f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=0.56
cc_32 VPB C1 0.00111502f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_33 VPB N_B1_M1006_g 0.0209765f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=0.56
cc_34 VPB N_B1_c_125_n 0.00236436f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_35 VPB N_A2_M1008_g 0.0209765f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=0.56
cc_36 VPB N_A2_c_160_n 0.00227301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A1_M1001_g 0.0249669f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=0.56
cc_38 VPB A1 0.0120881f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_39 VPB N_A1_c_197_n 0.00869351f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_40 VPB N_VPWR_c_222_n 0.0142261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_223_n 0.0049942f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.025
cc_42 VPB N_VPWR_c_224_n 0.0106587f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_43 VPB N_VPWR_c_225_n 0.0297238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_226_n 0.0105569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_227_n 0.00510476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_228_n 0.0140553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_229_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_230_n 0.0317393f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_221_n 0.0456197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_Y_c_276_n 7.43506e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB Y 0.0398112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_D1_M1002_g N_C1_M1003_g 0.0351687f $X=0.74 $Y=0.56 $X2=0 $Y2=0
cc_53 N_D1_M1007_g N_C1_M1004_g 0.0242684f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_54 D1 N_C1_M1004_g 0.00190382f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_55 N_D1_M1007_g C1 3.67424e-19 $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_56 N_D1_M1002_g C1 0.0041564f $X=0.74 $Y=0.56 $X2=0 $Y2=0
cc_57 D1 C1 0.0353271f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_58 D1 N_C1_c_87_n 7.6624e-19 $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_59 N_D1_c_55_n N_C1_c_87_n 0.0351687f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_60 D1 N_VPWR_M1007_s 0.00198669f $X=0.605 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_61 N_D1_M1007_g N_VPWR_c_222_n 0.00826526f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_62 N_D1_M1007_g N_VPWR_c_228_n 0.00360664f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_63 N_D1_M1007_g N_VPWR_c_221_n 0.00426085f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_64 D1 N_Y_M1007_d 0.00135505f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_65 N_D1_M1007_g N_Y_c_276_n 0.0141599f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_66 D1 N_Y_c_276_n 0.0157034f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_67 N_D1_c_55_n N_Y_c_276_n 3.22022e-19 $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_68 D1 N_Y_c_282_n 0.00106376f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_69 N_D1_M1007_g Y 0.00711205f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_70 N_D1_M1002_g Y 0.00405936f $X=0.74 $Y=0.56 $X2=0 $Y2=0
cc_71 D1 Y 0.0426598f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_72 N_D1_c_55_n Y 0.00690821f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_73 N_D1_M1002_g N_Y_c_275_n 0.00909066f $X=0.74 $Y=0.56 $X2=0 $Y2=0
cc_74 D1 N_Y_c_275_n 0.0134618f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_75 N_D1_c_55_n N_Y_c_275_n 0.00439402f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_76 N_D1_M1002_g N_VGND_c_354_n 0.0054895f $X=0.74 $Y=0.56 $X2=0 $Y2=0
cc_77 N_D1_M1002_g N_VGND_c_356_n 0.0108821f $X=0.74 $Y=0.56 $X2=0 $Y2=0
cc_78 N_C1_M1003_g N_B1_M1005_g 0.0250828f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_79 C1 N_B1_M1005_g 0.00931362f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_80 N_C1_M1004_g N_B1_M1006_g 0.034348f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_81 C1 N_B1_M1006_g 0.00111231f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_82 C1 N_B1_c_124_n 3.11466e-19 $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_83 N_C1_c_87_n N_B1_c_124_n 0.0168786f $X=1.19 $Y=1.16 $X2=0 $Y2=0
cc_84 N_C1_M1004_g N_B1_c_125_n 5.59388e-19 $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_85 C1 N_B1_c_125_n 0.0444609f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_86 N_C1_c_87_n N_B1_c_125_n 0.00150127f $X=1.19 $Y=1.16 $X2=0 $Y2=0
cc_87 C1 N_VPWR_M1004_d 0.00247112f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_88 N_C1_M1004_g N_VPWR_c_222_n 5.44914e-19 $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_89 N_C1_M1004_g N_VPWR_c_223_n 0.00302715f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_90 N_C1_M1004_g N_VPWR_c_228_n 0.00433717f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_91 N_C1_M1004_g N_VPWR_c_221_n 0.00617618f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_92 N_C1_M1004_g N_Y_c_290_n 0.0126428f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_93 C1 N_Y_c_290_n 0.021788f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_94 N_C1_c_87_n N_Y_c_290_n 5.76654e-19 $X=1.19 $Y=1.16 $X2=0 $Y2=0
cc_95 N_C1_M1003_g N_Y_c_275_n 0.00158098f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_96 C1 N_Y_c_275_n 0.0287849f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_97 C1 A_235_47# 0.00899777f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_98 N_C1_M1003_g N_VGND_c_354_n 0.00359186f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_99 C1 N_VGND_c_354_n 0.0207604f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_100 N_C1_M1003_g N_VGND_c_356_n 0.00542543f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_101 C1 N_VGND_c_356_n 0.0119505f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_102 N_B1_M1005_g N_A2_M1009_g 0.0161672f $X=1.64 $Y=0.56 $X2=0 $Y2=0
cc_103 N_B1_M1006_g N_A2_M1008_g 0.0252416f $X=1.64 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B1_c_125_n N_A2_M1008_g 8.73452e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B1_c_124_n N_A2_c_159_n 0.0152927f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B1_c_125_n N_A2_c_159_n 2.32847e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B1_M1006_g N_A2_c_160_n 0.00107501f $X=1.64 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B1_c_124_n N_A2_c_160_n 0.00198199f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_109 N_B1_c_125_n N_A2_c_160_n 0.0523216f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B1_M1006_g N_VPWR_c_223_n 0.0032033f $X=1.64 $Y=1.985 $X2=0 $Y2=0
cc_111 N_B1_M1006_g N_VPWR_c_230_n 0.00433717f $X=1.64 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B1_M1006_g N_VPWR_c_221_n 0.00642404f $X=1.64 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B1_c_125_n N_Y_M1006_d 0.00161675f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_M1006_g N_Y_c_290_n 0.0160687f $X=1.64 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B1_c_125_n N_Y_c_290_n 0.0116161f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B1_c_124_n N_Y_c_298_n 0.00272096f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B1_c_125_n N_Y_c_298_n 0.00376103f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_118 N_B1_c_124_n N_A_343_47#_c_331_n 0.00371445f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B1_c_125_n N_A_343_47#_c_331_n 0.0048014f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B1_M1005_g N_VGND_c_354_n 0.00585385f $X=1.64 $Y=0.56 $X2=0 $Y2=0
cc_121 N_B1_M1005_g N_VGND_c_356_n 0.0114525f $X=1.64 $Y=0.56 $X2=0 $Y2=0
cc_122 N_A2_M1009_g N_A1_M1000_g 0.0229885f $X=2.195 $Y=0.56 $X2=0 $Y2=0
cc_123 N_A2_c_160_n N_A1_M1000_g 0.00525794f $X=2.442 $Y=1.305 $X2=0 $Y2=0
cc_124 N_A2_M1008_g A1 2.15311e-19 $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A2_c_159_n A1 2.04949e-19 $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A2_c_160_n A1 0.0450995f $X=2.442 $Y=1.305 $X2=0 $Y2=0
cc_127 N_A2_M1008_g N_A1_c_197_n 0.0318348f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A2_c_159_n N_A1_c_197_n 0.0170516f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A2_M1008_g N_VPWR_c_225_n 0.00152974f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A2_M1008_g N_VPWR_c_230_n 0.00585385f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_131 A2 N_VPWR_c_230_n 0.0135336f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_132 N_A2_M1008_g N_VPWR_c_221_n 0.0113642f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_133 A2 N_VPWR_c_221_n 0.0125514f $X=2.445 $Y=2.125 $X2=0 $Y2=0
cc_134 N_A2_c_160_n N_Y_M1006_d 0.00202692f $X=2.442 $Y=1.305 $X2=0 $Y2=0
cc_135 N_A2_c_160_n N_Y_c_298_n 0.00695229f $X=2.442 $Y=1.305 $X2=0 $Y2=0
cc_136 A2 A_454_297# 0.0143594f $X=2.445 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_137 N_A2_c_160_n A_454_297# 0.00190855f $X=2.442 $Y=1.305 $X2=-0.19 $Y2=-0.24
cc_138 N_A2_c_160_n N_A_343_47#_c_331_n 0.00846891f $X=2.442 $Y=1.305 $X2=0
+ $Y2=0
cc_139 N_A2_M1009_g N_A_343_47#_c_329_n 0.0111755f $X=2.195 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A2_c_159_n N_A_343_47#_c_329_n 0.00106328f $X=2.285 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A2_c_160_n N_A_343_47#_c_329_n 0.0385903f $X=2.442 $Y=1.305 $X2=0 $Y2=0
cc_142 N_A2_M1009_g N_A_343_47#_c_330_n 5.62833e-19 $X=2.195 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A2_M1009_g N_VGND_c_353_n 0.00326685f $X=2.195 $Y=0.56 $X2=0 $Y2=0
cc_144 N_A2_M1009_g N_VGND_c_354_n 0.0042361f $X=2.195 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A2_M1009_g N_VGND_c_356_n 0.00617387f $X=2.195 $Y=0.56 $X2=0 $Y2=0
cc_146 A1 N_VPWR_M1001_d 0.00296264f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A1_M1001_g N_VPWR_c_225_n 0.0158096f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_148 A1 N_VPWR_c_225_n 0.0230817f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A1_c_197_n N_VPWR_c_225_n 0.00114781f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A1_M1001_g N_VPWR_c_230_n 0.00486043f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A1_M1001_g N_VPWR_c_221_n 0.00857998f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A1_M1000_g N_A_343_47#_c_329_n 0.0144721f $X=2.735 $Y=0.56 $X2=0 $Y2=0
cc_153 A1 N_A_343_47#_c_329_n 0.0258241f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A1_c_197_n N_A_343_47#_c_329_n 0.00212522f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A1_M1000_g N_A_343_47#_c_330_n 0.00561561f $X=2.735 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A1_M1000_g N_VGND_c_353_n 0.00433285f $X=2.735 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A1_M1000_g N_VGND_c_355_n 0.00414138f $X=2.735 $Y=0.56 $X2=0 $Y2=0
cc_158 N_A1_M1000_g N_VGND_c_356_n 0.00684473f $X=2.735 $Y=0.56 $X2=0 $Y2=0
cc_159 N_VPWR_c_221_n N_Y_M1007_d 0.00242341f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_160 N_VPWR_c_221_n N_Y_M1006_d 0.00426234f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_228_n N_Y_c_304_n 0.0140505f $X=1.21 $Y=2.72 $X2=0 $Y2=0
cc_162 N_VPWR_c_221_n N_Y_c_304_n 0.00897324f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_M1004_d N_Y_c_290_n 0.0109582f $X=1.175 $Y=1.485 $X2=0 $Y2=0
cc_164 N_VPWR_c_223_n N_Y_c_290_n 0.0167329f $X=1.375 $Y=2.34 $X2=0 $Y2=0
cc_165 N_VPWR_c_228_n N_Y_c_290_n 0.00247019f $X=1.21 $Y=2.72 $X2=0 $Y2=0
cc_166 N_VPWR_c_230_n N_Y_c_290_n 0.00268576f $X=2.785 $Y=2.72 $X2=0 $Y2=0
cc_167 N_VPWR_c_221_n N_Y_c_290_n 0.0108068f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_168 N_VPWR_c_230_n N_Y_c_311_n 0.0223083f $X=2.785 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_c_221_n N_Y_c_311_n 0.0132095f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_170 N_VPWR_M1007_s N_Y_c_276_n 0.00999205f $X=0.33 $Y=1.485 $X2=0 $Y2=0
cc_171 N_VPWR_c_222_n N_Y_c_276_n 0.019466f $X=0.455 $Y=2.34 $X2=0 $Y2=0
cc_172 N_VPWR_c_228_n N_Y_c_276_n 0.00218864f $X=1.21 $Y=2.72 $X2=0 $Y2=0
cc_173 N_VPWR_c_221_n N_Y_c_276_n 0.00525408f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_174 N_VPWR_c_222_n Y 0.00209642f $X=0.455 $Y=2.34 $X2=0 $Y2=0
cc_175 N_VPWR_c_226_n Y 0.00367525f $X=0.29 $Y=2.72 $X2=0 $Y2=0
cc_176 N_VPWR_c_221_n Y 0.00604532f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_177 N_VPWR_c_221_n A_454_297# 0.00484382f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_178 N_Y_c_275_n N_VGND_c_354_n 0.0406396f $X=0.525 $Y=0.4 $X2=0 $Y2=0
cc_179 N_Y_M1002_s N_VGND_c_356_n 0.00213418f $X=0.4 $Y=0.235 $X2=0 $Y2=0
cc_180 N_Y_c_275_n N_VGND_c_356_n 0.0230117f $X=0.525 $Y=0.4 $X2=0 $Y2=0
cc_181 A_163_47# N_VGND_c_356_n 0.00897657f $X=0.815 $Y=0.235 $X2=2.99 $Y2=0
cc_182 A_235_47# N_VGND_c_356_n 0.0104567f $X=1.175 $Y=0.235 $X2=1.19 $Y2=1.16
cc_183 N_A_343_47#_c_329_n N_VGND_M1009_d 0.00584429f $X=2.785 $Y=0.725
+ $X2=-0.19 $Y2=-0.24
cc_184 N_A_343_47#_c_329_n N_VGND_c_353_n 0.0212136f $X=2.785 $Y=0.725 $X2=0
+ $Y2=0
cc_185 N_A_343_47#_c_344_p N_VGND_c_354_n 0.0220464f $X=1.93 $Y=0.4 $X2=0 $Y2=0
cc_186 N_A_343_47#_c_329_n N_VGND_c_354_n 0.00292296f $X=2.785 $Y=0.725 $X2=0
+ $Y2=0
cc_187 N_A_343_47#_c_329_n N_VGND_c_355_n 0.00255018f $X=2.785 $Y=0.725 $X2=0
+ $Y2=0
cc_188 N_A_343_47#_c_330_n N_VGND_c_355_n 0.0208048f $X=2.95 $Y=0.4 $X2=0 $Y2=0
cc_189 N_A_343_47#_M1005_d N_VGND_c_356_n 0.00456992f $X=1.715 $Y=0.235 $X2=0
+ $Y2=0
cc_190 N_A_343_47#_M1000_d N_VGND_c_356_n 0.00213418f $X=2.81 $Y=0.235 $X2=0
+ $Y2=0
cc_191 N_A_343_47#_c_344_p N_VGND_c_356_n 0.0131491f $X=1.93 $Y=0.4 $X2=0 $Y2=0
cc_192 N_A_343_47#_c_329_n N_VGND_c_356_n 0.0103582f $X=2.785 $Y=0.725 $X2=0
+ $Y2=0
cc_193 N_A_343_47#_c_330_n N_VGND_c_356_n 0.0123922f $X=2.95 $Y=0.4 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a211oi_4.pxi.spice
* Created: Thu Aug 27 13:59:56 2020
* 
x_PM_SKY130_FD_SC_HD__A211OI_4%A2 N_A2_M1009_g N_A2_M16_noxref_g N_A2_M1018_g
+ N_A2_M17_noxref_g N_A2_M1025_g N_A2_M18_noxref_g N_A2_c_120_n N_A2_M1030_g
+ N_A2_M23_noxref_g N_A2_c_130_n N_A2_c_121_n N_A2_c_122_n A2 N_A2_c_123_n
+ N_A2_c_124_n A2 N_A2_c_125_n PM_SKY130_FD_SC_HD__A211OI_4%A2
x_PM_SKY130_FD_SC_HD__A211OI_4%A1 N_A1_M1013_g N_A1_M19_noxref_g N_A1_M1014_g
+ N_A1_M20_noxref_g N_A1_M1020_g N_A1_M21_noxref_g N_A1_M1024_g
+ N_A1_M22_noxref_g A1 N_A1_c_245_n N_A1_c_263_n N_A1_c_246_n
+ PM_SKY130_FD_SC_HD__A211OI_4%A1
x_PM_SKY130_FD_SC_HD__A211OI_4%B1 N_B1_c_310_n N_B1_M1002_g N_B1_M24_noxref_g
+ N_B1_M25_noxref_g N_B1_c_311_n N_B1_M1006_g N_B1_M26_noxref_g N_B1_c_312_n
+ N_B1_M1023_g N_B1_M1026_g N_B1_M31_noxref_g N_B1_c_348_p N_B1_c_313_n
+ N_B1_c_314_n N_B1_c_324_n N_B1_c_332_n N_B1_c_325_n N_B1_c_326_n B1
+ N_B1_c_315_n N_B1_c_316_n N_B1_c_317_n PM_SKY130_FD_SC_HD__A211OI_4%B1
x_PM_SKY130_FD_SC_HD__A211OI_4%C1 N_C1_M27_noxref_g N_C1_c_450_n N_C1_M1015_g
+ N_C1_M28_noxref_g N_C1_c_451_n N_C1_M1021_g N_C1_M29_noxref_g N_C1_c_452_n
+ N_C1_M1027_g N_C1_c_453_n N_C1_M1031_g N_C1_M30_noxref_g N_C1_c_454_n
+ N_C1_c_460_n C1 N_C1_c_455_n PM_SKY130_FD_SC_HD__A211OI_4%C1
x_PM_SKY130_FD_SC_HD__A211OI_4%noxref_7 N_noxref_7_M16_noxref_s
+ N_noxref_7_M17_noxref_d N_noxref_7_M19_noxref_d N_noxref_7_M21_noxref_d
+ N_noxref_7_M23_noxref_d N_noxref_7_M25_noxref_d N_noxref_7_M31_noxref_d
+ N_noxref_7_c_539_n N_noxref_7_c_540_n N_noxref_7_c_549_n N_noxref_7_c_588_p
+ N_noxref_7_c_553_n N_noxref_7_c_591_p N_noxref_7_c_555_n N_noxref_7_c_594_p
+ N_noxref_7_c_556_n N_noxref_7_c_558_n N_noxref_7_c_599_p N_noxref_7_c_541_n
+ N_noxref_7_c_559_n N_noxref_7_c_561_n N_noxref_7_c_562_n
+ PM_SKY130_FD_SC_HD__A211OI_4%noxref_7
x_PM_SKY130_FD_SC_HD__A211OI_4%VPWR N_VPWR_M16_noxref_d N_VPWR_M18_noxref_d
+ N_VPWR_M20_noxref_d N_VPWR_M22_noxref_d N_VPWR_c_634_n N_VPWR_c_635_n
+ N_VPWR_c_636_n N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n
+ N_VPWR_c_641_n N_VPWR_c_642_n N_VPWR_c_643_n VPWR N_VPWR_c_644_n
+ N_VPWR_c_645_n N_VPWR_c_633_n N_VPWR_c_647_n PM_SKY130_FD_SC_HD__A211OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A211OI_4%noxref_9 N_noxref_9_M24_noxref_d
+ N_noxref_9_M28_noxref_d N_noxref_9_c_749_n N_noxref_9_c_745_n
+ N_noxref_9_c_746_n PM_SKY130_FD_SC_HD__A211OI_4%noxref_9
x_PM_SKY130_FD_SC_HD__A211OI_4%Y N_Y_M1013_d N_Y_M1020_d N_Y_M1002_d N_Y_M1023_d
+ N_Y_M1021_d N_Y_M1031_d N_Y_M27_noxref_d N_Y_M29_noxref_d N_Y_c_800_n
+ N_Y_c_801_n N_Y_c_803_n N_Y_c_819_n N_Y_c_905_p N_Y_c_852_n N_Y_c_824_n
+ N_Y_c_912_p N_Y_c_829_n N_Y_c_794_n N_Y_c_804_n N_Y_c_806_n N_Y_c_839_n
+ N_Y_c_870_n N_Y_c_872_n N_Y_c_796_n N_Y_c_795_n Y N_Y_c_799_n
+ PM_SKY130_FD_SC_HD__A211OI_4%Y
x_PM_SKY130_FD_SC_HD__A211OI_4%VGND N_VGND_M1009_d N_VGND_M1018_d N_VGND_M1030_d
+ N_VGND_M1006_s N_VGND_M1015_s N_VGND_M1027_s N_VGND_M1026_s N_VGND_c_942_n
+ N_VGND_c_943_n N_VGND_c_944_n N_VGND_c_945_n N_VGND_c_946_n N_VGND_c_947_n
+ N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n N_VGND_c_952_n
+ N_VGND_c_953_n N_VGND_c_954_n VGND N_VGND_c_955_n N_VGND_c_956_n
+ N_VGND_c_957_n N_VGND_c_958_n N_VGND_c_959_n N_VGND_c_960_n N_VGND_c_961_n
+ N_VGND_c_962_n PM_SKY130_FD_SC_HD__A211OI_4%VGND
x_PM_SKY130_FD_SC_HD__A211OI_4%A_109_47# N_A_109_47#_M1009_s N_A_109_47#_M1025_s
+ N_A_109_47#_M1014_s N_A_109_47#_M1024_s N_A_109_47#_c_1068_n
+ N_A_109_47#_c_1074_n N_A_109_47#_c_1075_n N_A_109_47#_c_1077_n
+ N_A_109_47#_c_1078_n PM_SKY130_FD_SC_HD__A211OI_4%A_109_47#
cc_1 VNB N_A2_M1009_g 0.0243492f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A2_M16_noxref_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_3 VNB N_A2_M1018_g 0.0173626f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_4 VNB N_A2_M17_noxref_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_5 VNB N_A2_M1025_g 0.017802f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_6 VNB N_A2_M18_noxref_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_7 VNB N_A2_c_120_n 0.0164935f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.995
cc_8 VNB N_A2_c_121_n 0.00412892f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.16
cc_9 VNB N_A2_c_122_n 0.0185317f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.16
cc_10 VNB N_A2_c_123_n 0.0509684f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_11 VNB N_A2_c_124_n 0.0157817f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.33
cc_12 VNB N_A2_c_125_n 0.00216106f $X=-0.19 $Y=-0.24 $X2=1.385 $Y2=1.33
cc_13 VNB N_A1_M1013_g 0.017802f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_14 VNB N_A1_M19_noxref_g 4.64343e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_15 VNB N_A1_M1014_g 0.017506f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_16 VNB N_A1_M20_noxref_g 4.50136e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_17 VNB N_A1_M1020_g 0.017506f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_18 VNB N_A1_M21_noxref_g 4.5006e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_19 VNB N_A1_M1024_g 0.0177319f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.56
cc_20 VNB N_A1_M22_noxref_g 4.42713e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A1_c_245_n 0.00128095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A1_c_246_n 0.0617851f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_23 VNB N_B1_c_310_n 0.0168703f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_24 VNB N_B1_c_311_n 0.0165272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_B1_c_312_n 0.0161977f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_26 VNB N_B1_c_313_n 0.00332507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_B1_c_314_n 0.0224282f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.445
cc_28 VNB N_B1_c_315_n 0.0500449f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.33
cc_29 VNB N_B1_c_316_n 0.0187792f $X=-0.19 $Y=-0.24 $X2=1.165 $Y2=1.33
cc_30 VNB N_B1_c_317_n 0.00176906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_C1_c_450_n 0.0160696f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_32 VNB N_C1_c_451_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_C1_c_452_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_34 VNB N_C1_c_453_n 0.0161143f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_35 VNB N_C1_c_454_n 0.00215472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_C1_c_455_n 0.0655433f $X=-0.19 $Y=-0.24 $X2=1.22 $Y2=1.16
cc_37 VNB N_VPWR_c_633_n 0.30769f $X=-0.19 $Y=-0.24 $X2=1.165 $Y2=1.33
cc_38 VNB N_Y_c_794_n 0.00937344f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.33
cc_39 VNB N_Y_c_795_n 0.0219013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_942_n 0.0109754f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_41 VNB N_VGND_c_943_n 0.0185677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_944_n 0.00222423f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.325
cc_43 VNB N_VGND_c_945_n 0.0040921f $X=-0.19 $Y=-0.24 $X2=3.245 $Y2=1.535
cc_44 VNB N_VGND_c_946_n 0.0153014f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.445
cc_45 VNB N_VGND_c_947_n 3.27959e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_948_n 0.0111906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_949_n 3.03604e-19 $X=-0.19 $Y=-0.24 $X2=0.88 $Y2=1.16
cc_48 VNB N_VGND_c_950_n 3.05427e-19 $X=-0.19 $Y=-0.24 $X2=1.22 $Y2=1.16
cc_49 VNB N_VGND_c_951_n 0.0106585f $X=-0.19 $Y=-0.24 $X2=1.22 $Y2=1.16
cc_50 VNB N_VGND_c_952_n 0.0114478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_953_n 0.0537997f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.33
cc_52 VNB N_VGND_c_954_n 0.00323548f $X=-0.19 $Y=-0.24 $X2=0.88 $Y2=1.33
cc_53 VNB N_VGND_c_955_n 0.0147118f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.33
cc_54 VNB N_VGND_c_956_n 0.0109187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_957_n 0.0122674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_958_n 0.00333399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_959_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_960_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_961_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_962_n 0.350921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VPB N_A2_M16_noxref_g 0.0233062f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_62 VPB N_A2_M17_noxref_g 0.0177798f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_63 VPB N_A2_M18_noxref_g 0.0178048f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_64 VPB N_A2_M23_noxref_g 0.0169708f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_65 VPB N_A2_c_130_n 0.0147256f $X=-0.19 $Y=1.305 $X2=3.245 $Y2=1.535
cc_66 VPB N_A2_c_121_n 0.00227281f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.16
cc_67 VPB N_A2_c_122_n 0.00441099f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.16
cc_68 VPB N_A2_c_124_n 0.0141397f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.33
cc_69 VPB N_A2_c_125_n 0.00172186f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=1.33
cc_70 VPB N_A1_M19_noxref_g 0.0191776f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_71 VPB N_A1_M20_noxref_g 0.0189431f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_72 VPB N_A1_M21_noxref_g 0.0189419f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_73 VPB N_A1_M22_noxref_g 0.0191204f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B1_M24_noxref_g 0.0172006f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_75 VPB N_B1_M25_noxref_g 0.0171196f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_76 VPB N_B1_M26_noxref_g 0.0187667f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_77 VPB N_B1_M31_noxref_g 0.0223521f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=0.56
cc_78 VPB N_B1_c_313_n 4.1497e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_B1_c_314_n 0.00494045f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.445
cc_80 VPB N_B1_c_324_n 0.00238359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_B1_c_325_n 0.00143589f $X=-0.19 $Y=1.305 $X2=0.88 $Y2=1.16
cc_82 VPB N_B1_c_326_n 0.00234886f $X=-0.19 $Y=1.305 $X2=0.88 $Y2=1.16
cc_83 VPB N_B1_c_315_n 0.00996356f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.33
cc_84 VPB N_B1_c_317_n 0.00265396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_C1_M27_noxref_g 0.0188589f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_86 VPB N_C1_M28_noxref_g 0.0183752f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_87 VPB N_C1_M29_noxref_g 0.0186533f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.025
cc_88 VPB N_C1_M30_noxref_g 0.0192996f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=0.56
cc_89 VPB N_C1_c_460_n 0.00223318f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=1.535
cc_90 VPB N_C1_c_455_n 0.0124647f $X=-0.19 $Y=1.305 $X2=1.22 $Y2=1.16
cc_91 VPB N_noxref_7_c_539_n 0.0125686f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_92 VPB N_noxref_7_c_540_n 0.0144536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_noxref_7_c_541_n 0.00955326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_634_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_95 VPB N_VPWR_c_635_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_96 VPB N_VPWR_c_636_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_97 VPB N_VPWR_c_637_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=3.41 $Y2=0.56
cc_98 VPB N_VPWR_c_638_n 0.0109337f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_99 VPB N_VPWR_c_639_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_640_n 0.0109033f $X=-0.19 $Y=1.305 $X2=1.385 $Y2=1.535
cc_101 VPB N_VPWR_c_641_n 0.00436029f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.445
cc_102 VPB N_VPWR_c_642_n 0.0109033f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.16
cc_103 VPB N_VPWR_c_643_n 0.00436029f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.16
cc_104 VPB N_VPWR_c_644_n 0.0143745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_645_n 0.0912487f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.53
cc_106 VPB N_VPWR_c_633_n 0.0444431f $X=-0.19 $Y=1.305 $X2=1.165 $Y2=1.33
cc_107 VPB N_VPWR_c_647_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_noxref_9_c_745_n 0.00632438f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.295
cc_109 VPB N_noxref_9_c_746_n 0.00213042f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_110 VPB N_Y_c_796_n 0.00675691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_Y_c_795_n 0.00860934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB Y 0.00769973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_Y_c_799_n 0.00974655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 N_A2_M1025_g N_A1_M1013_g 0.0295534f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A2_M18_noxref_g N_A1_M19_noxref_g 0.0295534f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A2_c_130_n N_A1_M19_noxref_g 0.0107047f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_117 N_A2_c_130_n N_A1_M20_noxref_g 0.0107506f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_118 N_A2_c_130_n N_A1_M21_noxref_g 0.0107506f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_119 N_A2_c_120_n N_A1_M1024_g 0.028776f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A2_c_122_n N_A1_M1024_g 0.0218068f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A2_M23_noxref_g N_A1_M22_noxref_g 0.0458735f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A2_c_130_n N_A1_M22_noxref_g 0.0114935f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_123 N_A2_c_130_n N_A1_c_245_n 0.00873663f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_124 N_A2_c_123_n N_A1_c_245_n 3.00961e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A2_c_125_n N_A1_c_245_n 0.0138708f $X=1.385 $Y=1.33 $X2=0 $Y2=0
cc_126 N_A2_c_130_n N_A1_c_263_n 0.0886865f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_127 N_A2_c_121_n N_A1_c_263_n 0.015406f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A2_c_122_n N_A1_c_263_n 2.57681e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A2_c_130_n N_A1_c_246_n 0.00595574f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_130 N_A2_c_121_n N_A1_c_246_n 0.00562222f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A2_c_123_n N_A1_c_246_n 0.0295534f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A2_c_125_n N_A1_c_246_n 0.00160383f $X=1.385 $Y=1.33 $X2=0 $Y2=0
cc_133 N_A2_c_120_n N_B1_c_310_n 0.0281328f $X=3.41 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_134 N_A2_M23_noxref_g N_B1_M24_noxref_g 0.0281563f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A2_c_130_n N_B1_M24_noxref_g 9.54768e-19 $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_136 N_A2_c_130_n N_B1_c_332_n 0.00186069f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_137 N_A2_c_121_n N_B1_c_332_n 2.19649e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A2_c_121_n N_B1_c_315_n 0.00132623f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A2_c_122_n N_B1_c_315_n 0.0219965f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A2_M23_noxref_g N_B1_c_317_n 6.02781e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A2_c_130_n N_B1_c_317_n 0.00817198f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_142 N_A2_c_121_n N_B1_c_317_n 0.0359707f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A2_c_122_n N_B1_c_317_n 0.0010206f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A2_c_124_n N_noxref_7_M16_noxref_s 0.0028575f $X=1.09 $Y=1.33 $X2=-0.19
+ $Y2=-0.24
cc_145 N_A2_c_124_n N_noxref_7_M17_noxref_d 7.39973e-19 $X=1.09 $Y=1.33 $X2=0
+ $Y2=0
cc_146 N_A2_c_125_n N_noxref_7_M17_noxref_d 9.71905e-19 $X=1.385 $Y=1.33 $X2=0
+ $Y2=0
cc_147 N_A2_c_130_n N_noxref_7_M19_noxref_d 0.00166124f $X=3.245 $Y=1.535 $X2=0
+ $Y2=0
cc_148 N_A2_c_130_n N_noxref_7_M21_noxref_d 0.00166124f $X=3.245 $Y=1.535 $X2=0
+ $Y2=0
cc_149 N_A2_c_130_n N_noxref_7_M23_noxref_d 0.00143429f $X=3.245 $Y=1.535 $X2=0
+ $Y2=0
cc_150 N_A2_c_124_n N_noxref_7_c_539_n 0.0212345f $X=1.09 $Y=1.33 $X2=0 $Y2=0
cc_151 N_A2_M16_noxref_g N_noxref_7_c_549_n 0.0125846f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A2_M17_noxref_g N_noxref_7_c_549_n 0.0125846f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A2_c_123_n N_noxref_7_c_549_n 3.27531e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A2_c_124_n N_noxref_7_c_549_n 0.036224f $X=1.09 $Y=1.33 $X2=0 $Y2=0
cc_155 N_A2_M18_noxref_g N_noxref_7_c_553_n 0.0129515f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A2_c_125_n N_noxref_7_c_553_n 0.0342673f $X=1.385 $Y=1.33 $X2=0 $Y2=0
cc_157 N_A2_c_130_n N_noxref_7_c_555_n 0.0332445f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_158 N_A2_M23_noxref_g N_noxref_7_c_556_n 0.0129452f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A2_c_130_n N_noxref_7_c_556_n 0.0345375f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_160 N_A2_c_130_n N_noxref_7_c_558_n 0.00294201f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_161 N_A2_c_123_n N_noxref_7_c_559_n 3.64505e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A2_c_124_n N_noxref_7_c_559_n 0.0137945f $X=1.09 $Y=1.33 $X2=0 $Y2=0
cc_163 N_A2_c_130_n N_noxref_7_c_561_n 0.0127256f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_164 N_A2_c_130_n N_noxref_7_c_562_n 0.0127256f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_165 N_A2_c_124_n N_VPWR_M16_noxref_d 0.00172715f $X=1.09 $Y=1.33 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A2_c_130_n N_VPWR_M18_noxref_d 0.00166529f $X=3.245 $Y=1.535 $X2=0
+ $Y2=0
cc_167 N_A2_c_130_n N_VPWR_M20_noxref_d 0.00166529f $X=3.245 $Y=1.535 $X2=0
+ $Y2=0
cc_168 N_A2_c_130_n N_VPWR_M22_noxref_d 0.0016558f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_169 N_A2_M16_noxref_g N_VPWR_c_634_n 0.00834749f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A2_M17_noxref_g N_VPWR_c_634_n 0.00664421f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A2_M18_noxref_g N_VPWR_c_634_n 5.08801e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A2_M17_noxref_g N_VPWR_c_635_n 5.02907e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A2_M18_noxref_g N_VPWR_c_635_n 0.00640108f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A2_M23_noxref_g N_VPWR_c_637_n 0.00759476f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A2_M17_noxref_g N_VPWR_c_638_n 0.00339367f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A2_M18_noxref_g N_VPWR_c_638_n 0.00337001f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A2_M16_noxref_g N_VPWR_c_644_n 0.00339367f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A2_M23_noxref_g N_VPWR_c_645_n 0.00337001f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A2_M16_noxref_g N_VPWR_c_633_n 0.00489827f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A2_M17_noxref_g N_VPWR_c_633_n 0.00394406f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A2_M18_noxref_g N_VPWR_c_633_n 0.00390568f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A2_M23_noxref_g N_VPWR_c_633_n 0.00393288f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A2_c_130_n N_Y_c_800_n 0.0062004f $X=3.245 $Y=1.535 $X2=0 $Y2=0
cc_184 N_A2_c_120_n N_Y_c_801_n 0.0115989f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A2_c_122_n N_Y_c_801_n 0.00127448f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_c_120_n N_Y_c_803_n 4.57554e-19 $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A2_c_121_n N_Y_c_804_n 0.0212409f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A2_c_122_n N_Y_c_804_n 0.00127466f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A2_c_120_n N_Y_c_806_n 3.55166e-19 $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A2_M1009_g N_VGND_c_943_n 0.0036131f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A2_c_124_n N_VGND_c_943_n 0.0119939f $X=1.09 $Y=1.33 $X2=0 $Y2=0
cc_192 N_A2_M1009_g N_VGND_c_944_n 0.00122355f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A2_M1018_g N_VGND_c_944_n 0.00816829f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A2_M1025_g N_VGND_c_944_n 0.00277851f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A2_c_120_n N_VGND_c_945_n 0.00268723f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_M1025_g N_VGND_c_953_n 0.00418507f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A2_c_120_n N_VGND_c_953_n 0.00418549f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_M1009_g N_VGND_c_955_n 0.00583607f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A2_M1018_g N_VGND_c_955_n 0.00389579f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A2_M1009_g N_VGND_c_962_n 0.0114285f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A2_M1018_g N_VGND_c_962_n 0.00454817f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A2_M1025_g N_VGND_c_962_n 0.00569347f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A2_c_120_n N_VGND_c_962_n 0.00572071f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_M1018_g N_A_109_47#_c_1068_n 0.00977774f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A2_M1025_g N_A_109_47#_c_1068_n 0.010724f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A2_c_130_n N_A_109_47#_c_1068_n 0.0063014f $X=3.245 $Y=1.535 $X2=0
+ $Y2=0
cc_207 N_A2_c_123_n N_A_109_47#_c_1068_n 0.00195929f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A2_c_124_n N_A_109_47#_c_1068_n 0.0384914f $X=1.09 $Y=1.33 $X2=0 $Y2=0
cc_209 N_A2_c_125_n N_A_109_47#_c_1068_n 0.00247908f $X=1.385 $Y=1.33 $X2=0
+ $Y2=0
cc_210 N_A2_M1025_g N_A_109_47#_c_1074_n 0.00286712f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A2_M1018_g N_A_109_47#_c_1075_n 4.5955e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_212 N_A2_M1025_g N_A_109_47#_c_1075_n 0.00455129f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_213 N_A2_c_120_n N_A_109_47#_c_1077_n 0.00327517f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A2_c_123_n N_A_109_47#_c_1078_n 0.00199473f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A2_c_124_n N_A_109_47#_c_1078_n 0.0148737f $X=1.09 $Y=1.33 $X2=0 $Y2=0
cc_216 N_A1_M19_noxref_g N_noxref_7_c_553_n 0.0129515f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A1_M20_noxref_g N_noxref_7_c_555_n 0.0130325f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A1_M21_noxref_g N_noxref_7_c_555_n 0.0130325f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A1_M22_noxref_g N_noxref_7_c_556_n 0.0129515f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A1_M19_noxref_g N_VPWR_c_635_n 0.00640108f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A1_M20_noxref_g N_VPWR_c_635_n 5.02907e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A1_M19_noxref_g N_VPWR_c_636_n 5.02907e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A1_M20_noxref_g N_VPWR_c_636_n 0.00643498f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A1_M21_noxref_g N_VPWR_c_636_n 0.00643498f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A1_M22_noxref_g N_VPWR_c_636_n 5.02907e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A1_M21_noxref_g N_VPWR_c_637_n 5.02907e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A1_M22_noxref_g N_VPWR_c_637_n 0.00640108f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A1_M19_noxref_g N_VPWR_c_640_n 0.00337001f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A1_M20_noxref_g N_VPWR_c_640_n 0.00337001f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A1_M21_noxref_g N_VPWR_c_642_n 0.00337001f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_M22_noxref_g N_VPWR_c_642_n 0.00337001f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A1_M19_noxref_g N_VPWR_c_633_n 0.00390568f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_M20_noxref_g N_VPWR_c_633_n 0.00390568f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A1_M21_noxref_g N_VPWR_c_633_n 0.00390568f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A1_M22_noxref_g N_VPWR_c_633_n 0.00390568f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A1_M1013_g N_Y_c_800_n 0.00275946f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A1_M1014_g N_Y_c_800_n 0.00889421f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_238 N_A1_M1020_g N_Y_c_800_n 0.00889421f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_239 N_A1_M1024_g N_Y_c_800_n 0.00960368f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_240 N_A1_c_245_n N_Y_c_800_n 3.52947e-19 $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A1_c_263_n N_Y_c_800_n 0.0751905f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A1_c_246_n N_Y_c_800_n 0.00589357f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A1_M1013_g N_VGND_c_953_n 0.00357877f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_244 N_A1_M1014_g N_VGND_c_953_n 0.00357877f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_245 N_A1_M1020_g N_VGND_c_953_n 0.00357877f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A1_M1024_g N_VGND_c_953_n 0.00357877f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A1_M1013_g N_VGND_c_962_n 0.00525237f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A1_M1014_g N_VGND_c_962_n 0.00522516f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A1_M1020_g N_VGND_c_962_n 0.00522516f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A1_M1024_g N_VGND_c_962_n 0.00525237f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_251 N_A1_M1013_g N_A_109_47#_c_1077_n 0.0110389f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A1_M1014_g N_A_109_47#_c_1077_n 0.00970685f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A1_M1020_g N_A_109_47#_c_1077_n 0.00970685f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A1_M1024_g N_A_109_47#_c_1077_n 0.00970685f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A1_c_245_n N_A_109_47#_c_1077_n 0.0033735f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_M26_noxref_g N_C1_M27_noxref_g 0.0536525f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_B1_c_312_n N_C1_c_450_n 0.0123011f $X=4.745 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B1_c_324_n N_C1_M29_noxref_g 0.00272354f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_259 N_B1_c_316_n N_C1_c_453_n 0.0253187f $X=6.852 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B1_M31_noxref_g N_C1_M30_noxref_g 0.0528792f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_261 N_B1_c_324_n N_C1_M30_noxref_g 0.00979653f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_262 N_B1_c_325_n N_C1_M30_noxref_g 0.00154686f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_263 N_B1_c_326_n N_C1_M30_noxref_g 0.0020707f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_264 N_B1_c_348_p N_C1_c_454_n 0.0161108f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_265 N_B1_c_324_n N_C1_c_454_n 0.0116052f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_266 N_B1_c_315_n N_C1_c_454_n 0.00185061f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B1_c_313_n N_C1_c_460_n 0.0185481f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B1_c_324_n N_C1_c_460_n 0.0135717f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_269 N_B1_c_325_n N_C1_c_460_n 0.00280085f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_270 N_B1_c_326_n N_C1_c_460_n 0.01337f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_271 N_B1_c_348_p N_C1_c_455_n 2.52572e-19 $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_c_313_n N_C1_c_455_n 0.00351952f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_273 N_B1_c_314_n N_C1_c_455_n 0.0216302f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B1_c_315_n N_C1_c_455_n 0.0233896f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_275 N_B1_c_324_n N_noxref_7_M25_noxref_d 0.00108324f $X=6.53 $Y=1.53 $X2=0
+ $Y2=0
cc_276 N_B1_c_317_n N_noxref_7_M25_noxref_d 0.00152787f $X=4.46 $Y=1.325 $X2=0
+ $Y2=0
cc_277 N_B1_M24_noxref_g N_noxref_7_c_541_n 0.0103545f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_278 N_B1_M25_noxref_g N_noxref_7_c_541_n 0.00861238f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_279 N_B1_M26_noxref_g N_noxref_7_c_541_n 0.00881116f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_B1_M31_noxref_g N_noxref_7_c_541_n 0.00889686f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_B1_c_332_n N_noxref_7_c_541_n 0.00198712f $X=4.06 $Y=1.53 $X2=0 $Y2=0
cc_282 N_B1_c_317_n N_noxref_7_c_541_n 0.00153958f $X=4.46 $Y=1.325 $X2=0 $Y2=0
cc_283 N_B1_M24_noxref_g N_VPWR_c_637_n 0.00110007f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B1_M24_noxref_g N_VPWR_c_645_n 0.00357877f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_285 N_B1_M25_noxref_g N_VPWR_c_645_n 0.00357877f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_286 N_B1_M26_noxref_g N_VPWR_c_645_n 0.00357877f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_287 N_B1_M31_noxref_g N_VPWR_c_645_n 0.00357877f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_288 N_B1_M24_noxref_g N_VPWR_c_633_n 0.00525237f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_289 N_B1_M25_noxref_g N_VPWR_c_633_n 0.00522516f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_290 N_B1_M26_noxref_g N_VPWR_c_633_n 0.00531933f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_291 N_B1_M31_noxref_g N_VPWR_c_633_n 0.00630671f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_292 N_B1_c_332_n N_noxref_9_M24_noxref_d 0.00166705f $X=4.06 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_293 N_B1_c_317_n N_noxref_9_M24_noxref_d 0.00110785f $X=4.46 $Y=1.325
+ $X2=-0.19 $Y2=-0.24
cc_294 N_B1_M24_noxref_g N_noxref_9_c_749_n 0.00421954f $X=3.83 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_B1_M25_noxref_g N_noxref_9_c_749_n 0.0119464f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_B1_M26_noxref_g N_noxref_9_c_749_n 0.00663528f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_B1_c_348_p N_noxref_9_c_749_n 0.00189129f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_298 N_B1_c_324_n N_noxref_9_c_749_n 0.00803351f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_299 N_B1_c_332_n N_noxref_9_c_749_n 0.00519502f $X=4.06 $Y=1.53 $X2=0 $Y2=0
cc_300 N_B1_c_315_n N_noxref_9_c_749_n 0.00143028f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_301 N_B1_c_317_n N_noxref_9_c_749_n 0.0304533f $X=4.46 $Y=1.325 $X2=0 $Y2=0
cc_302 N_B1_M26_noxref_g N_noxref_9_c_745_n 2.69506e-19 $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_B1_c_324_n N_noxref_9_c_745_n 0.0507522f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_304 N_B1_M25_noxref_g N_noxref_9_c_746_n 0.00141078f $X=4.25 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_B1_M26_noxref_g N_noxref_9_c_746_n 0.0188666f $X=4.67 $Y=1.985 $X2=0
+ $Y2=0
cc_306 N_B1_c_348_p N_noxref_9_c_746_n 0.00886294f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_307 N_B1_c_324_n N_noxref_9_c_746_n 0.0232691f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_308 N_B1_c_332_n N_noxref_9_c_746_n 0.00106885f $X=4.06 $Y=1.53 $X2=0 $Y2=0
cc_309 N_B1_c_315_n N_noxref_9_c_746_n 0.00256547f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_310 N_B1_c_317_n N_noxref_9_c_746_n 0.011957f $X=4.46 $Y=1.325 $X2=0 $Y2=0
cc_311 N_B1_c_324_n N_Y_M29_noxref_d 6.70552e-19 $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_312 N_B1_c_310_n N_Y_c_801_n 0.00832889f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B1_c_332_n N_Y_c_801_n 3.37147e-19 $X=4.06 $Y=1.53 $X2=0 $Y2=0
cc_314 N_B1_c_317_n N_Y_c_801_n 0.00918679f $X=4.46 $Y=1.325 $X2=0 $Y2=0
cc_315 N_B1_c_310_n N_Y_c_803_n 0.00468937f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B1_c_311_n N_Y_c_819_n 0.0115999f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B1_c_312_n N_Y_c_819_n 0.0122125f $X=4.745 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_324_n N_Y_c_819_n 0.00174752f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_319 N_B1_c_315_n N_Y_c_819_n 0.00268078f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_320 N_B1_c_317_n N_Y_c_819_n 0.03541f $X=4.46 $Y=1.325 $X2=0 $Y2=0
cc_321 N_B1_M31_noxref_g N_Y_c_824_n 0.00963234f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_322 N_B1_c_313_n N_Y_c_824_n 0.0034881f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_323 N_B1_c_324_n N_Y_c_824_n 0.016947f $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_324 N_B1_c_325_n N_Y_c_824_n 0.00928386f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_325 N_B1_c_326_n N_Y_c_824_n 0.00728805f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_326 N_B1_c_324_n N_Y_c_829_n 9.92915e-19 $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_327 N_B1_c_313_n N_Y_c_794_n 0.0235262f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_328 N_B1_c_314_n N_Y_c_794_n 0.00144581f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_329 N_B1_c_325_n N_Y_c_794_n 0.00198287f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_330 N_B1_c_316_n N_Y_c_794_n 0.0123625f $X=6.852 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B1_c_310_n N_Y_c_806_n 0.00242778f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B1_c_324_n N_Y_c_806_n 5.08128e-19 $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_333 N_B1_c_332_n N_Y_c_806_n 7.20097e-19 $X=4.06 $Y=1.53 $X2=0 $Y2=0
cc_334 N_B1_c_315_n N_Y_c_806_n 0.00403832f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_335 N_B1_c_317_n N_Y_c_806_n 0.0235246f $X=4.46 $Y=1.325 $X2=0 $Y2=0
cc_336 N_B1_c_324_n N_Y_c_839_n 9.96425e-19 $X=6.53 $Y=1.53 $X2=0 $Y2=0
cc_337 N_B1_M31_noxref_g N_Y_c_796_n 0.00646907f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_338 N_B1_c_325_n N_Y_c_796_n 0.00468212f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_339 N_B1_c_326_n N_Y_c_796_n 0.00570118f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_340 N_B1_M31_noxref_g N_Y_c_795_n 0.00369184f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_341 N_B1_c_313_n N_Y_c_795_n 0.0248551f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_342 N_B1_c_314_n N_Y_c_795_n 0.00763345f $X=6.85 $Y=1.16 $X2=0 $Y2=0
cc_343 N_B1_c_325_n N_Y_c_795_n 0.00201895f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_344 N_B1_c_326_n N_Y_c_795_n 0.00655305f $X=6.675 $Y=1.53 $X2=0 $Y2=0
cc_345 N_B1_c_316_n N_Y_c_795_n 0.005786f $X=6.852 $Y=0.995 $X2=0 $Y2=0
cc_346 N_B1_M31_noxref_g Y 0.0078069f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_347 N_B1_M31_noxref_g N_Y_c_799_n 0.00567077f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_348 N_B1_c_324_n noxref_12 2.11753e-19 $X=6.53 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_349 N_B1_c_325_n noxref_12 0.00287969f $X=6.675 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_350 N_B1_c_326_n noxref_12 0.00297068f $X=6.675 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_351 N_B1_c_310_n N_VGND_c_945_n 0.00145354f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_352 N_B1_c_310_n N_VGND_c_946_n 0.00420025f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_353 N_B1_c_311_n N_VGND_c_946_n 0.00351072f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_354 N_B1_c_310_n N_VGND_c_947_n 4.62158e-19 $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_355 N_B1_c_311_n N_VGND_c_947_n 0.00656161f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_356 N_B1_c_312_n N_VGND_c_947_n 0.00627278f $X=4.745 $Y=0.995 $X2=0 $Y2=0
cc_357 N_B1_c_312_n N_VGND_c_948_n 0.00351072f $X=4.745 $Y=0.995 $X2=0 $Y2=0
cc_358 N_B1_c_312_n N_VGND_c_949_n 5.03945e-19 $X=4.745 $Y=0.995 $X2=0 $Y2=0
cc_359 N_B1_c_316_n N_VGND_c_950_n 0.00105539f $X=6.852 $Y=0.995 $X2=0 $Y2=0
cc_360 N_B1_c_316_n N_VGND_c_952_n 0.00849116f $X=6.852 $Y=0.995 $X2=0 $Y2=0
cc_361 N_B1_c_316_n N_VGND_c_957_n 0.00365142f $X=6.852 $Y=0.995 $X2=0 $Y2=0
cc_362 N_B1_c_310_n N_VGND_c_962_n 0.00584714f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_363 N_B1_c_311_n N_VGND_c_962_n 0.00420947f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_364 N_B1_c_312_n N_VGND_c_962_n 0.00408624f $X=4.745 $Y=0.995 $X2=0 $Y2=0
cc_365 N_B1_c_316_n N_VGND_c_962_n 0.00428413f $X=6.852 $Y=0.995 $X2=0 $Y2=0
cc_366 N_C1_M27_noxref_g N_noxref_7_c_541_n 0.0129515f $X=5.12 $Y=1.985 $X2=0
+ $Y2=0
cc_367 N_C1_M28_noxref_g N_noxref_7_c_541_n 0.0112707f $X=5.55 $Y=1.985 $X2=0
+ $Y2=0
cc_368 N_C1_M29_noxref_g N_noxref_7_c_541_n 0.0114193f $X=5.98 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_C1_M30_noxref_g N_noxref_7_c_541_n 0.0115734f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_C1_M27_noxref_g N_VPWR_c_645_n 0.00357877f $X=5.12 $Y=1.985 $X2=0 $Y2=0
cc_371 N_C1_M28_noxref_g N_VPWR_c_645_n 0.00357877f $X=5.55 $Y=1.985 $X2=0 $Y2=0
cc_372 N_C1_M29_noxref_g N_VPWR_c_645_n 0.00357877f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_373 N_C1_M30_noxref_g N_VPWR_c_645_n 0.00357877f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_374 N_C1_M27_noxref_g N_VPWR_c_633_n 0.00539468f $X=5.12 $Y=1.985 $X2=0 $Y2=0
cc_375 N_C1_M28_noxref_g N_VPWR_c_633_n 0.00531884f $X=5.55 $Y=1.985 $X2=0 $Y2=0
cc_376 N_C1_M29_noxref_g N_VPWR_c_633_n 0.00537207f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_377 N_C1_M30_noxref_g N_VPWR_c_633_n 0.00547202f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_378 N_C1_M27_noxref_g N_noxref_9_c_745_n 0.014111f $X=5.12 $Y=1.985 $X2=0
+ $Y2=0
cc_379 N_C1_M28_noxref_g N_noxref_9_c_745_n 0.0109926f $X=5.55 $Y=1.985 $X2=0
+ $Y2=0
cc_380 N_C1_M29_noxref_g N_noxref_9_c_745_n 0.00451953f $X=5.98 $Y=1.985 $X2=0
+ $Y2=0
cc_381 N_C1_c_454_n N_noxref_9_c_745_n 0.0650168f $X=6.13 $Y=1.155 $X2=0 $Y2=0
cc_382 N_C1_c_460_n N_noxref_9_c_745_n 0.0180537f $X=6.185 $Y=1.16 $X2=0 $Y2=0
cc_383 N_C1_c_455_n N_noxref_9_c_745_n 0.00553579f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_384 N_C1_M27_noxref_g N_noxref_9_c_746_n 0.00613333f $X=5.12 $Y=1.985 $X2=0
+ $Y2=0
cc_385 N_C1_c_460_n N_Y_M29_noxref_d 0.00474778f $X=6.185 $Y=1.16 $X2=0 $Y2=0
cc_386 N_C1_c_450_n N_Y_c_852_n 0.0112545f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_387 N_C1_c_451_n N_Y_c_852_n 0.0112545f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_388 N_C1_c_454_n N_Y_c_852_n 0.0397307f $X=6.13 $Y=1.155 $X2=0 $Y2=0
cc_389 N_C1_c_455_n N_Y_c_852_n 0.00229737f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_390 N_C1_M27_noxref_g N_Y_c_824_n 0.00332425f $X=5.12 $Y=1.985 $X2=0 $Y2=0
cc_391 N_C1_M28_noxref_g N_Y_c_824_n 0.00971281f $X=5.55 $Y=1.985 $X2=0 $Y2=0
cc_392 N_C1_M29_noxref_g N_Y_c_824_n 0.0108104f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_393 N_C1_M30_noxref_g N_Y_c_824_n 0.0105097f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_394 N_C1_c_454_n N_Y_c_824_n 0.00145459f $X=6.13 $Y=1.155 $X2=0 $Y2=0
cc_395 N_C1_c_460_n N_Y_c_824_n 0.0128459f $X=6.185 $Y=1.16 $X2=0 $Y2=0
cc_396 N_C1_c_455_n N_Y_c_824_n 3.95205e-19 $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_397 N_C1_c_452_n N_Y_c_829_n 0.011457f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_398 N_C1_c_454_n N_Y_c_829_n 0.0138108f $X=6.13 $Y=1.155 $X2=0 $Y2=0
cc_399 N_C1_c_460_n N_Y_c_829_n 0.0149229f $X=6.185 $Y=1.16 $X2=0 $Y2=0
cc_400 N_C1_c_455_n N_Y_c_829_n 0.00213112f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_401 N_C1_c_453_n N_Y_c_794_n 0.0126398f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_402 N_C1_c_454_n N_Y_c_839_n 0.00332969f $X=6.13 $Y=1.155 $X2=0 $Y2=0
cc_403 N_C1_c_455_n N_Y_c_839_n 3.42634e-19 $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_404 N_C1_c_454_n N_Y_c_870_n 0.0126553f $X=6.13 $Y=1.155 $X2=0 $Y2=0
cc_405 N_C1_c_455_n N_Y_c_870_n 0.00231294f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_406 N_C1_c_453_n N_Y_c_872_n 0.00357123f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_407 N_C1_M30_noxref_g N_Y_c_796_n 0.00110866f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_408 N_C1_c_450_n N_VGND_c_947_n 5.0063e-19 $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_409 N_C1_c_450_n N_VGND_c_948_n 0.00338189f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_410 N_C1_c_450_n N_VGND_c_949_n 0.00647313f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_411 N_C1_c_451_n N_VGND_c_949_n 0.00644706f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_412 N_C1_c_452_n N_VGND_c_949_n 5.02907e-19 $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_413 N_C1_c_451_n N_VGND_c_950_n 5.02907e-19 $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_414 N_C1_c_452_n N_VGND_c_950_n 0.00643498f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_415 N_C1_c_453_n N_VGND_c_950_n 0.00788135f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_416 N_C1_c_453_n N_VGND_c_952_n 0.00103379f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_417 N_C1_c_451_n N_VGND_c_956_n 0.00338189f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_418 N_C1_c_452_n N_VGND_c_956_n 0.00337001f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_419 N_C1_c_453_n N_VGND_c_957_n 0.00337001f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_420 N_C1_c_450_n N_VGND_c_962_n 0.00396432f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_421 N_C1_c_451_n N_VGND_c_962_n 0.00392481f $X=5.59 $Y=0.995 $X2=0 $Y2=0
cc_422 N_C1_c_452_n N_VGND_c_962_n 0.00390568f $X=6.01 $Y=0.995 $X2=0 $Y2=0
cc_423 N_C1_c_453_n N_VGND_c_962_n 0.00400203f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_424 N_noxref_7_c_549_n N_VPWR_M16_noxref_d 0.00320329f $X=1.015 $Y=1.94
+ $X2=-0.19 $Y2=1.305
cc_425 N_noxref_7_c_553_n N_VPWR_M18_noxref_d 0.00331224f $X=1.855 $Y=1.95 $X2=0
+ $Y2=0
cc_426 N_noxref_7_c_555_n N_VPWR_M20_noxref_d 0.00320354f $X=2.695 $Y=1.95 $X2=0
+ $Y2=0
cc_427 N_noxref_7_c_556_n N_VPWR_M22_noxref_d 0.00327888f $X=3.535 $Y=1.95 $X2=0
+ $Y2=0
cc_428 N_noxref_7_c_549_n N_VPWR_c_634_n 0.0165403f $X=1.015 $Y=1.94 $X2=0 $Y2=0
cc_429 N_noxref_7_c_553_n N_VPWR_c_635_n 0.0165079f $X=1.855 $Y=1.95 $X2=0 $Y2=0
cc_430 N_noxref_7_c_555_n N_VPWR_c_636_n 0.0165079f $X=2.695 $Y=1.95 $X2=0 $Y2=0
cc_431 N_noxref_7_c_556_n N_VPWR_c_637_n 0.0165079f $X=3.535 $Y=1.95 $X2=0 $Y2=0
cc_432 N_noxref_7_c_549_n N_VPWR_c_638_n 0.00250343f $X=1.015 $Y=1.94 $X2=0
+ $Y2=0
cc_433 N_noxref_7_c_588_p N_VPWR_c_638_n 0.0113839f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_434 N_noxref_7_c_553_n N_VPWR_c_638_n 0.00263532f $X=1.855 $Y=1.95 $X2=0
+ $Y2=0
cc_435 N_noxref_7_c_553_n N_VPWR_c_640_n 0.00263532f $X=1.855 $Y=1.95 $X2=0
+ $Y2=0
cc_436 N_noxref_7_c_591_p N_VPWR_c_640_n 0.0113839f $X=1.94 $Y=2.3 $X2=0 $Y2=0
cc_437 N_noxref_7_c_555_n N_VPWR_c_640_n 0.00263532f $X=2.695 $Y=1.95 $X2=0
+ $Y2=0
cc_438 N_noxref_7_c_555_n N_VPWR_c_642_n 0.00263532f $X=2.695 $Y=1.95 $X2=0
+ $Y2=0
cc_439 N_noxref_7_c_594_p N_VPWR_c_642_n 0.0113839f $X=2.78 $Y=2.3 $X2=0 $Y2=0
cc_440 N_noxref_7_c_556_n N_VPWR_c_642_n 0.00263532f $X=3.535 $Y=1.95 $X2=0
+ $Y2=0
cc_441 N_noxref_7_c_540_n N_VPWR_c_644_n 0.0172654f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_442 N_noxref_7_c_549_n N_VPWR_c_644_n 0.00250343f $X=1.015 $Y=1.94 $X2=0
+ $Y2=0
cc_443 N_noxref_7_c_556_n N_VPWR_c_645_n 0.00263532f $X=3.535 $Y=1.95 $X2=0
+ $Y2=0
cc_444 N_noxref_7_c_599_p N_VPWR_c_645_n 0.0114548f $X=3.62 $Y=2.255 $X2=0 $Y2=0
cc_445 N_noxref_7_c_541_n N_VPWR_c_645_n 0.200564f $X=7.1 $Y=2.34 $X2=0 $Y2=0
cc_446 N_noxref_7_M16_noxref_s N_VPWR_c_633_n 0.00226392f $X=0.135 $Y=1.485
+ $X2=0 $Y2=0
cc_447 N_noxref_7_M17_noxref_d N_VPWR_c_633_n 0.00247944f $X=0.965 $Y=1.485
+ $X2=0 $Y2=0
cc_448 N_noxref_7_M19_noxref_d N_VPWR_c_633_n 0.00246541f $X=1.805 $Y=1.485
+ $X2=0 $Y2=0
cc_449 N_noxref_7_M21_noxref_d N_VPWR_c_633_n 0.00246541f $X=2.645 $Y=1.485
+ $X2=0 $Y2=0
cc_450 N_noxref_7_M23_noxref_d N_VPWR_c_633_n 0.00231679f $X=3.485 $Y=1.485
+ $X2=0 $Y2=0
cc_451 N_noxref_7_M25_noxref_d N_VPWR_c_633_n 0.00215227f $X=4.325 $Y=1.485
+ $X2=0 $Y2=0
cc_452 N_noxref_7_M31_noxref_d N_VPWR_c_633_n 0.00209344f $X=6.965 $Y=1.485
+ $X2=0 $Y2=0
cc_453 N_noxref_7_c_540_n N_VPWR_c_633_n 0.00954719f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_454 N_noxref_7_c_549_n N_VPWR_c_633_n 0.0100872f $X=1.015 $Y=1.94 $X2=0 $Y2=0
cc_455 N_noxref_7_c_588_p N_VPWR_c_633_n 0.00646745f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_456 N_noxref_7_c_553_n N_VPWR_c_633_n 0.0103305f $X=1.855 $Y=1.95 $X2=0 $Y2=0
cc_457 N_noxref_7_c_591_p N_VPWR_c_633_n 0.00646745f $X=1.94 $Y=2.3 $X2=0 $Y2=0
cc_458 N_noxref_7_c_555_n N_VPWR_c_633_n 0.0103305f $X=2.695 $Y=1.95 $X2=0 $Y2=0
cc_459 N_noxref_7_c_594_p N_VPWR_c_633_n 0.00646745f $X=2.78 $Y=2.3 $X2=0 $Y2=0
cc_460 N_noxref_7_c_556_n N_VPWR_c_633_n 0.0103305f $X=3.535 $Y=1.95 $X2=0 $Y2=0
cc_461 N_noxref_7_c_599_p N_VPWR_c_633_n 0.00653402f $X=3.62 $Y=2.255 $X2=0
+ $Y2=0
cc_462 N_noxref_7_c_541_n N_VPWR_c_633_n 0.12763f $X=7.1 $Y=2.34 $X2=0 $Y2=0
cc_463 N_noxref_7_c_541_n N_noxref_9_M24_noxref_d 0.0031348f $X=7.1 $Y=2.34
+ $X2=-0.19 $Y2=1.305
cc_464 N_noxref_7_c_541_n N_noxref_9_M28_noxref_d 0.00334977f $X=7.1 $Y=2.34
+ $X2=0 $Y2=0
cc_465 N_noxref_7_M25_noxref_d N_noxref_9_c_749_n 0.00345664f $X=4.325 $Y=1.485
+ $X2=0 $Y2=0
cc_466 N_noxref_7_c_541_n N_noxref_9_c_749_n 0.0370815f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_467 N_noxref_7_c_541_n N_noxref_9_c_745_n 0.00576787f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_468 N_noxref_7_c_541_n N_noxref_9_c_746_n 0.016595f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_469 N_noxref_7_c_541_n noxref_10 0.00440165f $X=7.1 $Y=2.34 $X2=-0.19
+ $Y2=1.305
cc_470 N_noxref_7_c_541_n N_Y_M27_noxref_d 0.00334977f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_471 N_noxref_7_c_541_n N_Y_M29_noxref_d 0.00375335f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_472 N_noxref_7_c_541_n N_Y_c_824_n 0.0897932f $X=7.1 $Y=2.34 $X2=0 $Y2=0
cc_473 N_noxref_7_M31_noxref_d N_Y_c_796_n 0.00242325f $X=6.965 $Y=1.485 $X2=0
+ $Y2=0
cc_474 N_noxref_7_M31_noxref_d Y 8.67893e-19 $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_475 N_noxref_7_M31_noxref_d N_Y_c_799_n 0.00312578f $X=6.965 $Y=1.485 $X2=0
+ $Y2=0
cc_476 N_noxref_7_c_541_n N_Y_c_799_n 0.0219024f $X=7.1 $Y=2.34 $X2=0 $Y2=0
cc_477 N_noxref_7_c_541_n noxref_12 0.0039288f $X=7.1 $Y=2.34 $X2=-0.19
+ $Y2=1.305
cc_478 N_VPWR_c_633_n N_noxref_9_M24_noxref_d 0.00216833f $X=7.13 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_479 N_VPWR_c_633_n N_noxref_9_M28_noxref_d 0.00224864f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_633_n noxref_10 0.00240926f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_481 N_VPWR_c_633_n N_Y_M27_noxref_d 0.00224864f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_482 N_VPWR_c_633_n N_Y_M29_noxref_d 0.00240926f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_c_633_n N_Y_c_799_n 9.82724e-19 $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_484 N_VPWR_c_633_n noxref_12 0.00248956f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_485 N_noxref_9_c_745_n noxref_10 0.00174389f $X=5.765 $Y=1.61 $X2=-0.19
+ $Y2=1.305
cc_486 N_noxref_9_c_746_n noxref_10 0.0056067f $X=4.77 $Y=1.57 $X2=-0.19
+ $Y2=1.305
cc_487 N_noxref_9_c_745_n N_Y_M27_noxref_d 0.00179007f $X=5.765 $Y=1.61 $X2=0
+ $Y2=0
cc_488 N_noxref_9_c_746_n N_Y_c_819_n 0.00283531f $X=4.77 $Y=1.57 $X2=0 $Y2=0
cc_489 N_noxref_9_M28_noxref_d N_Y_c_824_n 0.00327822f $X=5.625 $Y=1.485 $X2=0
+ $Y2=0
cc_490 N_noxref_9_c_745_n N_Y_c_824_n 0.0384307f $X=5.765 $Y=1.61 $X2=0 $Y2=0
cc_491 N_noxref_9_c_746_n N_Y_c_824_n 0.0127836f $X=4.77 $Y=1.57 $X2=0 $Y2=0
cc_492 N_noxref_9_c_745_n N_Y_c_839_n 0.00246739f $X=5.765 $Y=1.61 $X2=0 $Y2=0
cc_493 N_noxref_9_c_746_n N_Y_c_839_n 0.00100183f $X=4.77 $Y=1.57 $X2=0 $Y2=0
cc_494 N_Y_c_824_n noxref_12 0.00429548f $X=6.93 $Y=1.975 $X2=-0.19 $Y2=-0.24
cc_495 N_Y_c_801_n N_VGND_M1030_d 0.00665097f $X=3.875 $Y=0.78 $X2=0 $Y2=0
cc_496 N_Y_c_819_n N_VGND_M1006_s 0.00323842f $X=4.875 $Y=0.74 $X2=0 $Y2=0
cc_497 N_Y_c_852_n N_VGND_M1015_s 0.00308951f $X=5.715 $Y=0.745 $X2=0 $Y2=0
cc_498 N_Y_c_829_n N_VGND_M1027_s 0.00169165f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_499 N_Y_c_872_n N_VGND_M1027_s 0.00133935f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_500 N_Y_c_794_n N_VGND_M1026_s 0.00594168f $X=7.105 $Y=0.72 $X2=0 $Y2=0
cc_501 N_Y_c_795_n N_VGND_M1026_s 0.00104353f $X=7.102 $Y=1.495 $X2=0 $Y2=0
cc_502 N_Y_c_801_n N_VGND_c_945_n 0.012114f $X=3.875 $Y=0.78 $X2=0 $Y2=0
cc_503 N_Y_c_801_n N_VGND_c_946_n 0.00211912f $X=3.875 $Y=0.78 $X2=0 $Y2=0
cc_504 N_Y_c_803_n N_VGND_c_946_n 0.01976f $X=4.06 $Y=0.42 $X2=0 $Y2=0
cc_505 N_Y_c_819_n N_VGND_c_946_n 0.00264265f $X=4.875 $Y=0.74 $X2=0 $Y2=0
cc_506 N_Y_c_819_n N_VGND_c_947_n 0.0163189f $X=4.875 $Y=0.74 $X2=0 $Y2=0
cc_507 N_Y_c_819_n N_VGND_c_948_n 0.0027458f $X=4.875 $Y=0.74 $X2=0 $Y2=0
cc_508 N_Y_c_905_p N_VGND_c_948_n 0.0114803f $X=4.96 $Y=0.42 $X2=0 $Y2=0
cc_509 N_Y_c_852_n N_VGND_c_948_n 0.00253904f $X=5.715 $Y=0.745 $X2=0 $Y2=0
cc_510 N_Y_c_852_n N_VGND_c_949_n 0.0154525f $X=5.715 $Y=0.745 $X2=0 $Y2=0
cc_511 N_Y_c_829_n N_VGND_c_950_n 0.0161789f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_512 N_Y_c_794_n N_VGND_c_952_n 0.0238522f $X=7.105 $Y=0.72 $X2=0 $Y2=0
cc_513 N_Y_c_801_n N_VGND_c_953_n 0.00212504f $X=3.875 $Y=0.78 $X2=0 $Y2=0
cc_514 N_Y_c_852_n N_VGND_c_956_n 0.00253904f $X=5.715 $Y=0.745 $X2=0 $Y2=0
cc_515 N_Y_c_912_p N_VGND_c_956_n 0.0113089f $X=5.8 $Y=0.42 $X2=0 $Y2=0
cc_516 N_Y_c_829_n N_VGND_c_956_n 0.00260639f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_517 N_Y_c_794_n N_VGND_c_957_n 0.00856645f $X=7.105 $Y=0.72 $X2=0 $Y2=0
cc_518 N_Y_M1013_d N_VGND_c_962_n 0.00216833f $X=1.805 $Y=0.235 $X2=0 $Y2=0
cc_519 N_Y_M1020_d N_VGND_c_962_n 0.00216833f $X=2.645 $Y=0.235 $X2=0 $Y2=0
cc_520 N_Y_M1002_d N_VGND_c_962_n 0.00281385f $X=3.905 $Y=0.235 $X2=0 $Y2=0
cc_521 N_Y_M1023_d N_VGND_c_962_n 0.00252936f $X=4.82 $Y=0.235 $X2=0 $Y2=0
cc_522 N_Y_M1021_d N_VGND_c_962_n 0.00247241f $X=5.665 $Y=0.235 $X2=0 $Y2=0
cc_523 N_Y_M1031_d N_VGND_c_962_n 0.00318969f $X=6.505 $Y=0.235 $X2=0 $Y2=0
cc_524 N_Y_c_801_n N_VGND_c_962_n 0.00863387f $X=3.875 $Y=0.78 $X2=0 $Y2=0
cc_525 N_Y_c_803_n N_VGND_c_962_n 0.0120072f $X=4.06 $Y=0.42 $X2=0 $Y2=0
cc_526 N_Y_c_819_n N_VGND_c_962_n 0.0104634f $X=4.875 $Y=0.74 $X2=0 $Y2=0
cc_527 N_Y_c_905_p N_VGND_c_962_n 0.0064465f $X=4.96 $Y=0.42 $X2=0 $Y2=0
cc_528 N_Y_c_852_n N_VGND_c_962_n 0.0101296f $X=5.715 $Y=0.745 $X2=0 $Y2=0
cc_529 N_Y_c_912_p N_VGND_c_962_n 0.00645162f $X=5.8 $Y=0.42 $X2=0 $Y2=0
cc_530 N_Y_c_829_n N_VGND_c_962_n 0.00587314f $X=6.23 $Y=0.74 $X2=0 $Y2=0
cc_531 N_Y_c_794_n N_VGND_c_962_n 0.0161063f $X=7.105 $Y=0.72 $X2=0 $Y2=0
cc_532 N_Y_c_800_n N_A_109_47#_M1014_s 0.00307484f $X=3.235 $Y=0.77 $X2=0 $Y2=0
cc_533 N_Y_c_800_n N_A_109_47#_M1024_s 0.00335846f $X=3.235 $Y=0.77 $X2=0 $Y2=0
cc_534 N_Y_c_804_n N_A_109_47#_M1024_s 9.51e-19 $X=3.33 $Y=0.77 $X2=0 $Y2=0
cc_535 N_Y_M1013_d N_A_109_47#_c_1077_n 0.00306229f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_536 N_Y_M1020_d N_A_109_47#_c_1077_n 0.00306229f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_537 N_Y_c_800_n N_A_109_47#_c_1077_n 0.0770667f $X=3.235 $Y=0.77 $X2=0 $Y2=0
cc_538 N_Y_c_801_n N_A_109_47#_c_1077_n 0.00178381f $X=3.875 $Y=0.78 $X2=0 $Y2=0
cc_539 N_VGND_c_962_n N_A_109_47#_M1009_s 0.00352549f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_540 N_VGND_c_962_n N_A_109_47#_M1025_s 0.00215206f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_962_n N_A_109_47#_M1014_s 0.00215227f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_542 N_VGND_c_962_n N_A_109_47#_M1024_s 0.00212015f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_M1018_d N_A_109_47#_c_1068_n 0.00306545f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_544 N_VGND_c_944_n N_A_109_47#_c_1068_n 0.0130903f $X=1.1 $Y=0.36 $X2=0 $Y2=0
cc_545 N_VGND_c_953_n N_A_109_47#_c_1068_n 0.00211912f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_546 N_VGND_c_955_n N_A_109_47#_c_1068_n 0.00224973f $X=0.95 $Y=0 $X2=0 $Y2=0
cc_547 N_VGND_c_962_n N_A_109_47#_c_1068_n 0.00895942f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_548 N_VGND_c_953_n N_A_109_47#_c_1074_n 0.0151511f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_549 N_VGND_c_962_n N_A_109_47#_c_1074_n 0.00939123f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_550 N_VGND_c_953_n N_A_109_47#_c_1077_n 0.098072f $X=3.535 $Y=0 $X2=0 $Y2=0
cc_551 N_VGND_c_962_n N_A_109_47#_c_1077_n 0.0628764f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_955_n N_A_109_47#_c_1078_n 0.00434645f $X=0.95 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_962_n N_A_109_47#_c_1078_n 0.00655826f $X=7.13 $Y=0 $X2=0 $Y2=0

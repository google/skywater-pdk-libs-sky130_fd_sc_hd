* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
M1000 VGND a_505_21# a_439_47# VNB nshort w=420000u l=150000u
+  ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u
M1001 a_76_199# A0 a_218_374# VPB phighvt w=420000u l=150000u
+  ad=3.864e+11p pd=2.68e+06u as=1.533e+11p ps=1.57e+06u
M1002 VPWR a_505_21# a_535_374# VPB phighvt w=420000u l=150000u
+  ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_218_374# S VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_218_47# S VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1005 a_76_199# A1 a_218_47# VNB nshort w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1006 a_535_374# A1 a_76_199# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_76_199# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1008 a_505_21# S VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1009 a_505_21# S VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1010 VGND a_76_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1011 a_439_47# A0 a_76_199# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

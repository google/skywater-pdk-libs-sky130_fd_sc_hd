* File: sky130_fd_sc_hd__o41ai_4.pxi.spice
* Created: Tue Sep  1 19:26:52 2020
* 
x_PM_SKY130_FD_SC_HD__O41AI_4%B1 N_B1_M1020_g N_B1_M1003_g N_B1_M1028_g
+ N_B1_M1006_g N_B1_M1030_g N_B1_M1031_g N_B1_c_173_n N_B1_M1038_g N_B1_M1036_g
+ B1 B1 B1 B1 PM_SKY130_FD_SC_HD__O41AI_4%B1
x_PM_SKY130_FD_SC_HD__O41AI_4%A4 N_A4_c_244_n N_A4_M1010_g N_A4_M1014_g
+ N_A4_M1013_g N_A4_M1025_g N_A4_M1021_g N_A4_M1026_g N_A4_c_249_n N_A4_M1024_g
+ N_A4_M1035_g A4 A4 A4 A4 PM_SKY130_FD_SC_HD__O41AI_4%A4
x_PM_SKY130_FD_SC_HD__O41AI_4%A3 N_A3_M1017_g N_A3_M1001_g N_A3_M1022_g
+ N_A3_M1015_g N_A3_M1029_g N_A3_M1019_g N_A3_M1032_g N_A3_M1037_g A3 A3 A3 A3
+ N_A3_c_348_n N_A3_c_349_n PM_SKY130_FD_SC_HD__O41AI_4%A3
x_PM_SKY130_FD_SC_HD__O41AI_4%A2 N_A2_M1000_g N_A2_M1002_g N_A2_M1004_g
+ N_A2_M1027_g N_A2_M1005_g N_A2_M1033_g N_A2_M1011_g N_A2_M1039_g A2 A2 A2 A2
+ N_A2_c_441_n N_A2_c_442_n PM_SKY130_FD_SC_HD__O41AI_4%A2
x_PM_SKY130_FD_SC_HD__O41AI_4%A1 N_A1_M1008_g N_A1_M1007_g N_A1_M1009_g
+ N_A1_M1016_g N_A1_M1012_g N_A1_M1023_g N_A1_M1018_g N_A1_M1034_g A1 A1 A1 A1
+ N_A1_c_542_n A1 PM_SKY130_FD_SC_HD__O41AI_4%A1
x_PM_SKY130_FD_SC_HD__O41AI_4%VPWR N_VPWR_M1003_s N_VPWR_M1006_s N_VPWR_M1036_s
+ N_VPWR_M1007_s N_VPWR_M1023_s N_VPWR_c_622_n N_VPWR_c_623_n N_VPWR_c_624_n
+ N_VPWR_c_625_n N_VPWR_c_626_n N_VPWR_c_627_n N_VPWR_c_628_n N_VPWR_c_629_n
+ N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_632_n N_VPWR_c_633_n VPWR
+ N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_621_n N_VPWR_c_637_n
+ PM_SKY130_FD_SC_HD__O41AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O41AI_4%Y N_Y_M1020_s N_Y_M1030_s N_Y_M1003_d N_Y_M1031_d
+ N_Y_M1014_s N_Y_M1026_s N_Y_c_750_n N_Y_c_790_n N_Y_c_753_n N_Y_c_798_n
+ N_Y_c_754_n N_Y_c_755_n Y Y Y Y Y Y N_Y_c_760_n N_Y_c_761_n N_Y_c_752_n
+ N_Y_c_784_n N_Y_c_787_n PM_SKY130_FD_SC_HD__O41AI_4%Y
x_PM_SKY130_FD_SC_HD__O41AI_4%A_467_297# N_A_467_297#_M1014_d
+ N_A_467_297#_M1025_d N_A_467_297#_M1035_d N_A_467_297#_M1015_s
+ N_A_467_297#_M1037_s N_A_467_297#_c_848_n N_A_467_297#_c_856_n
+ N_A_467_297#_c_849_n N_A_467_297#_c_902_n N_A_467_297#_c_858_n
+ N_A_467_297#_c_850_n N_A_467_297#_c_851_n N_A_467_297#_c_865_n
+ N_A_467_297#_c_852_n N_A_467_297#_c_853_n N_A_467_297#_c_894_n
+ N_A_467_297#_c_854_n PM_SKY130_FD_SC_HD__O41AI_4%A_467_297#
x_PM_SKY130_FD_SC_HD__O41AI_4%A_885_297# N_A_885_297#_M1001_d
+ N_A_885_297#_M1019_d N_A_885_297#_M1002_d N_A_885_297#_M1033_d
+ N_A_885_297#_c_920_n N_A_885_297#_c_921_n N_A_885_297#_c_923_n
+ N_A_885_297#_c_949_n N_A_885_297#_c_919_n N_A_885_297#_c_956_p
+ N_A_885_297#_c_926_n N_A_885_297#_c_959_p N_A_885_297#_c_940_n
+ N_A_885_297#_c_942_n PM_SKY130_FD_SC_HD__O41AI_4%A_885_297#
x_PM_SKY130_FD_SC_HD__O41AI_4%A_1243_297# N_A_1243_297#_M1002_s
+ N_A_1243_297#_M1027_s N_A_1243_297#_M1039_s N_A_1243_297#_M1016_d
+ N_A_1243_297#_M1034_d N_A_1243_297#_c_960_n N_A_1243_297#_c_961_n
+ N_A_1243_297#_c_962_n N_A_1243_297#_c_980_n N_A_1243_297#_c_963_n
+ N_A_1243_297#_c_988_n N_A_1243_297#_c_964_n N_A_1243_297#_c_1003_n
+ N_A_1243_297#_c_965_n N_A_1243_297#_c_966_n N_A_1243_297#_c_967_n
+ N_A_1243_297#_c_968_n N_A_1243_297#_c_969_n
+ PM_SKY130_FD_SC_HD__O41AI_4%A_1243_297#
x_PM_SKY130_FD_SC_HD__O41AI_4%A_27_47# N_A_27_47#_M1020_d N_A_27_47#_M1028_d
+ N_A_27_47#_M1038_d N_A_27_47#_M1010_d N_A_27_47#_M1013_d N_A_27_47#_M1024_d
+ N_A_27_47#_M1022_s N_A_27_47#_M1032_s N_A_27_47#_M1000_s N_A_27_47#_M1004_s
+ N_A_27_47#_M1011_s N_A_27_47#_M1009_s N_A_27_47#_M1018_s N_A_27_47#_c_1045_n
+ N_A_27_47#_c_1046_n N_A_27_47#_c_1047_n N_A_27_47#_c_1079_n
+ N_A_27_47#_c_1077_n N_A_27_47#_c_1048_n N_A_27_47#_c_1049_n
+ N_A_27_47#_c_1089_n N_A_27_47#_c_1050_n N_A_27_47#_c_1097_n
+ N_A_27_47#_c_1051_n N_A_27_47#_c_1111_n N_A_27_47#_c_1052_n
+ N_A_27_47#_c_1053_n N_A_27_47#_c_1054_n N_A_27_47#_c_1055_n
+ N_A_27_47#_c_1056_n N_A_27_47#_c_1137_n N_A_27_47#_c_1057_n
+ N_A_27_47#_c_1145_n N_A_27_47#_c_1058_n N_A_27_47#_c_1163_n
+ N_A_27_47#_c_1059_n N_A_27_47#_c_1060_n N_A_27_47#_c_1061_n
+ N_A_27_47#_c_1062_n N_A_27_47#_c_1063_n N_A_27_47#_c_1064_n
+ N_A_27_47#_c_1065_n N_A_27_47#_c_1066_n N_A_27_47#_c_1067_n
+ N_A_27_47#_c_1068_n PM_SKY130_FD_SC_HD__O41AI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O41AI_4%VGND N_VGND_M1010_s N_VGND_M1021_s N_VGND_M1017_d
+ N_VGND_M1029_d N_VGND_M1000_d N_VGND_M1005_d N_VGND_M1008_d N_VGND_M1012_d
+ N_VGND_c_1272_n N_VGND_c_1273_n N_VGND_c_1274_n N_VGND_c_1275_n
+ N_VGND_c_1276_n N_VGND_c_1277_n N_VGND_c_1278_n N_VGND_c_1279_n
+ N_VGND_c_1280_n N_VGND_c_1281_n N_VGND_c_1282_n N_VGND_c_1283_n
+ N_VGND_c_1284_n N_VGND_c_1285_n N_VGND_c_1286_n N_VGND_c_1287_n
+ N_VGND_c_1288_n N_VGND_c_1289_n N_VGND_c_1290_n N_VGND_c_1291_n
+ N_VGND_c_1292_n N_VGND_c_1293_n N_VGND_c_1294_n VGND N_VGND_c_1295_n
+ N_VGND_c_1296_n N_VGND_c_1297_n PM_SKY130_FD_SC_HD__O41AI_4%VGND
cc_1 VNB N_B1_M1020_g 0.0229701f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_B1_M1028_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_B1_M1006_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_4 VNB N_B1_M1030_g 0.0172834f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_5 VNB N_B1_M1031_g 4.49859e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_6 VNB N_B1_c_173_n 0.0878075f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.025
cc_7 VNB N_B1_M1038_g 0.0209309f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_8 VNB N_B1_M1036_g 5.34616e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_9 VNB B1 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_10 VNB N_A4_c_244_n 0.0196825f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.015
cc_11 VNB N_A4_M1013_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_12 VNB N_A4_M1025_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_13 VNB N_A4_M1021_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_14 VNB N_A4_M1026_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_15 VNB N_A4_c_249_n 0.0793088f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A4_M1024_g 0.0175639f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_17 VNB N_A4_M1035_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_18 VNB A4 0.00371738f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_19 VNB N_A3_M1017_g 0.0175639f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_A3_M1001_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_21 VNB N_A3_M1022_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_22 VNB N_A3_M1015_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_23 VNB N_A3_M1029_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_24 VNB N_A3_M1019_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_25 VNB N_A3_M1032_g 0.0238771f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_26 VNB N_A3_M1037_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_27 VNB N_A3_c_348_n 0.0582256f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_28 VNB N_A3_c_349_n 0.0315688f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_29 VNB N_A2_M1000_g 0.0238771f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_30 VNB N_A2_M1002_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_31 VNB N_A2_M1004_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_32 VNB N_A2_M1027_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_33 VNB N_A2_M1005_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_34 VNB N_A2_M1033_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_35 VNB N_A2_M1011_g 0.0175639f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_36 VNB N_A2_M1039_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_37 VNB N_A2_c_441_n 0.00640919f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_38 VNB N_A2_c_442_n 0.0734508f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_39 VNB N_A1_M1008_g 0.0175639f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_40 VNB N_A1_M1007_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_41 VNB N_A1_M1009_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_42 VNB N_A1_M1016_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_43 VNB N_A1_M1012_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_44 VNB N_A1_M1023_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_45 VNB N_A1_M1018_g 0.0238771f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_46 VNB N_A1_M1034_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_47 VNB A1 0.0254859f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_48 VNB N_A1_c_542_n 0.0760363f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_49 VNB N_VPWR_c_621_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_750_n 0.00745062f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_51 VNB Y 0.00995045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_752_n 0.00378775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_27_47#_c_1045_n 0.00929764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_27_47#_c_1046_n 0.0185818f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_55 VNB N_A_27_47#_c_1047_n 0.0110516f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_56 VNB N_A_27_47#_c_1048_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_57 VNB N_A_27_47#_c_1049_n 0.00163327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_27_47#_c_1050_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_27_47#_c_1051_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_27_47#_c_1052_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_27_47#_c_1053_n 0.00360197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_27_47#_c_1054_n 0.00942896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_27_47#_c_1055_n 0.0035283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_27_47#_c_1056_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_27_47#_c_1057_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_27_47#_c_1058_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_27_47#_c_1059_n 0.0116174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_27_47#_c_1060_n 0.0181379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_27_47#_c_1061_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_27_47#_c_1062_n 0.00496586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_27_47#_c_1063_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_27_47#_c_1064_n 0.00204484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_27_47#_c_1065_n 0.00270871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_27_47#_c_1066_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_27_47#_c_1067_n 0.00365945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_27_47#_c_1068_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1272_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_78 VNB N_VGND_c_1273_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_79 VNB N_VGND_c_1274_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_80 VNB N_VGND_c_1275_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1276_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_82 VNB N_VGND_c_1277_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_83 VNB N_VGND_c_1278_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.16
cc_84 VNB N_VGND_c_1279_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1280_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1281_n 0.0659631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1282_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1283_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1284_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1285_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1286_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1287_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1288_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1289_n 0.0295085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1290_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1291_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1292_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1293_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1294_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1295_n 0.0224294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1296_n 0.478686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1297_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VPB N_B1_M1003_g 0.0263683f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_104 VPB N_B1_M1006_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_105 VPB N_B1_M1031_g 0.0191788f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_106 VPB N_B1_c_173_n 0.00817555f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.025
cc_107 VPB N_B1_M1036_g 0.0231694f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_108 VPB N_A4_M1014_g 0.0225954f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_109 VPB N_A4_M1025_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_110 VPB N_A4_M1026_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_111 VPB N_A4_c_249_n 0.00750268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A4_M1035_g 0.0197272f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_113 VPB N_A3_M1001_g 0.0194911f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_114 VPB N_A3_M1015_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_115 VPB N_A3_M1019_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_116 VPB N_A3_M1037_g 0.0267067f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_117 VPB N_A2_M1002_g 0.0267067f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_118 VPB N_A2_M1027_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_119 VPB N_A2_M1033_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_120 VPB N_A2_M1039_g 0.0194853f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_121 VPB N_A1_M1007_g 0.0194853f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_122 VPB N_A1_M1016_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_123 VPB N_A1_M1023_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_124 VPB N_A1_M1034_g 0.0267067f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_125 VPB N_VPWR_c_622_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_623_n 0.0462623f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_127 VPB N_VPWR_c_624_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_625_n 0.0108807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_626_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_627_n 0.00410835f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_131 VPB N_VPWR_c_628_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_629_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_630_n 0.145051f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_134 VPB N_VPWR_c_631_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_135 VPB N_VPWR_c_632_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_136 VPB N_VPWR_c_633_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_137 VPB N_VPWR_c_634_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_635_n 0.0229574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_621_n 0.0614248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_637_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_Y_c_753_n 0.0044278f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.295
cc_142 VPB N_Y_c_754_n 0.0140549f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_143 VPB N_Y_c_755_n 0.00223815f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_144 VPB Y 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB Y 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB Y 0.00399002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB Y 0.00335687f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_148 VPB N_Y_c_760_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_Y_c_761_n 8.47385e-19 $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.175
cc_150 VPB N_A_467_297#_c_848_n 0.0050955f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_151 VPB N_A_467_297#_c_849_n 0.00181858f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.295
cc_152 VPB N_A_467_297#_c_850_n 0.00289964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_467_297#_c_851_n 0.00292689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_467_297#_c_852_n 0.00559623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_467_297#_c_853_n 0.00485985f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_156 VPB N_A_467_297#_c_854_n 0.00223815f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_157 VPB N_A_885_297#_c_919_n 0.0109117f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_158 VPB N_A_1243_297#_c_960_n 0.00485985f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_159 VPB N_A_1243_297#_c_961_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_1243_297#_c_962_n 0.00405856f $X=-0.19 $Y=1.305 $X2=1.31
+ $Y2=1.295
cc_161 VPB N_A_1243_297#_c_963_n 0.00218965f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_162 VPB N_A_1243_297#_c_964_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0.61
+ $Y2=1.105
cc_163 VPB N_A_1243_297#_c_965_n 0.0117183f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_164 VPB N_A_1243_297#_c_966_n 0.032376f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_165 VPB N_A_1243_297#_c_967_n 0.00223815f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_166 VPB N_A_1243_297#_c_968_n 0.0036674f $X=-0.19 $Y=1.305 $X2=0.235
+ $Y2=1.175
cc_167 VPB N_A_1243_297#_c_969_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 N_B1_M1038_g N_A4_c_249_n 0.00520634f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_169 N_B1_M1003_g N_VPWR_c_623_n 0.00410837f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_170 N_B1_c_173_n N_VPWR_c_623_n 0.00562759f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_171 B1 N_VPWR_c_623_n 0.0194886f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_172 N_B1_M1006_g N_VPWR_c_624_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B1_M1031_g N_VPWR_c_624_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B1_M1036_g N_VPWR_c_625_n 0.00321269f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_175 N_B1_M1003_g N_VPWR_c_628_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B1_M1006_g N_VPWR_c_628_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B1_M1031_g N_VPWR_c_634_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_178 N_B1_M1036_g N_VPWR_c_634_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_179 N_B1_M1003_g N_VPWR_c_621_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B1_M1006_g N_VPWR_c_621_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B1_M1031_g N_VPWR_c_621_n 0.00950154f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B1_M1036_g N_VPWR_c_621_n 0.0108276f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_M1020_g N_Y_c_750_n 0.00398755f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_184 N_B1_M1028_g N_Y_c_750_n 0.0112239f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_185 N_B1_M1030_g N_Y_c_750_n 0.0112239f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_186 N_B1_c_173_n N_Y_c_750_n 0.0062366f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_187 N_B1_M1038_g N_Y_c_750_n 0.0148982f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_188 B1 N_Y_c_750_n 0.0875307f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_189 N_B1_M1003_g Y 0.00276634f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B1_M1006_g Y 0.00135419f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_191 N_B1_c_173_n Y 0.00206439f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_192 B1 Y 0.026643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_193 N_B1_M1031_g Y 0.00135419f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B1_c_173_n Y 0.00206439f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_195 N_B1_M1036_g Y 0.00135419f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_196 B1 Y 0.026643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_197 N_B1_M1038_g Y 0.015255f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_198 B1 Y 0.016453f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_199 N_B1_M1006_g N_Y_c_760_n 0.0107189f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B1_M1031_g N_Y_c_760_n 0.0107189f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_201 N_B1_c_173_n N_Y_c_760_n 0.00198252f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_202 B1 N_Y_c_760_n 0.0359514f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_203 N_B1_M1036_g N_Y_c_761_n 0.0140198f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_204 B1 N_Y_c_761_n 9.95686e-19 $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_205 N_B1_M1003_g N_Y_c_784_n 0.0095746f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B1_M1006_g N_Y_c_784_n 0.0106215f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B1_M1031_g N_Y_c_784_n 7.66249e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_M1006_g N_Y_c_787_n 7.66249e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1031_g N_Y_c_787_n 0.0106215f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_M1036_g N_Y_c_787_n 0.0156353f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1036_g N_A_467_297#_c_848_n 0.00112495f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_B1_M1020_g N_A_27_47#_c_1046_n 4.62458e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_213 N_B1_c_173_n N_A_27_47#_c_1046_n 0.00581864f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_214 B1 N_A_27_47#_c_1046_n 0.0194124f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_215 N_B1_M1020_g N_A_27_47#_c_1047_n 0.0103313f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_216 N_B1_M1028_g N_A_27_47#_c_1047_n 0.00866705f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_217 N_B1_M1030_g N_A_27_47#_c_1047_n 0.00866705f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_218 N_B1_M1038_g N_A_27_47#_c_1047_n 0.00866705f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_219 B1 N_A_27_47#_c_1047_n 0.00349599f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_220 N_B1_M1038_g N_A_27_47#_c_1077_n 0.00325806f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_221 N_B1_M1038_g N_A_27_47#_c_1049_n 6.50799e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_222 N_B1_M1020_g N_VGND_c_1281_n 0.00357877f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_223 N_B1_M1028_g N_VGND_c_1281_n 0.00357877f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_224 N_B1_M1030_g N_VGND_c_1281_n 0.00357877f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_225 N_B1_M1038_g N_VGND_c_1281_n 0.00357877f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_226 N_B1_M1020_g N_VGND_c_1296_n 0.00617937f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_227 N_B1_M1028_g N_VGND_c_1296_n 0.00522516f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_228 N_B1_M1030_g N_VGND_c_1296_n 0.00522516f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_229 N_B1_M1038_g N_VGND_c_1296_n 0.00655123f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A4_M1024_g N_A3_M1017_g 0.0149322f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A4_M1035_g N_A3_M1001_g 0.0149322f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A4_c_249_n A3 2.3095e-19 $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_233 A4 A3 0.0118208f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_234 N_A4_c_249_n N_A3_c_348_n 0.0149322f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_235 A4 N_A3_c_348_n 0.00161014f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_236 N_A4_M1014_g N_VPWR_c_625_n 0.00229957f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A4_M1014_g N_VPWR_c_630_n 0.00357877f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A4_M1025_g N_VPWR_c_630_n 0.00357877f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A4_M1026_g N_VPWR_c_630_n 0.00357877f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A4_M1035_g N_VPWR_c_630_n 0.00357877f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A4_M1014_g N_VPWR_c_621_n 0.00655123f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A4_M1025_g N_VPWR_c_621_n 0.00522516f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A4_M1026_g N_VPWR_c_621_n 0.00522516f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A4_M1035_g N_VPWR_c_621_n 0.00525237f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A4_M1014_g N_Y_c_790_n 0.0115312f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A4_M1025_g N_Y_c_790_n 0.00688691f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A4_M1026_g N_Y_c_790_n 5.34018e-19 $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A4_M1025_g N_Y_c_753_n 0.0107189f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A4_M1026_g N_Y_c_753_n 0.0120586f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A4_c_249_n N_Y_c_753_n 0.00404321f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_251 N_A4_M1035_g N_Y_c_753_n 0.00263685f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_252 A4 N_Y_c_753_n 0.0625945f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_253 N_A4_M1025_g N_Y_c_798_n 5.34018e-19 $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_254 N_A4_M1026_g N_Y_c_798_n 0.00688691f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A4_M1035_g N_Y_c_798_n 0.00570839f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A4_M1014_g N_Y_c_754_n 0.0128219f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A4_c_249_n N_Y_c_754_n 0.00582639f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_258 A4 N_Y_c_754_n 0.0259352f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_259 N_A4_M1014_g N_Y_c_755_n 0.0013397f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A4_M1025_g N_Y_c_755_n 0.0013397f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A4_c_249_n N_Y_c_755_n 0.00206069f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_262 A4 N_Y_c_755_n 0.026643f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_263 N_A4_c_244_n Y 0.00245645f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A4_M1014_g Y 0.00328446f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A4_c_249_n Y 0.00436648f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_266 A4 Y 0.0151254f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_267 N_A4_c_244_n N_Y_c_752_n 6.0652e-19 $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A4_M1014_g N_A_467_297#_c_856_n 0.0112878f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A4_M1025_g N_A_467_297#_c_856_n 0.0112878f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A4_M1026_g N_A_467_297#_c_858_n 0.0112437f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A4_M1035_g N_A_467_297#_c_858_n 0.0112878f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A4_M1035_g N_A_467_297#_c_850_n 3.16391e-19 $X=3.93 $Y=1.985 $X2=0
+ $Y2=0
cc_273 N_A4_c_244_n N_A_27_47#_c_1079_n 0.00244813f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A4_c_244_n N_A_27_47#_c_1077_n 0.00411304f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A4_M1013_g N_A_27_47#_c_1077_n 5.16591e-19 $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_276 N_A4_c_244_n N_A_27_47#_c_1048_n 0.00850187f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A4_M1013_g N_A_27_47#_c_1048_n 0.00845772f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A4_c_249_n N_A_27_47#_c_1048_n 0.00205431f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_279 A4 N_A_27_47#_c_1048_n 0.0359512f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_280 N_A4_c_244_n N_A_27_47#_c_1049_n 0.00126526f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A4_c_249_n N_A_27_47#_c_1049_n 0.00627033f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_282 A4 N_A_27_47#_c_1049_n 0.0222017f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_283 N_A4_c_244_n N_A_27_47#_c_1089_n 5.77985e-19 $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A4_M1013_g N_A_27_47#_c_1089_n 0.00655349f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A4_M1021_g N_A_27_47#_c_1089_n 0.00655349f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A4_M1024_g N_A_27_47#_c_1089_n 5.77985e-19 $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A4_M1021_g N_A_27_47#_c_1050_n 0.00850187f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A4_c_249_n N_A_27_47#_c_1050_n 0.00205431f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_289 N_A4_M1024_g N_A_27_47#_c_1050_n 0.00850187f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_290 A4 N_A_27_47#_c_1050_n 0.0359512f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_291 N_A4_M1021_g N_A_27_47#_c_1097_n 5.77985e-19 $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A4_M1024_g N_A_27_47#_c_1097_n 0.00655349f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A4_M1013_g N_A_27_47#_c_1061_n 0.00110555f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A4_M1021_g N_A_27_47#_c_1061_n 0.00110555f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_295 N_A4_c_249_n N_A_27_47#_c_1061_n 0.00213429f $X=3.93 $Y=1.025 $X2=0 $Y2=0
cc_296 A4 N_A_27_47#_c_1061_n 0.0265408f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_297 N_A4_M1024_g N_A_27_47#_c_1062_n 0.00110056f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_298 A4 N_A_27_47#_c_1062_n 0.00357912f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_299 N_A4_c_244_n N_VGND_c_1272_n 0.00268723f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A4_M1013_g N_VGND_c_1272_n 0.00146448f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_301 N_A4_M1021_g N_VGND_c_1273_n 0.00146448f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_302 N_A4_M1024_g N_VGND_c_1273_n 0.00146448f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_303 N_A4_c_244_n N_VGND_c_1281_n 0.00422898f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A4_M1013_g N_VGND_c_1283_n 0.00424416f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A4_M1021_g N_VGND_c_1283_n 0.00424416f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A4_M1024_g N_VGND_c_1285_n 0.00424416f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A4_c_244_n N_VGND_c_1296_n 0.00707121f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A4_M1013_g N_VGND_c_1296_n 0.00573607f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A4_M1021_g N_VGND_c_1296_n 0.00573607f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A4_M1024_g N_VGND_c_1296_n 0.00576327f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_311 A3 N_A2_c_441_n 0.0162228f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_312 N_A3_c_349_n N_A2_c_441_n 0.00187335f $X=5.815 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A3_c_349_n N_A2_c_442_n 0.0104238f $X=5.815 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A3_M1001_g N_VPWR_c_630_n 0.00539841f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A3_M1015_g N_VPWR_c_630_n 0.00357877f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A3_M1019_g N_VPWR_c_630_n 0.00357877f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A3_M1037_g N_VPWR_c_630_n 0.00357877f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A3_M1001_g N_VPWR_c_621_n 0.00961452f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A3_M1015_g N_VPWR_c_621_n 0.00522516f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A3_M1019_g N_VPWR_c_621_n 0.00522516f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A3_M1037_g N_VPWR_c_621_n 0.00660224f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A3_M1001_g N_A_467_297#_c_851_n 0.0128171f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A3_M1015_g N_A_467_297#_c_851_n 0.0106747f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_324 A3 N_A_467_297#_c_851_n 0.0356421f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_325 N_A3_c_348_n N_A_467_297#_c_851_n 0.00198252f $X=5.685 $Y=1.16 $X2=0
+ $Y2=0
cc_326 N_A3_M1001_g N_A_467_297#_c_865_n 4.50937e-19 $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_327 N_A3_M1015_g N_A_467_297#_c_865_n 0.0071026f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A3_M1019_g N_A_467_297#_c_865_n 0.00688691f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A3_M1037_g N_A_467_297#_c_865_n 5.34018e-19 $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_330 N_A3_M1019_g N_A_467_297#_c_852_n 0.0107189f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A3_M1037_g N_A_467_297#_c_852_n 0.0123922f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_332 A3 N_A_467_297#_c_852_n 0.062283f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_333 N_A3_c_348_n N_A_467_297#_c_852_n 0.00198252f $X=5.685 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A3_c_349_n N_A_467_297#_c_852_n 0.00687658f $X=5.815 $Y=1.16 $X2=0
+ $Y2=0
cc_335 N_A3_M1019_g N_A_467_297#_c_853_n 5.34018e-19 $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A3_M1037_g N_A_467_297#_c_853_n 0.00688691f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A3_M1015_g N_A_467_297#_c_854_n 0.0013397f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A3_M1019_g N_A_467_297#_c_854_n 0.0013397f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_339 A3 N_A_467_297#_c_854_n 0.026643f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_340 N_A3_c_348_n N_A_467_297#_c_854_n 0.00206069f $X=5.685 $Y=1.16 $X2=0
+ $Y2=0
cc_341 N_A3_M1001_g N_A_885_297#_c_920_n 0.0057144f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A3_M1015_g N_A_885_297#_c_921_n 0.0112878f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_343 N_A3_M1019_g N_A_885_297#_c_921_n 0.0112878f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A3_M1001_g N_A_885_297#_c_923_n 0.00200125f $X=4.35 $Y=1.985 $X2=0
+ $Y2=0
cc_345 N_A3_M1037_g N_A_885_297#_c_919_n 0.0133908f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A3_M1037_g N_A_1243_297#_c_962_n 4.1126e-19 $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_347 N_A3_M1017_g N_A_27_47#_c_1097_n 0.00655349f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A3_M1022_g N_A_27_47#_c_1097_n 5.77985e-19 $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A3_M1017_g N_A_27_47#_c_1051_n 0.00844712f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A3_M1022_g N_A_27_47#_c_1051_n 0.00850187f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_351 A3 N_A_27_47#_c_1051_n 0.0356419f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_352 N_A3_c_348_n N_A_27_47#_c_1051_n 0.00205431f $X=5.685 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A3_M1017_g N_A_27_47#_c_1111_n 5.77985e-19 $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A3_M1022_g N_A_27_47#_c_1111_n 0.00655349f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A3_M1029_g N_A_27_47#_c_1111_n 0.00655349f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A3_M1032_g N_A_27_47#_c_1111_n 5.77985e-19 $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A3_M1029_g N_A_27_47#_c_1052_n 0.00850187f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A3_M1032_g N_A_27_47#_c_1052_n 0.00850187f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_359 A3 N_A_27_47#_c_1052_n 0.0359512f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_360 N_A3_c_348_n N_A_27_47#_c_1052_n 0.00205431f $X=5.685 $Y=1.16 $X2=0 $Y2=0
cc_361 N_A3_M1029_g N_A_27_47#_c_1053_n 5.77985e-19 $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A3_M1032_g N_A_27_47#_c_1053_n 0.00655349f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A3_c_349_n N_A_27_47#_c_1054_n 0.00114284f $X=5.815 $Y=1.16 $X2=0 $Y2=0
cc_364 N_A3_M1017_g N_A_27_47#_c_1062_n 0.00147648f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A3_M1022_g N_A_27_47#_c_1063_n 0.00110555f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A3_M1029_g N_A_27_47#_c_1063_n 0.00110555f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_367 A3 N_A_27_47#_c_1063_n 0.0265408f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_368 N_A3_c_348_n N_A_27_47#_c_1063_n 0.00213429f $X=5.685 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A3_M1032_g N_A_27_47#_c_1064_n 0.00134339f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_370 A3 N_A_27_47#_c_1064_n 0.0262291f $X=5.69 $Y=1.105 $X2=0 $Y2=0
cc_371 N_A3_c_349_n N_A_27_47#_c_1064_n 0.00712258f $X=5.815 $Y=1.16 $X2=0 $Y2=0
cc_372 N_A3_M1017_g N_VGND_c_1274_n 0.00146448f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_373 N_A3_M1022_g N_VGND_c_1274_n 0.00146448f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_374 N_A3_M1029_g N_VGND_c_1275_n 0.00146448f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_375 N_A3_M1032_g N_VGND_c_1275_n 0.00268723f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_376 N_A3_M1017_g N_VGND_c_1285_n 0.00424416f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A3_M1022_g N_VGND_c_1287_n 0.00424416f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_378 N_A3_M1029_g N_VGND_c_1287_n 0.00424416f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_379 N_A3_M1032_g N_VGND_c_1289_n 0.00424416f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_380 N_A3_M1017_g N_VGND_c_1296_n 0.00576327f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_381 N_A3_M1022_g N_VGND_c_1296_n 0.00573607f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_382 N_A3_M1029_g N_VGND_c_1296_n 0.00573607f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_383 N_A3_M1032_g N_VGND_c_1296_n 0.00706214f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_384 N_A2_M1011_g N_A1_M1008_g 0.0139989f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_385 N_A2_M1039_g N_A1_M1007_g 0.0165165f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_386 N_A2_c_441_n A1 0.0138625f $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A2_c_442_n A1 2.463e-19 $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_388 N_A2_c_441_n N_A1_c_542_n 2.463e-19 $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A2_c_442_n N_A1_c_542_n 0.0184699f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A2_M1002_g N_VPWR_c_630_n 0.00357877f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_391 N_A2_M1027_g N_VPWR_c_630_n 0.00357877f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A2_M1033_g N_VPWR_c_630_n 0.00357877f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A2_M1039_g N_VPWR_c_630_n 0.00541359f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A2_M1002_g N_VPWR_c_621_n 0.00660224f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_395 N_A2_M1027_g N_VPWR_c_621_n 0.00522516f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_396 N_A2_M1033_g N_VPWR_c_621_n 0.00522516f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A2_M1039_g N_VPWR_c_621_n 0.00965151f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_398 N_A2_M1002_g N_A_467_297#_c_852_n 4.1126e-19 $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_399 N_A2_M1002_g N_A_885_297#_c_919_n 0.0133908f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A2_M1027_g N_A_885_297#_c_926_n 0.0112437f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_401 N_A2_M1033_g N_A_885_297#_c_926_n 0.0112878f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A2_M1002_g N_A_1243_297#_c_960_n 0.00688691f $X=6.55 $Y=1.985 $X2=0
+ $Y2=0
cc_403 N_A2_M1027_g N_A_1243_297#_c_960_n 5.34018e-19 $X=6.97 $Y=1.985 $X2=0
+ $Y2=0
cc_404 N_A2_M1002_g N_A_1243_297#_c_961_n 0.0107189f $X=6.55 $Y=1.985 $X2=0
+ $Y2=0
cc_405 N_A2_M1027_g N_A_1243_297#_c_961_n 0.0107189f $X=6.97 $Y=1.985 $X2=0
+ $Y2=0
cc_406 N_A2_c_441_n N_A_1243_297#_c_961_n 0.0359514f $X=7.775 $Y=1.16 $X2=0
+ $Y2=0
cc_407 N_A2_c_442_n N_A_1243_297#_c_961_n 0.00198252f $X=7.81 $Y=1.16 $X2=0
+ $Y2=0
cc_408 N_A2_M1002_g N_A_1243_297#_c_962_n 0.00167331f $X=6.55 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A2_c_441_n N_A_1243_297#_c_962_n 0.0275081f $X=7.775 $Y=1.16 $X2=0
+ $Y2=0
cc_410 N_A2_c_442_n N_A_1243_297#_c_962_n 0.00251862f $X=7.81 $Y=1.16 $X2=0
+ $Y2=0
cc_411 N_A2_M1002_g N_A_1243_297#_c_980_n 5.34018e-19 $X=6.55 $Y=1.985 $X2=0
+ $Y2=0
cc_412 N_A2_M1027_g N_A_1243_297#_c_980_n 0.00688691f $X=6.97 $Y=1.985 $X2=0
+ $Y2=0
cc_413 N_A2_M1033_g N_A_1243_297#_c_980_n 0.00688691f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_414 N_A2_M1039_g N_A_1243_297#_c_980_n 5.34018e-19 $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_415 N_A2_M1033_g N_A_1243_297#_c_963_n 0.0107189f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_A2_M1039_g N_A_1243_297#_c_963_n 0.0107189f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_417 N_A2_c_441_n N_A_1243_297#_c_963_n 0.0359514f $X=7.775 $Y=1.16 $X2=0
+ $Y2=0
cc_418 N_A2_c_442_n N_A_1243_297#_c_963_n 0.00198252f $X=7.81 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A2_M1033_g N_A_1243_297#_c_988_n 5.84415e-19 $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A2_M1039_g N_A_1243_297#_c_988_n 0.0102534f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_421 N_A2_M1027_g N_A_1243_297#_c_967_n 0.0013397f $X=6.97 $Y=1.985 $X2=0
+ $Y2=0
cc_422 N_A2_M1033_g N_A_1243_297#_c_967_n 0.0013397f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_423 N_A2_c_441_n N_A_1243_297#_c_967_n 0.026643f $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_424 N_A2_c_442_n N_A_1243_297#_c_967_n 0.00206069f $X=7.81 $Y=1.16 $X2=0
+ $Y2=0
cc_425 N_A2_M1039_g N_A_1243_297#_c_968_n 0.00134394f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_A2_c_441_n N_A_1243_297#_c_968_n 0.00679601f $X=7.775 $Y=1.16 $X2=0
+ $Y2=0
cc_427 N_A2_c_442_n N_A_1243_297#_c_968_n 0.00126157f $X=7.81 $Y=1.16 $X2=0
+ $Y2=0
cc_428 N_A2_c_441_n N_A_27_47#_c_1054_n 3.43563e-19 $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_429 N_A2_M1000_g N_A_27_47#_c_1055_n 0.00650773f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_430 N_A2_M1004_g N_A_27_47#_c_1055_n 5.76511e-19 $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_431 N_A2_M1000_g N_A_27_47#_c_1056_n 0.00850187f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_432 N_A2_M1004_g N_A_27_47#_c_1056_n 0.00850187f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_433 N_A2_c_441_n N_A_27_47#_c_1056_n 0.0359512f $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_434 N_A2_c_442_n N_A_27_47#_c_1056_n 0.00205431f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_435 N_A2_M1000_g N_A_27_47#_c_1137_n 5.76511e-19 $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_436 N_A2_M1004_g N_A_27_47#_c_1137_n 0.00650773f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_437 N_A2_M1005_g N_A_27_47#_c_1137_n 0.00650773f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_438 N_A2_M1011_g N_A_27_47#_c_1137_n 5.76511e-19 $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_439 N_A2_M1005_g N_A_27_47#_c_1057_n 0.00850187f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_440 N_A2_M1011_g N_A_27_47#_c_1057_n 0.00850187f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_441 N_A2_c_441_n N_A_27_47#_c_1057_n 0.0359512f $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_442 N_A2_c_442_n N_A_27_47#_c_1057_n 0.00205431f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A2_M1005_g N_A_27_47#_c_1145_n 5.76511e-19 $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_444 N_A2_M1011_g N_A_27_47#_c_1145_n 0.00650773f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_445 N_A2_M1000_g N_A_27_47#_c_1065_n 0.00134325f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_446 N_A2_c_441_n N_A_27_47#_c_1065_n 0.0273875f $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_447 N_A2_c_442_n N_A_27_47#_c_1065_n 0.00260793f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_448 N_A2_M1004_g N_A_27_47#_c_1066_n 0.00110541f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_449 N_A2_M1005_g N_A_27_47#_c_1066_n 0.00110541f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_450 N_A2_c_441_n N_A_27_47#_c_1066_n 0.0265235f $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_451 N_A2_c_442_n N_A_27_47#_c_1066_n 0.00213376f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_452 N_A2_M1011_g N_A_27_47#_c_1067_n 0.00110042f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_453 N_A2_c_441_n N_A_27_47#_c_1067_n 0.00676573f $X=7.775 $Y=1.16 $X2=0 $Y2=0
cc_454 N_A2_c_442_n N_A_27_47#_c_1067_n 0.00130397f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_455 N_A2_M1000_g N_VGND_c_1276_n 0.00268723f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_456 N_A2_M1004_g N_VGND_c_1276_n 0.00146448f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_457 N_A2_M1004_g N_VGND_c_1277_n 0.00424619f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_458 N_A2_M1005_g N_VGND_c_1277_n 0.00424619f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_459 N_A2_M1005_g N_VGND_c_1278_n 0.00146448f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_460 N_A2_M1011_g N_VGND_c_1278_n 0.00146448f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_461 N_A2_M1000_g N_VGND_c_1289_n 0.00424619f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_462 N_A2_M1011_g N_VGND_c_1291_n 0.00424619f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_463 N_A2_M1000_g N_VGND_c_1296_n 0.00706231f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_464 N_A2_M1004_g N_VGND_c_1296_n 0.00573624f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_465 N_A2_M1005_g N_VGND_c_1296_n 0.00573624f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_466 N_A2_M1011_g N_VGND_c_1296_n 0.00576344f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_467 N_A1_M1007_g N_VPWR_c_626_n 0.00268723f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_468 N_A1_M1016_g N_VPWR_c_626_n 0.00146448f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_469 N_A1_M1023_g N_VPWR_c_627_n 0.00146448f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_470 N_A1_M1034_g N_VPWR_c_627_n 0.00268723f $X=9.49 $Y=1.985 $X2=0 $Y2=0
cc_471 N_A1_M1007_g N_VPWR_c_630_n 0.00541359f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_472 N_A1_M1016_g N_VPWR_c_632_n 0.00541359f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_473 N_A1_M1023_g N_VPWR_c_632_n 0.00541359f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_474 N_A1_M1034_g N_VPWR_c_635_n 0.00541359f $X=9.49 $Y=1.985 $X2=0 $Y2=0
cc_475 N_A1_M1007_g N_VPWR_c_621_n 0.00952874f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_476 N_A1_M1016_g N_VPWR_c_621_n 0.00950154f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_477 N_A1_M1023_g N_VPWR_c_621_n 0.00950154f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_478 N_A1_M1034_g N_VPWR_c_621_n 0.0105778f $X=9.49 $Y=1.985 $X2=0 $Y2=0
cc_479 N_A1_M1007_g N_A_1243_297#_c_988_n 0.0106215f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_480 N_A1_M1016_g N_A_1243_297#_c_988_n 7.66249e-19 $X=8.65 $Y=1.985 $X2=0
+ $Y2=0
cc_481 N_A1_M1007_g N_A_1243_297#_c_964_n 0.0107189f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_482 N_A1_M1016_g N_A_1243_297#_c_964_n 0.0107189f $X=8.65 $Y=1.985 $X2=0
+ $Y2=0
cc_483 A1 N_A_1243_297#_c_964_n 0.0359514f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_484 N_A1_c_542_n N_A_1243_297#_c_964_n 0.00198252f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_485 N_A1_M1007_g N_A_1243_297#_c_1003_n 7.66249e-19 $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_486 N_A1_M1016_g N_A_1243_297#_c_1003_n 0.0106215f $X=8.65 $Y=1.985 $X2=0
+ $Y2=0
cc_487 N_A1_M1023_g N_A_1243_297#_c_1003_n 0.0106215f $X=9.07 $Y=1.985 $X2=0
+ $Y2=0
cc_488 N_A1_M1034_g N_A_1243_297#_c_1003_n 7.66249e-19 $X=9.49 $Y=1.985 $X2=0
+ $Y2=0
cc_489 N_A1_M1023_g N_A_1243_297#_c_965_n 0.0107189f $X=9.07 $Y=1.985 $X2=0
+ $Y2=0
cc_490 N_A1_M1034_g N_A_1243_297#_c_965_n 0.0124067f $X=9.49 $Y=1.985 $X2=0
+ $Y2=0
cc_491 A1 N_A_1243_297#_c_965_n 0.0633629f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_492 N_A1_c_542_n N_A_1243_297#_c_965_n 0.0050791f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_493 N_A1_M1023_g N_A_1243_297#_c_966_n 7.66249e-19 $X=9.07 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_A1_M1034_g N_A_1243_297#_c_966_n 0.0106215f $X=9.49 $Y=1.985 $X2=0
+ $Y2=0
cc_495 N_A1_M1007_g N_A_1243_297#_c_968_n 0.00134394f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_496 A1 N_A_1243_297#_c_968_n 0.00231112f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_497 N_A1_M1016_g N_A_1243_297#_c_969_n 0.00135419f $X=8.65 $Y=1.985 $X2=0
+ $Y2=0
cc_498 N_A1_M1023_g N_A_1243_297#_c_969_n 0.00135419f $X=9.07 $Y=1.985 $X2=0
+ $Y2=0
cc_499 A1 N_A_1243_297#_c_969_n 0.026643f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_500 N_A1_c_542_n N_A_1243_297#_c_969_n 0.00206439f $X=9.535 $Y=1.16 $X2=0
+ $Y2=0
cc_501 N_A1_M1008_g N_A_27_47#_c_1145_n 0.00650773f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_502 N_A1_M1009_g N_A_27_47#_c_1145_n 5.76511e-19 $X=8.65 $Y=0.56 $X2=0 $Y2=0
cc_503 N_A1_M1008_g N_A_27_47#_c_1058_n 0.00850187f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_504 N_A1_M1009_g N_A_27_47#_c_1058_n 0.00850187f $X=8.65 $Y=0.56 $X2=0 $Y2=0
cc_505 A1 N_A_27_47#_c_1058_n 0.0359512f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_506 N_A1_c_542_n N_A_27_47#_c_1058_n 0.00205431f $X=9.535 $Y=1.16 $X2=0 $Y2=0
cc_507 N_A1_M1008_g N_A_27_47#_c_1163_n 5.76511e-19 $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_508 N_A1_M1009_g N_A_27_47#_c_1163_n 0.00650773f $X=8.65 $Y=0.56 $X2=0 $Y2=0
cc_509 N_A1_M1012_g N_A_27_47#_c_1163_n 0.00650773f $X=9.07 $Y=0.56 $X2=0 $Y2=0
cc_510 N_A1_M1018_g N_A_27_47#_c_1163_n 5.76511e-19 $X=9.49 $Y=0.56 $X2=0 $Y2=0
cc_511 N_A1_M1012_g N_A_27_47#_c_1059_n 0.00850187f $X=9.07 $Y=0.56 $X2=0 $Y2=0
cc_512 N_A1_M1018_g N_A_27_47#_c_1059_n 0.00976982f $X=9.49 $Y=0.56 $X2=0 $Y2=0
cc_513 A1 N_A_27_47#_c_1059_n 0.063242f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_514 N_A1_c_542_n N_A_27_47#_c_1059_n 0.00525496f $X=9.535 $Y=1.16 $X2=0 $Y2=0
cc_515 N_A1_M1012_g N_A_27_47#_c_1060_n 5.76511e-19 $X=9.07 $Y=0.56 $X2=0 $Y2=0
cc_516 N_A1_M1018_g N_A_27_47#_c_1060_n 0.00650773f $X=9.49 $Y=0.56 $X2=0 $Y2=0
cc_517 N_A1_M1008_g N_A_27_47#_c_1067_n 0.00110042f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_518 A1 N_A_27_47#_c_1067_n 0.00230134f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_519 N_A1_M1009_g N_A_27_47#_c_1068_n 0.00110541f $X=8.65 $Y=0.56 $X2=0 $Y2=0
cc_520 N_A1_M1012_g N_A_27_47#_c_1068_n 0.00110541f $X=9.07 $Y=0.56 $X2=0 $Y2=0
cc_521 A1 N_A_27_47#_c_1068_n 0.0265235f $X=9.85 $Y=1.105 $X2=0 $Y2=0
cc_522 N_A1_c_542_n N_A_27_47#_c_1068_n 0.00213376f $X=9.535 $Y=1.16 $X2=0 $Y2=0
cc_523 N_A1_M1008_g N_VGND_c_1279_n 0.00146448f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_524 N_A1_M1009_g N_VGND_c_1279_n 0.00146448f $X=8.65 $Y=0.56 $X2=0 $Y2=0
cc_525 N_A1_M1012_g N_VGND_c_1280_n 0.00146448f $X=9.07 $Y=0.56 $X2=0 $Y2=0
cc_526 N_A1_M1018_g N_VGND_c_1280_n 0.00268723f $X=9.49 $Y=0.56 $X2=0 $Y2=0
cc_527 N_A1_M1008_g N_VGND_c_1291_n 0.00424619f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_528 N_A1_M1009_g N_VGND_c_1293_n 0.00424619f $X=8.65 $Y=0.56 $X2=0 $Y2=0
cc_529 N_A1_M1012_g N_VGND_c_1293_n 0.00424619f $X=9.07 $Y=0.56 $X2=0 $Y2=0
cc_530 N_A1_M1018_g N_VGND_c_1295_n 0.00424619f $X=9.49 $Y=0.56 $X2=0 $Y2=0
cc_531 N_A1_M1008_g N_VGND_c_1296_n 0.00576344f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_532 N_A1_M1009_g N_VGND_c_1296_n 0.00573624f $X=8.65 $Y=0.56 $X2=0 $Y2=0
cc_533 N_A1_M1012_g N_VGND_c_1296_n 0.00573624f $X=9.07 $Y=0.56 $X2=0 $Y2=0
cc_534 N_A1_M1018_g N_VGND_c_1296_n 0.00681247f $X=9.49 $Y=0.56 $X2=0 $Y2=0
cc_535 N_VPWR_c_621_n N_Y_M1003_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_536 N_VPWR_c_621_n N_Y_M1031_d 0.00215201f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_537 N_VPWR_c_621_n N_Y_M1014_s 0.00216833f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_538 N_VPWR_c_621_n N_Y_M1026_s 0.00216833f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_c_623_n Y 0.00873275f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_540 N_VPWR_M1036_s Y 0.00299357f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_541 N_VPWR_c_625_n Y 0.0175453f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_542 N_VPWR_M1006_s N_Y_c_760_n 0.00185611f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_543 N_VPWR_c_624_n N_Y_c_760_n 0.0104788f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_544 N_VPWR_c_625_n N_Y_c_761_n 5.07258e-19 $X=1.94 $Y=2 $X2=0 $Y2=0
cc_545 N_VPWR_c_628_n N_Y_c_784_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_546 N_VPWR_c_621_n N_Y_c_784_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_547 N_VPWR_c_634_n N_Y_c_787_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_548 N_VPWR_c_621_n N_Y_c_787_n 0.0122217f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_549 N_VPWR_c_621_n N_A_467_297#_M1014_d 0.00209324f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_550 N_VPWR_c_621_n N_A_467_297#_M1025_d 0.0021521f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_621_n N_A_467_297#_M1035_d 0.00385313f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_621_n N_A_467_297#_M1015_s 0.00216833f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_621_n N_A_467_297#_M1037_s 0.00210147f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_625_n N_A_467_297#_c_848_n 0.033926f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_555 N_VPWR_c_630_n N_A_467_297#_c_856_n 0.0358391f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_621_n N_A_467_297#_c_856_n 0.0234424f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_625_n N_A_467_297#_c_849_n 0.0136295f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_558 N_VPWR_c_630_n N_A_467_297#_c_849_n 0.0173913f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_621_n N_A_467_297#_c_849_n 0.00962794f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_630_n N_A_467_297#_c_858_n 0.0473059f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_621_n N_A_467_297#_c_858_n 0.0299894f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_630_n N_A_467_297#_c_894_n 0.0114668f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_621_n N_A_467_297#_c_894_n 0.006547f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_564 N_VPWR_c_621_n N_A_885_297#_M1001_d 0.00215206f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_565 N_VPWR_c_621_n N_A_885_297#_M1019_d 0.0021521f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_621_n N_A_885_297#_M1002_d 0.0021521f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_621_n N_A_885_297#_M1033_d 0.00385313f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_630_n N_A_885_297#_c_921_n 0.0358391f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_621_n N_A_885_297#_c_921_n 0.0234424f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_630_n N_A_885_297#_c_923_n 0.0152535f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_621_n N_A_885_297#_c_923_n 0.00941307f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_630_n N_A_885_297#_c_919_n 0.0690823f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_621_n N_A_885_297#_c_919_n 0.04281f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_574 N_VPWR_c_630_n N_A_885_297#_c_926_n 0.0473059f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_621_n N_A_885_297#_c_926_n 0.0299789f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_630_n N_A_885_297#_c_940_n 0.0114668f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_621_n N_A_885_297#_c_940_n 0.00653655f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_630_n N_A_885_297#_c_942_n 0.0114668f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_621_n N_A_885_297#_c_942_n 0.00653655f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_580 N_VPWR_c_621_n N_A_1243_297#_M1002_s 0.00210147f $X=9.89 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_581 N_VPWR_c_621_n N_A_1243_297#_M1027_s 0.00216833f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_621_n N_A_1243_297#_M1039_s 0.00215201f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_621_n N_A_1243_297#_M1016_d 0.00215201f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_584 N_VPWR_c_621_n N_A_1243_297#_M1034_d 0.00225715f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_630_n N_A_1243_297#_c_988_n 0.0189039f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_621_n N_A_1243_297#_c_988_n 0.0122217f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_587 N_VPWR_M1007_s N_A_1243_297#_c_964_n 0.00185611f $X=8.305 $Y=1.485 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_626_n N_A_1243_297#_c_964_n 0.0104788f $X=8.44 $Y=2 $X2=0 $Y2=0
cc_589 N_VPWR_c_632_n N_A_1243_297#_c_1003_n 0.0189039f $X=9.195 $Y=2.72 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_621_n N_A_1243_297#_c_1003_n 0.0122217f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_591 N_VPWR_M1023_s N_A_1243_297#_c_965_n 0.00185611f $X=9.145 $Y=1.485 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_627_n N_A_1243_297#_c_965_n 0.0104788f $X=9.28 $Y=2 $X2=0 $Y2=0
cc_593 N_VPWR_c_635_n N_A_1243_297#_c_966_n 0.0210107f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_621_n N_A_1243_297#_c_966_n 0.0124268f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_623_n N_A_27_47#_c_1046_n 7.91944e-19 $X=0.26 $Y=1.66 $X2=0
+ $Y2=0
cc_596 N_Y_c_754_n N_A_467_297#_M1014_d 0.00272914f $X=2.715 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_597 N_Y_c_753_n N_A_467_297#_M1025_d 0.00165831f $X=3.555 $Y=1.53 $X2=0 $Y2=0
cc_598 N_Y_c_754_n N_A_467_297#_c_848_n 0.0198097f $X=2.715 $Y=1.53 $X2=0 $Y2=0
cc_599 N_Y_c_787_n N_A_467_297#_c_848_n 0.00146999f $X=1.52 $Y=1.66 $X2=0 $Y2=0
cc_600 N_Y_M1014_s N_A_467_297#_c_856_n 0.00312348f $X=2.745 $Y=1.485 $X2=0
+ $Y2=0
cc_601 N_Y_c_790_n N_A_467_297#_c_856_n 0.015949f $X=2.88 $Y=1.66 $X2=0 $Y2=0
cc_602 N_Y_c_753_n N_A_467_297#_c_902_n 0.0126919f $X=3.555 $Y=1.53 $X2=0 $Y2=0
cc_603 N_Y_M1026_s N_A_467_297#_c_858_n 0.00312348f $X=3.585 $Y=1.485 $X2=0
+ $Y2=0
cc_604 N_Y_c_798_n N_A_467_297#_c_858_n 0.015949f $X=3.72 $Y=1.66 $X2=0 $Y2=0
cc_605 N_Y_c_753_n N_A_467_297#_c_850_n 0.00902116f $X=3.555 $Y=1.53 $X2=0 $Y2=0
cc_606 N_Y_c_750_n N_A_27_47#_M1028_d 0.00162207f $X=1.87 $Y=0.77 $X2=0 $Y2=0
cc_607 N_Y_c_752_n N_A_27_47#_M1038_d 0.00318776f $X=2.015 $Y=0.905 $X2=0 $Y2=0
cc_608 N_Y_c_750_n N_A_27_47#_c_1046_n 0.0120147f $X=1.87 $Y=0.77 $X2=0 $Y2=0
cc_609 N_Y_M1020_s N_A_27_47#_c_1047_n 0.00305599f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_610 N_Y_M1030_s N_A_27_47#_c_1047_n 0.00305599f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_611 N_Y_c_750_n N_A_27_47#_c_1047_n 0.0666979f $X=1.87 $Y=0.77 $X2=0 $Y2=0
cc_612 N_Y_c_752_n N_A_27_47#_c_1047_n 0.0229034f $X=2.015 $Y=0.905 $X2=0 $Y2=0
cc_613 N_Y_c_752_n N_A_27_47#_c_1077_n 0.00788354f $X=2.015 $Y=0.905 $X2=0 $Y2=0
cc_614 N_Y_c_752_n N_A_27_47#_c_1049_n 0.0144435f $X=2.015 $Y=0.905 $X2=0 $Y2=0
cc_615 N_Y_M1020_s N_VGND_c_1296_n 0.00216833f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_616 N_Y_M1030_s N_VGND_c_1296_n 0.00216833f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_617 N_A_467_297#_c_851_n N_A_885_297#_M1001_d 0.00165831f $X=4.815 $Y=1.53
+ $X2=-0.19 $Y2=1.305
cc_618 N_A_467_297#_c_852_n N_A_885_297#_M1019_d 0.00165831f $X=5.655 $Y=1.53
+ $X2=0 $Y2=0
cc_619 N_A_467_297#_c_851_n N_A_885_297#_c_920_n 0.0148589f $X=4.815 $Y=1.53
+ $X2=0 $Y2=0
cc_620 N_A_467_297#_M1015_s N_A_885_297#_c_921_n 0.00312348f $X=4.845 $Y=1.485
+ $X2=0 $Y2=0
cc_621 N_A_467_297#_c_865_n N_A_885_297#_c_921_n 0.015949f $X=4.98 $Y=1.66 $X2=0
+ $Y2=0
cc_622 N_A_467_297#_c_852_n N_A_885_297#_c_949_n 0.0126919f $X=5.655 $Y=1.53
+ $X2=0 $Y2=0
cc_623 N_A_467_297#_M1037_s N_A_885_297#_c_919_n 0.00480843f $X=5.685 $Y=1.485
+ $X2=0 $Y2=0
cc_624 N_A_467_297#_c_853_n N_A_885_297#_c_919_n 0.0205836f $X=5.82 $Y=1.66
+ $X2=0 $Y2=0
cc_625 N_A_467_297#_c_853_n N_A_1243_297#_c_960_n 0.0391942f $X=5.82 $Y=1.66
+ $X2=0 $Y2=0
cc_626 N_A_467_297#_c_852_n N_A_1243_297#_c_962_n 0.0147157f $X=5.655 $Y=1.53
+ $X2=0 $Y2=0
cc_627 N_A_467_297#_c_850_n N_A_27_47#_c_1062_n 0.00708581f $X=4.14 $Y=1.615
+ $X2=0 $Y2=0
cc_628 N_A_467_297#_c_851_n N_A_27_47#_c_1062_n 0.00274641f $X=4.815 $Y=1.53
+ $X2=0 $Y2=0
cc_629 N_A_467_297#_c_852_n N_A_27_47#_c_1064_n 2.06363e-19 $X=5.655 $Y=1.53
+ $X2=0 $Y2=0
cc_630 N_A_885_297#_c_919_n N_A_1243_297#_M1002_s 0.00480843f $X=6.675 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_631 N_A_885_297#_c_926_n N_A_1243_297#_M1027_s 0.00312348f $X=7.515 $Y=2.38
+ $X2=0 $Y2=0
cc_632 N_A_885_297#_c_919_n N_A_1243_297#_c_960_n 0.0205836f $X=6.675 $Y=2.38
+ $X2=0 $Y2=0
cc_633 N_A_885_297#_M1002_d N_A_1243_297#_c_961_n 0.00165831f $X=6.625 $Y=1.485
+ $X2=0 $Y2=0
cc_634 N_A_885_297#_c_956_p N_A_1243_297#_c_961_n 0.0126919f $X=6.76 $Y=1.95
+ $X2=0 $Y2=0
cc_635 N_A_885_297#_c_926_n N_A_1243_297#_c_980_n 0.015949f $X=7.515 $Y=2.38
+ $X2=0 $Y2=0
cc_636 N_A_885_297#_M1033_d N_A_1243_297#_c_963_n 0.00165831f $X=7.465 $Y=1.485
+ $X2=0 $Y2=0
cc_637 N_A_885_297#_c_959_p N_A_1243_297#_c_963_n 0.0126919f $X=7.6 $Y=1.95
+ $X2=0 $Y2=0
cc_638 N_A_1243_297#_c_968_n N_A_27_47#_c_1067_n 0.00895629f $X=8.02 $Y=1.53
+ $X2=0 $Y2=0
cc_639 N_A_27_47#_c_1048_n N_VGND_M1010_s 0.00169589f $X=3.135 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_640 N_A_27_47#_c_1050_n N_VGND_M1021_s 0.00169589f $X=3.975 $Y=0.82 $X2=0
+ $Y2=0
cc_641 N_A_27_47#_c_1051_n N_VGND_M1017_d 0.00169589f $X=4.815 $Y=0.82 $X2=0
+ $Y2=0
cc_642 N_A_27_47#_c_1052_n N_VGND_M1029_d 0.00169589f $X=5.655 $Y=0.82 $X2=0
+ $Y2=0
cc_643 N_A_27_47#_c_1056_n N_VGND_M1000_d 0.00169589f $X=7.015 $Y=0.82 $X2=0
+ $Y2=0
cc_644 N_A_27_47#_c_1057_n N_VGND_M1005_d 0.00169589f $X=7.855 $Y=0.82 $X2=0
+ $Y2=0
cc_645 N_A_27_47#_c_1058_n N_VGND_M1008_d 0.00169589f $X=8.695 $Y=0.82 $X2=0
+ $Y2=0
cc_646 N_A_27_47#_c_1059_n N_VGND_M1012_d 0.00169589f $X=9.535 $Y=0.82 $X2=0
+ $Y2=0
cc_647 N_A_27_47#_c_1048_n N_VGND_c_1272_n 0.0111177f $X=3.135 $Y=0.82 $X2=0
+ $Y2=0
cc_648 N_A_27_47#_c_1050_n N_VGND_c_1273_n 0.0111177f $X=3.975 $Y=0.82 $X2=0
+ $Y2=0
cc_649 N_A_27_47#_c_1051_n N_VGND_c_1274_n 0.0111177f $X=4.815 $Y=0.82 $X2=0
+ $Y2=0
cc_650 N_A_27_47#_c_1052_n N_VGND_c_1275_n 0.0111177f $X=5.655 $Y=0.82 $X2=0
+ $Y2=0
cc_651 N_A_27_47#_c_1056_n N_VGND_c_1276_n 0.0111177f $X=7.015 $Y=0.82 $X2=0
+ $Y2=0
cc_652 N_A_27_47#_c_1056_n N_VGND_c_1277_n 0.00193763f $X=7.015 $Y=0.82 $X2=0
+ $Y2=0
cc_653 N_A_27_47#_c_1137_n N_VGND_c_1277_n 0.0182681f $X=7.18 $Y=0.38 $X2=0
+ $Y2=0
cc_654 N_A_27_47#_c_1057_n N_VGND_c_1277_n 0.00193763f $X=7.855 $Y=0.82 $X2=0
+ $Y2=0
cc_655 N_A_27_47#_c_1057_n N_VGND_c_1278_n 0.0111177f $X=7.855 $Y=0.82 $X2=0
+ $Y2=0
cc_656 N_A_27_47#_c_1058_n N_VGND_c_1279_n 0.0111177f $X=8.695 $Y=0.82 $X2=0
+ $Y2=0
cc_657 N_A_27_47#_c_1059_n N_VGND_c_1280_n 0.0111177f $X=9.535 $Y=0.82 $X2=0
+ $Y2=0
cc_658 N_A_27_47#_c_1045_n N_VGND_c_1281_n 0.0180491f $X=0.215 $Y=0.465 $X2=0
+ $Y2=0
cc_659 N_A_27_47#_c_1047_n N_VGND_c_1281_n 0.114888f $X=2.35 $Y=0.36 $X2=0 $Y2=0
cc_660 N_A_27_47#_c_1079_n N_VGND_c_1281_n 0.0172052f $X=2.487 $Y=0.465 $X2=0
+ $Y2=0
cc_661 N_A_27_47#_c_1048_n N_VGND_c_1281_n 0.00193763f $X=3.135 $Y=0.82 $X2=0
+ $Y2=0
cc_662 N_A_27_47#_c_1048_n N_VGND_c_1283_n 0.00193763f $X=3.135 $Y=0.82 $X2=0
+ $Y2=0
cc_663 N_A_27_47#_c_1089_n N_VGND_c_1283_n 0.0188551f $X=3.3 $Y=0.38 $X2=0 $Y2=0
cc_664 N_A_27_47#_c_1050_n N_VGND_c_1283_n 0.00193763f $X=3.975 $Y=0.82 $X2=0
+ $Y2=0
cc_665 N_A_27_47#_c_1050_n N_VGND_c_1285_n 0.00193763f $X=3.975 $Y=0.82 $X2=0
+ $Y2=0
cc_666 N_A_27_47#_c_1097_n N_VGND_c_1285_n 0.0188551f $X=4.14 $Y=0.38 $X2=0
+ $Y2=0
cc_667 N_A_27_47#_c_1051_n N_VGND_c_1285_n 0.00193763f $X=4.815 $Y=0.82 $X2=0
+ $Y2=0
cc_668 N_A_27_47#_c_1051_n N_VGND_c_1287_n 0.00193763f $X=4.815 $Y=0.82 $X2=0
+ $Y2=0
cc_669 N_A_27_47#_c_1111_n N_VGND_c_1287_n 0.0188551f $X=4.98 $Y=0.38 $X2=0
+ $Y2=0
cc_670 N_A_27_47#_c_1052_n N_VGND_c_1287_n 0.00193763f $X=5.655 $Y=0.82 $X2=0
+ $Y2=0
cc_671 N_A_27_47#_c_1052_n N_VGND_c_1289_n 0.00193763f $X=5.655 $Y=0.82 $X2=0
+ $Y2=0
cc_672 N_A_27_47#_c_1053_n N_VGND_c_1289_n 0.0209752f $X=5.82 $Y=0.38 $X2=0
+ $Y2=0
cc_673 N_A_27_47#_c_1054_n N_VGND_c_1289_n 0.00282615f $X=6.175 $Y=0.82 $X2=0
+ $Y2=0
cc_674 N_A_27_47#_c_1055_n N_VGND_c_1289_n 0.020318f $X=6.34 $Y=0.38 $X2=0 $Y2=0
cc_675 N_A_27_47#_c_1056_n N_VGND_c_1289_n 0.00193763f $X=7.015 $Y=0.82 $X2=0
+ $Y2=0
cc_676 N_A_27_47#_c_1057_n N_VGND_c_1291_n 0.00193763f $X=7.855 $Y=0.82 $X2=0
+ $Y2=0
cc_677 N_A_27_47#_c_1145_n N_VGND_c_1291_n 0.0182681f $X=8.02 $Y=0.38 $X2=0
+ $Y2=0
cc_678 N_A_27_47#_c_1058_n N_VGND_c_1291_n 0.00193763f $X=8.695 $Y=0.82 $X2=0
+ $Y2=0
cc_679 N_A_27_47#_c_1058_n N_VGND_c_1293_n 0.00193763f $X=8.695 $Y=0.82 $X2=0
+ $Y2=0
cc_680 N_A_27_47#_c_1163_n N_VGND_c_1293_n 0.0182681f $X=8.86 $Y=0.38 $X2=0
+ $Y2=0
cc_681 N_A_27_47#_c_1059_n N_VGND_c_1293_n 0.00193763f $X=9.535 $Y=0.82 $X2=0
+ $Y2=0
cc_682 N_A_27_47#_c_1059_n N_VGND_c_1295_n 0.00193763f $X=9.535 $Y=0.82 $X2=0
+ $Y2=0
cc_683 N_A_27_47#_c_1060_n N_VGND_c_1295_n 0.0202909f $X=9.7 $Y=0.38 $X2=0 $Y2=0
cc_684 N_A_27_47#_M1020_d N_VGND_c_1296_n 0.00209324f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_685 N_A_27_47#_M1028_d N_VGND_c_1296_n 0.00215227f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_686 N_A_27_47#_M1038_d N_VGND_c_1296_n 0.00209344f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_687 N_A_27_47#_M1010_d N_VGND_c_1296_n 0.0020932f $X=2.335 $Y=0.235 $X2=0
+ $Y2=0
cc_688 N_A_27_47#_M1013_d N_VGND_c_1296_n 0.00215201f $X=3.165 $Y=0.235 $X2=0
+ $Y2=0
cc_689 N_A_27_47#_M1024_d N_VGND_c_1296_n 0.00215201f $X=4.005 $Y=0.235 $X2=0
+ $Y2=0
cc_690 N_A_27_47#_M1022_s N_VGND_c_1296_n 0.00215201f $X=4.845 $Y=0.235 $X2=0
+ $Y2=0
cc_691 N_A_27_47#_M1032_s N_VGND_c_1296_n 0.00209319f $X=5.685 $Y=0.235 $X2=0
+ $Y2=0
cc_692 N_A_27_47#_M1000_s N_VGND_c_1296_n 0.0020946f $X=6.215 $Y=0.235 $X2=0
+ $Y2=0
cc_693 N_A_27_47#_M1004_s N_VGND_c_1296_n 0.00215347f $X=7.045 $Y=0.235 $X2=0
+ $Y2=0
cc_694 N_A_27_47#_M1011_s N_VGND_c_1296_n 0.00215347f $X=7.885 $Y=0.235 $X2=0
+ $Y2=0
cc_695 N_A_27_47#_M1009_s N_VGND_c_1296_n 0.00215347f $X=8.725 $Y=0.235 $X2=0
+ $Y2=0
cc_696 N_A_27_47#_M1018_s N_VGND_c_1296_n 0.00225867f $X=9.565 $Y=0.235 $X2=0
+ $Y2=0
cc_697 N_A_27_47#_c_1045_n N_VGND_c_1296_n 0.0100013f $X=0.215 $Y=0.465 $X2=0
+ $Y2=0
cc_698 N_A_27_47#_c_1047_n N_VGND_c_1296_n 0.0719952f $X=2.35 $Y=0.36 $X2=0
+ $Y2=0
cc_699 N_A_27_47#_c_1079_n N_VGND_c_1296_n 0.0103686f $X=2.487 $Y=0.465 $X2=0
+ $Y2=0
cc_700 N_A_27_47#_c_1048_n N_VGND_c_1296_n 0.00828806f $X=3.135 $Y=0.82 $X2=0
+ $Y2=0
cc_701 N_A_27_47#_c_1089_n N_VGND_c_1296_n 0.0122069f $X=3.3 $Y=0.38 $X2=0 $Y2=0
cc_702 N_A_27_47#_c_1050_n N_VGND_c_1296_n 0.00828806f $X=3.975 $Y=0.82 $X2=0
+ $Y2=0
cc_703 N_A_27_47#_c_1097_n N_VGND_c_1296_n 0.0122069f $X=4.14 $Y=0.38 $X2=0
+ $Y2=0
cc_704 N_A_27_47#_c_1051_n N_VGND_c_1296_n 0.00828806f $X=4.815 $Y=0.82 $X2=0
+ $Y2=0
cc_705 N_A_27_47#_c_1111_n N_VGND_c_1296_n 0.0122069f $X=4.98 $Y=0.38 $X2=0
+ $Y2=0
cc_706 N_A_27_47#_c_1052_n N_VGND_c_1296_n 0.00828806f $X=5.655 $Y=0.82 $X2=0
+ $Y2=0
cc_707 N_A_27_47#_c_1053_n N_VGND_c_1296_n 0.0124119f $X=5.82 $Y=0.38 $X2=0
+ $Y2=0
cc_708 N_A_27_47#_c_1054_n N_VGND_c_1296_n 0.00497105f $X=6.175 $Y=0.82 $X2=0
+ $Y2=0
cc_709 N_A_27_47#_c_1055_n N_VGND_c_1296_n 0.0123792f $X=6.34 $Y=0.38 $X2=0
+ $Y2=0
cc_710 N_A_27_47#_c_1056_n N_VGND_c_1296_n 0.00828806f $X=7.015 $Y=0.82 $X2=0
+ $Y2=0
cc_711 N_A_27_47#_c_1137_n N_VGND_c_1296_n 0.0121741f $X=7.18 $Y=0.38 $X2=0
+ $Y2=0
cc_712 N_A_27_47#_c_1057_n N_VGND_c_1296_n 0.00828806f $X=7.855 $Y=0.82 $X2=0
+ $Y2=0
cc_713 N_A_27_47#_c_1145_n N_VGND_c_1296_n 0.0121741f $X=8.02 $Y=0.38 $X2=0
+ $Y2=0
cc_714 N_A_27_47#_c_1058_n N_VGND_c_1296_n 0.00828806f $X=8.695 $Y=0.82 $X2=0
+ $Y2=0
cc_715 N_A_27_47#_c_1163_n N_VGND_c_1296_n 0.0121741f $X=8.86 $Y=0.38 $X2=0
+ $Y2=0
cc_716 N_A_27_47#_c_1059_n N_VGND_c_1296_n 0.00828806f $X=9.535 $Y=0.82 $X2=0
+ $Y2=0
cc_717 N_A_27_47#_c_1060_n N_VGND_c_1296_n 0.0123792f $X=9.7 $Y=0.38 $X2=0 $Y2=0

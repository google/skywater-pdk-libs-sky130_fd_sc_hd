* File: sky130_fd_sc_hd__bufbuf_8.pxi.spice
* Created: Thu Aug 27 14:10:21 2020
* 
x_PM_SKY130_FD_SC_HD__BUFBUF_8%A N_A_M1022_g N_A_M1018_g A N_A_c_142_n
+ PM_SKY130_FD_SC_HD__BUFBUF_8%A
x_PM_SKY130_FD_SC_HD__BUFBUF_8%A_27_47# N_A_27_47#_M1022_s N_A_27_47#_M1018_s
+ N_A_27_47#_M1007_g N_A_27_47#_M1023_g N_A_27_47#_c_170_n N_A_27_47#_c_177_n
+ N_A_27_47#_c_171_n N_A_27_47#_c_172_n N_A_27_47#_c_178_n N_A_27_47#_c_179_n
+ N_A_27_47#_c_173_n N_A_27_47#_c_174_n N_A_27_47#_c_175_n
+ PM_SKY130_FD_SC_HD__BUFBUF_8%A_27_47#
x_PM_SKY130_FD_SC_HD__BUFBUF_8%A_206_47# N_A_206_47#_M1007_d N_A_206_47#_M1023_d
+ N_A_206_47#_M1002_g N_A_206_47#_M1016_g N_A_206_47#_M1008_g
+ N_A_206_47#_M1020_g N_A_206_47#_M1025_g N_A_206_47#_M1021_g
+ N_A_206_47#_c_253_n N_A_206_47#_c_244_n N_A_206_47#_c_245_n
+ N_A_206_47#_c_246_n N_A_206_47#_c_254_n N_A_206_47#_c_247_n
+ N_A_206_47#_c_248_n N_A_206_47#_c_249_n PM_SKY130_FD_SC_HD__BUFBUF_8%A_206_47#
x_PM_SKY130_FD_SC_HD__BUFBUF_8%A_318_47# N_A_318_47#_M1002_d N_A_318_47#_M1008_d
+ N_A_318_47#_M1016_s N_A_318_47#_M1020_s N_A_318_47#_M1001_g
+ N_A_318_47#_M1000_g N_A_318_47#_M1003_g N_A_318_47#_M1006_g
+ N_A_318_47#_M1004_g N_A_318_47#_M1009_g N_A_318_47#_M1005_g
+ N_A_318_47#_M1010_g N_A_318_47#_M1011_g N_A_318_47#_M1015_g
+ N_A_318_47#_M1012_g N_A_318_47#_M1017_g N_A_318_47#_M1013_g
+ N_A_318_47#_M1019_g N_A_318_47#_M1014_g N_A_318_47#_M1024_g
+ N_A_318_47#_c_358_n N_A_318_47#_c_375_n N_A_318_47#_c_359_n
+ N_A_318_47#_c_360_n N_A_318_47#_c_376_n N_A_318_47#_c_377_n
+ N_A_318_47#_c_402_n N_A_318_47#_c_405_n N_A_318_47#_c_361_n
+ N_A_318_47#_c_362_n N_A_318_47#_c_363_n N_A_318_47#_c_364_n
+ N_A_318_47#_c_379_n N_A_318_47#_c_365_n N_A_318_47#_c_366_n
+ PM_SKY130_FD_SC_HD__BUFBUF_8%A_318_47#
x_PM_SKY130_FD_SC_HD__BUFBUF_8%VPWR N_VPWR_M1018_d N_VPWR_M1016_d N_VPWR_M1021_d
+ N_VPWR_M1006_d N_VPWR_M1010_d N_VPWR_M1017_d N_VPWR_M1024_d N_VPWR_c_581_n
+ N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n
+ N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n N_VPWR_c_591_n
+ N_VPWR_c_592_n N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n N_VPWR_c_596_n
+ N_VPWR_c_597_n N_VPWR_c_598_n VPWR N_VPWR_c_599_n N_VPWR_c_600_n
+ N_VPWR_c_580_n N_VPWR_c_602_n N_VPWR_c_603_n PM_SKY130_FD_SC_HD__BUFBUF_8%VPWR
x_PM_SKY130_FD_SC_HD__BUFBUF_8%X N_X_M1001_d N_X_M1004_d N_X_M1011_d N_X_M1013_d
+ N_X_M1000_s N_X_M1009_s N_X_M1015_s N_X_M1019_s N_X_c_703_n N_X_c_704_n
+ N_X_c_684_n N_X_c_685_n N_X_c_693_n N_X_c_694_n N_X_c_731_n N_X_c_735_n
+ N_X_c_686_n N_X_c_695_n N_X_c_747_n N_X_c_751_n N_X_c_687_n N_X_c_696_n
+ N_X_c_763_n N_X_c_766_n N_X_c_688_n N_X_c_697_n N_X_c_689_n N_X_c_698_n
+ N_X_c_690_n N_X_c_699_n N_X_c_691_n N_X_c_700_n X X
+ PM_SKY130_FD_SC_HD__BUFBUF_8%X
x_PM_SKY130_FD_SC_HD__BUFBUF_8%VGND N_VGND_M1022_d N_VGND_M1002_s N_VGND_M1025_s
+ N_VGND_M1003_s N_VGND_M1005_s N_VGND_M1012_s N_VGND_M1014_s N_VGND_c_847_n
+ N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n N_VGND_c_852_n
+ N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n N_VGND_c_857_n
+ N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n N_VGND_c_862_n
+ N_VGND_c_863_n N_VGND_c_864_n VGND N_VGND_c_865_n N_VGND_c_866_n
+ N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n PM_SKY130_FD_SC_HD__BUFBUF_8%VGND
cc_1 VNB N_A_M1022_g 0.0365152f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_142_n 0.0382658f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_47#_c_170_n 0.0188691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_c_171_n 0.00168076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_172_n 0.00952728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_173_n 0.00752922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_174_n 0.0240805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_175_n 0.0200736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_206_47#_M1002_g 0.0215628f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_11 VNB N_A_206_47#_M1016_g 5.45489e-19 $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_12 VNB N_A_206_47#_M1008_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_206_47#_M1020_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_206_47#_M1025_g 0.0175122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_206_47#_M1021_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_206_47#_c_244_n 0.00535692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_206_47#_c_245_n 0.0194792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_206_47#_c_246_n 0.00655664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_206_47#_c_247_n 7.03049e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_206_47#_c_248_n 0.00238516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_206_47#_c_249_n 0.0498731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_318_47#_M1001_g 0.0176384f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_23 VNB N_A_318_47#_M1000_g 4.62868e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_318_47#_M1003_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_318_47#_M1006_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_318_47#_M1004_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_318_47#_M1009_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_318_47#_M1005_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_318_47#_M1010_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_318_47#_M1011_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_318_47#_M1015_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_318_47#_M1012_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_318_47#_M1017_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_318_47#_M1013_g 0.0172996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_318_47#_M1019_g 4.50112e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_318_47#_M1014_g 0.0210056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_318_47#_M1024_g 5.05833e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_318_47#_c_358_n 0.00443915f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_318_47#_c_359_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_318_47#_c_360_n 0.00437286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_318_47#_c_361_n 0.00354558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_318_47#_c_362_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_318_47#_c_363_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_318_47#_c_364_n 0.00345692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_318_47#_c_365_n 0.0013705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_318_47#_c_366_n 0.129098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VPWR_c_580_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_684_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_X_c_685_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_X_c_686_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_X_c_687_n 0.00308894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_X_c_688_n 0.0176068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_X_c_689_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_X_c_690_n 0.00222994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_X_c_691_n 0.00308159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB X 0.0251467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_847_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_848_n 0.0334581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_849_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_850_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_851_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_852_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_853_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_854_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_855_n 0.0168651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_856_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_857_n 0.0174747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_858_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_859_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_860_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_861_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_862_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_863_n 0.0168468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_864_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_865_n 0.0173377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_866_n 0.0159811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_867_n 0.34545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_868_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_869_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VPB N_A_M1018_g 0.0270892f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.805
cc_81 VPB N_A_c_142_n 0.00905856f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_82 VPB N_A_27_47#_M1023_g 0.0253519f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_83 VPB N_A_27_47#_c_177_n 0.0247548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_178_n 8.47385e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_179_n 0.00916145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_173_n 0.00599891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_27_47#_c_174_n 0.00499463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_206_47#_M1016_g 0.023984f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_89 VPB N_A_206_47#_M1020_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_206_47#_M1021_g 0.0194268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_206_47#_c_253_n 0.0082657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_206_47#_c_254_n 0.0019845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_206_47#_c_247_n 0.00515443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_318_47#_M1000_g 0.0196632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_318_47#_M1006_g 0.0191654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_318_47#_M1009_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_318_47#_M1010_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_318_47#_M1015_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_318_47#_M1017_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_318_47#_M1019_g 0.0191828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_318_47#_M1024_g 0.0233343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_318_47#_c_375_n 0.00772239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_318_47#_c_376_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_318_47#_c_377_n 0.00444397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_318_47#_c_362_n 0.00301948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_318_47#_c_379_n 0.00360324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_581_n 0.0138494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_582_n 0.0339308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_583_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_584_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_585_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_586_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_587_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_588_n 0.00416524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_589_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_590_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_591_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_592_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_593_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_594_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_595_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_596_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_597_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_598_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_599_n 0.0193829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_600_n 0.0174178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_580_n 0.073988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_602_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_603_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_X_c_693_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_X_c_694_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_X_c_695_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_X_c_696_n 0.00309768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_X_c_697_n 0.00317615f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_X_c_698_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_X_c_699_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_X_c_700_n 0.00309026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB X 0.00876037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB X 0.0236103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 N_A_M1018_g N_A_27_47#_M1023_g 0.0219942f $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_141 N_A_M1022_g N_A_27_47#_c_170_n 0.00852486f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_M1018_g N_A_27_47#_c_177_n 0.00823618f $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_143 N_A_M1022_g N_A_27_47#_c_171_n 0.00951801f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_144 A N_A_27_47#_c_171_n 9.95686e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A_M1022_g N_A_27_47#_c_172_n 0.00432116f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_146 A N_A_27_47#_c_172_n 0.0254341f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A_c_142_n N_A_27_47#_c_172_n 0.00729231f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_M1018_g N_A_27_47#_c_178_n 0.0115545f $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_149 A N_A_27_47#_c_178_n 9.95686e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A_M1018_g N_A_27_47#_c_179_n 0.00167422f $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_151 A N_A_27_47#_c_179_n 0.02566f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A_c_142_n N_A_27_47#_c_179_n 0.00705182f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_M1022_g N_A_27_47#_c_173_n 0.0081897f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_154 A N_A_27_47#_c_173_n 0.0161599f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_c_142_n N_A_27_47#_c_174_n 0.0157425f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_M1022_g N_A_27_47#_c_175_n 0.0229168f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A_M1022_g N_A_206_47#_c_246_n 6.25469e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_M1018_g N_A_206_47#_c_254_n 6.64196e-19 $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_159 N_A_M1018_g N_VPWR_c_581_n 0.0026193f $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_160 N_A_M1018_g N_VPWR_c_599_n 0.00411454f $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_161 N_A_M1018_g N_VPWR_c_580_n 0.00474973f $X=0.47 $Y=1.805 $X2=0 $Y2=0
cc_162 N_A_M1022_g N_VGND_c_847_n 0.00278284f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_M1022_g N_VGND_c_865_n 0.00424619f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_M1022_g N_VGND_c_867_n 0.00694488f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_27_47#_M1023_g N_A_206_47#_c_253_n 0.00949196f $X=0.955 $Y=1.985
+ $X2=0 $Y2=0
cc_166 N_A_27_47#_c_173_n N_A_206_47#_c_244_n 0.013229f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_174_n N_A_206_47#_c_244_n 0.00184284f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_175_n N_A_206_47#_c_244_n 0.00264865f $X=0.947 $Y=0.995
+ $X2=0 $Y2=0
cc_169 N_A_27_47#_c_170_n N_A_206_47#_c_246_n 0.00470936f $X=0.26 $Y=0.47 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_173_n N_A_206_47#_c_246_n 0.00878707f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_174_n N_A_206_47#_c_246_n 0.0010811f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_175_n N_A_206_47#_c_246_n 0.00856287f $X=0.947 $Y=0.995
+ $X2=0 $Y2=0
cc_173 N_A_27_47#_M1023_g N_A_206_47#_c_254_n 0.00352886f $X=0.955 $Y=1.985
+ $X2=0 $Y2=0
cc_174 N_A_27_47#_c_177_n N_A_206_47#_c_254_n 0.00469532f $X=0.26 $Y=1.63 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_173_n N_A_206_47#_c_254_n 0.00695096f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_174_n N_A_206_47#_c_254_n 0.00102817f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_M1023_g N_A_206_47#_c_247_n 0.003729f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_173_n N_A_206_47#_c_247_n 0.0129861f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_174_n N_A_206_47#_c_247_n 0.00115087f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_173_n N_A_206_47#_c_248_n 0.0172594f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_174_n N_A_206_47#_c_248_n 0.00480542f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_173_n N_VPWR_M1018_d 0.00417893f $X=0.955 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_183 N_A_27_47#_M1023_g N_VPWR_c_581_n 0.0126293f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_177_n N_VPWR_c_581_n 0.0153501f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_178_n N_VPWR_c_581_n 6.14392e-19 $X=0.61 $Y=1.53 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_173_n N_VPWR_c_581_n 0.0138849f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_47#_M1023_g N_VPWR_c_582_n 0.00541359f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_177_n N_VPWR_c_599_n 0.00780663f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_189 N_A_27_47#_M1023_g N_VPWR_c_580_n 0.0124033f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_177_n N_VPWR_c_580_n 0.010413f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_173_n N_VGND_M1022_d 0.00371268f $X=0.955 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_192 N_A_27_47#_c_171_n N_VGND_c_847_n 8.13279e-19 $X=0.61 $Y=0.82 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_173_n N_VGND_c_847_n 0.0133682f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_175_n N_VGND_c_847_n 0.00530447f $X=0.947 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_173_n N_VGND_c_848_n 2.28683e-19 $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_175_n N_VGND_c_848_n 0.00541562f $X=0.947 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_170_n N_VGND_c_865_n 0.0203493f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_171_n N_VGND_c_865_n 0.00230723f $X=0.61 $Y=0.82 $X2=0 $Y2=0
cc_199 N_A_27_47#_M1022_s N_VGND_c_867_n 0.00210264f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_170_n N_VGND_c_867_n 0.0124514f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_171_n N_VGND_c_867_n 0.00386518f $X=0.61 $Y=0.82 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_173_n N_VGND_c_867_n 0.00111682f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_175_n N_VGND_c_867_n 0.0112121f $X=0.947 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_206_47#_M1025_g N_A_318_47#_M1001_g 0.021435f $X=2.765 $Y=0.56 $X2=0
+ $Y2=0
cc_205 N_A_206_47#_M1021_g N_A_318_47#_M1000_g 0.021435f $X=2.765 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_206_47#_M1002_g N_A_318_47#_c_358_n 0.00636826f $X=1.925 $Y=0.56
+ $X2=0 $Y2=0
cc_207 N_A_206_47#_M1008_g N_A_318_47#_c_358_n 5.23702e-19 $X=2.345 $Y=0.56
+ $X2=0 $Y2=0
cc_208 N_A_206_47#_c_246_n N_A_318_47#_c_358_n 0.0399373f $X=1.165 $Y=0.4 $X2=0
+ $Y2=0
cc_209 N_A_206_47#_M1016_g N_A_318_47#_c_375_n 0.0102729f $X=1.925 $Y=1.985
+ $X2=0 $Y2=0
cc_210 N_A_206_47#_M1020_g N_A_318_47#_c_375_n 6.98608e-19 $X=2.345 $Y=1.985
+ $X2=0 $Y2=0
cc_211 N_A_206_47#_c_254_n N_A_318_47#_c_375_n 0.0714571f $X=1.165 $Y=1.63 $X2=0
+ $Y2=0
cc_212 N_A_206_47#_M1002_g N_A_318_47#_c_359_n 0.00850187f $X=1.925 $Y=0.56
+ $X2=0 $Y2=0
cc_213 N_A_206_47#_M1008_g N_A_318_47#_c_359_n 0.00850187f $X=2.345 $Y=0.56
+ $X2=0 $Y2=0
cc_214 N_A_206_47#_c_245_n N_A_318_47#_c_359_n 0.0596152f $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_215 N_A_206_47#_c_249_n N_A_318_47#_c_359_n 0.00205431f $X=2.765 $Y=1.16
+ $X2=0 $Y2=0
cc_216 N_A_206_47#_M1002_g N_A_318_47#_c_360_n 0.00126794f $X=1.925 $Y=0.56
+ $X2=0 $Y2=0
cc_217 N_A_206_47#_c_245_n N_A_318_47#_c_360_n 0.0278128f $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_218 N_A_206_47#_c_246_n N_A_318_47#_c_360_n 0.0147614f $X=1.165 $Y=0.4 $X2=0
+ $Y2=0
cc_219 N_A_206_47#_M1016_g N_A_318_47#_c_376_n 0.0107189f $X=1.925 $Y=1.985
+ $X2=0 $Y2=0
cc_220 N_A_206_47#_M1020_g N_A_318_47#_c_376_n 0.0107189f $X=2.345 $Y=1.985
+ $X2=0 $Y2=0
cc_221 N_A_206_47#_c_245_n N_A_318_47#_c_376_n 0.0596157f $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_222 N_A_206_47#_c_249_n N_A_318_47#_c_376_n 0.00198252f $X=2.765 $Y=1.16
+ $X2=0 $Y2=0
cc_223 N_A_206_47#_M1016_g N_A_318_47#_c_377_n 0.00168781f $X=1.925 $Y=1.985
+ $X2=0 $Y2=0
cc_224 N_A_206_47#_c_245_n N_A_318_47#_c_377_n 0.0279329f $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_225 N_A_206_47#_c_247_n N_A_318_47#_c_377_n 0.0146634f $X=1.19 $Y=1.545 $X2=0
+ $Y2=0
cc_226 N_A_206_47#_M1002_g N_A_318_47#_c_402_n 5.24491e-19 $X=1.925 $Y=0.56
+ $X2=0 $Y2=0
cc_227 N_A_206_47#_M1008_g N_A_318_47#_c_402_n 0.00647394f $X=2.345 $Y=0.56
+ $X2=0 $Y2=0
cc_228 N_A_206_47#_M1025_g N_A_318_47#_c_402_n 0.00647394f $X=2.765 $Y=0.56
+ $X2=0 $Y2=0
cc_229 N_A_206_47#_M1016_g N_A_318_47#_c_405_n 6.99397e-19 $X=1.925 $Y=1.985
+ $X2=0 $Y2=0
cc_230 N_A_206_47#_M1020_g N_A_318_47#_c_405_n 0.0103785f $X=2.345 $Y=1.985
+ $X2=0 $Y2=0
cc_231 N_A_206_47#_M1021_g N_A_318_47#_c_405_n 0.0103785f $X=2.765 $Y=1.985
+ $X2=0 $Y2=0
cc_232 N_A_206_47#_M1025_g N_A_318_47#_c_361_n 0.00412488f $X=2.765 $Y=0.56
+ $X2=0 $Y2=0
cc_233 N_A_206_47#_c_249_n N_A_318_47#_c_362_n 0.00407173f $X=2.765 $Y=1.16
+ $X2=0 $Y2=0
cc_234 N_A_206_47#_M1008_g N_A_318_47#_c_364_n 0.00123754f $X=2.345 $Y=0.56
+ $X2=0 $Y2=0
cc_235 N_A_206_47#_M1025_g N_A_318_47#_c_364_n 0.0107176f $X=2.765 $Y=0.56 $X2=0
+ $Y2=0
cc_236 N_A_206_47#_c_249_n N_A_318_47#_c_364_n 0.00205431f $X=2.765 $Y=1.16
+ $X2=0 $Y2=0
cc_237 N_A_206_47#_M1020_g N_A_318_47#_c_379_n 0.00139111f $X=2.345 $Y=1.985
+ $X2=0 $Y2=0
cc_238 N_A_206_47#_M1021_g N_A_318_47#_c_379_n 0.0131306f $X=2.765 $Y=1.985
+ $X2=0 $Y2=0
cc_239 N_A_206_47#_c_249_n N_A_318_47#_c_379_n 0.00198252f $X=2.765 $Y=1.16
+ $X2=0 $Y2=0
cc_240 N_A_206_47#_c_245_n N_A_318_47#_c_365_n 0.0176501f $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_241 N_A_206_47#_c_249_n N_A_318_47#_c_365_n 0.00200384f $X=2.765 $Y=1.16
+ $X2=0 $Y2=0
cc_242 N_A_206_47#_c_249_n N_A_318_47#_c_366_n 0.021435f $X=2.765 $Y=1.16 $X2=0
+ $Y2=0
cc_243 N_A_206_47#_c_253_n N_VPWR_c_581_n 0.0395707f $X=1.165 $Y=2.31 $X2=0
+ $Y2=0
cc_244 N_A_206_47#_M1016_g N_VPWR_c_582_n 0.00541359f $X=1.925 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_A_206_47#_c_253_n N_VPWR_c_582_n 0.0246229f $X=1.165 $Y=2.31 $X2=0
+ $Y2=0
cc_246 N_A_206_47#_M1016_g N_VPWR_c_583_n 0.0027696f $X=1.925 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_206_47#_M1020_g N_VPWR_c_583_n 0.00154685f $X=2.345 $Y=1.985 $X2=0
+ $Y2=0
cc_248 N_A_206_47#_M1021_g N_VPWR_c_584_n 0.00154685f $X=2.765 $Y=1.985 $X2=0
+ $Y2=0
cc_249 N_A_206_47#_M1020_g N_VPWR_c_589_n 0.00541359f $X=2.345 $Y=1.985 $X2=0
+ $Y2=0
cc_250 N_A_206_47#_M1021_g N_VPWR_c_589_n 0.00541359f $X=2.765 $Y=1.985 $X2=0
+ $Y2=0
cc_251 N_A_206_47#_M1023_d N_VPWR_c_580_n 0.00209319f $X=1.03 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_206_47#_M1016_g N_VPWR_c_580_n 0.0108276f $X=1.925 $Y=1.985 $X2=0
+ $Y2=0
cc_253 N_A_206_47#_M1020_g N_VPWR_c_580_n 0.00950154f $X=2.345 $Y=1.985 $X2=0
+ $Y2=0
cc_254 N_A_206_47#_M1021_g N_VPWR_c_580_n 0.00952874f $X=2.765 $Y=1.985 $X2=0
+ $Y2=0
cc_255 N_A_206_47#_c_253_n N_VPWR_c_580_n 0.0143524f $X=1.165 $Y=2.31 $X2=0
+ $Y2=0
cc_256 N_A_206_47#_M1025_g N_X_c_703_n 5.23702e-19 $X=2.765 $Y=0.56 $X2=0 $Y2=0
cc_257 N_A_206_47#_M1021_g N_X_c_704_n 6.98608e-19 $X=2.765 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_206_47#_c_246_n N_VGND_c_847_n 0.0177486f $X=1.165 $Y=0.4 $X2=0 $Y2=0
cc_259 N_A_206_47#_M1002_g N_VGND_c_848_n 0.00424619f $X=1.925 $Y=0.56 $X2=0
+ $Y2=0
cc_260 N_A_206_47#_c_246_n N_VGND_c_848_n 0.0237276f $X=1.165 $Y=0.4 $X2=0 $Y2=0
cc_261 N_A_206_47#_M1002_g N_VGND_c_849_n 0.00268723f $X=1.925 $Y=0.56 $X2=0
+ $Y2=0
cc_262 N_A_206_47#_M1008_g N_VGND_c_849_n 0.00146448f $X=2.345 $Y=0.56 $X2=0
+ $Y2=0
cc_263 N_A_206_47#_M1025_g N_VGND_c_850_n 0.00146448f $X=2.765 $Y=0.56 $X2=0
+ $Y2=0
cc_264 N_A_206_47#_M1008_g N_VGND_c_855_n 0.00423644f $X=2.345 $Y=0.56 $X2=0
+ $Y2=0
cc_265 N_A_206_47#_M1025_g N_VGND_c_855_n 0.00423644f $X=2.765 $Y=0.56 $X2=0
+ $Y2=0
cc_266 N_A_206_47#_M1007_d N_VGND_c_867_n 0.0020946f $X=1.03 $Y=0.235 $X2=0
+ $Y2=0
cc_267 N_A_206_47#_M1002_g N_VGND_c_867_n 0.00706231f $X=1.925 $Y=0.56 $X2=0
+ $Y2=0
cc_268 N_A_206_47#_M1008_g N_VGND_c_867_n 0.00575105f $X=2.345 $Y=0.56 $X2=0
+ $Y2=0
cc_269 N_A_206_47#_M1025_g N_VGND_c_867_n 0.00577825f $X=2.765 $Y=0.56 $X2=0
+ $Y2=0
cc_270 N_A_206_47#_c_246_n N_VGND_c_867_n 0.0142792f $X=1.165 $Y=0.4 $X2=0 $Y2=0
cc_271 N_A_318_47#_c_376_n N_VPWR_M1016_d 0.00165831f $X=2.39 $Y=1.53 $X2=0
+ $Y2=0
cc_272 N_A_318_47#_c_379_n N_VPWR_M1021_d 0.00187252f $X=2.975 $Y=1.53 $X2=0
+ $Y2=0
cc_273 N_A_318_47#_c_375_n N_VPWR_c_582_n 0.0210382f $X=1.715 $Y=1.63 $X2=0
+ $Y2=0
cc_274 N_A_318_47#_c_376_n N_VPWR_c_583_n 0.0126919f $X=2.39 $Y=1.53 $X2=0 $Y2=0
cc_275 N_A_318_47#_M1000_g N_VPWR_c_584_n 0.00154685f $X=3.185 $Y=1.985 $X2=0
+ $Y2=0
cc_276 N_A_318_47#_c_379_n N_VPWR_c_584_n 0.0126919f $X=2.975 $Y=1.53 $X2=0
+ $Y2=0
cc_277 N_A_318_47#_M1006_g N_VPWR_c_585_n 0.00146448f $X=3.605 $Y=1.985 $X2=0
+ $Y2=0
cc_278 N_A_318_47#_M1009_g N_VPWR_c_585_n 0.00146448f $X=4.025 $Y=1.985 $X2=0
+ $Y2=0
cc_279 N_A_318_47#_M1010_g N_VPWR_c_586_n 0.00146448f $X=4.445 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A_318_47#_M1015_g N_VPWR_c_586_n 0.00146448f $X=4.865 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_A_318_47#_M1017_g N_VPWR_c_587_n 0.00146448f $X=5.285 $Y=1.985 $X2=0
+ $Y2=0
cc_282 N_A_318_47#_M1019_g N_VPWR_c_587_n 0.00146448f $X=5.705 $Y=1.985 $X2=0
+ $Y2=0
cc_283 N_A_318_47#_M1024_g N_VPWR_c_588_n 0.00316354f $X=6.125 $Y=1.985 $X2=0
+ $Y2=0
cc_284 N_A_318_47#_c_405_n N_VPWR_c_589_n 0.0189039f $X=2.555 $Y=1.63 $X2=0
+ $Y2=0
cc_285 N_A_318_47#_M1000_g N_VPWR_c_591_n 0.00541359f $X=3.185 $Y=1.985 $X2=0
+ $Y2=0
cc_286 N_A_318_47#_M1006_g N_VPWR_c_591_n 0.00541359f $X=3.605 $Y=1.985 $X2=0
+ $Y2=0
cc_287 N_A_318_47#_M1009_g N_VPWR_c_593_n 0.00541359f $X=4.025 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_318_47#_M1010_g N_VPWR_c_593_n 0.00541359f $X=4.445 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_A_318_47#_M1015_g N_VPWR_c_595_n 0.00541359f $X=4.865 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_A_318_47#_M1017_g N_VPWR_c_595_n 0.00541359f $X=5.285 $Y=1.985 $X2=0
+ $Y2=0
cc_291 N_A_318_47#_M1019_g N_VPWR_c_597_n 0.00541359f $X=5.705 $Y=1.985 $X2=0
+ $Y2=0
cc_292 N_A_318_47#_M1024_g N_VPWR_c_597_n 0.00541359f $X=6.125 $Y=1.985 $X2=0
+ $Y2=0
cc_293 N_A_318_47#_M1016_s N_VPWR_c_580_n 0.00209319f $X=1.59 $Y=1.485 $X2=0
+ $Y2=0
cc_294 N_A_318_47#_M1020_s N_VPWR_c_580_n 0.00215201f $X=2.42 $Y=1.485 $X2=0
+ $Y2=0
cc_295 N_A_318_47#_M1000_g N_VPWR_c_580_n 0.00952874f $X=3.185 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_318_47#_M1006_g N_VPWR_c_580_n 0.00950154f $X=3.605 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_A_318_47#_M1009_g N_VPWR_c_580_n 0.00950154f $X=4.025 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_318_47#_M1010_g N_VPWR_c_580_n 0.00950154f $X=4.445 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A_318_47#_M1015_g N_VPWR_c_580_n 0.00950154f $X=4.865 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_A_318_47#_M1017_g N_VPWR_c_580_n 0.00950154f $X=5.285 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A_318_47#_M1019_g N_VPWR_c_580_n 0.00950154f $X=5.705 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_A_318_47#_M1024_g N_VPWR_c_580_n 0.0106471f $X=6.125 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_318_47#_c_375_n N_VPWR_c_580_n 0.0124268f $X=1.715 $Y=1.63 $X2=0
+ $Y2=0
cc_304 N_A_318_47#_c_405_n N_VPWR_c_580_n 0.0122217f $X=2.555 $Y=1.63 $X2=0
+ $Y2=0
cc_305 N_A_318_47#_M1001_g N_X_c_703_n 0.00636826f $X=3.185 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A_318_47#_M1003_g N_X_c_703_n 0.00636826f $X=3.605 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A_318_47#_M1004_g N_X_c_703_n 5.23702e-19 $X=4.025 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A_318_47#_c_402_n N_X_c_703_n 0.00518536f $X=2.555 $Y=0.4 $X2=0 $Y2=0
cc_309 N_A_318_47#_M1000_g N_X_c_704_n 0.0102729f $X=3.185 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_318_47#_M1006_g N_X_c_704_n 0.0106215f $X=3.605 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A_318_47#_M1009_g N_X_c_704_n 7.66249e-19 $X=4.025 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A_318_47#_c_405_n N_X_c_704_n 0.00518536f $X=2.555 $Y=1.63 $X2=0 $Y2=0
cc_313 N_A_318_47#_M1003_g N_X_c_684_n 0.00850187f $X=3.605 $Y=0.56 $X2=0 $Y2=0
cc_314 N_A_318_47#_M1004_g N_X_c_684_n 0.00850187f $X=4.025 $Y=0.56 $X2=0 $Y2=0
cc_315 N_A_318_47#_c_363_n N_X_c_684_n 0.0359512f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_318_47#_c_366_n N_X_c_684_n 0.00205431f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_318_47#_M1001_g N_X_c_685_n 0.00240257f $X=3.185 $Y=0.56 $X2=0 $Y2=0
cc_318 N_A_318_47#_M1003_g N_X_c_685_n 0.00109384f $X=3.605 $Y=0.56 $X2=0 $Y2=0
cc_319 N_A_318_47#_c_363_n N_X_c_685_n 0.0265235f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_318_47#_c_364_n N_X_c_685_n 0.00795337f $X=2.975 $Y=0.82 $X2=0 $Y2=0
cc_321 N_A_318_47#_c_366_n N_X_c_685_n 0.00213376f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A_318_47#_M1006_g N_X_c_693_n 0.0107189f $X=3.605 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_318_47#_M1009_g N_X_c_693_n 0.0107189f $X=4.025 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A_318_47#_c_363_n N_X_c_693_n 0.0359514f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_318_47#_c_366_n N_X_c_693_n 0.00198252f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A_318_47#_M1000_g N_X_c_694_n 0.00265135f $X=3.185 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A_318_47#_M1006_g N_X_c_694_n 0.00134262f $X=3.605 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_318_47#_c_363_n N_X_c_694_n 0.026643f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_318_47#_c_379_n N_X_c_694_n 0.0088897f $X=2.975 $Y=1.53 $X2=0 $Y2=0
cc_330 N_A_318_47#_c_366_n N_X_c_694_n 0.00206439f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_318_47#_M1003_g N_X_c_731_n 5.23702e-19 $X=3.605 $Y=0.56 $X2=0 $Y2=0
cc_332 N_A_318_47#_M1004_g N_X_c_731_n 0.00636826f $X=4.025 $Y=0.56 $X2=0 $Y2=0
cc_333 N_A_318_47#_M1005_g N_X_c_731_n 0.00636826f $X=4.445 $Y=0.56 $X2=0 $Y2=0
cc_334 N_A_318_47#_M1011_g N_X_c_731_n 5.23702e-19 $X=4.865 $Y=0.56 $X2=0 $Y2=0
cc_335 N_A_318_47#_M1006_g N_X_c_735_n 7.66249e-19 $X=3.605 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_318_47#_M1009_g N_X_c_735_n 0.0106215f $X=4.025 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_318_47#_M1010_g N_X_c_735_n 0.0106215f $X=4.445 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A_318_47#_M1015_g N_X_c_735_n 7.66249e-19 $X=4.865 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A_318_47#_M1005_g N_X_c_686_n 0.00850187f $X=4.445 $Y=0.56 $X2=0 $Y2=0
cc_340 N_A_318_47#_M1011_g N_X_c_686_n 0.00850187f $X=4.865 $Y=0.56 $X2=0 $Y2=0
cc_341 N_A_318_47#_c_363_n N_X_c_686_n 0.0359512f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_342 N_A_318_47#_c_366_n N_X_c_686_n 0.00205431f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_318_47#_M1010_g N_X_c_695_n 0.0107189f $X=4.445 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A_318_47#_M1015_g N_X_c_695_n 0.0107189f $X=4.865 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A_318_47#_c_363_n N_X_c_695_n 0.0359514f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A_318_47#_c_366_n N_X_c_695_n 0.00198252f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A_318_47#_M1005_g N_X_c_747_n 5.23702e-19 $X=4.445 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A_318_47#_M1011_g N_X_c_747_n 0.00636826f $X=4.865 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A_318_47#_M1012_g N_X_c_747_n 0.00636826f $X=5.285 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A_318_47#_M1013_g N_X_c_747_n 5.23702e-19 $X=5.705 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A_318_47#_M1010_g N_X_c_751_n 7.66249e-19 $X=4.445 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A_318_47#_M1015_g N_X_c_751_n 0.0106215f $X=4.865 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A_318_47#_M1017_g N_X_c_751_n 0.0106215f $X=5.285 $Y=1.985 $X2=0 $Y2=0
cc_354 N_A_318_47#_M1019_g N_X_c_751_n 7.66249e-19 $X=5.705 $Y=1.985 $X2=0 $Y2=0
cc_355 N_A_318_47#_M1012_g N_X_c_687_n 0.00850187f $X=5.285 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_318_47#_M1013_g N_X_c_687_n 0.00985957f $X=5.705 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_318_47#_c_363_n N_X_c_687_n 0.00820272f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_358 N_A_318_47#_c_366_n N_X_c_687_n 0.00243099f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_359 N_A_318_47#_M1017_g N_X_c_696_n 0.0107189f $X=5.285 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A_318_47#_M1019_g N_X_c_696_n 0.0120766f $X=5.705 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A_318_47#_c_363_n N_X_c_696_n 0.00820272f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_362 N_A_318_47#_c_366_n N_X_c_696_n 0.00233927f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_363 N_A_318_47#_M1012_g N_X_c_763_n 5.23702e-19 $X=5.285 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A_318_47#_M1013_g N_X_c_763_n 0.00636826f $X=5.705 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A_318_47#_M1014_g N_X_c_763_n 0.0109928f $X=6.125 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A_318_47#_M1017_g N_X_c_766_n 7.66249e-19 $X=5.285 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A_318_47#_M1019_g N_X_c_766_n 0.0106215f $X=5.705 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A_318_47#_M1024_g N_X_c_766_n 0.0167471f $X=6.125 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A_318_47#_M1014_g N_X_c_688_n 0.0118401f $X=6.125 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_318_47#_M1024_g N_X_c_697_n 0.0140571f $X=6.125 $Y=1.985 $X2=0 $Y2=0
cc_371 N_A_318_47#_M1004_g N_X_c_689_n 0.00110541f $X=4.025 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_318_47#_M1005_g N_X_c_689_n 0.00110541f $X=4.445 $Y=0.56 $X2=0 $Y2=0
cc_373 N_A_318_47#_c_363_n N_X_c_689_n 0.0265235f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_318_47#_c_366_n N_X_c_689_n 0.00213376f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_375 N_A_318_47#_M1009_g N_X_c_698_n 0.00135419f $X=4.025 $Y=1.985 $X2=0 $Y2=0
cc_376 N_A_318_47#_M1010_g N_X_c_698_n 0.00135419f $X=4.445 $Y=1.985 $X2=0 $Y2=0
cc_377 N_A_318_47#_c_363_n N_X_c_698_n 0.026643f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_378 N_A_318_47#_c_366_n N_X_c_698_n 0.00206439f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A_318_47#_M1011_g N_X_c_690_n 0.00110541f $X=4.865 $Y=0.56 $X2=0 $Y2=0
cc_380 N_A_318_47#_M1012_g N_X_c_690_n 0.00110541f $X=5.285 $Y=0.56 $X2=0 $Y2=0
cc_381 N_A_318_47#_c_363_n N_X_c_690_n 0.0265235f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_382 N_A_318_47#_c_366_n N_X_c_690_n 0.00213376f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_318_47#_M1015_g N_X_c_699_n 0.00135419f $X=4.865 $Y=1.985 $X2=0 $Y2=0
cc_384 N_A_318_47#_M1017_g N_X_c_699_n 0.00135419f $X=5.285 $Y=1.985 $X2=0 $Y2=0
cc_385 N_A_318_47#_c_363_n N_X_c_699_n 0.026643f $X=5.015 $Y=1.16 $X2=0 $Y2=0
cc_386 N_A_318_47#_c_366_n N_X_c_699_n 0.00206439f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A_318_47#_M1013_g N_X_c_691_n 0.00141219f $X=5.705 $Y=0.56 $X2=0 $Y2=0
cc_388 N_A_318_47#_M1014_g N_X_c_691_n 0.00141219f $X=6.125 $Y=0.56 $X2=0 $Y2=0
cc_389 N_A_318_47#_c_366_n N_X_c_691_n 0.00264592f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A_318_47#_M1019_g N_X_c_700_n 0.00167056f $X=5.705 $Y=1.985 $X2=0 $Y2=0
cc_391 N_A_318_47#_M1024_g N_X_c_700_n 0.00167056f $X=6.125 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A_318_47#_c_366_n N_X_c_700_n 0.00256174f $X=6.125 $Y=1.16 $X2=0 $Y2=0
cc_393 N_A_318_47#_M1014_g X 0.0207748f $X=6.125 $Y=0.56 $X2=0 $Y2=0
cc_394 N_A_318_47#_c_359_n N_VGND_M1002_s 0.00162006f $X=2.39 $Y=0.82 $X2=0
+ $Y2=0
cc_395 N_A_318_47#_c_364_n N_VGND_M1025_s 0.00186748f $X=2.975 $Y=0.82 $X2=0
+ $Y2=0
cc_396 N_A_318_47#_c_358_n N_VGND_c_848_n 0.020318f $X=1.715 $Y=0.4 $X2=0 $Y2=0
cc_397 N_A_318_47#_c_359_n N_VGND_c_848_n 0.00193763f $X=2.39 $Y=0.82 $X2=0
+ $Y2=0
cc_398 N_A_318_47#_c_359_n N_VGND_c_849_n 0.0122414f $X=2.39 $Y=0.82 $X2=0 $Y2=0
cc_399 N_A_318_47#_M1001_g N_VGND_c_850_n 0.00146448f $X=3.185 $Y=0.56 $X2=0
+ $Y2=0
cc_400 N_A_318_47#_c_364_n N_VGND_c_850_n 0.0122414f $X=2.975 $Y=0.82 $X2=0
+ $Y2=0
cc_401 N_A_318_47#_M1003_g N_VGND_c_851_n 0.00146448f $X=3.605 $Y=0.56 $X2=0
+ $Y2=0
cc_402 N_A_318_47#_M1004_g N_VGND_c_851_n 0.00146448f $X=4.025 $Y=0.56 $X2=0
+ $Y2=0
cc_403 N_A_318_47#_M1005_g N_VGND_c_852_n 0.00146448f $X=4.445 $Y=0.56 $X2=0
+ $Y2=0
cc_404 N_A_318_47#_M1011_g N_VGND_c_852_n 0.00146448f $X=4.865 $Y=0.56 $X2=0
+ $Y2=0
cc_405 N_A_318_47#_M1012_g N_VGND_c_853_n 0.00146448f $X=5.285 $Y=0.56 $X2=0
+ $Y2=0
cc_406 N_A_318_47#_M1013_g N_VGND_c_853_n 0.00146448f $X=5.705 $Y=0.56 $X2=0
+ $Y2=0
cc_407 N_A_318_47#_M1014_g N_VGND_c_854_n 0.00316354f $X=6.125 $Y=0.56 $X2=0
+ $Y2=0
cc_408 N_A_318_47#_c_359_n N_VGND_c_855_n 0.00390702f $X=2.39 $Y=0.82 $X2=0
+ $Y2=0
cc_409 N_A_318_47#_c_402_n N_VGND_c_855_n 0.0179571f $X=2.555 $Y=0.4 $X2=0 $Y2=0
cc_410 N_A_318_47#_M1001_g N_VGND_c_857_n 0.00541562f $X=3.185 $Y=0.56 $X2=0
+ $Y2=0
cc_411 N_A_318_47#_M1003_g N_VGND_c_857_n 0.00424619f $X=3.605 $Y=0.56 $X2=0
+ $Y2=0
cc_412 N_A_318_47#_M1004_g N_VGND_c_859_n 0.00424619f $X=4.025 $Y=0.56 $X2=0
+ $Y2=0
cc_413 N_A_318_47#_M1005_g N_VGND_c_859_n 0.00424619f $X=4.445 $Y=0.56 $X2=0
+ $Y2=0
cc_414 N_A_318_47#_M1011_g N_VGND_c_861_n 0.00424619f $X=4.865 $Y=0.56 $X2=0
+ $Y2=0
cc_415 N_A_318_47#_M1012_g N_VGND_c_861_n 0.00424619f $X=5.285 $Y=0.56 $X2=0
+ $Y2=0
cc_416 N_A_318_47#_M1013_g N_VGND_c_863_n 0.00424619f $X=5.705 $Y=0.56 $X2=0
+ $Y2=0
cc_417 N_A_318_47#_M1014_g N_VGND_c_863_n 0.00424619f $X=6.125 $Y=0.56 $X2=0
+ $Y2=0
cc_418 N_A_318_47#_M1002_d N_VGND_c_867_n 0.0020946f $X=1.59 $Y=0.235 $X2=0
+ $Y2=0
cc_419 N_A_318_47#_M1008_d N_VGND_c_867_n 0.00215347f $X=2.42 $Y=0.235 $X2=0
+ $Y2=0
cc_420 N_A_318_47#_M1001_g N_VGND_c_867_n 0.00952891f $X=3.185 $Y=0.56 $X2=0
+ $Y2=0
cc_421 N_A_318_47#_M1003_g N_VGND_c_867_n 0.00573624f $X=3.605 $Y=0.56 $X2=0
+ $Y2=0
cc_422 N_A_318_47#_M1004_g N_VGND_c_867_n 0.00573624f $X=4.025 $Y=0.56 $X2=0
+ $Y2=0
cc_423 N_A_318_47#_M1005_g N_VGND_c_867_n 0.00573624f $X=4.445 $Y=0.56 $X2=0
+ $Y2=0
cc_424 N_A_318_47#_M1011_g N_VGND_c_867_n 0.00573624f $X=4.865 $Y=0.56 $X2=0
+ $Y2=0
cc_425 N_A_318_47#_M1012_g N_VGND_c_867_n 0.00573624f $X=5.285 $Y=0.56 $X2=0
+ $Y2=0
cc_426 N_A_318_47#_M1013_g N_VGND_c_867_n 0.00573624f $X=5.705 $Y=0.56 $X2=0
+ $Y2=0
cc_427 N_A_318_47#_M1014_g N_VGND_c_867_n 0.0068818f $X=6.125 $Y=0.56 $X2=0
+ $Y2=0
cc_428 N_A_318_47#_c_358_n N_VGND_c_867_n 0.0123792f $X=1.715 $Y=0.4 $X2=0 $Y2=0
cc_429 N_A_318_47#_c_359_n N_VGND_c_867_n 0.012122f $X=2.39 $Y=0.82 $X2=0 $Y2=0
cc_430 N_A_318_47#_c_402_n N_VGND_c_867_n 0.0120759f $X=2.555 $Y=0.4 $X2=0 $Y2=0
cc_431 N_A_318_47#_c_364_n N_VGND_c_867_n 6.28727e-19 $X=2.975 $Y=0.82 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_580_n N_X_M1000_s 0.00215201f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_433 N_VPWR_c_580_n N_X_M1009_s 0.00215201f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_434 N_VPWR_c_580_n N_X_M1015_s 0.00215201f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_435 N_VPWR_c_580_n N_X_M1019_s 0.00215201f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_436 N_VPWR_c_591_n N_X_c_704_n 0.0189039f $X=3.73 $Y=2.72 $X2=0 $Y2=0
cc_437 N_VPWR_c_580_n N_X_c_704_n 0.0122217f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_438 N_VPWR_M1006_d N_X_c_693_n 0.00185611f $X=3.68 $Y=1.485 $X2=0 $Y2=0
cc_439 N_VPWR_c_585_n N_X_c_693_n 0.0104788f $X=3.815 $Y=2 $X2=0 $Y2=0
cc_440 N_VPWR_c_593_n N_X_c_735_n 0.0189039f $X=4.57 $Y=2.72 $X2=0 $Y2=0
cc_441 N_VPWR_c_580_n N_X_c_735_n 0.0122217f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_442 N_VPWR_M1010_d N_X_c_695_n 0.00185611f $X=4.52 $Y=1.485 $X2=0 $Y2=0
cc_443 N_VPWR_c_586_n N_X_c_695_n 0.0104788f $X=4.655 $Y=2 $X2=0 $Y2=0
cc_444 N_VPWR_c_595_n N_X_c_751_n 0.0189039f $X=5.41 $Y=2.72 $X2=0 $Y2=0
cc_445 N_VPWR_c_580_n N_X_c_751_n 0.0122217f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_M1017_d N_X_c_696_n 0.00185611f $X=5.36 $Y=1.485 $X2=0 $Y2=0
cc_447 N_VPWR_c_587_n N_X_c_696_n 0.0104788f $X=5.495 $Y=2 $X2=0 $Y2=0
cc_448 N_VPWR_c_597_n N_X_c_766_n 0.0189039f $X=6.25 $Y=2.72 $X2=0 $Y2=0
cc_449 N_VPWR_c_580_n N_X_c_766_n 0.0122217f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_M1024_d N_X_c_697_n 0.0028854f $X=6.2 $Y=1.485 $X2=0 $Y2=0
cc_451 N_VPWR_c_588_n N_X_c_697_n 0.0108818f $X=6.335 $Y=2 $X2=0 $Y2=0
cc_452 N_VPWR_M1024_d X 0.00130765f $X=6.2 $Y=1.485 $X2=0 $Y2=0
cc_453 N_X_c_684_n N_VGND_M1003_s 0.00162006f $X=4.07 $Y=0.82 $X2=0 $Y2=0
cc_454 N_X_c_686_n N_VGND_M1005_s 0.00162006f $X=4.91 $Y=0.82 $X2=0 $Y2=0
cc_455 N_X_c_687_n N_VGND_M1012_s 0.00162006f $X=5.75 $Y=0.82 $X2=0 $Y2=0
cc_456 N_X_c_688_n N_VGND_M1014_s 0.00311553f $X=6.435 $Y=0.82 $X2=0 $Y2=0
cc_457 N_X_c_684_n N_VGND_c_851_n 0.0122414f $X=4.07 $Y=0.82 $X2=0 $Y2=0
cc_458 N_X_c_686_n N_VGND_c_852_n 0.0122414f $X=4.91 $Y=0.82 $X2=0 $Y2=0
cc_459 N_X_c_687_n N_VGND_c_853_n 0.0122414f $X=5.75 $Y=0.82 $X2=0 $Y2=0
cc_460 N_X_c_688_n N_VGND_c_854_n 0.0127122f $X=6.435 $Y=0.82 $X2=0 $Y2=0
cc_461 N_X_c_703_n N_VGND_c_857_n 0.0182681f $X=3.395 $Y=0.4 $X2=0 $Y2=0
cc_462 N_X_c_684_n N_VGND_c_857_n 0.00193763f $X=4.07 $Y=0.82 $X2=0 $Y2=0
cc_463 N_X_c_684_n N_VGND_c_859_n 0.00193763f $X=4.07 $Y=0.82 $X2=0 $Y2=0
cc_464 N_X_c_731_n N_VGND_c_859_n 0.0182681f $X=4.235 $Y=0.4 $X2=0 $Y2=0
cc_465 N_X_c_686_n N_VGND_c_859_n 0.00193763f $X=4.91 $Y=0.82 $X2=0 $Y2=0
cc_466 N_X_c_686_n N_VGND_c_861_n 0.00193763f $X=4.91 $Y=0.82 $X2=0 $Y2=0
cc_467 N_X_c_747_n N_VGND_c_861_n 0.0182681f $X=5.075 $Y=0.4 $X2=0 $Y2=0
cc_468 N_X_c_687_n N_VGND_c_861_n 0.00193763f $X=5.75 $Y=0.82 $X2=0 $Y2=0
cc_469 N_X_c_687_n N_VGND_c_863_n 0.00193763f $X=5.75 $Y=0.82 $X2=0 $Y2=0
cc_470 N_X_c_763_n N_VGND_c_863_n 0.0182681f $X=5.915 $Y=0.4 $X2=0 $Y2=0
cc_471 N_X_c_688_n N_VGND_c_863_n 0.00193763f $X=6.435 $Y=0.82 $X2=0 $Y2=0
cc_472 N_X_c_688_n N_VGND_c_866_n 0.00652531f $X=6.435 $Y=0.82 $X2=0 $Y2=0
cc_473 N_X_M1001_d N_VGND_c_867_n 0.00215347f $X=3.26 $Y=0.235 $X2=0 $Y2=0
cc_474 N_X_M1004_d N_VGND_c_867_n 0.00215347f $X=4.1 $Y=0.235 $X2=0 $Y2=0
cc_475 N_X_M1011_d N_VGND_c_867_n 0.00215347f $X=4.94 $Y=0.235 $X2=0 $Y2=0
cc_476 N_X_M1013_d N_VGND_c_867_n 0.00215347f $X=5.78 $Y=0.235 $X2=0 $Y2=0
cc_477 N_X_c_703_n N_VGND_c_867_n 0.0121741f $X=3.395 $Y=0.4 $X2=0 $Y2=0
cc_478 N_X_c_684_n N_VGND_c_867_n 0.00825759f $X=4.07 $Y=0.82 $X2=0 $Y2=0
cc_479 N_X_c_731_n N_VGND_c_867_n 0.0121741f $X=4.235 $Y=0.4 $X2=0 $Y2=0
cc_480 N_X_c_686_n N_VGND_c_867_n 0.00825759f $X=4.91 $Y=0.82 $X2=0 $Y2=0
cc_481 N_X_c_747_n N_VGND_c_867_n 0.0121741f $X=5.075 $Y=0.4 $X2=0 $Y2=0
cc_482 N_X_c_687_n N_VGND_c_867_n 0.00825759f $X=5.75 $Y=0.82 $X2=0 $Y2=0
cc_483 N_X_c_763_n N_VGND_c_867_n 0.0121741f $X=5.915 $Y=0.4 $X2=0 $Y2=0
cc_484 N_X_c_688_n N_VGND_c_867_n 0.0154886f $X=6.435 $Y=0.82 $X2=0 $Y2=0

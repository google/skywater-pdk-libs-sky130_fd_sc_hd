* File: sky130_fd_sc_hd__a21o_2.spice
* Created: Tue Sep  1 18:52:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21o_2.pex.spice"
.subckt sky130_fd_sc_hd__a21o_2  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_X_M1003_d N_A_80_199#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1003_d N_A_80_199#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.1105 PD=0.93 PS=0.99 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_A_80_199#_M1001_d N_B1_M1001_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1625 AS=0.1105 PD=1.15 PS=0.99 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75001.1
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1006 A_458_47# N_A1_M1006_g N_A_80_199#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.1625 PD=1.03 PS=1.15 NRD=24.912 NRS=40.608 M=1 R=4.33333
+ SA=75001.8 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_458_47# VNB NSHORT L=0.15 W=0.65 AD=0.17225
+ AS=0.1235 PD=1.83 PS=1.03 NRD=0 NRS=24.912 M=1 R=4.33333 SA=75002.3 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1004_d N_A_80_199#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1004_d N_A_80_199#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_386_297#_M1002_d N_B1_M1002_g N_A_80_199#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_386_297#_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1575 AS=0.14 PD=1.315 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_386_297#_M1008_d N_A2_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1575 PD=2.52 PS=1.315 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a21o_2.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
M1000 Z A a_204_309# VPB phighvt w=1e+06u l=150000u
+  ad=5.193e+11p pd=5.08e+06u as=5.238e+11p ps=4.96e+06u
M1001 a_204_309# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR TE_B a_204_309# VPB phighvt w=940000u l=150000u
+  ad=5.24375e+11p pd=4.93e+06u as=0p ps=0u
M1003 a_214_120# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=5.586e+11p pd=5.63e+06u as=2.834e+11p ps=3.2e+06u
M1004 a_204_309# TE_B VPWR VPB phighvt w=940000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_27_47# a_214_120# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR TE_B a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1007 a_214_120# A Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1008 VGND TE_B a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1009 Z A a_214_120# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

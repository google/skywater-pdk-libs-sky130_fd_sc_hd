* File: sky130_fd_sc_hd__buf_1.spice.SKY130_FD_SC_HD__BUF_1.pxi
* Created: Thu Aug 27 14:09:37 2020
* 
x_PM_SKY130_FD_SC_HD__BUF_1%A N_A_c_37_n N_A_c_38_n N_A_M1003_g N_A_M1000_g
+ N_A_c_41_n N_A_c_42_n A PM_SKY130_FD_SC_HD__BUF_1%A
x_PM_SKY130_FD_SC_HD__BUF_1%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1000_s
+ N_A_27_47#_M1001_g N_A_27_47#_M1002_g N_A_27_47#_c_109_p N_A_27_47#_c_131_p
+ N_A_27_47#_c_72_n N_A_27_47#_c_73_n N_A_27_47#_c_78_n N_A_27_47#_c_79_n
+ N_A_27_47#_c_80_n N_A_27_47#_c_74_n N_A_27_47#_c_75_n N_A_27_47#_c_76_n
+ PM_SKY130_FD_SC_HD__BUF_1%A_27_47#
x_PM_SKY130_FD_SC_HD__BUF_1%VPWR N_VPWR_M1000_d N_VPWR_c_139_n VPWR VPWR
+ N_VPWR_c_140_n N_VPWR_c_141_n N_VPWR_c_138_n N_VPWR_c_143_n
+ PM_SKY130_FD_SC_HD__BUF_1%VPWR
x_PM_SKY130_FD_SC_HD__BUF_1%X N_X_M1001_d N_X_M1002_d N_X_c_163_n N_X_c_160_n
+ N_X_c_161_n X X X PM_SKY130_FD_SC_HD__BUF_1%X
x_PM_SKY130_FD_SC_HD__BUF_1%VGND N_VGND_M1003_d N_VGND_c_184_n VGND VGND
+ N_VGND_c_185_n VGND N_VGND_c_186_n N_VGND_c_187_n N_VGND_c_188_n
+ PM_SKY130_FD_SC_HD__BUF_1%VGND
cc_1 VNB N_A_c_37_n 0.0488646f $X=-0.19 $Y=-0.24 $X2=0.44 $Y2=1.325
cc_2 VNB N_A_c_38_n 0.0179813f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.83
cc_3 VNB A 0.016387f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1001_g 0.0289578f $X=-0.19 $Y=-0.24 $X2=0.455 $Y2=1.5
cc_5 VNB N_A_27_47#_c_72_n 0.004553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_73_n 0.00316029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_74_n 0.00160894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_75_n 0.0188254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_76_n 0.00216225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VPWR_c_138_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_X_c_160_n 0.0257842f $X=-0.19 $Y=-0.24 $X2=0.455 $Y2=1.62
cc_12 VNB N_X_c_161_n 0.00808244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB X 0.0145716f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=1.16
cc_14 VNB N_VGND_c_184_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.62
cc_15 VNB N_VGND_c_185_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_186_n 0.0153759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_187_n 0.10585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_188_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VPB N_A_c_37_n 0.00828629f $X=-0.19 $Y=1.305 $X2=0.44 $Y2=1.325
cc_20 VPB N_A_c_41_n 0.0136328f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.5
cc_21 VPB N_A_c_42_n 0.0273733f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.62
cc_22 VPB A 0.00599714f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_23 VPB N_A_27_47#_M1002_g 0.0288767f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_24 VPB N_A_27_47#_c_78_n 0.00437821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_A_27_47#_c_79_n 0.00777514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_27_47#_c_80_n 0.00135348f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_27_47#_c_74_n 6.84768e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_27_47#_c_75_n 0.00891828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_139_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.62
cc_30 VPB N_VPWR_c_140_n 0.0161285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_141_n 0.0152818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_138_n 0.0448622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_143_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_X_c_163_n 0.010634f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.5
cc_35 VPB N_X_c_160_n 0.0120491f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.62
cc_36 VPB X 0.0297138f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_37 N_A_c_37_n N_A_27_47#_M1001_g 0.003841f $X=0.44 $Y=1.325 $X2=0 $Y2=0
cc_38 N_A_c_38_n N_A_27_47#_M1001_g 0.0209393f $X=0.47 $Y=0.83 $X2=0 $Y2=0
cc_39 N_A_c_41_n N_A_27_47#_M1002_g 0.00368068f $X=0.455 $Y=1.5 $X2=0 $Y2=0
cc_40 N_A_c_42_n N_A_27_47#_M1002_g 0.016665f $X=0.455 $Y=1.62 $X2=0 $Y2=0
cc_41 N_A_c_37_n N_A_27_47#_c_72_n 0.00107654f $X=0.44 $Y=1.325 $X2=0 $Y2=0
cc_42 N_A_c_38_n N_A_27_47#_c_72_n 0.0150007f $X=0.47 $Y=0.83 $X2=0 $Y2=0
cc_43 A N_A_27_47#_c_72_n 0.00712115f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_44 N_A_c_37_n N_A_27_47#_c_73_n 0.00127129f $X=0.44 $Y=1.325 $X2=0 $Y2=0
cc_45 A N_A_27_47#_c_73_n 0.0143207f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_46 N_A_c_37_n N_A_27_47#_c_78_n 3.11379e-19 $X=0.44 $Y=1.325 $X2=0 $Y2=0
cc_47 N_A_c_42_n N_A_27_47#_c_78_n 0.0189812f $X=0.455 $Y=1.62 $X2=0 $Y2=0
cc_48 A N_A_27_47#_c_78_n 0.00700834f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_49 N_A_c_37_n N_A_27_47#_c_79_n 0.00130855f $X=0.44 $Y=1.325 $X2=0 $Y2=0
cc_50 A N_A_27_47#_c_79_n 0.0154136f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_51 N_A_c_42_n N_A_27_47#_c_80_n 7.5643e-19 $X=0.455 $Y=1.62 $X2=0 $Y2=0
cc_52 N_A_c_41_n N_A_27_47#_c_74_n 0.00318841f $X=0.455 $Y=1.5 $X2=0 $Y2=0
cc_53 N_A_c_37_n N_A_27_47#_c_75_n 0.0204881f $X=0.44 $Y=1.325 $X2=0 $Y2=0
cc_54 A N_A_27_47#_c_75_n 3.0111e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A_c_37_n N_A_27_47#_c_76_n 0.00318841f $X=0.44 $Y=1.325 $X2=0 $Y2=0
cc_56 N_A_c_38_n N_A_27_47#_c_76_n 0.00318324f $X=0.47 $Y=0.83 $X2=0 $Y2=0
cc_57 A N_A_27_47#_c_76_n 0.0231805f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_42_n N_VPWR_c_139_n 0.0118915f $X=0.455 $Y=1.62 $X2=0 $Y2=0
cc_59 N_A_c_42_n N_VPWR_c_140_n 0.00505556f $X=0.455 $Y=1.62 $X2=0 $Y2=0
cc_60 N_A_c_42_n N_VPWR_c_138_n 0.00946027f $X=0.455 $Y=1.62 $X2=0 $Y2=0
cc_61 N_A_c_38_n N_VGND_c_184_n 0.00787353f $X=0.47 $Y=0.83 $X2=0 $Y2=0
cc_62 N_A_c_38_n N_VGND_c_185_n 0.00367706f $X=0.47 $Y=0.83 $X2=0 $Y2=0
cc_63 N_A_c_38_n N_VGND_c_187_n 0.00526324f $X=0.47 $Y=0.83 $X2=0 $Y2=0
cc_64 N_A_27_47#_c_78_n N_VPWR_M1000_d 0.00190738f $X=0.67 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_27_47#_M1002_g N_VPWR_c_139_n 0.0118404f $X=0.91 $Y=2.09 $X2=0 $Y2=0
cc_66 N_A_27_47#_c_78_n N_VPWR_c_139_n 0.0169772f $X=0.67 $Y=1.62 $X2=0 $Y2=0
cc_67 N_A_27_47#_c_74_n N_VPWR_c_139_n 4.75835e-19 $X=0.86 $Y=1.225 $X2=0 $Y2=0
cc_68 N_A_27_47#_c_75_n N_VPWR_c_139_n 3.47424e-19 $X=0.86 $Y=1.225 $X2=0 $Y2=0
cc_69 N_A_27_47#_c_109_p N_VPWR_c_140_n 0.012308f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_70 N_A_27_47#_M1002_g N_VPWR_c_141_n 0.00505556f $X=0.91 $Y=2.09 $X2=0 $Y2=0
cc_71 N_A_27_47#_M1000_s N_VPWR_c_138_n 0.00490516f $X=0.135 $Y=1.695 $X2=0
+ $Y2=0
cc_72 N_A_27_47#_M1002_g N_VPWR_c_138_n 0.00946027f $X=0.91 $Y=2.09 $X2=0 $Y2=0
cc_73 N_A_27_47#_c_109_p N_VPWR_c_138_n 0.00685509f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_74 N_A_27_47#_M1002_g N_X_c_163_n 0.00347811f $X=0.91 $Y=2.09 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_78_n N_X_c_163_n 0.0108135f $X=0.67 $Y=1.62 $X2=0 $Y2=0
cc_76 N_A_27_47#_M1001_g N_X_c_160_n 0.00638849f $X=0.91 $Y=0.495 $X2=0 $Y2=0
cc_77 N_A_27_47#_M1002_g N_X_c_160_n 0.0036109f $X=0.91 $Y=2.09 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_72_n N_X_c_160_n 0.00248131f $X=0.67 $Y=0.72 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_78_n N_X_c_160_n 0.00136803f $X=0.67 $Y=1.62 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_80_n N_X_c_160_n 0.0072356f $X=0.755 $Y=1.535 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_74_n N_X_c_160_n 0.0245674f $X=0.86 $Y=1.225 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_75_n N_X_c_160_n 0.00754311f $X=0.86 $Y=1.225 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_76_n N_X_c_160_n 0.0127597f $X=0.807 $Y=1.06 $X2=0 $Y2=0
cc_84 N_A_27_47#_M1001_g N_X_c_161_n 0.00222896f $X=0.91 $Y=0.495 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_72_n N_X_c_161_n 0.00484499f $X=0.67 $Y=0.72 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_72_n N_VGND_M1003_d 0.00183491f $X=0.67 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_27_47#_M1001_g N_VGND_c_184_n 0.00801602f $X=0.91 $Y=0.495 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_72_n N_VGND_c_184_n 0.0159274f $X=0.67 $Y=0.72 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_74_n N_VGND_c_184_n 3.89729e-19 $X=0.86 $Y=1.225 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_75_n N_VGND_c_184_n 2.8407e-19 $X=0.86 $Y=1.225 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_131_p N_VGND_c_185_n 0.01143f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_72_n N_VGND_c_185_n 0.00260015f $X=0.67 $Y=0.72 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1001_g N_VGND_c_186_n 0.00505556f $X=0.91 $Y=0.495 $X2=0 $Y2=0
cc_94 N_A_27_47#_M1003_s N_VGND_c_187_n 0.00369894f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_M1001_g N_VGND_c_187_n 0.00957284f $X=0.91 $Y=0.495 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_131_p N_VGND_c_187_n 0.00643448f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_72_n N_VGND_c_187_n 0.00595413f $X=0.67 $Y=0.72 $X2=0 $Y2=0
cc_98 N_VPWR_c_138_n N_X_M1002_d 0.00348182f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_99 N_VPWR_c_141_n X 0.0183559f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_100 N_VPWR_c_138_n X 0.0103212f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_101 X N_VGND_c_186_n 0.0178913f $X=1.055 $Y=0.425 $X2=0 $Y2=0
cc_102 N_X_M1001_d N_VGND_c_187_n 0.00387172f $X=0.985 $Y=0.235 $X2=0 $Y2=0
cc_103 X N_VGND_c_187_n 0.00991282f $X=1.055 $Y=0.425 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__maj3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
M1000 a_441_47# B a_47_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.226e+11p ps=2.74e+06u
M1001 a_285_47# A VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=6.1335e+11p ps=5.72e+06u
M1002 a_47_47# B a_285_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_285_369# A VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=9.168e+11p ps=7.56e+06u
M1004 VPWR A a_129_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1005 a_47_47# B a_285_369# VPB phighvt w=640000u l=150000u
+  ad=3.392e+11p pd=3.62e+06u as=0p ps=0u
M1006 VPWR a_47_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 X a_47_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_129_47# C a_47_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 a_129_369# C a_47_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C a_441_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1011 VGND C a_441_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_47_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1013 VGND A a_129_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_441_369# B a_47_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_47_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


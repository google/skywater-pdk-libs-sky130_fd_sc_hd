* File: sky130_fd_sc_hd__or3b_4.spice.pex
* Created: Thu Aug 27 14:43:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR3B_4%C_N 3 7 9 10 17
c28 3 0 1.41829e-19 $X=0.47 $Y=0.445
r29 14 17 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r31 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r33 5 7 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=2.01
r34 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r35 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_4%A_176_21# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 38 46 47 48 52 56 62 65 67 69 70 78
c147 36 0 2.84877e-20 $X=2.215 $Y=1.985
r148 72 74 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.955 $Y=1.16
+ $X2=1.375 $Y2=1.16
r149 64 70 1.17118 $w=2.05e-07 $l=1.1e-07 $layer=LI1_cond $X=3.952 $Y=0.825
+ $X2=3.952 $Y2=0.715
r150 64 65 74.9313 $w=2.03e-07 $l=1.385e-06 $layer=LI1_cond $X=3.952 $Y=0.825
+ $X2=3.952 $Y2=2.21
r151 60 70 8.64332 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.787 $Y=0.715
+ $X2=3.952 $Y2=0.715
r152 60 69 7.27802 $w=2.18e-07 $l=1.27e-07 $layer=LI1_cond $X=3.787 $Y=0.715
+ $X2=3.66 $Y2=0.715
r153 60 62 6.10117 $w=2.53e-07 $l=1.35e-07 $layer=LI1_cond $X=3.787 $Y=0.605
+ $X2=3.787 $Y2=0.47
r154 56 65 6.82152 $w=2.15e-07 $l=1.49543e-07 $layer=LI1_cond $X=3.85 $Y=2.317
+ $X2=3.952 $Y2=2.21
r155 56 58 5.62821 $w=2.13e-07 $l=1.05e-07 $layer=LI1_cond $X=3.85 $Y=2.317
+ $X2=3.745 $Y2=2.317
r156 55 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=0.74
+ $X2=2.845 $Y2=0.74
r157 55 69 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.93 $Y=0.74
+ $X2=3.66 $Y2=0.74
r158 50 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.655
+ $X2=2.845 $Y2=0.74
r159 50 52 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.845 $Y=0.655
+ $X2=2.845 $Y2=0.47
r160 49 66 1.35458 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=2.4 $Y=0.74
+ $X2=2.297 $Y2=0.74
r161 48 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.74
+ $X2=2.845 $Y2=0.74
r162 48 49 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.76 $Y=0.74
+ $X2=2.4 $Y2=0.74
r163 46 66 9.83255 $w=1.89e-07 $l=1.58272e-07 $layer=LI1_cond $X=2.28 $Y=0.89
+ $X2=2.297 $Y2=0.74
r164 46 47 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.28 $Y=0.89
+ $X2=2.28 $Y2=1.075
r165 45 78 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.12 $Y=1.16
+ $X2=2.215 $Y2=1.16
r166 45 76 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=2.12 $Y=1.16
+ $X2=1.795 $Y2=1.16
r167 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.12
+ $Y=1.16 $X2=2.12 $Y2=1.16
r168 41 76 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.44 $Y=1.16
+ $X2=1.795 $Y2=1.16
r169 41 74 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.44 $Y=1.16
+ $X2=1.375 $Y2=1.16
r170 40 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.44 $Y=1.16
+ $X2=2.12 $Y2=1.16
r171 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.44
+ $Y=1.16 $X2=1.44 $Y2=1.16
r172 38 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.195 $Y=1.16
+ $X2=2.28 $Y2=1.075
r173 38 44 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.195 $Y=1.16
+ $X2=2.12 $Y2=1.16
r174 34 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.325
+ $X2=2.215 $Y2=1.16
r175 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.215 $Y=1.325
+ $X2=2.215 $Y2=1.985
r176 31 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=0.995
+ $X2=2.215 $Y2=1.16
r177 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.215 $Y=0.995
+ $X2=2.215 $Y2=0.56
r178 27 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.325
+ $X2=1.795 $Y2=1.16
r179 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.795 $Y=1.325
+ $X2=1.795 $Y2=1.985
r180 24 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=0.995
+ $X2=1.795 $Y2=1.16
r181 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.795 $Y=0.995
+ $X2=1.795 $Y2=0.56
r182 20 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.16
r183 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.985
r184 17 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=1.16
r185 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=0.56
r186 13 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.16
r187 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.985
r188 10 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.16
r189 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r190 3 58 600 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=1.485 $X2=3.745 $Y2=2.295
r191 2 62 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=3.61
+ $Y=0.235 $X2=3.745 $Y2=0.47
r192 1 52 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.235 $X2=2.845 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_4%A 1 3 6 8 10 11 13
r47 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.635
+ $Y=1.16 $X2=2.635 $Y2=1.16
r48 8 13 3.72017 $w=2.83e-07 $l=9.2e-08 $layer=LI1_cond $X=2.627 $Y=1.557
+ $X2=2.535 $Y2=1.557
r49 8 10 15.2875 $w=1.83e-07 $l=2.55e-07 $layer=LI1_cond $X=2.627 $Y=1.415
+ $X2=2.627 $Y2=1.16
r50 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.325
+ $X2=2.635 $Y2=1.16
r51 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.635 $Y=1.325
+ $X2=2.635 $Y2=1.985
r52 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=0.995
+ $X2=2.635 $Y2=1.16
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.635 $Y=0.995
+ $X2=2.635 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_4%B 3 6 8 9 13 14 15
c41 14 0 2.84877e-20 $X=3.115 $Y=1.16
r42 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.16
+ $X2=3.115 $Y2=1.325
r43 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.16
+ $X2=3.115 $Y2=0.995
r44 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.115
+ $Y=1.16 $X2=3.115 $Y2=1.16
r45 8 9 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=3.045 $Y=1.19
+ $X2=3.045 $Y2=1.53
r46 8 14 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=3.045 $Y=1.19 $X2=3.045
+ $Y2=1.16
r47 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.055 $Y=1.985
+ $X2=3.055 $Y2=1.325
r48 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.055 $Y=0.56
+ $X2=3.055 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_4%A_27_47# 1 2 9 12 16 18 19 20 23 24 27 30 32
+ 34 35 39
r98 35 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.16
+ $X2=3.595 $Y2=1.325
r99 35 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.16
+ $X2=3.595 $Y2=0.995
r100 34 37 7.0829 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=1.16
+ $X2=3.535 $Y2=1.325
r101 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.595
+ $Y=1.16 $X2=3.595 $Y2=1.16
r102 27 37 27.3079 $w=2.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.505 $Y=1.87
+ $X2=3.505 $Y2=1.325
r103 25 32 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.765 $Y=1.955
+ $X2=0.68 $Y2=1.925
r104 24 27 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.39 $Y=1.955
+ $X2=3.505 $Y2=1.87
r105 24 25 171.257 $w=1.68e-07 $l=2.625e-06 $layer=LI1_cond $X=3.39 $Y=1.955
+ $X2=0.765 $Y2=1.955
r106 23 32 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.68 $Y=1.81
+ $X2=0.68 $Y2=1.925
r107 22 23 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=0.68 $Y=0.905
+ $X2=0.68 $Y2=1.81
r108 21 30 1.45362 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.925
+ $X2=0.215 $Y2=1.925
r109 20 32 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=1.925
+ $X2=0.68 $Y2=1.925
r110 20 21 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.595 $Y=1.925
+ $X2=0.345 $Y2=1.925
r111 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.68 $Y2=0.905
r112 18 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.345 $Y2=0.82
r113 14 19 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.345 $Y2=0.82
r114 14 16 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.215 $Y2=0.455
r115 12 40 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.535 $Y=1.985
+ $X2=3.535 $Y2=1.325
r116 9 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.535 $Y=0.56
+ $X2=3.535 $Y2=0.995
r117 2 30 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.8 $X2=0.26 $Y2=1.975
r118 1 16 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_4%VPWR 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r66 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r67 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 42 52 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 39 51 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.595 $Y=2.72
+ $X2=2.425 $Y2=2.72
r72 39 41 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=2.595 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r74 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r75 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r76 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=2.72
+ $X2=1.585 $Y2=2.72
r77 35 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.75 $Y=2.72 $X2=2.07
+ $Y2=2.72
r78 34 51 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.425 $Y2=2.72
r79 34 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 30 45 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.91 $Y=2.72 $X2=0.73
+ $Y2=2.72
r84 30 32 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=2.72
+ $X2=1.585 $Y2=2.72
r86 29 32 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.42 $Y=2.72 $X2=1.15
+ $Y2=2.72
r87 24 45 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=0.73
+ $Y2=2.72
r88 24 26 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=0.23
+ $Y2=2.72
r89 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 18 51 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=2.635
+ $X2=2.425 $Y2=2.72
r92 18 20 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.425 $Y=2.635
+ $X2=2.425 $Y2=2.295
r93 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=2.635
+ $X2=1.585 $Y2=2.72
r94 14 16 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.585 $Y=2.635
+ $X2=1.585 $Y2=2.295
r95 10 45 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r96 10 12 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.295
r97 3 20 600 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.485 $X2=2.425 $Y2=2.295
r98 2 16 600 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.485 $X2=1.585 $Y2=2.295
r99 1 12 600 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.8 $X2=0.745 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_4%X 1 2 3 4 14 17 19 22 23 24 26 29
c66 23 0 1.41829e-19 $X=1.132 $Y=0.82
r67 29 32 33.9667 $w=2.83e-07 $l=8.4e-07 $layer=LI1_cond $X=2.005 $Y=1.557
+ $X2=1.165 $Y2=1.557
r68 26 28 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.972 $Y=0.42
+ $X2=1.972 $Y2=0.585
r69 24 32 2.4262 $w=2.83e-07 $l=6e-08 $layer=LI1_cond $X=1.105 $Y=1.557
+ $X2=1.165 $Y2=1.557
r70 22 28 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=1.94 $Y2=0.585
r71 20 23 2.76166 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.33 $Y=0.82
+ $X2=1.132 $Y2=0.82
r72 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.855 $Y=0.82
+ $X2=1.94 $Y2=0.735
r73 19 20 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.855 $Y=0.82
+ $X2=1.33 $Y2=0.82
r74 15 23 3.70735 $w=2.5e-07 $l=1.0015e-07 $layer=LI1_cond $X=1.165 $Y=0.735
+ $X2=1.132 $Y2=0.82
r75 15 17 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=0.735
+ $X2=1.165 $Y2=0.395
r76 14 24 7.39867 $w=2.85e-07 $l=1.79538e-07 $layer=LI1_cond $X=1.02 $Y=1.415
+ $X2=1.105 $Y2=1.557
r77 13 23 3.70735 $w=2.5e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.02 $Y=0.905
+ $X2=1.132 $Y2=0.82
r78 13 14 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.02 $Y=0.905
+ $X2=1.02 $Y2=1.415
r79 4 29 600 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.485 $X2=2.005 $Y2=1.615
r80 3 32 600 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.615
r81 2 26 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.87
+ $Y=0.235 $X2=2.005 $Y2=0.42
r82 1 17 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.235 $X2=1.165 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_4%VGND 1 2 3 4 17 21 25 29 32 33 35 36 38 39 40
+ 53 54 57 60
r82 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r83 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r84 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r85 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r86 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r87 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r88 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r89 45 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r90 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r91 42 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.705
+ $Y2=0
r92 42 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=1.15
+ $Y2=0
r93 40 58 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r94 40 60 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r95 38 50 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.99
+ $Y2=0
r96 38 39 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.295
+ $Y2=0
r97 37 53 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.49 $Y=0 $X2=3.91
+ $Y2=0
r98 37 39 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.49 $Y=0 $X2=3.295
+ $Y2=0
r99 35 47 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.07
+ $Y2=0
r100 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.425
+ $Y2=0
r101 34 50 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.99
+ $Y2=0
r102 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.425
+ $Y2=0
r103 32 44 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.5 $Y=0 $X2=1.15
+ $Y2=0
r104 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=0 $X2=1.585
+ $Y2=0
r105 31 47 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=2.07
+ $Y2=0
r106 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.585
+ $Y2=0
r107 27 39 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0
r108 27 29 9.30819 $w=3.88e-07 $l=3.15e-07 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0.4
r109 23 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0
r110 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0.4
r111 19 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.585 $Y2=0
r112 19 21 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.585 $Y=0.085
+ $X2=1.585 $Y2=0.4
r113 15 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r114 15 17 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.4
r115 4 29 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.265 $Y2=0.4
r116 3 25 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.235 $X2=2.425 $Y2=0.4
r117 2 21 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.585 $Y2=0.4
r118 1 17 182 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.705 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__and4b_1.spice.SKY130_FD_SC_HD__AND4B_1.pxi
* Created: Thu Aug 27 14:08:41 2020
* 
x_PM_SKY130_FD_SC_HD__AND4B_1%A_N N_A_N_M1008_g N_A_N_M1005_g A_N A_N
+ N_A_N_c_80_n PM_SKY130_FD_SC_HD__AND4B_1%A_N
x_PM_SKY130_FD_SC_HD__AND4B_1%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1005_s
+ N_A_27_47#_c_111_n N_A_27_47#_M1010_g N_A_27_47#_c_112_n N_A_27_47#_c_113_n
+ N_A_27_47#_M1003_g N_A_27_47#_c_178_p N_A_27_47#_c_120_n N_A_27_47#_c_114_n
+ N_A_27_47#_c_115_n N_A_27_47#_c_121_n N_A_27_47#_c_122_n N_A_27_47#_c_116_n
+ N_A_27_47#_c_123_n N_A_27_47#_c_117_n PM_SKY130_FD_SC_HD__AND4B_1%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4B_1%B N_B_M1006_g N_B_M1004_g B B B B N_B_c_190_n
+ PM_SKY130_FD_SC_HD__AND4B_1%B
x_PM_SKY130_FD_SC_HD__AND4B_1%C N_C_M1002_g N_C_M1001_g C C C C N_C_c_228_n
+ PM_SKY130_FD_SC_HD__AND4B_1%C
x_PM_SKY130_FD_SC_HD__AND4B_1%D N_D_M1009_g N_D_M1011_g D D D N_D_c_266_n
+ PM_SKY130_FD_SC_HD__AND4B_1%D
x_PM_SKY130_FD_SC_HD__AND4B_1%A_193_413# N_A_193_413#_M1003_s
+ N_A_193_413#_M1010_d N_A_193_413#_M1001_d N_A_193_413#_M1007_g
+ N_A_193_413#_M1000_g N_A_193_413#_c_306_n N_A_193_413#_c_312_n
+ N_A_193_413#_c_313_n N_A_193_413#_c_314_n N_A_193_413#_c_315_n
+ N_A_193_413#_c_316_n N_A_193_413#_c_322_n N_A_193_413#_c_317_n
+ N_A_193_413#_c_318_n N_A_193_413#_c_307_n N_A_193_413#_c_308_n
+ N_A_193_413#_c_309_n PM_SKY130_FD_SC_HD__AND4B_1%A_193_413#
x_PM_SKY130_FD_SC_HD__AND4B_1%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_M1011_d
+ N_VPWR_c_400_n N_VPWR_c_401_n VPWR N_VPWR_c_402_n N_VPWR_c_403_n
+ N_VPWR_c_404_n N_VPWR_c_399_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n
+ N_VPWR_c_409_n PM_SKY130_FD_SC_HD__AND4B_1%VPWR
x_PM_SKY130_FD_SC_HD__AND4B_1%X N_X_M1007_d N_X_M1000_d N_X_c_459_n N_X_c_461_n
+ N_X_c_460_n X X X N_X_c_463_n PM_SKY130_FD_SC_HD__AND4B_1%X
x_PM_SKY130_FD_SC_HD__AND4B_1%VGND N_VGND_M1008_d N_VGND_M1009_d N_VGND_c_479_n
+ N_VGND_c_480_n VGND N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n
+ N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n PM_SKY130_FD_SC_HD__AND4B_1%VGND
cc_1 VNB N_A_N_M1008_g 0.0403072f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.0172275f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A_N_c_80_n 0.036838f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_47#_c_111_n 0.0433735f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_5 VNB N_A_27_47#_c_112_n 0.0358152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_113_n 0.0169127f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_7 VNB N_A_27_47#_c_114_n 0.00644367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_115_n 0.00818302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_116_n 0.00317446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_117_n 0.00221925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_M1004_g 0.0361509f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_12 VNB B 0.00330189f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_13 VNB N_B_c_190_n 0.0223034f $X=-0.19 $Y=-0.24 $X2=0.267 $Y2=1.53
cc_14 VNB N_C_M1002_g 0.0284736f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_15 VNB C 0.00432191f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_C_c_228_n 0.0208562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_M1009_g 0.0264844f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB D 0.00964293f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_D_c_266_n 0.0205332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_193_413#_c_306_n 0.00814249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_193_413#_c_307_n 0.00247125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_193_413#_c_308_n 0.0238065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_193_413#_c_309_n 0.020172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_399_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_459_n 0.020416f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_26 VNB N_X_c_460_n 0.0224947f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_27 VNB N_VGND_c_479_n 0.00557802f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_28 VNB N_VGND_c_480_n 0.00276554f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_29 VNB N_VGND_c_481_n 0.0151229f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_30 VNB N_VGND_c_482_n 0.052683f $X=-0.19 $Y=-0.24 $X2=0.267 $Y2=1.53
cc_31 VNB N_VGND_c_483_n 0.018123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_484_n 0.206027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_485_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_486_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_A_N_M1005_g 0.0614435f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_36 VPB A_N 0.0203025f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_37 VPB N_A_N_c_80_n 0.0101167f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_38 VPB N_A_27_47#_c_111_n 0.00669282f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_39 VPB N_A_27_47#_M1010_g 0.0550489f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_40 VPB N_A_27_47#_c_120_n 0.00220604f $X=-0.19 $Y=1.305 $X2=0.267 $Y2=1.53
cc_41 VPB N_A_27_47#_c_121_n 0.00786997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_122_n 0.00841734f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_123_n 0.00931061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_117_n 4.82126e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B_M1006_g 0.0545611f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_46 VPB B 0.00435974f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_47 VPB N_B_c_190_n 0.0165518f $X=-0.19 $Y=1.305 $X2=0.267 $Y2=1.53
cc_48 VPB N_C_M1001_g 0.05509f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_49 VPB C 0.00450837f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_50 VPB N_C_c_228_n 0.00453948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_D_M1011_g 0.0471738f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_52 VPB D 0.00663196f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_53 VPB N_D_c_266_n 0.00449071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_193_413#_M1000_g 0.0217459f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_55 VPB N_A_193_413#_c_306_n 0.0114802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_193_413#_c_312_n 4.33886e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_193_413#_c_313_n 0.0263913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_193_413#_c_314_n 3.38187e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_193_413#_c_315_n 0.00385753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_193_413#_c_316_n 0.00107927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_193_413#_c_317_n 0.00210916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_193_413#_c_318_n 0.00286967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_193_413#_c_307_n 2.26104e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_193_413#_c_308_n 0.00510782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_400_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_401_n 0.00231197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_402_n 0.0151914f $X=-0.19 $Y=1.305 $X2=0.267 $Y2=1.53
cc_68 VPB N_VPWR_c_403_n 0.014199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_404_n 0.0157545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_399_n 0.0453489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_406_n 0.00436502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_407_n 0.0178771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_408_n 0.0121841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_409_n 0.00522141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_X_c_461_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_76 VPB N_X_c_460_n 0.00876896f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_77 VPB N_X_c_463_n 0.0322452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 N_A_N_M1008_g N_A_27_47#_c_111_n 0.00821899f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_79 A_N N_A_27_47#_c_111_n 2.78759e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A_N_c_80_n N_A_27_47#_c_111_n 0.0202235f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_N_M1005_g N_A_27_47#_M1010_g 0.0381875f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_82 N_A_N_M1005_g N_A_27_47#_c_120_n 0.00268857f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_83 N_A_N_M1008_g N_A_27_47#_c_114_n 0.0161999f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_84 A_N N_A_27_47#_c_114_n 0.00807147f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_85 N_A_N_c_80_n N_A_27_47#_c_114_n 3.50292e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_86 A_N N_A_27_47#_c_115_n 0.0153899f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_N_c_80_n N_A_27_47#_c_115_n 0.00135787f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_N_M1005_g N_A_27_47#_c_121_n 0.0154869f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_89 A_N N_A_27_47#_c_121_n 0.00829866f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_90 A_N N_A_27_47#_c_122_n 0.0162852f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_91 N_A_N_c_80_n N_A_27_47#_c_122_n 6.55167e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_N_M1008_g N_A_27_47#_c_116_n 0.0039865f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_N_M1005_g N_A_27_47#_c_123_n 0.00616503f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_94 A_N N_A_27_47#_c_123_n 0.0253512f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_95 A_N N_A_27_47#_c_117_n 0.0252802f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_N_c_80_n N_A_27_47#_c_117_n 0.00237414f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_N_M1008_g N_A_193_413#_c_306_n 0.00189977f $X=0.47 $Y=0.445 $X2=0
+ $Y2=0
cc_98 N_A_N_M1008_g N_A_193_413#_c_322_n 0.00162248f $X=0.47 $Y=0.445 $X2=0
+ $Y2=0
cc_99 N_A_N_M1005_g N_VPWR_c_400_n 0.00898724f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_100 N_A_N_M1005_g N_VPWR_c_402_n 0.00347311f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_101 N_A_N_M1005_g N_VPWR_c_399_n 0.00503562f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_102 N_A_N_M1008_g N_VGND_c_479_n 0.00947303f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A_N_M1008_g N_VGND_c_481_n 0.00341689f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_N_M1008_g N_VGND_c_484_n 0.00493711f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_111_n N_B_M1004_g 0.00259332f $X=0.89 $Y=1.325 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_113_n N_B_M1004_g 0.0481451f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_113_n B 0.00259364f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_111_n N_B_c_190_n 0.00439184f $X=0.89 $Y=1.325 $X2=0 $Y2=0
cc_109 N_A_27_47#_M1010_g N_B_c_190_n 0.023308f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_112_n N_B_c_190_n 0.00350435f $X=1.335 $Y=0.805 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_111_n N_A_193_413#_c_306_n 0.00454513f $X=0.89 $Y=1.325
+ $X2=0 $Y2=0
cc_112 N_A_27_47#_M1010_g N_A_193_413#_c_306_n 0.00502314f $X=0.89 $Y=2.275
+ $X2=0 $Y2=0
cc_113 N_A_27_47#_c_112_n N_A_193_413#_c_306_n 0.0138926f $X=1.335 $Y=0.805
+ $X2=0 $Y2=0
cc_114 N_A_27_47#_c_113_n N_A_193_413#_c_306_n 0.00254183f $X=1.41 $Y=0.73 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_114_n N_A_193_413#_c_306_n 0.00826266f $X=0.63 $Y=0.74 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_121_n N_A_193_413#_c_306_n 0.00149659f $X=0.63 $Y=1.93 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_116_n N_A_193_413#_c_306_n 0.00750984f $X=0.715 $Y=0.995
+ $X2=0 $Y2=0
cc_118 N_A_27_47#_c_123_n N_A_193_413#_c_306_n 0.0236604f $X=0.715 $Y=1.845
+ $X2=0 $Y2=0
cc_119 N_A_27_47#_c_117_n N_A_193_413#_c_306_n 0.0248826f $X=0.895 $Y=1.16 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_M1010_g N_A_193_413#_c_312_n 0.00564962f $X=0.89 $Y=2.275
+ $X2=0 $Y2=0
cc_121 N_A_27_47#_c_112_n N_A_193_413#_c_322_n 0.00225284f $X=1.335 $Y=0.805
+ $X2=0 $Y2=0
cc_122 N_A_27_47#_M1010_g N_A_193_413#_c_317_n 0.0023712f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_121_n N_A_193_413#_c_317_n 0.00785419f $X=0.63 $Y=1.93 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_M1010_g N_VPWR_c_400_n 0.0104697f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_121_n N_VPWR_c_400_n 0.0183339f $X=0.63 $Y=1.93 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_120_n N_VPWR_c_402_n 0.0118773f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_121_n N_VPWR_c_402_n 0.002454f $X=0.63 $Y=1.93 $X2=0 $Y2=0
cc_128 N_A_27_47#_M1005_s N_VPWR_c_399_n 0.00356395f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_M1010_g N_VPWR_c_399_n 0.0084266f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_120_n N_VPWR_c_399_n 0.00664644f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_121_n N_VPWR_c_399_n 0.00517911f $X=0.63 $Y=1.93 $X2=0 $Y2=0
cc_132 N_A_27_47#_M1010_g N_VPWR_c_407_n 0.0046653f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_133 N_A_27_47#_M1010_g N_VPWR_c_408_n 9.75794e-19 $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_114_n N_VGND_M1008_d 0.00183923f $X=0.63 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_27_47#_c_111_n N_VGND_c_479_n 0.00103651f $X=0.89 $Y=1.325 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_c_113_n N_VGND_c_479_n 0.00276694f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_114_n N_VGND_c_479_n 0.0179795f $X=0.63 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_117_n N_VGND_c_479_n 0.00157757f $X=0.895 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_c_178_p N_VGND_c_481_n 0.0118061f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_114_n N_VGND_c_481_n 0.00273399f $X=0.63 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_111_n N_VGND_c_482_n 0.00419046f $X=0.89 $Y=1.325 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_c_112_n N_VGND_c_482_n 6.44498e-19 $X=1.335 $Y=0.805 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_c_113_n N_VGND_c_482_n 0.00585385f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_144 N_A_27_47#_M1008_s N_VGND_c_484_n 0.00352789f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_111_n N_VGND_c_484_n 0.00578911f $X=0.89 $Y=1.325 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_113_n N_VGND_c_484_n 0.0119273f $X=1.41 $Y=0.73 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_178_p N_VGND_c_484_n 0.00663203f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_114_n N_VGND_c_484_n 0.00544343f $X=0.63 $Y=0.74 $X2=0 $Y2=0
cc_149 N_B_M1004_g N_C_M1002_g 0.029948f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_150 B N_C_M1002_g 5.45207e-19 $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_151 N_B_M1006_g N_C_M1001_g 0.0139464f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_152 B N_C_M1001_g 9.46813e-19 $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_153 N_B_c_190_n N_C_M1001_g 0.00254887f $X=1.77 $Y=1.27 $X2=0 $Y2=0
cc_154 N_B_M1006_g C 7.90751e-19 $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_155 N_B_M1004_g C 0.00677686f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_156 B C 0.0804026f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_157 N_B_M1004_g N_C_c_228_n 0.0181019f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_158 B N_C_c_228_n 3.5867e-19 $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_159 N_B_M1004_g N_A_193_413#_c_306_n 8.15967e-19 $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_160 B N_A_193_413#_c_306_n 0.0696125f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_161 N_B_c_190_n N_A_193_413#_c_306_n 0.00941695f $X=1.77 $Y=1.27 $X2=0 $Y2=0
cc_162 N_B_M1006_g N_A_193_413#_c_312_n 0.00653277f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_163 N_B_M1006_g N_A_193_413#_c_313_n 0.0159719f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_164 B N_A_193_413#_c_313_n 0.0220118f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_165 N_B_c_190_n N_A_193_413#_c_313_n 0.00218571f $X=1.77 $Y=1.27 $X2=0 $Y2=0
cc_166 N_B_M1006_g N_VPWR_c_400_n 9.59561e-19 $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_167 N_B_M1006_g N_VPWR_c_399_n 0.00450838f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_168 N_B_M1006_g N_VPWR_c_407_n 0.00343969f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_169 N_B_M1006_g N_VPWR_c_408_n 0.00975543f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_170 N_B_M1004_g N_VGND_c_482_n 0.00449772f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_171 B N_VGND_c_482_n 0.00798731f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_172 N_B_M1004_g N_VGND_c_484_n 0.00715864f $X=1.77 $Y=0.445 $X2=0 $Y2=0
cc_173 B N_VGND_c_484_n 0.00921996f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_174 B A_297_47# 0.00129203f $X=1.525 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_175 N_C_M1002_g N_D_M1009_g 0.0374912f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_176 C N_D_M1009_g 0.00158447f $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_177 N_C_M1001_g N_D_M1011_g 0.0343885f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_178 C N_D_M1011_g 3.3807e-19 $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_179 N_C_M1002_g D 0.00680155f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_180 C D 0.0740266f $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_181 C N_D_c_266_n 3.35477e-19 $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_182 N_C_c_228_n N_D_c_266_n 0.0202262f $X=2.21 $Y=1.16 $X2=0 $Y2=0
cc_183 N_C_M1001_g N_A_193_413#_c_313_n 0.0147503f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_184 C N_A_193_413#_c_313_n 0.0209083f $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_185 N_C_c_228_n N_A_193_413#_c_313_n 3.89084e-19 $X=2.21 $Y=1.16 $X2=0 $Y2=0
cc_186 N_C_M1001_g N_A_193_413#_c_314_n 0.00439741f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_187 N_C_M1001_g N_VPWR_c_403_n 0.00343969f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_188 N_C_M1001_g N_VPWR_c_399_n 0.0041399f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_189 N_C_M1001_g N_VPWR_c_408_n 0.00847709f $X=2.27 $Y=2.275 $X2=0 $Y2=0
cc_190 N_C_M1002_g N_VGND_c_480_n 0.00204992f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_191 C N_VGND_c_480_n 0.00148293f $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_192 N_C_M1002_g N_VGND_c_482_n 0.00456292f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_193 C N_VGND_c_482_n 0.0079878f $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_194 N_C_M1002_g N_VGND_c_484_n 0.0075516f $X=2.27 $Y=0.445 $X2=0 $Y2=0
cc_195 C N_VGND_c_484_n 0.00889453f $X=2.03 $Y=0.425 $X2=0 $Y2=0
cc_196 C A_369_47# 0.00374224f $X=2.03 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_197 N_D_M1011_g N_A_193_413#_M1000_g 0.033628f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_198 D N_A_193_413#_M1000_g 9.78277e-19 $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_199 N_D_M1011_g N_A_193_413#_c_314_n 6.38571e-19 $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_200 N_D_M1011_g N_A_193_413#_c_315_n 0.0124544f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_201 D N_A_193_413#_c_315_n 0.0160658f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_202 N_D_c_266_n N_A_193_413#_c_315_n 2.05349e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_203 N_D_M1011_g N_A_193_413#_c_316_n 0.00489639f $X=2.735 $Y=2.275 $X2=0
+ $Y2=0
cc_204 D N_A_193_413#_c_316_n 0.0291205f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_205 D N_A_193_413#_c_318_n 0.0110373f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_206 D N_A_193_413#_c_307_n 0.0256593f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_207 N_D_c_266_n N_A_193_413#_c_307_n 0.00175898f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_208 D N_A_193_413#_c_308_n 3.78352e-19 $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_209 N_D_c_266_n N_A_193_413#_c_308_n 0.0203238f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_210 N_D_M1009_g N_A_193_413#_c_309_n 0.0233641f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_211 D N_A_193_413#_c_309_n 0.0027953f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_212 N_D_M1011_g N_VPWR_c_401_n 0.00172637f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_213 N_D_M1011_g N_VPWR_c_403_n 0.00430148f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_214 N_D_M1011_g N_VPWR_c_399_n 0.00592266f $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_215 N_D_M1011_g N_VPWR_c_408_n 5.46734e-19 $X=2.735 $Y=2.275 $X2=0 $Y2=0
cc_216 N_D_M1009_g N_X_c_459_n 8.37986e-19 $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_217 D N_X_c_459_n 0.00558165f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_218 D N_X_c_460_n 0.00615197f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_219 N_D_M1009_g N_VGND_c_480_n 0.00959191f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_220 D N_VGND_c_480_n 0.00336096f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_221 N_D_M1009_g N_VGND_c_482_n 0.0034272f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_222 D N_VGND_c_482_n 0.00485239f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_223 N_D_M1009_g N_VGND_c_484_n 0.00412264f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_224 D N_VGND_c_484_n 0.00767675f $X=2.5 $Y=0.765 $X2=0 $Y2=0
cc_225 N_A_193_413#_c_315_n N_VPWR_M1011_d 0.00620895f $X=2.995 $Y=1.96 $X2=0
+ $Y2=0
cc_226 N_A_193_413#_c_316_n N_VPWR_M1011_d 0.00386409f $X=3.08 $Y=1.875 $X2=0
+ $Y2=0
cc_227 N_A_193_413#_c_312_n N_VPWR_c_400_n 0.0127254f $X=1.235 $Y=2.3 $X2=0
+ $Y2=0
cc_228 N_A_193_413#_M1000_g N_VPWR_c_401_n 0.00722566f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_193_413#_c_315_n N_VPWR_c_401_n 0.0182012f $X=2.995 $Y=1.96 $X2=0
+ $Y2=0
cc_230 N_A_193_413#_c_313_n N_VPWR_c_403_n 0.00337363f $X=2.44 $Y=1.96 $X2=0
+ $Y2=0
cc_231 N_A_193_413#_c_314_n N_VPWR_c_403_n 0.0114872f $X=2.525 $Y=2.3 $X2=0
+ $Y2=0
cc_232 N_A_193_413#_c_315_n N_VPWR_c_403_n 0.00306482f $X=2.995 $Y=1.96 $X2=0
+ $Y2=0
cc_233 N_A_193_413#_M1000_g N_VPWR_c_404_n 0.00539353f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_193_413#_c_315_n N_VPWR_c_404_n 3.95781e-19 $X=2.995 $Y=1.96 $X2=0
+ $Y2=0
cc_235 N_A_193_413#_M1010_d N_VPWR_c_399_n 0.0107282f $X=0.965 $Y=2.065 $X2=0
+ $Y2=0
cc_236 N_A_193_413#_M1001_d N_VPWR_c_399_n 0.0031023f $X=2.345 $Y=2.065 $X2=0
+ $Y2=0
cc_237 N_A_193_413#_M1000_g N_VPWR_c_399_n 0.0096554f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_193_413#_c_312_n N_VPWR_c_399_n 0.00646998f $X=1.235 $Y=2.3 $X2=0
+ $Y2=0
cc_239 N_A_193_413#_c_313_n N_VPWR_c_399_n 0.0139338f $X=2.44 $Y=1.96 $X2=0
+ $Y2=0
cc_240 N_A_193_413#_c_314_n N_VPWR_c_399_n 0.00644606f $X=2.525 $Y=2.3 $X2=0
+ $Y2=0
cc_241 N_A_193_413#_c_315_n N_VPWR_c_399_n 0.00680748f $X=2.995 $Y=1.96 $X2=0
+ $Y2=0
cc_242 N_A_193_413#_c_312_n N_VPWR_c_407_n 0.0118139f $X=1.235 $Y=2.3 $X2=0
+ $Y2=0
cc_243 N_A_193_413#_c_313_n N_VPWR_c_407_n 0.00371004f $X=2.44 $Y=1.96 $X2=0
+ $Y2=0
cc_244 N_A_193_413#_c_312_n N_VPWR_c_408_n 0.0145995f $X=1.235 $Y=2.3 $X2=0
+ $Y2=0
cc_245 N_A_193_413#_c_313_n N_VPWR_c_408_n 0.0445621f $X=2.44 $Y=1.96 $X2=0
+ $Y2=0
cc_246 N_A_193_413#_c_314_n N_VPWR_c_408_n 0.0156363f $X=2.525 $Y=2.3 $X2=0
+ $Y2=0
cc_247 N_A_193_413#_c_309_n N_X_c_459_n 0.0098106f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_193_413#_M1000_g N_X_c_460_n 0.00335436f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_193_413#_c_316_n N_X_c_460_n 0.00879353f $X=3.08 $Y=1.875 $X2=0 $Y2=0
cc_250 N_A_193_413#_c_307_n N_X_c_460_n 0.0243303f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_193_413#_c_308_n N_X_c_460_n 0.00753767f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A_193_413#_c_309_n N_X_c_460_n 0.00320939f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_193_413#_c_322_n N_VGND_c_479_n 0.0128716f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_254 N_A_193_413#_c_307_n N_VGND_c_480_n 0.00303163f $X=3.17 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A_193_413#_c_308_n N_VGND_c_480_n 8.59493e-19 $X=3.17 $Y=1.16 $X2=0
+ $Y2=0
cc_256 N_A_193_413#_c_309_n N_VGND_c_480_n 0.00417809f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A_193_413#_c_322_n N_VGND_c_482_n 0.0143957f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_258 N_A_193_413#_c_309_n N_VGND_c_483_n 0.00541489f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_193_413#_M1003_s N_VGND_c_484_n 0.00244967f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_260 N_A_193_413#_c_322_n N_VGND_c_484_n 0.00874023f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_261 N_A_193_413#_c_309_n N_VGND_c_484_n 0.0107167f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_399_n N_X_M1000_d 0.00387172f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_263 N_VPWR_c_404_n N_X_c_463_n 0.018001f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_264 N_VPWR_c_399_n N_X_c_463_n 0.00993603f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_265 N_X_c_459_n N_VGND_c_483_n 0.0172615f $X=3.51 $Y=0.805 $X2=0 $Y2=0
cc_266 N_X_M1007_d N_VGND_c_484_n 0.00211564f $X=3.285 $Y=0.235 $X2=0 $Y2=0
cc_267 N_X_c_459_n N_VGND_c_484_n 0.012566f $X=3.51 $Y=0.805 $X2=0 $Y2=0
cc_268 N_VGND_c_484_n A_297_47# 0.00309773f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_269 N_VGND_c_484_n A_369_47# 0.00925104f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_270 N_VGND_c_484_n A_469_47# 0.00782994f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o221ai_1.pxi.spice
* Created: Thu Aug 27 14:37:09 2020
* 
x_PM_SKY130_FD_SC_HD__O221AI_1%C1 N_C1_c_55_n N_C1_M1008_g N_C1_c_56_n
+ N_C1_M1002_g C1 N_C1_c_57_n PM_SKY130_FD_SC_HD__O221AI_1%C1
x_PM_SKY130_FD_SC_HD__O221AI_1%B1 N_B1_M1006_g N_B1_M1003_g B1 N_B1_c_80_n
+ N_B1_c_81_n N_B1_c_82_n PM_SKY130_FD_SC_HD__O221AI_1%B1
x_PM_SKY130_FD_SC_HD__O221AI_1%B2 N_B2_M1005_g N_B2_M1000_g B2 N_B2_c_111_n
+ N_B2_c_112_n PM_SKY130_FD_SC_HD__O221AI_1%B2
x_PM_SKY130_FD_SC_HD__O221AI_1%A2 N_A2_c_147_n N_A2_M1001_g N_A2_M1007_g
+ N_A2_c_148_n N_A2_c_149_n N_A2_c_150_n N_A2_c_154_n A2
+ PM_SKY130_FD_SC_HD__O221AI_1%A2
x_PM_SKY130_FD_SC_HD__O221AI_1%A1 N_A1_c_193_n N_A1_M1004_g N_A1_M1009_g A1
+ N_A1_c_195_n PM_SKY130_FD_SC_HD__O221AI_1%A1
x_PM_SKY130_FD_SC_HD__O221AI_1%Y N_Y_M1008_s N_Y_M1002_s N_Y_M1005_d N_Y_c_219_n
+ N_Y_c_223_n N_Y_c_224_n N_Y_c_220_n N_Y_c_221_n N_Y_c_232_n N_Y_c_222_n
+ N_Y_c_241_n N_Y_c_256_p Y Y PM_SKY130_FD_SC_HD__O221AI_1%Y
x_PM_SKY130_FD_SC_HD__O221AI_1%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_c_280_n
+ N_VPWR_c_281_n VPWR N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n
+ N_VPWR_c_279_n PM_SKY130_FD_SC_HD__O221AI_1%VPWR
x_PM_SKY130_FD_SC_HD__O221AI_1%A_109_47# N_A_109_47#_M1008_d N_A_109_47#_M1006_d
+ N_A_109_47#_c_326_n PM_SKY130_FD_SC_HD__O221AI_1%A_109_47#
x_PM_SKY130_FD_SC_HD__O221AI_1%A_213_123# N_A_213_123#_M1006_s
+ N_A_213_123#_M1000_d N_A_213_123#_M1004_d N_A_213_123#_c_340_n
+ N_A_213_123#_c_341_n N_A_213_123#_c_342_n N_A_213_123#_c_349_n
+ PM_SKY130_FD_SC_HD__O221AI_1%A_213_123#
x_PM_SKY130_FD_SC_HD__O221AI_1%VGND N_VGND_M1001_d N_VGND_c_383_n VGND
+ N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n
+ PM_SKY130_FD_SC_HD__O221AI_1%VGND
cc_1 VNB N_C1_c_55_n 0.0251668f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_C1_c_56_n 0.0319478f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_3 VNB N_C1_c_57_n 0.013208f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_4 VNB N_B1_c_80_n 0.0279788f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_5 VNB N_B1_c_81_n 0.00334141f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_6 VNB N_B1_c_82_n 0.0201382f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_7 VNB B2 0.0059886f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB N_B2_c_111_n 0.0185644f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_9 VNB N_B2_c_112_n 0.0172889f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_10 VNB N_A2_c_147_n 0.0172889f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_11 VNB N_A2_c_148_n 5.9128e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_149_n 0.00330957f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_13 VNB N_A2_c_150_n 0.0195476f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_14 VNB N_A1_c_193_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_15 VNB A1 0.00957755f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_A1_c_195_n 0.0358799f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_17 VNB N_Y_c_219_n 0.011033f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_18 VNB N_Y_c_220_n 0.00197206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_221_n 0.00810425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_222_n 0.00977255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_279_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_109_47#_c_326_n 0.0105337f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_23 VNB N_A_213_123#_c_340_n 0.00258612f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_24 VNB N_A_213_123#_c_341_n 0.00767792f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.16
cc_25 VNB N_A_213_123#_c_342_n 0.016608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_383_n 0.0046757f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_27 VNB N_VGND_c_384_n 0.0626928f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_28 VNB N_VGND_c_385_n 0.0173701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_386_n 0.182957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_387_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_C1_c_56_n 0.00589404f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.325
cc_32 VPB N_C1_M1002_g 0.0285599f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_33 VPB N_C1_c_57_n 0.00220476f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_34 VPB N_B1_M1003_g 0.0221077f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_35 VPB N_B1_c_80_n 0.00606202f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_36 VPB N_B1_c_81_n 0.00129527f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_37 VPB N_B2_M1005_g 0.0205458f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_38 VPB B2 0.00202192f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_39 VPB N_B2_c_111_n 0.00394553f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_40 VPB N_A2_M1007_g 0.0182281f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_41 VPB N_A2_c_148_n 0.00302356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A2_c_150_n 0.00589507f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_43 VPB N_A2_c_154_n 0.00333901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A1_M1009_g 0.0245333f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_45 VPB N_A1_c_195_n 0.010169f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_46 VPB N_Y_c_223_n 0.00939401f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_47 VPB N_Y_c_224_n 0.0294554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_Y_c_222_n 0.00447382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_280_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_281_n 0.0463797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_282_n 0.0159927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_283_n 0.0410358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_284_n 0.0156238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_279_n 0.0430098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_C1_c_56_n N_B1_c_80_n 0.00459621f $X=0.49 $Y=1.325 $X2=0 $Y2=0
cc_56 N_C1_c_56_n N_Y_c_223_n 0.00277415f $X=0.49 $Y=1.325 $X2=0 $Y2=0
cc_57 N_C1_c_57_n N_Y_c_223_n 0.0235546f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_58 N_C1_c_55_n N_Y_c_220_n 0.0131586f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_59 N_C1_c_57_n N_Y_c_220_n 0.00689596f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_60 N_C1_c_56_n N_Y_c_221_n 0.0022807f $X=0.49 $Y=1.325 $X2=0 $Y2=0
cc_61 N_C1_c_57_n N_Y_c_221_n 0.0212593f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_62 N_C1_M1002_g N_Y_c_232_n 0.0176964f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_63 N_C1_c_57_n N_Y_c_232_n 0.00546771f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_64 N_C1_c_55_n N_Y_c_222_n 0.00725552f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_65 N_C1_c_56_n N_Y_c_222_n 0.0096204f $X=0.49 $Y=1.325 $X2=0 $Y2=0
cc_66 N_C1_c_57_n N_Y_c_222_n 0.0253963f $X=0.38 $Y=1.16 $X2=0 $Y2=0
cc_67 N_C1_M1002_g N_VPWR_c_282_n 0.00526846f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_68 N_C1_M1002_g N_VPWR_c_284_n 0.0131577f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_69 N_C1_M1002_g N_VPWR_c_279_n 0.00978613f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_70 N_C1_c_55_n N_A_109_47#_c_326_n 0.00471569f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_71 N_C1_c_55_n N_A_213_123#_c_340_n 7.52591e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_72 N_C1_c_55_n N_VGND_c_384_n 0.00414876f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_73 N_C1_c_55_n N_VGND_c_386_n 0.00805596f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_74 N_B1_M1003_g N_B2_M1005_g 0.0421451f $X=1.4 $Y=1.985 $X2=0 $Y2=0
cc_75 N_B1_c_80_n B2 0.0026179f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B1_c_81_n B2 0.0270001f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B1_c_80_n N_B2_c_111_n 0.0421451f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B1_c_81_n N_B2_c_111_n 2.48845e-19 $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B1_c_82_n N_B2_c_112_n 0.0269334f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B1_M1003_g N_Y_c_222_n 0.00424932f $X=1.4 $Y=1.985 $X2=0 $Y2=0
cc_81 N_B1_c_80_n N_Y_c_222_n 9.59576e-19 $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B1_c_81_n N_Y_c_222_n 0.0265744f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B1_c_82_n N_Y_c_222_n 0.00352102f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_84 N_B1_M1003_g N_Y_c_241_n 0.0203375f $X=1.4 $Y=1.985 $X2=0 $Y2=0
cc_85 N_B1_c_80_n N_Y_c_241_n 0.00414942f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B1_c_81_n N_Y_c_241_n 0.0241806f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B1_M1003_g Y 0.00303841f $X=1.4 $Y=1.985 $X2=0 $Y2=0
cc_88 N_B1_M1003_g N_VPWR_c_283_n 0.00526846f $X=1.4 $Y=1.985 $X2=0 $Y2=0
cc_89 N_B1_M1003_g N_VPWR_c_284_n 0.014984f $X=1.4 $Y=1.985 $X2=0 $Y2=0
cc_90 N_B1_M1003_g N_VPWR_c_279_n 0.00883818f $X=1.4 $Y=1.985 $X2=0 $Y2=0
cc_91 N_B1_c_82_n N_A_109_47#_c_326_n 0.0100597f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B1_c_80_n N_A_213_123#_c_340_n 0.00413873f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B1_c_81_n N_A_213_123#_c_340_n 0.0239752f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B1_c_82_n N_A_213_123#_c_340_n 0.0104059f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B1_c_82_n N_VGND_c_384_n 0.00368123f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B1_c_82_n N_VGND_c_386_n 0.00665061f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B2_c_112_n N_A2_c_147_n 0.0218722f $X=1.85 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_98 N_B2_M1005_g N_A2_M1007_g 0.0164192f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_99 N_B2_M1005_g N_A2_c_148_n 0.002036f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_100 B2 N_A2_c_148_n 0.0036494f $X=1.705 $Y=1.105 $X2=0 $Y2=0
cc_101 B2 N_A2_c_149_n 0.0132014f $X=1.705 $Y=1.105 $X2=0 $Y2=0
cc_102 N_B2_c_111_n N_A2_c_149_n 5.64036e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_103 B2 N_A2_c_150_n 0.00105031f $X=1.705 $Y=1.105 $X2=0 $Y2=0
cc_104 N_B2_c_111_n N_A2_c_150_n 0.0209307f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B2_M1005_g N_A2_c_154_n 7.27201e-19 $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B2_M1005_g N_Y_c_241_n 0.00361313f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_107 B2 N_Y_c_241_n 0.0140494f $X=1.705 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B2_M1005_g Y 0.0228649f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_109 B2 Y 0.0176866f $X=1.705 $Y=1.105 $X2=0 $Y2=0
cc_110 N_B2_c_111_n Y 0.00274012f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_111 N_B2_M1005_g N_VPWR_c_283_n 0.0038803f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B2_M1005_g N_VPWR_c_284_n 0.00276282f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B2_M1005_g N_VPWR_c_279_n 0.00632068f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B2_c_112_n N_A_109_47#_c_326_n 0.00249547f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_115 B2 N_A_213_123#_c_340_n 0.0273492f $X=1.705 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B2_c_112_n N_A_213_123#_c_340_n 0.00972005f $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_117 B2 N_A_213_123#_c_349_n 0.00294124f $X=1.705 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B2_c_111_n N_A_213_123#_c_349_n 9.04308e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B2_c_112_n N_A_213_123#_c_349_n 9.65579e-19 $X=1.85 $Y=0.995 $X2=0
+ $Y2=0
cc_120 N_B2_c_112_n N_VGND_c_384_n 0.00414876f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B2_c_112_n N_VGND_c_386_n 0.00600769f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A2_c_147_n N_A1_c_193_n 0.0275845f $X=2.33 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_123 N_A2_M1007_g N_A1_M1009_g 0.0473146f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A2_c_154_n N_A1_M1009_g 0.00153496f $X=2.57 $Y=1.615 $X2=0 $Y2=0
cc_125 N_A2_c_148_n A1 0.00228278f $X=2.4 $Y=1.445 $X2=0 $Y2=0
cc_126 N_A2_c_149_n A1 0.0137887f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A2_c_150_n A1 2.26845e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A2_c_148_n N_A1_c_195_n 0.0036734f $X=2.4 $Y=1.445 $X2=0 $Y2=0
cc_129 N_A2_c_149_n N_A1_c_195_n 5.53273e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A2_c_150_n N_A1_c_195_n 0.0473146f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A2_M1007_g Y 0.00974911f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A2_c_149_n Y 0.00268175f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A2_c_150_n Y 9.94463e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A2_c_154_n N_VPWR_c_281_n 0.00642006f $X=2.57 $Y=1.615 $X2=0 $Y2=0
cc_135 N_A2_M1007_g N_VPWR_c_283_n 0.00585385f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_136 A2 N_VPWR_c_283_n 0.00781264f $X=2.485 $Y=1.785 $X2=0 $Y2=0
cc_137 N_A2_M1007_g N_VPWR_c_279_n 0.0110996f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_138 A2 N_VPWR_c_279_n 0.00776711f $X=2.485 $Y=1.785 $X2=0 $Y2=0
cc_139 N_A2_c_154_n A_493_297# 2.83863e-19 $X=2.57 $Y=1.615 $X2=-0.19 $Y2=-0.24
cc_140 A2 A_493_297# 0.00459627f $X=2.485 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_141 N_A2_c_147_n N_A_213_123#_c_341_n 0.0124263f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A2_c_149_n N_A_213_123#_c_341_n 0.0139391f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A2_c_150_n N_A_213_123#_c_341_n 0.00152291f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A2_c_154_n N_A_213_123#_c_341_n 0.00437253f $X=2.57 $Y=1.615 $X2=0
+ $Y2=0
cc_145 N_A2_c_147_n N_A_213_123#_c_342_n 5.19775e-19 $X=2.33 $Y=0.995 $X2=0
+ $Y2=0
cc_146 N_A2_c_149_n N_A_213_123#_c_349_n 0.00293317f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A2_c_150_n N_A_213_123#_c_349_n 5.40128e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_147_n N_VGND_c_383_n 0.00268723f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_147_n N_VGND_c_384_n 0.00433717f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A2_c_147_n N_VGND_c_386_n 0.00612585f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_M1009_g N_VPWR_c_281_n 0.00518824f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_152 A1 N_VPWR_c_281_n 0.0202856f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A1_c_195_n N_VPWR_c_281_n 0.00551671f $X=2.935 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A1_M1009_g N_VPWR_c_283_n 0.00585385f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A1_M1009_g N_VPWR_c_279_n 0.0114326f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A1_c_193_n N_A_213_123#_c_341_n 0.00944054f $X=2.75 $Y=0.995 $X2=0
+ $Y2=0
cc_157 A1 N_A_213_123#_c_341_n 0.0276659f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A1_c_195_n N_A_213_123#_c_341_n 0.00664911f $X=2.935 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A1_c_193_n N_A_213_123#_c_342_n 0.00594411f $X=2.75 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A1_c_193_n N_VGND_c_383_n 0.00268723f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A1_c_193_n N_VGND_c_385_n 0.00421028f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A1_c_193_n N_VGND_c_386_n 0.00663995f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_163 N_Y_c_232_n N_VPWR_M1002_d 3.68853e-19 $X=0.635 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_164 N_Y_c_222_n N_VPWR_M1002_d 2.88346e-19 $X=0.737 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_165 N_Y_c_241_n N_VPWR_M1002_d 0.017061f $X=1.735 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_166 N_Y_c_256_p N_VPWR_M1002_d 0.00335069f $X=0.737 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_167 N_Y_c_224_n N_VPWR_c_282_n 0.0194075f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_168 Y N_VPWR_c_283_n 0.0335667f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_169 N_Y_c_232_n N_VPWR_c_284_n 0.00207535f $X=0.635 $Y=1.6 $X2=0 $Y2=0
cc_170 N_Y_c_241_n N_VPWR_c_284_n 0.0363263f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_171 N_Y_c_256_p N_VPWR_c_284_n 0.018393f $X=0.737 $Y=1.6 $X2=0 $Y2=0
cc_172 Y N_VPWR_c_284_n 0.0246f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_173 N_Y_M1002_s N_VPWR_c_279_n 0.00399293f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_174 N_Y_M1005_d N_VPWR_c_279_n 0.00605065f $X=1.865 $Y=1.485 $X2=0 $Y2=0
cc_175 N_Y_c_224_n N_VPWR_c_279_n 0.0107063f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_176 Y N_VPWR_c_279_n 0.018974f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_177 N_Y_c_241_n A_295_297# 0.00628361f $X=1.735 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_178 N_Y_c_220_n N_A_109_47#_M1008_d 0.00337828f $X=0.635 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_179 N_Y_c_222_n N_A_109_47#_M1008_d 8.9915e-19 $X=0.737 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_180 N_Y_c_220_n N_A_109_47#_c_326_n 0.0200608f $X=0.635 $Y=0.735 $X2=0 $Y2=0
cc_181 N_Y_c_220_n N_A_213_123#_c_340_n 0.0166778f $X=0.635 $Y=0.735 $X2=0 $Y2=0
cc_182 N_Y_c_241_n N_A_213_123#_c_340_n 0.00263868f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_183 Y N_A_213_123#_c_349_n 0.00442842f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_184 N_Y_c_219_n N_VGND_c_384_n 0.0102332f $X=0.215 $Y=0.645 $X2=0 $Y2=0
cc_185 N_Y_c_220_n N_VGND_c_384_n 0.00239565f $X=0.635 $Y=0.735 $X2=0 $Y2=0
cc_186 N_Y_M1008_s N_VGND_c_386_n 0.00237941f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_187 N_Y_c_219_n N_VGND_c_386_n 0.00923165f $X=0.215 $Y=0.645 $X2=0 $Y2=0
cc_188 N_Y_c_220_n N_VGND_c_386_n 0.00439354f $X=0.635 $Y=0.735 $X2=0 $Y2=0
cc_189 N_VPWR_c_279_n A_295_297# 0.0102589f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_190 N_VPWR_c_279_n A_493_297# 0.00170476f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_191 N_A_109_47#_c_326_n N_A_213_123#_M1006_s 0.0045726f $X=1.61 $Y=0.39
+ $X2=-0.19 $Y2=-0.24
cc_192 N_A_109_47#_M1006_d N_A_213_123#_c_340_n 0.00327018f $X=1.475 $Y=0.235
+ $X2=0 $Y2=0
cc_193 N_A_109_47#_c_326_n N_A_213_123#_c_340_n 0.0404059f $X=1.61 $Y=0.39 $X2=0
+ $Y2=0
cc_194 N_A_109_47#_c_326_n N_VGND_c_384_n 0.0557511f $X=1.61 $Y=0.39 $X2=0 $Y2=0
cc_195 N_A_109_47#_M1008_d N_VGND_c_386_n 0.0021262f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_196 N_A_109_47#_M1006_d N_VGND_c_386_n 0.00218617f $X=1.475 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_A_109_47#_c_326_n N_VGND_c_386_n 0.0443103f $X=1.61 $Y=0.39 $X2=0 $Y2=0
cc_198 N_A_213_123#_c_341_n N_VGND_M1001_d 0.00427606f $X=2.795 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_199 N_A_213_123#_c_341_n N_VGND_c_383_n 0.012114f $X=2.795 $Y=0.78 $X2=0
+ $Y2=0
cc_200 N_A_213_123#_c_340_n N_VGND_c_384_n 0.00239565f $X=1.945 $Y=0.735 $X2=0
+ $Y2=0
cc_201 N_A_213_123#_c_341_n N_VGND_c_384_n 0.00284679f $X=2.795 $Y=0.78 $X2=0
+ $Y2=0
cc_202 N_A_213_123#_c_349_n N_VGND_c_384_n 0.0155299f $X=2.03 $Y=0.66 $X2=0
+ $Y2=0
cc_203 N_A_213_123#_c_341_n N_VGND_c_385_n 0.00211912f $X=2.795 $Y=0.78 $X2=0
+ $Y2=0
cc_204 N_A_213_123#_c_342_n N_VGND_c_385_n 0.01858f $X=2.96 $Y=0.39 $X2=0 $Y2=0
cc_205 N_A_213_123#_M1006_s N_VGND_c_386_n 0.0020511f $X=1.065 $Y=0.615 $X2=0
+ $Y2=0
cc_206 N_A_213_123#_M1000_d N_VGND_c_386_n 0.0032344f $X=1.895 $Y=0.235 $X2=0
+ $Y2=0
cc_207 N_A_213_123#_M1004_d N_VGND_c_386_n 0.00210425f $X=2.825 $Y=0.235 $X2=0
+ $Y2=0
cc_208 N_A_213_123#_c_340_n N_VGND_c_386_n 0.00558585f $X=1.945 $Y=0.735 $X2=0
+ $Y2=0
cc_209 N_A_213_123#_c_341_n N_VGND_c_386_n 0.0101818f $X=2.795 $Y=0.78 $X2=0
+ $Y2=0
cc_210 N_A_213_123#_c_342_n N_VGND_c_386_n 0.0125989f $X=2.96 $Y=0.39 $X2=0
+ $Y2=0
cc_211 N_A_213_123#_c_349_n N_VGND_c_386_n 0.0103304f $X=2.03 $Y=0.66 $X2=0
+ $Y2=0

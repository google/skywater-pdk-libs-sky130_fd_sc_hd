* File: sky130_fd_sc_hd__o21ba_1.pex.spice
* Created: Tue Sep  1 19:21:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21BA_1%A_79_199# 1 2 9 13 15 17 20 25 26 30 31 33
+ 37
c80 26 0 1.5038e-19 $X=0.595 $Y=1.16
r81 31 33 0.474307 $w=5.78e-07 $l=2.3e-08 $layer=LI1_cond $X=2.412 $Y=1.745
+ $X2=2.435 $Y2=1.745
r82 29 31 9.42427 $w=5.78e-07 $l=4.57e-07 $layer=LI1_cond $X=1.955 $Y=1.745
+ $X2=2.412 $Y2=1.745
r83 29 30 8.37612 $w=5.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.745
+ $X2=1.87 $Y2=1.745
r84 26 38 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=1.325
r85 26 37 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.562 $Y=1.16
+ $X2=0.562 $Y2=0.995
r86 25 28 6.13995 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.685 $Y=1.16
+ $X2=0.685 $Y2=1.325
r87 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r88 18 29 8.09873 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=1.955 $Y=1.455
+ $X2=1.955 $Y2=1.745
r89 18 20 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.955 $Y=1.455
+ $X2=1.955 $Y2=0.57
r90 17 30 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.86 $Y=1.95
+ $X2=1.87 $Y2=1.95
r91 15 17 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.727 $Y=1.865
+ $X2=0.86 $Y2=1.95
r92 15 28 23.4837 $w=2.63e-07 $l=5.4e-07 $layer=LI1_cond $X=0.727 $Y=1.865
+ $X2=0.727 $Y2=1.325
r93 13 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.55 $Y=0.56
+ $X2=0.55 $Y2=0.995
r94 9 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r95 2 33 300 $w=1.7e-07 $l=5.64137e-07 $layer=licon1_PDIFF $count=2 $X=2.24
+ $Y=1.485 $X2=2.435 $Y2=1.96
r96 2 33 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.485 $X2=2.435 $Y2=1.62
r97 1 20 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.235 $X2=1.955 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%B1_N 3 6 8 11 13
c34 6 0 1.93433e-19 $X=1.035 $Y=1.695
r35 11 14 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.16
+ $X2=1.115 $Y2=1.325
r36 11 13 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.16
+ $X2=1.115 $Y2=0.995
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=1.16 $X2=1.135 $Y2=1.16
r38 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.035 $Y=1.695
+ $X2=1.035 $Y2=1.325
r39 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.035 $Y=0.675
+ $X2=1.035 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%A_222_93# 1 2 7 9 12 14 15 16 20 25 28
r54 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.615
+ $Y=1.16 $X2=1.615 $Y2=1.16
r55 23 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.615 $Y=1.525
+ $X2=1.615 $Y2=1.16
r56 22 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.615 $Y=0.825
+ $X2=1.615 $Y2=1.16
r57 21 28 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.33 $Y=0.74
+ $X2=1.245 $Y2=0.66
r58 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.53 $Y=0.74
+ $X2=1.615 $Y2=0.825
r59 20 21 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.53 $Y=0.74 $X2=1.33
+ $Y2=0.74
r60 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.53 $Y=1.61
+ $X2=1.615 $Y2=1.525
r61 16 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.53 $Y=1.61
+ $X2=1.245 $Y2=1.61
r62 14 26 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=2.09 $Y=1.16
+ $X2=1.615 $Y2=1.16
r63 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.09 $Y=1.16
+ $X2=2.165 $Y2=1.16
r64 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=1.325
+ $X2=2.165 $Y2=1.16
r65 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.165 $Y=1.325
+ $X2=2.165 $Y2=1.985
r66 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=1.16
r67 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=0.56
r68 2 18 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.485 $X2=1.245 $Y2=1.61
r69 1 28 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.465 $X2=1.245 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%A2 3 6 8 11 13
r34 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.16
+ $X2=2.585 $Y2=1.325
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.16
+ $X2=2.585 $Y2=0.995
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=1.16 $X2=2.585 $Y2=1.16
r37 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.645 $Y=1.985
+ $X2=2.645 $Y2=1.325
r38 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.645 $Y=0.56
+ $X2=2.645 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%A1 3 7 8 11 13
r26 11 14 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.16
+ $X2=3.105 $Y2=1.325
r27 11 13 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.16
+ $X2=3.105 $Y2=0.995
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.115
+ $Y=1.16 $X2=3.115 $Y2=1.16
r29 8 12 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.45 $Y=1.18
+ $X2=3.115 $Y2=1.18
r30 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.065 $Y=0.56
+ $X2=3.065 $Y2=0.995
r31 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.005 $Y=1.985
+ $X2=3.005 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%X 1 2 10 15 16 17
c19 17 0 1.12617e-19 $X=0.23 $Y=2.21
c20 15 0 8.0816e-20 $X=0.26 $Y=1.645
r21 17 22 3.89797 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=0.255 $Y=2.21
+ $X2=0.255 $Y2=2.325
r22 15 16 6.33887 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=1.645
+ $X2=0.255 $Y2=1.48
r23 13 17 18.9814 $w=3.38e-07 $l=5.6e-07 $layer=LI1_cond $X=0.255 $Y=1.65
+ $X2=0.255 $Y2=2.21
r24 13 15 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.255 $Y=1.65
+ $X2=0.255 $Y2=1.645
r25 12 16 29.602 $w=2.53e-07 $l=6.55e-07 $layer=LI1_cond $X=0.212 $Y=0.825
+ $X2=0.212 $Y2=1.48
r26 10 12 6.27783 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=0.66
+ $X2=0.265 $Y2=0.825
r27 2 22 400 $w=1.7e-07 $l=9.00333e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.325
r28 2 15 400 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.645
r29 1 10 182 $w=1.7e-07 $l=4.83477e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.235 $X2=0.34 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%VPWR 1 2 3 12 16 20 25 26 27 29 34 44 45 48
+ 51
r51 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 42 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 42 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.08 $Y=2.72
+ $X2=1.915 $Y2=2.72
r58 39 41 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.08 $Y=2.72 $X2=2.99
+ $Y2=2.72
r59 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 38 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 35 48 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=0.8 $Y2=2.72
r63 35 37 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.005 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=2.72
+ $X2=1.915 $Y2=2.72
r65 34 37 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.75 $Y=2.72
+ $X2=1.61 $Y2=2.72
r66 29 48 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.8 $Y2=2.72
r67 29 31 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 27 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 25 41 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.05 $Y=2.72 $X2=2.99
+ $Y2=2.72
r71 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=2.72
+ $X2=3.215 $Y2=2.72
r72 24 44 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.38 $Y=2.72 $X2=3.45
+ $Y2=2.72
r73 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=2.72
+ $X2=3.215 $Y2=2.72
r74 20 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.215 $Y=1.62
+ $X2=3.215 $Y2=2.3
r75 18 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.635
+ $X2=3.215 $Y2=2.72
r76 18 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.215 $Y=2.635
+ $X2=3.215 $Y2=2.3
r77 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=2.635
+ $X2=1.915 $Y2=2.72
r78 14 16 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.915 $Y=2.635
+ $X2=1.915 $Y2=2.3
r79 10 48 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=2.635 $X2=0.8
+ $Y2=2.72
r80 10 12 9.69739 $w=4.08e-07 $l=3.45e-07 $layer=LI1_cond $X=0.8 $Y=2.635
+ $X2=0.8 $Y2=2.29
r81 3 23 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.485 $X2=3.215 $Y2=2.3
r82 3 20 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.485 $X2=3.215 $Y2=1.62
r83 2 16 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.485 $X2=1.915 $Y2=2.3
r84 1 12 600 $w=1.7e-07 $l=9.06146e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.76 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%VGND 1 2 9 13 16 17 19 20 21 34 35
c45 9 0 1.5038e-19 $X=0.795 $Y=0.66
r46 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r47 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r48 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r49 29 32 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r50 28 31 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r51 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r52 25 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r53 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r54 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r55 19 31 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.77 $Y=0 $X2=2.53
+ $Y2=0
r56 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0 $X2=2.855
+ $Y2=0
r57 18 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=3.45
+ $Y2=0
r58 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0 $X2=2.855
+ $Y2=0
r59 16 24 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.69
+ $Y2=0
r60 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.795
+ $Y2=0
r61 15 28 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.15
+ $Y2=0
r62 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.795
+ $Y2=0
r63 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r64 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.39
r65 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r66 7 9 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.66
r67 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.235 $X2=2.855 $Y2=0.39
r68 1 9 182 $w=1.7e-07 $l=5.02867e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.235 $X2=0.795 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_1%A_448_47# 1 2 9 11 12 15
r28 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.275 $Y=0.735
+ $X2=3.275 $Y2=0.39
r29 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.11 $Y=0.82
+ $X2=3.275 $Y2=0.735
r30 11 12 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.11 $Y=0.82 $X2=2.6
+ $Y2=0.82
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.435 $Y=0.735
+ $X2=2.6 $Y2=0.82
r32 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.435 $Y=0.735
+ $X2=2.435 $Y2=0.39
r33 2 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.235 $X2=3.275 $Y2=0.39
r34 1 9 91 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=2 $X=2.24
+ $Y=0.235 $X2=2.435 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__or2_1.spice.SKY130_FD_SC_HD__OR2_1.pxi
* Created: Thu Aug 27 14:42:34 2020
* 
x_PM_SKY130_FD_SC_HD__OR2_1%B N_B_M1003_g N_B_M1004_g B B N_B_c_41_n
+ PM_SKY130_FD_SC_HD__OR2_1%B
x_PM_SKY130_FD_SC_HD__OR2_1%A N_A_M1000_g N_A_M1002_g A A N_A_c_69_n
+ PM_SKY130_FD_SC_HD__OR2_1%A
x_PM_SKY130_FD_SC_HD__OR2_1%A_68_297# N_A_68_297#_M1003_d N_A_68_297#_M1004_s
+ N_A_68_297#_M1001_g N_A_68_297#_M1005_g N_A_68_297#_c_104_n
+ N_A_68_297#_c_124_n N_A_68_297#_c_110_n N_A_68_297#_c_105_n
+ N_A_68_297#_c_106_n N_A_68_297#_c_120_n N_A_68_297#_c_107_n
+ PM_SKY130_FD_SC_HD__OR2_1%A_68_297#
x_PM_SKY130_FD_SC_HD__OR2_1%VPWR N_VPWR_M1002_d N_VPWR_c_162_n VPWR
+ N_VPWR_c_163_n N_VPWR_c_164_n N_VPWR_c_161_n N_VPWR_c_166_n
+ PM_SKY130_FD_SC_HD__OR2_1%VPWR
x_PM_SKY130_FD_SC_HD__OR2_1%X N_X_M1001_d N_X_M1005_d N_X_c_181_n X X
+ PM_SKY130_FD_SC_HD__OR2_1%X
x_PM_SKY130_FD_SC_HD__OR2_1%VGND N_VGND_M1003_s N_VGND_M1000_d N_VGND_c_206_n
+ N_VGND_c_207_n N_VGND_c_208_n N_VGND_c_209_n N_VGND_c_210_n VGND
+ N_VGND_c_211_n N_VGND_c_212_n PM_SKY130_FD_SC_HD__OR2_1%VGND
cc_1 VNB N_B_M1003_g 0.0331172f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.445
cc_2 VNB B 0.0261495f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B_c_41_n 0.0393495f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.16
cc_4 VNB N_A_M1000_g 0.0285171f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.445
cc_5 VNB A 0.00450205f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_6 VNB N_A_c_69_n 0.0206472f $X=-0.19 $Y=-0.24 $X2=0.415 $Y2=1.16
cc_7 VNB N_A_68_297#_c_104_n 0.00420445f $X=-0.19 $Y=-0.24 $X2=0.415 $Y2=1.16
cc_8 VNB N_A_68_297#_c_105_n 9.29423e-19 $X=-0.19 $Y=-0.24 $X2=0.322 $Y2=0.85
cc_9 VNB N_A_68_297#_c_106_n 0.0280668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_68_297#_c_107_n 0.0202332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_VPWR_c_161_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.16
cc_12 VNB N_X_c_181_n 0.0333687f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_13 VNB X 0.02761f $X=-0.19 $Y=-0.24 $X2=0.415 $Y2=1.16
cc_14 VNB N_VGND_c_206_n 0.0144081f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.695
cc_15 VNB N_VGND_c_207_n 0.0185f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_16 VNB N_VGND_c_208_n 0.00493424f $X=-0.19 $Y=-0.24 $X2=0.415 $Y2=1.16
cc_17 VNB N_VGND_c_209_n 0.0193288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_210_n 0.00410625f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.16
cc_19 VNB N_VGND_c_211_n 0.0250559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_212_n 0.149265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_B_M1004_g 0.0272481f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.695
cc_22 VPB B 0.00782337f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_23 VPB N_B_c_41_n 0.0115141f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_24 VPB N_A_M1002_g 0.0206595f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.695
cc_25 VPB A 0.00167213f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_26 VPB N_A_c_69_n 0.0045414f $X=-0.19 $Y=1.305 $X2=0.415 $Y2=1.16
cc_27 VPB N_A_68_297#_M1005_g 0.0254771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_68_297#_c_104_n 0.00160812f $X=-0.19 $Y=1.305 $X2=0.415 $Y2=1.16
cc_29 VPB N_A_68_297#_c_110_n 0.0175009f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.16
cc_30 VPB N_A_68_297#_c_105_n 0.00146985f $X=-0.19 $Y=1.305 $X2=0.322 $Y2=0.85
cc_31 VPB N_A_68_297#_c_106_n 0.00684409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_162_n 0.0215687f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.695
cc_33 VPB N_VPWR_c_163_n 0.0385795f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_34 VPB N_VPWR_c_164_n 0.0223354f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.16
cc_35 VPB N_VPWR_c_161_n 0.0829129f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_36 VPB N_VPWR_c_166_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB X 0.0263845f $X=-0.19 $Y=1.305 $X2=0.415 $Y2=1.16
cc_38 VPB X 0.0318853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 N_B_M1003_g N_A_M1000_g 0.0223994f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_40 N_B_M1004_g N_A_M1002_g 0.0318915f $X=0.675 $Y=1.695 $X2=0 $Y2=0
cc_41 N_B_M1003_g A 2.11082e-19 $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_42 N_B_c_41_n A 3.17146e-19 $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_43 N_B_c_41_n N_A_c_69_n 0.0318915f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_44 N_B_M1003_g N_A_68_297#_c_104_n 0.0117741f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_45 N_B_M1004_g N_A_68_297#_c_104_n 0.00820962f $X=0.675 $Y=1.695 $X2=0 $Y2=0
cc_46 B N_A_68_297#_c_104_n 0.0411416f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_47 N_B_c_41_n N_A_68_297#_c_104_n 0.00980993f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_48 N_B_M1004_g N_A_68_297#_c_110_n 0.0174028f $X=0.675 $Y=1.695 $X2=0 $Y2=0
cc_49 B N_A_68_297#_c_110_n 0.0188518f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_50 N_B_c_41_n N_A_68_297#_c_110_n 0.00488703f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_51 N_B_M1003_g N_A_68_297#_c_120_n 0.00364962f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_52 N_B_M1004_g N_VPWR_c_163_n 0.00327927f $X=0.675 $Y=1.695 $X2=0 $Y2=0
cc_53 N_B_M1004_g N_VPWR_c_161_n 0.00417489f $X=0.675 $Y=1.695 $X2=0 $Y2=0
cc_54 B N_VGND_c_206_n 0.00162397f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_55 N_B_M1003_g N_VGND_c_207_n 0.00448362f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_56 B N_VGND_c_207_n 0.0206591f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_B_c_41_n N_VGND_c_207_n 0.00110332f $X=0.675 $Y=1.16 $X2=0 $Y2=0
cc_58 N_B_M1003_g N_VGND_c_209_n 0.00556805f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_59 N_B_M1003_g N_VGND_c_212_n 0.010966f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_60 B N_VGND_c_212_n 0.00417208f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_A_68_297#_M1005_g 0.0193785f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_A_68_297#_c_104_n 0.0104173f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_63 A N_A_68_297#_c_104_n 0.0413542f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_64 N_A_M1002_g N_A_68_297#_c_124_n 0.0158541f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_65 A N_A_68_297#_c_124_n 0.0182242f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_66 N_A_c_69_n N_A_68_297#_c_124_n 7.21566e-19 $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_A_68_297#_c_110_n 9.32062e-19 $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_68 N_A_M1002_g N_A_68_297#_c_105_n 8.77094e-19 $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_69 A N_A_68_297#_c_105_n 0.0183661f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_70 N_A_c_69_n N_A_68_297#_c_105_n 3.45798e-19 $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_69_n N_A_68_297#_c_106_n 0.0199989f $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_A_68_297#_c_107_n 0.0173675f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_73 A N_A_68_297#_c_107_n 0.00454052f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_74 N_A_M1002_g N_VPWR_c_162_n 0.00404488f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_75 N_A_M1002_g N_VPWR_c_163_n 0.00327927f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_76 N_A_M1002_g N_VPWR_c_161_n 0.00417489f $X=1.035 $Y=1.695 $X2=0 $Y2=0
cc_77 N_A_M1000_g N_X_c_181_n 8.74927e-19 $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_78 A N_X_c_181_n 0.0031434f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_79 A X 0.00569575f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_80 A N_VGND_M1000_d 0.00243754f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_M1000_g N_VGND_c_208_n 0.00453377f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_82 A N_VGND_c_208_n 0.0080166f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_83 N_A_c_69_n N_VGND_c_208_n 2.29546e-19 $X=1.095 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_M1000_g N_VGND_c_209_n 0.00585385f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_M1000_g N_VGND_c_212_n 0.0077776f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_86 A N_VGND_c_212_n 0.00654989f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_87 N_A_68_297#_c_124_n A_150_297# 0.00473129f $X=1.525 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_68_297#_c_110_n A_150_297# 0.00144354f $X=0.84 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_68_297#_c_124_n N_VPWR_M1002_d 0.00769283f $X=1.525 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_90 N_A_68_297#_M1005_g N_VPWR_c_162_n 0.014753f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_68_297#_c_124_n N_VPWR_c_162_n 0.0201472f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A_68_297#_M1005_g N_VPWR_c_164_n 0.0046653f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_68_297#_M1005_g N_VPWR_c_161_n 0.00915924f $X=1.52 $Y=1.985 $X2=0
+ $Y2=0
cc_94 N_A_68_297#_c_124_n N_X_M1005_d 0.00236185f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A_68_297#_c_105_n N_X_c_181_n 0.00844569f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_68_297#_c_106_n N_X_c_181_n 0.00409566f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_68_297#_c_107_n N_X_c_181_n 0.00857784f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A_68_297#_M1005_g X 0.00780242f $X=1.52 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_68_297#_c_124_n X 0.0144304f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_100 N_A_68_297#_c_105_n X 0.038181f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_68_297#_c_106_n X 0.00826352f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_68_297#_c_107_n X 0.00270973f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_68_297#_c_124_n X 0.00364128f $X=1.525 $Y=1.58 $X2=0 $Y2=0
cc_104 N_A_68_297#_c_106_n X 0.0026095f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_68_297#_c_107_n N_VGND_c_208_n 0.0028487f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_A_68_297#_c_120_n N_VGND_c_209_n 0.0147354f $X=0.825 $Y=0.43 $X2=0
+ $Y2=0
cc_107 N_A_68_297#_c_107_n N_VGND_c_211_n 0.00539883f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_108 N_A_68_297#_M1003_d N_VGND_c_212_n 0.00250238f $X=0.69 $Y=0.235 $X2=0
+ $Y2=0
cc_109 N_A_68_297#_c_120_n N_VGND_c_212_n 0.010419f $X=0.825 $Y=0.43 $X2=0 $Y2=0
cc_110 N_A_68_297#_c_107_n N_VGND_c_212_n 0.0107909f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_111 N_VPWR_c_161_n N_X_M1005_d 0.00452756f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_112 N_VPWR_c_162_n X 3.8678e-19 $X=1.31 $Y=1.92 $X2=0 $Y2=0
cc_113 N_VPWR_c_164_n X 0.0375063f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_114 N_VPWR_c_161_n X 0.0205064f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_115 N_X_c_181_n N_VGND_c_211_n 0.0408267f $X=2.022 $Y=0.54 $X2=0 $Y2=0
cc_116 N_X_M1001_d N_VGND_c_212_n 0.00209344f $X=1.595 $Y=0.235 $X2=0 $Y2=0
cc_117 N_X_c_181_n N_VGND_c_212_n 0.0233535f $X=2.022 $Y=0.54 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__mux2i_2.spice.SKY130_FD_SC_HD__MUX2I_2.pxi
* Created: Thu Aug 27 14:28:02 2020
* 
x_PM_SKY130_FD_SC_HD__MUX2I_2%S N_S_c_82_n N_S_M1016_g N_S_M1010_g N_S_c_83_n
+ N_S_M1004_g N_S_M1000_g N_S_c_84_n N_S_M1009_g N_S_M1001_g S S N_S_c_86_n
+ PM_SKY130_FD_SC_HD__MUX2I_2%S
x_PM_SKY130_FD_SC_HD__MUX2I_2%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1010_s
+ N_A_27_47#_M1008_g N_A_27_47#_M1011_g N_A_27_47#_M1013_g N_A_27_47#_M1014_g
+ N_A_27_47#_c_151_n N_A_27_47#_c_170_n N_A_27_47#_c_158_n N_A_27_47#_c_177_n
+ N_A_27_47#_c_152_n N_A_27_47#_c_159_n N_A_27_47#_c_160_n N_A_27_47#_c_161_n
+ N_A_27_47#_c_180_n N_A_27_47#_c_153_n N_A_27_47#_c_154_n
+ PM_SKY130_FD_SC_HD__MUX2I_2%A_27_47#
x_PM_SKY130_FD_SC_HD__MUX2I_2%A0 N_A0_c_244_n N_A0_M1002_g N_A0_M1003_g
+ N_A0_c_245_n N_A0_M1005_g N_A0_M1012_g A0 A0 A0 N_A0_c_247_n N_A0_c_248_n
+ PM_SKY130_FD_SC_HD__MUX2I_2%A0
x_PM_SKY130_FD_SC_HD__MUX2I_2%A1 N_A1_c_299_n N_A1_M1006_g N_A1_M1007_g
+ N_A1_c_300_n N_A1_M1017_g N_A1_M1015_g A1 A1 N_A1_c_301_n N_A1_c_302_n
+ PM_SKY130_FD_SC_HD__MUX2I_2%A1
x_PM_SKY130_FD_SC_HD__MUX2I_2%VPWR N_VPWR_M1010_d N_VPWR_M1001_d N_VPWR_M1014_d
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_351_n VPWR N_VPWR_c_352_n N_VPWR_c_353_n
+ N_VPWR_c_344_n N_VPWR_c_355_n PM_SKY130_FD_SC_HD__MUX2I_2%VPWR
x_PM_SKY130_FD_SC_HD__MUX2I_2%A_193_297# N_A_193_297#_M1000_s
+ N_A_193_297#_M1003_d N_A_193_297#_c_416_n N_A_193_297#_c_419_n
+ N_A_193_297#_c_420_n N_A_193_297#_c_434_n N_A_193_297#_c_415_n
+ PM_SKY130_FD_SC_HD__MUX2I_2%A_193_297#
x_PM_SKY130_FD_SC_HD__MUX2I_2%A_361_297# N_A_361_297#_M1011_s
+ N_A_361_297#_M1007_s N_A_361_297#_c_469_n N_A_361_297#_c_465_n
+ N_A_361_297#_c_463_n N_A_361_297#_c_464_n
+ PM_SKY130_FD_SC_HD__MUX2I_2%A_361_297#
x_PM_SKY130_FD_SC_HD__MUX2I_2%Y N_Y_M1002_d N_Y_M1005_d N_Y_M1017_d N_Y_M1003_s
+ N_Y_M1012_s N_Y_M1015_d N_Y_c_499_n Y Y N_Y_c_503_n Y Y
+ PM_SKY130_FD_SC_HD__MUX2I_2%Y
x_PM_SKY130_FD_SC_HD__MUX2I_2%VGND N_VGND_M1016_d N_VGND_M1009_s N_VGND_M1013_s
+ N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n N_VGND_c_557_n N_VGND_c_558_n
+ N_VGND_c_559_n N_VGND_c_560_n VGND N_VGND_c_561_n N_VGND_c_562_n
+ N_VGND_c_563_n N_VGND_c_564_n PM_SKY130_FD_SC_HD__MUX2I_2%VGND
x_PM_SKY130_FD_SC_HD__MUX2I_2%A_193_47# N_A_193_47#_M1004_d N_A_193_47#_M1006_s
+ N_A_193_47#_c_629_n N_A_193_47#_c_630_n N_A_193_47#_c_631_n
+ N_A_193_47#_c_632_n N_A_193_47#_c_633_n PM_SKY130_FD_SC_HD__MUX2I_2%A_193_47#
x_PM_SKY130_FD_SC_HD__MUX2I_2%A_361_47# N_A_361_47#_M1008_d N_A_361_47#_M1002_s
+ N_A_361_47#_c_717_n N_A_361_47#_c_695_n N_A_361_47#_c_696_n
+ N_A_361_47#_c_697_n PM_SKY130_FD_SC_HD__MUX2I_2%A_361_47#
cc_1 VNB N_S_c_82_n 0.0189749f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_S_c_83_n 0.0157864f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_S_c_84_n 0.0157144f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB S 0.00140974f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_5 VNB N_S_c_86_n 0.0512782f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_6 VNB N_A_27_47#_M1008_g 0.0171828f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_7 VNB N_A_27_47#_M1013_g 0.0227686f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_8 VNB N_A_27_47#_c_151_n 0.027241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_152_n 0.01296f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.85
cc_10 VNB N_A_27_47#_c_153_n 0.00229698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_154_n 0.0296451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A0_c_244_n 0.0212161f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_A0_c_245_n 0.016268f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_14 VNB A0 0.00185106f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_15 VNB N_A0_c_247_n 0.0473557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A0_c_248_n 0.0297862f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_17 VNB N_A1_c_299_n 0.0158472f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_18 VNB N_A1_c_300_n 0.0196132f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_19 VNB N_A1_c_301_n 0.0501319f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_20 VNB N_A1_c_302_n 0.00251523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_344_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_499_n 0.00990813f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_23 VNB Y 0.0350897f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_24 VNB N_VGND_c_554_n 4.10862e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_25 VNB N_VGND_c_555_n 0.00247096f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_26 VNB N_VGND_c_556_n 0.00411685f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_27 VNB N_VGND_c_557_n 0.0167892f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_28 VNB N_VGND_c_558_n 0.00356594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_559_n 0.0152839f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_30 VNB N_VGND_c_560_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_561_n 0.0154495f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_32 VNB N_VGND_c_562_n 0.0647519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_563_n 0.259129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_564_n 0.00423302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_47#_c_629_n 0.0189307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_47#_c_630_n 0.00311847f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_37 VNB N_A_193_47#_c_631_n 0.00634489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_c_632_n 0.0029815f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_39 VNB N_A_193_47#_c_633_n 0.00210775f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_40 VNB N_A_361_47#_c_695_n 9.62668e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_41 VNB N_A_361_47#_c_696_n 9.23525e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_361_47#_c_697_n 0.00980739f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_43 VPB N_S_M1010_g 0.0217492f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_S_M1000_g 0.0182511f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_45 VPB N_S_M1001_g 0.0169285f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_46 VPB S 8.43337e-19 $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_47 VPB N_S_c_86_n 0.00799888f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_48 VPB N_A_27_47#_M1011_g 0.0185382f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_49 VPB N_A_27_47#_M1014_g 0.0259828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_151_n 0.00903094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_158_n 0.00325282f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_52 VPB N_A_27_47#_c_159_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_160_n 0.0128993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_161_n 0.0169831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_153_n 0.00316123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_154_n 0.0050694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A0_M1003_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_58 VPB N_A0_M1012_g 0.0192809f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_59 VPB N_A0_c_248_n 0.00607782f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_60 VPB N_A1_M1007_g 0.0193168f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_A1_M1015_g 0.0223888f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_A1_c_301_n 0.014288f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_63 VPB N_A1_c_302_n 0.00326631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_345_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_65 VPB N_VPWR_c_346_n 3.15634e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_66 VPB N_VPWR_c_347_n 0.00851371f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_67 VPB N_VPWR_c_348_n 0.0124848f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_68 VPB N_VPWR_c_349_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_350_n 0.0145058f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_70 VPB N_VPWR_c_351_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_352_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_72 VPB N_VPWR_c_353_n 0.0624642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_344_n 0.0467416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_355_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_193_297#_c_415_n 0.00583938f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_76 VPB N_A_361_297#_c_463_n 0.00609927f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_77 VPB N_A_361_297#_c_464_n 0.00182633f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_78 VPB Y 0.0367183f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_79 VPB Y 0.00218948f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_80 VPB N_Y_c_503_n 0.00762094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 N_S_c_84_n N_A_27_47#_M1008_g 0.0138377f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_82 N_S_M1001_g N_A_27_47#_M1011_g 0.0435283f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_83 N_S_c_82_n N_A_27_47#_c_151_n 0.00708648f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_84 N_S_M1010_g N_A_27_47#_c_151_n 0.00603009f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_85 S N_A_27_47#_c_151_n 0.0341606f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_86 N_S_c_86_n N_A_27_47#_c_151_n 0.00922146f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_87 N_S_M1010_g N_A_27_47#_c_170_n 0.0169771f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_88 N_S_M1000_g N_A_27_47#_c_170_n 0.0180709f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_89 N_S_M1001_g N_A_27_47#_c_170_n 0.00701627f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_90 S N_A_27_47#_c_170_n 0.0235323f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_91 N_S_c_86_n N_A_27_47#_c_170_n 0.00301158f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_92 N_S_M1000_g N_A_27_47#_c_158_n 0.0029474f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 N_S_M1001_g N_A_27_47#_c_158_n 0.00334921f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_94 S N_A_27_47#_c_177_n 0.00624934f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_95 N_S_c_86_n N_A_27_47#_c_177_n 0.0115245f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_96 N_S_M1010_g N_A_27_47#_c_161_n 0.0144508f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_97 N_S_c_86_n N_A_27_47#_c_180_n 5.75762e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_98 N_S_c_86_n N_A_27_47#_c_154_n 0.0171028f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_99 N_S_M1010_g N_VPWR_c_345_n 0.00874453f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_100 N_S_M1000_g N_VPWR_c_345_n 0.00850568f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_101 N_S_M1001_g N_VPWR_c_345_n 0.00110281f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_102 N_S_M1000_g N_VPWR_c_346_n 0.00110281f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_103 N_S_M1001_g N_VPWR_c_346_n 0.00816739f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_104 N_S_M1000_g N_VPWR_c_348_n 0.00436751f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_105 N_S_M1001_g N_VPWR_c_348_n 0.00348405f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_106 N_S_M1010_g N_VPWR_c_352_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_S_M1010_g N_VPWR_c_344_n 0.008846f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_108 N_S_M1000_g N_VPWR_c_344_n 0.00702003f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_109 N_S_M1001_g N_VPWR_c_344_n 0.00414556f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_110 N_S_M1010_g N_A_193_297#_c_416_n 5.24915e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_111 N_S_M1000_g N_A_193_297#_c_416_n 0.00447395f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_112 N_S_M1001_g N_A_193_297#_c_416_n 0.00975793f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_113 N_S_M1001_g N_A_193_297#_c_419_n 0.0034207f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_114 N_S_M1001_g N_A_193_297#_c_420_n 6.60451e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_115 S N_VGND_M1016_d 0.00249482f $X=0.61 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_116 N_S_c_82_n N_VGND_c_554_n 0.0124497f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_117 N_S_c_83_n N_VGND_c_554_n 0.0101604f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_118 N_S_c_84_n N_VGND_c_554_n 0.00137663f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_119 S N_VGND_c_554_n 0.0143427f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_120 N_S_c_86_n N_VGND_c_554_n 3.90313e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_121 N_S_c_84_n N_VGND_c_555_n 0.00157006f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_122 N_S_c_83_n N_VGND_c_557_n 0.00505556f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_123 N_S_c_84_n N_VGND_c_557_n 0.00563907f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_124 N_S_c_82_n N_VGND_c_561_n 0.0046653f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_125 N_S_c_82_n N_VGND_c_563_n 0.00895857f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_126 N_S_c_83_n N_VGND_c_563_n 0.00858194f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_127 N_S_c_84_n N_VGND_c_563_n 0.00613461f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_128 S N_VGND_c_563_n 8.77277e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_129 N_S_c_84_n N_A_193_47#_c_629_n 0.00239247f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_130 N_S_c_83_n N_A_193_47#_c_630_n 0.00408989f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_131 N_S_c_84_n N_A_193_47#_c_630_n 0.0025566f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_132 S N_A_193_47#_c_630_n 0.00758543f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_133 N_S_c_86_n N_A_193_47#_c_630_n 0.00252992f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_134 N_S_c_83_n N_A_193_47#_c_633_n 6.21302e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_135 N_S_c_84_n N_A_193_47#_c_633_n 0.00450329f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_136 S N_A_193_47#_c_633_n 0.00434984f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_137 N_S_c_86_n N_A_193_47#_c_633_n 0.00269478f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_180_n A0 0.00694836f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_154_n A0 9.19871e-19 $X=2.15 $Y=1.175 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1013_g N_A0_c_247_n 0.0177662f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_180_n N_A0_c_247_n 2.76827e-19 $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_170_n N_VPWR_M1010_d 0.00452837f $X=1.225 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A_27_47#_c_170_n N_VPWR_c_345_n 0.00643049f $X=1.225 $Y=1.58 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_M1011_g N_VPWR_c_346_n 0.00688248f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_M1014_g N_VPWR_c_346_n 4.79856e-19 $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_M1014_g N_VPWR_c_347_n 0.00311793f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_M1011_g N_VPWR_c_350_n 0.00417846f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_M1014_g N_VPWR_c_350_n 0.00433859f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_160_n N_VPWR_c_352_n 0.0177247f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_150 N_A_27_47#_M1010_s N_VPWR_c_344_n 0.00382897f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_M1011_g N_VPWR_c_344_n 0.00627998f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_M1014_g N_VPWR_c_344_n 0.00713033f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_160_n N_VPWR_c_344_n 0.00987844f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_170_n N_A_193_297#_M1000_s 0.0040413f $X=1.225 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_155 N_A_27_47#_M1011_g N_A_193_297#_c_416_n 0.00606173f $X=1.73 $Y=1.985
+ $X2=0 $Y2=0
cc_156 N_A_27_47#_c_170_n N_A_193_297#_c_416_n 0.0244519f $X=1.225 $Y=1.58 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_161_n N_A_193_297#_c_416_n 0.00436842f $X=0.215 $Y=2.135
+ $X2=0 $Y2=0
cc_158 N_A_27_47#_c_153_n N_A_193_297#_c_416_n 0.00493725f $X=1.655 $Y=1.2 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_M1011_g N_A_193_297#_c_419_n 0.00449992f $X=1.73 $Y=1.985
+ $X2=0 $Y2=0
cc_160 N_A_27_47#_M1014_g N_A_193_297#_c_419_n 9.29105e-19 $X=2.15 $Y=1.985
+ $X2=0 $Y2=0
cc_161 N_A_27_47#_M1011_g N_A_193_297#_c_420_n 0.00337042f $X=1.73 $Y=1.985
+ $X2=0 $Y2=0
cc_162 N_A_27_47#_c_153_n N_A_193_297#_c_420_n 0.0106017f $X=1.655 $Y=1.2 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_M1011_g N_A_193_297#_c_415_n 0.00702893f $X=1.73 $Y=1.985
+ $X2=0 $Y2=0
cc_164 N_A_27_47#_M1014_g N_A_193_297#_c_415_n 0.0143493f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_180_n N_A_193_297#_c_415_n 0.01543f $X=1.82 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_154_n N_A_193_297#_c_415_n 0.0019787f $X=2.15 $Y=1.175 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_M1011_g N_A_361_297#_c_465_n 0.00402742f $X=1.73 $Y=1.985
+ $X2=0 $Y2=0
cc_168 N_A_27_47#_M1014_g N_A_361_297#_c_465_n 0.010267f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_M1014_g N_A_361_297#_c_463_n 0.0118711f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_M1014_g N_A_361_297#_c_464_n 0.00138752f $X=2.15 $Y=1.985
+ $X2=0 $Y2=0
cc_171 N_A_27_47#_M1008_g N_VGND_c_555_n 0.0106535f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1013_g N_VGND_c_555_n 8.5303e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_180_n N_VGND_c_555_n 0.00158864f $X=1.82 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_153_n N_VGND_c_555_n 0.00821347f $X=1.655 $Y=1.2 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_154_n N_VGND_c_555_n 3.34217e-19 $X=2.15 $Y=1.175 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1013_g N_VGND_c_556_n 0.0030732f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1008_g N_VGND_c_559_n 0.0046653f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A_27_47#_M1013_g N_VGND_c_559_n 0.00439206f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_152_n N_VGND_c_561_n 0.0112151f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1016_s N_VGND_c_563_n 0.00394021f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1008_g N_VGND_c_563_n 0.00443939f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1013_g N_VGND_c_563_n 0.00689604f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_152_n N_VGND_c_563_n 0.00939877f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1008_g N_A_193_47#_c_629_n 0.00435566f $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_M1013_g N_A_193_47#_c_629_n 0.00251177f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_177_n N_A_193_47#_c_629_n 0.00387656f $X=1.395 $Y=1.24 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_180_n N_A_193_47#_c_629_n 0.011031f $X=1.82 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_153_n N_A_193_47#_c_629_n 0.00714923f $X=1.655 $Y=1.2 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_154_n N_A_193_47#_c_629_n 0.00259044f $X=2.15 $Y=1.175 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1008_g N_A_193_47#_c_630_n 2.13938e-19 $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_170_n N_A_193_47#_c_630_n 0.00479736f $X=1.225 $Y=1.58 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_177_n N_A_193_47#_c_630_n 0.00277842f $X=1.395 $Y=1.24 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1008_g N_A_193_47#_c_633_n 3.04786e-19 $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_170_n N_A_193_47#_c_633_n 0.00337433f $X=1.225 $Y=1.58 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_177_n N_A_193_47#_c_633_n 0.00145554f $X=1.395 $Y=1.24 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_M1008_g N_A_361_47#_c_695_n 9.44612e-19 $X=1.73 $Y=0.56 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_180_n N_A_361_47#_c_695_n 0.00859309f $X=1.82 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_154_n N_A_361_47#_c_695_n 0.00209037f $X=2.15 $Y=1.175 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_M1013_g N_A_361_47#_c_697_n 0.0145901f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_200 N_A0_c_245_n N_A1_c_299_n 0.0231532f $X=3.51 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_201 N_A0_M1012_g N_A1_M1007_g 0.0414912f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_202 A0 N_A1_c_301_n 0.00129358f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A0_c_248_n N_A1_c_301_n 0.0189538f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A0_c_248_n N_A1_c_302_n 0.00117539f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A0_M1003_g N_VPWR_c_347_n 0.00285342f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A0_M1003_g N_VPWR_c_353_n 0.00366111f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A0_M1012_g N_VPWR_c_353_n 0.00366111f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A0_M1003_g N_VPWR_c_344_n 0.00656615f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A0_M1012_g N_VPWR_c_344_n 0.00536271f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A0_M1003_g N_A_193_297#_c_434_n 0.00350536f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A0_M1012_g N_A_193_297#_c_434_n 0.00531718f $X=3.51 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A0_c_248_n N_A_193_297#_c_434_n 0.00208572f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A0_M1003_g N_A_193_297#_c_415_n 0.00978883f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_214 A0 N_A_193_297#_c_415_n 0.0503682f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_215 N_A0_c_247_n N_A_193_297#_c_415_n 0.0117023f $X=3.015 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A0_M1003_g N_A_361_297#_c_469_n 0.0125459f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A0_M1012_g N_A_361_297#_c_469_n 0.0127111f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_218 A0 N_A_361_297#_c_469_n 0.00216392f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_219 N_A0_M1003_g N_A_361_297#_c_464_n 0.00339149f $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A0_c_244_n N_Y_c_499_n 0.00830822f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A0_c_245_n N_Y_c_499_n 0.00914927f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_222 A0 N_Y_c_499_n 9.08118e-19 $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_223 N_A0_M1003_g Y 0.00789149f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A0_M1012_g Y 0.00789149f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A0_c_244_n N_VGND_c_556_n 0.00241512f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A0_c_244_n N_VGND_c_562_n 0.00366111f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A0_c_245_n N_VGND_c_562_n 0.00366111f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A0_c_244_n N_VGND_c_563_n 0.00650956f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A0_c_245_n N_VGND_c_563_n 0.00530612f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A0_c_244_n N_A_193_47#_c_629_n 0.00167352f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A0_c_245_n N_A_193_47#_c_629_n 0.00455389f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_232 A0 N_A_193_47#_c_629_n 0.0270209f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A0_c_247_n N_A_193_47#_c_629_n 0.0136728f $X=3.015 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A0_c_248_n N_A_193_47#_c_629_n 0.00319156f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A0_c_245_n N_A_193_47#_c_631_n 0.00135525f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A0_c_245_n N_A_193_47#_c_632_n 0.00141163f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A0_c_244_n N_A_361_47#_c_696_n 0.00478547f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A0_c_245_n N_A_361_47#_c_696_n 0.0040908f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A0_c_248_n N_A_361_47#_c_696_n 0.00218833f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A0_c_244_n N_A_361_47#_c_697_n 0.00889719f $X=3.09 $Y=0.995 $X2=0 $Y2=0
cc_241 A0 N_A_361_47#_c_697_n 0.0624906f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_242 N_A0_c_247_n N_A_361_47#_c_697_n 0.012914f $X=3.015 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A1_M1007_g N_VPWR_c_353_n 0.00366111f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A1_M1015_g N_VPWR_c_353_n 0.00366111f $X=4.395 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A1_M1007_g N_VPWR_c_344_n 0.00537647f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A1_M1015_g N_VPWR_c_344_n 0.00634973f $X=4.395 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A1_M1007_g N_A_193_297#_c_434_n 0.00105222f $X=3.97 $Y=1.985 $X2=0
+ $Y2=0
cc_248 N_A1_M1007_g N_A_361_297#_c_469_n 0.0130945f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A1_M1015_g N_A_361_297#_c_469_n 0.00377055f $X=4.395 $Y=1.985 $X2=0
+ $Y2=0
cc_250 N_A1_c_301_n N_A_361_297#_c_469_n 0.00230667f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A1_c_302_n N_A_361_297#_c_469_n 0.0014153f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A1_c_302_n N_Y_M1015_d 0.00371992f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A1_c_299_n N_Y_c_499_n 0.00798178f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_300_n N_Y_c_499_n 0.0132534f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_301_n N_Y_c_499_n 0.00265292f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A1_c_302_n N_Y_c_499_n 0.0080624f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A1_c_300_n Y 0.0133829f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A1_M1015_g Y 0.0172805f $X=4.395 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A1_c_301_n Y 0.00949568f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A1_c_302_n Y 0.047363f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A1_M1007_g Y 0.00792292f $X=3.97 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A1_M1015_g Y 0.00964912f $X=4.395 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A1_c_302_n Y 0.00617293f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A1_c_299_n N_VGND_c_562_n 0.00366111f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A1_c_300_n N_VGND_c_562_n 0.00366111f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A1_c_299_n N_VGND_c_563_n 0.00527136f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A1_c_300_n N_VGND_c_563_n 0.00643087f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A1_c_299_n N_A_193_47#_c_631_n 0.00651291f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A1_c_300_n N_A_193_47#_c_631_n 4.34273e-19 $X=4.395 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A1_c_299_n N_A_193_47#_c_632_n 0.0113598f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_c_300_n N_A_193_47#_c_632_n 0.00587593f $X=4.395 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A1_c_301_n N_A_193_47#_c_632_n 0.00357711f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A1_c_302_n N_A_193_47#_c_632_n 0.00224159f $X=4.55 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A1_c_299_n N_A_361_47#_c_696_n 3.55919e-19 $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_275 N_VPWR_c_344_n N_A_193_297#_M1000_s 0.00347015f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_276 N_VPWR_c_344_n N_A_193_297#_M1003_d 0.00219239f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_M1001_d N_A_193_297#_c_416_n 0.00413587f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_346_n N_A_193_297#_c_416_n 0.0117417f $X=1.52 $Y=2.34 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_348_n N_A_193_297#_c_416_n 0.00524457f $X=1.355 $Y=2.72 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_350_n N_A_193_297#_c_416_n 7.30294e-19 $X=2.275 $Y=2.72 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_344_n N_A_193_297#_c_416_n 0.0131723f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_282 N_VPWR_M1001_d N_A_193_297#_c_419_n 0.00196174f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_283 N_VPWR_M1001_d N_A_193_297#_c_420_n 0.00182267f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_284 N_VPWR_M1014_d N_A_193_297#_c_415_n 0.00659088f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_344_n N_A_361_297#_M1011_s 0.00385308f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_286 N_VPWR_c_344_n N_A_361_297#_M1007_s 0.00223299f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_350_n N_A_361_297#_c_465_n 0.0133351f $X=2.275 $Y=2.72 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_344_n N_A_361_297#_c_465_n 0.00851918f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_289 N_VPWR_M1014_d N_A_361_297#_c_463_n 0.00499382f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_347_n N_A_361_297#_c_463_n 0.0190091f $X=2.36 $Y=2.34 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_350_n N_A_361_297#_c_463_n 0.0023677f $X=2.275 $Y=2.72 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_353_n N_A_361_297#_c_463_n 0.0029367f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_344_n N_A_361_297#_c_463_n 0.0104748f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_344_n N_Y_M1003_s 0.00211652f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_295 N_VPWR_c_344_n N_Y_M1012_s 0.00250095f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_c_344_n N_Y_M1015_d 0.0037321f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_c_347_n Y 0.0134692f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_298 N_VPWR_c_353_n Y 0.0918031f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_299 N_VPWR_c_344_n Y 0.0708847f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_300 N_VPWR_c_353_n N_Y_c_503_n 0.0126008f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_c_344_n N_Y_c_503_n 0.00848438f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_302 N_A_193_297#_c_415_n N_A_361_297#_M1011_s 0.00369598f $X=3.135 $Y=1.605
+ $X2=-0.19 $Y2=1.305
cc_303 N_A_193_297#_M1003_d N_A_361_297#_c_469_n 0.00328697f $X=3.165 $Y=1.485
+ $X2=0 $Y2=0
cc_304 N_A_193_297#_c_434_n N_A_361_297#_c_469_n 0.0138241f $X=3.3 $Y=1.63 $X2=0
+ $Y2=0
cc_305 N_A_193_297#_c_415_n N_A_361_297#_c_469_n 0.00991501f $X=3.135 $Y=1.605
+ $X2=0 $Y2=0
cc_306 N_A_193_297#_c_416_n N_A_361_297#_c_465_n 0.0145256f $X=1.565 $Y=1.92
+ $X2=0 $Y2=0
cc_307 N_A_193_297#_c_415_n N_A_361_297#_c_465_n 0.0108445f $X=3.135 $Y=1.605
+ $X2=0 $Y2=0
cc_308 N_A_193_297#_c_415_n N_A_361_297#_c_463_n 0.0546462f $X=3.135 $Y=1.605
+ $X2=0 $Y2=0
cc_309 N_A_193_297#_c_415_n N_Y_M1003_s 0.00491846f $X=3.135 $Y=1.605 $X2=0
+ $Y2=0
cc_310 N_A_193_297#_M1003_d Y 0.00325828f $X=3.165 $Y=1.485 $X2=0 $Y2=0
cc_311 N_A_193_297#_c_415_n N_A_193_47#_c_629_n 0.0110369f $X=3.135 $Y=1.605
+ $X2=0 $Y2=0
cc_312 N_A_193_297#_c_415_n N_A_361_47#_c_695_n 6.39736e-19 $X=3.135 $Y=1.605
+ $X2=0 $Y2=0
cc_313 N_A_193_297#_c_415_n N_A_361_47#_c_697_n 0.00600989f $X=3.135 $Y=1.605
+ $X2=0 $Y2=0
cc_314 N_A_361_297#_c_469_n N_Y_M1003_s 0.00156706f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_315 N_A_361_297#_c_464_n N_Y_M1003_s 0.00476462f $X=2.885 $Y=1.96 $X2=0 $Y2=0
cc_316 N_A_361_297#_c_469_n N_Y_M1012_s 0.00948762f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_317 N_A_361_297#_c_469_n Y 0.00693589f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_318 N_A_361_297#_M1007_s Y 0.00336272f $X=4.045 $Y=1.485 $X2=0 $Y2=0
cc_319 N_A_361_297#_c_464_n Y 0.0832255f $X=2.885 $Y=1.96 $X2=0 $Y2=0
cc_320 N_Y_c_499_n N_VGND_c_556_n 0.0100248f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_321 N_Y_c_499_n N_VGND_c_562_n 0.104172f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_322 N_Y_M1002_d N_VGND_c_563_n 0.00173965f $X=2.755 $Y=0.235 $X2=0 $Y2=0
cc_323 N_Y_M1005_d N_VGND_c_563_n 0.00202839f $X=3.585 $Y=0.235 $X2=0 $Y2=0
cc_324 N_Y_M1017_d N_VGND_c_563_n 0.00374041f $X=4.47 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_c_499_n N_VGND_c_563_n 0.0534042f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_326 N_Y_c_499_n N_A_193_47#_M1006_s 0.00329612f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_327 N_Y_M1005_d N_A_193_47#_c_629_n 0.0016435f $X=3.585 $Y=0.235 $X2=0 $Y2=0
cc_328 N_Y_c_499_n N_A_193_47#_c_629_n 0.00972835f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_329 N_Y_M1005_d N_A_193_47#_c_631_n 8.99988e-19 $X=3.585 $Y=0.235 $X2=0 $Y2=0
cc_330 N_Y_c_499_n N_A_193_47#_c_631_n 0.00242641f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_331 N_Y_c_499_n N_A_193_47#_c_632_n 0.0198172f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_332 Y N_A_193_47#_c_632_n 0.00599706f $X=4.75 $Y=1.785 $X2=0 $Y2=0
cc_333 N_Y_c_499_n N_A_361_47#_M1002_s 0.00313852f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_334 N_Y_c_499_n N_A_361_47#_c_696_n 0.0124572f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_335 N_Y_M1002_d N_A_361_47#_c_697_n 0.0032442f $X=2.755 $Y=0.235 $X2=0 $Y2=0
cc_336 N_Y_c_499_n N_A_361_47#_c_697_n 0.0139901f $X=4.805 $Y=0.38 $X2=0 $Y2=0
cc_337 N_VGND_c_563_n N_A_193_47#_M1004_d 0.00375977f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_338 N_VGND_c_563_n N_A_193_47#_M1006_s 0.00217386f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_M1009_s N_A_193_47#_c_629_n 6.81311e-19 $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_340 N_VGND_c_555_n N_A_193_47#_c_629_n 0.0131229f $X=1.52 $Y=0.38 $X2=0 $Y2=0
cc_341 N_VGND_c_556_n N_A_193_47#_c_629_n 8.4091e-19 $X=2.36 $Y=0.38 $X2=0 $Y2=0
cc_342 N_VGND_c_563_n N_A_193_47#_c_629_n 0.114455f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_555_n N_A_193_47#_c_630_n 0.0011828f $X=1.52 $Y=0.38 $X2=0 $Y2=0
cc_344 N_VGND_c_563_n N_A_193_47#_c_630_n 0.0148873f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_345 N_VGND_c_563_n N_A_193_47#_c_631_n 0.0146444f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_555_n N_A_193_47#_c_633_n 0.0118123f $X=1.52 $Y=0.38 $X2=0 $Y2=0
cc_347 N_VGND_c_557_n N_A_193_47#_c_633_n 0.00439594f $X=1.435 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_563_n N_A_193_47#_c_633_n 0.00311968f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_563_n N_A_361_47#_M1008_d 0.00232941f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_350 N_VGND_c_563_n N_A_361_47#_M1002_s 0.00179951f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_559_n N_A_361_47#_c_717_n 0.00899783f $X=2.275 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_563_n N_A_361_47#_c_717_n 0.00300001f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_555_n N_A_361_47#_c_695_n 0.00701214f $X=1.52 $Y=0.38 $X2=0
+ $Y2=0
cc_354 N_VGND_M1013_s N_A_361_47#_c_697_n 0.00319634f $X=2.225 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_VGND_c_556_n N_A_361_47#_c_697_n 0.0102463f $X=2.36 $Y=0.38 $X2=0 $Y2=0
cc_356 N_VGND_c_559_n N_A_361_47#_c_697_n 0.00271438f $X=2.275 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_562_n N_A_361_47#_c_697_n 0.00399916f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_563_n N_A_361_47#_c_697_n 0.0069082f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_359 N_A_193_47#_c_629_n N_A_361_47#_M1008_d 6.95505e-19 $X=3.79 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_360 N_A_193_47#_c_629_n N_A_361_47#_c_695_n 0.00918232f $X=3.79 $Y=0.85 $X2=0
+ $Y2=0
cc_361 N_A_193_47#_c_633_n N_A_361_47#_c_695_n 2.83204e-19 $X=1.1 $Y=0.74 $X2=0
+ $Y2=0
cc_362 N_A_193_47#_c_629_n N_A_361_47#_c_696_n 0.0128528f $X=3.79 $Y=0.85 $X2=0
+ $Y2=0
cc_363 N_A_193_47#_c_631_n N_A_361_47#_c_696_n 0.00122289f $X=3.935 $Y=0.85
+ $X2=0 $Y2=0
cc_364 N_A_193_47#_c_632_n N_A_361_47#_c_696_n 0.00513096f $X=3.935 $Y=0.85
+ $X2=0 $Y2=0
cc_365 N_A_193_47#_c_629_n N_A_361_47#_c_697_n 0.0389669f $X=3.79 $Y=0.85 $X2=0
+ $Y2=0

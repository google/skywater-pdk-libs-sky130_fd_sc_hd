# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlygate4sd1_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.555000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 0.255000 2.700000 0.825000 ;
        RECT 2.440000 1.495000 2.700000 2.465000 ;
        RECT 2.530000 0.825000 2.700000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.550000  0.085000 0.765000 0.545000 ;
        RECT 1.910000  0.085000 2.240000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 0.550000 2.175000 0.765000 2.635000 ;
        RECT 1.910000 1.915000 2.270000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.785000 0.895000 2.005000 ;
      RECT 0.085000 2.005000 0.380000 2.465000 ;
      RECT 0.095000 0.255000 0.380000 0.715000 ;
      RECT 0.095000 0.715000 0.895000 0.885000 ;
      RECT 0.725000 0.885000 0.895000 0.995000 ;
      RECT 0.725000 0.995000 0.980000 1.325000 ;
      RECT 0.725000 1.325000 0.895000 1.785000 ;
      RECT 0.935000 0.255000 1.320000 0.545000 ;
      RECT 0.935000 2.175000 1.320000 2.465000 ;
      RECT 1.150000 0.545000 1.320000 1.075000 ;
      RECT 1.150000 1.075000 1.900000 1.275000 ;
      RECT 1.150000 1.275000 1.320000 2.175000 ;
      RECT 1.515000 0.255000 1.740000 0.735000 ;
      RECT 1.515000 0.735000 2.240000 0.905000 ;
      RECT 1.515000 1.575000 2.240000 1.745000 ;
      RECT 1.515000 1.745000 1.740000 2.430000 ;
      RECT 2.070000 0.905000 2.240000 0.995000 ;
      RECT 2.070000 0.995000 2.360000 1.325000 ;
      RECT 2.070000 1.325000 2.240000 1.575000 ;
  END
END sky130_fd_sc_hd__dlygate4sd1_1

* File: sky130_fd_sc_hd__o22ai_2.spice.pex
* Created: Thu Aug 27 14:37:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O22AI_2%B1 1 3 6 8 10 13 15 21 22
r41 20 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.82 $Y=1.16 $X2=0.91
+ $Y2=1.16
r42 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.82
+ $Y=1.16 $X2=0.82 $Y2=1.16
r43 17 20 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.82 $Y2=1.16
r44 15 21 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.18
+ $X2=0.82 $Y2=1.18
r45 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r46 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r47 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r48 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r49 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r51 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%B2 1 3 6 8 10 13 15 21 22
r48 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.76
+ $Y=1.16 $X2=1.76 $Y2=1.16
r49 19 21 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.75 $Y=1.16 $X2=1.76
+ $Y2=1.16
r50 17 19 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.75 $Y2=1.16
r51 15 22 0.466005 $w=7.68e-07 $l=3e-08 $layer=LI1_cond $X=1.54 $Y=1.19 $X2=1.54
+ $Y2=1.16
r52 11 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r54 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325 $X2=1.33
+ $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995 $X2=1.33
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%A2 1 3 6 8 10 13 15 22
r52 20 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.06 $Y=1.16 $X2=3.15
+ $Y2=1.16
r53 17 20 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.73 $Y=1.16
+ $X2=3.06 $Y2=1.16
r54 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.06
+ $Y=1.16 $X2=3.06 $Y2=1.16
r55 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.16
r56 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.985
r57 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=1.16
r58 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=0.56
r59 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.16
r60 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.73 $Y=1.325 $X2=2.73
+ $Y2=1.985
r61 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=0.995
+ $X2=2.73 $Y2=1.16
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.73 $Y=0.995 $X2=2.73
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%A1 1 3 6 8 10 13 15 21
r42 19 21 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=3.99 $Y=1.16 $X2=4
+ $Y2=1.16
r43 17 19 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.57 $Y=1.16
+ $X2=3.99 $Y2=1.16
r44 15 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4 $Y=1.16
+ $X2=4 $Y2=1.16
r45 11 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.16
r46 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.985
r47 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=0.995
+ $X2=3.99 $Y2=1.16
r48 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.99 $Y=0.995
+ $X2=3.99 $Y2=0.56
r49 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.57 $Y=1.325 $X2=3.57
+ $Y2=1.985
r51 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=0.995
+ $X2=3.57 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.57 $Y=0.995 $X2=3.57
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%A_27_297# 1 2 3 10 12 14 16 17 18 22
r36 20 22 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.96 $Y=2.295
+ $X2=1.96 $Y2=1.96
r37 19 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.38
+ $X2=1.12 $Y2=2.38
r38 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.835 $Y=2.38
+ $X2=1.96 $Y2=2.295
r39 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=2.38
+ $X2=1.245 $Y2=2.38
r40 17 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.295
+ $X2=1.12 $Y2=2.38
r41 16 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=1.54
r42 16 17 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=2.295
r43 15 25 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r44 14 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=1.12 $Y2=1.54
r45 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=0.405 $Y2=1.54
r46 10 25 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r47 10 12 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r48 3 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.96
r49 2 29 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r50 2 27 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r51 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r52 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r55 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r57 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r58 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 28 31 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 27 30 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 25 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r64 25 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 20 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r66 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 16 30 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.655 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.655 $Y=2.72
+ $X2=3.78 $Y2=2.72
r71 15 33 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.905 $Y=2.72
+ $X2=4.37 $Y2=2.72
r72 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.905 $Y=2.72
+ $X2=3.78 $Y2=2.72
r73 11 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=2.635
+ $X2=3.78 $Y2=2.72
r74 11 13 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.78 $Y=2.635
+ $X2=3.78 $Y2=1.96
r75 7 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r76 7 9 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=1.96
r77 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.645
+ $Y=1.485 $X2=3.78 $Y2=1.96
r78 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%Y 1 2 3 4 17 19 26 29 30 33 36 37 41 44
r75 41 44 1.23232 $w=1.78e-07 $l=2e-08 $layer=LI1_cond $X=2.095 $Y=1.535
+ $X2=2.075 $Y2=1.535
r76 37 41 6.62226 $w=1.8e-07 $l=1.22e-07 $layer=LI1_cond $X=2.217 $Y=1.535
+ $X2=2.095 $Y2=1.535
r77 37 44 2.03333 $w=1.78e-07 $l=3.3e-08 $layer=LI1_cond $X=2.042 $Y=1.535
+ $X2=2.075 $Y2=1.535
r78 34 37 20.6138 $w=3.08e-07 $l=5.4e-07 $layer=LI1_cond $X=2.217 $Y=0.905
+ $X2=2.217 $Y2=1.445
r79 31 37 23.2293 $w=1.78e-07 $l=3.77e-07 $layer=LI1_cond $X=1.665 $Y=1.535
+ $X2=2.042 $Y2=1.535
r80 31 33 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=1.535
+ $X2=1.54 $Y2=1.535
r81 28 30 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=0.775
+ $X2=1.705 $Y2=0.775
r82 28 29 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=0.775
+ $X2=1.375 $Y2=0.775
r83 26 29 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=0.865 $Y=0.815
+ $X2=1.375 $Y2=0.815
r84 24 26 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=0.775
+ $X2=0.865 $Y2=0.775
r85 20 37 6.62226 $w=1.8e-07 $l=1.23e-07 $layer=LI1_cond $X=2.34 $Y=1.535
+ $X2=2.217 $Y2=1.535
r86 19 36 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.815 $Y=1.535
+ $X2=2.94 $Y2=1.535
r87 19 20 29.2677 $w=1.78e-07 $l=4.75e-07 $layer=LI1_cond $X=2.815 $Y=1.535
+ $X2=2.34 $Y2=1.535
r88 17 34 7.02594 $w=1.8e-07 $l=1.60823e-07 $layer=LI1_cond $X=2.095 $Y=0.815
+ $X2=2.217 $Y2=0.905
r89 17 30 24.0303 $w=1.78e-07 $l=3.9e-07 $layer=LI1_cond $X=2.095 $Y=0.815
+ $X2=1.705 $Y2=0.815
r90 4 36 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.485 $X2=2.94 $Y2=1.62
r91 3 33 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.62
r92 2 28 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.73
r93 1 24 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%A_475_297# 1 2 3 12 14 15 16 17 18 20 22
r36 20 29 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.202 $Y=1.625
+ $X2=4.202 $Y2=1.54
r37 20 22 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=4.202 $Y=1.625
+ $X2=4.202 $Y2=2.3
r38 19 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=1.54
+ $X2=3.36 $Y2=1.54
r39 18 29 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.075 $Y=1.54
+ $X2=4.202 $Y2=1.54
r40 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.075 $Y=1.54
+ $X2=3.485 $Y2=1.54
r41 17 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=2.295
+ $X2=3.36 $Y2=2.38
r42 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=1.625
+ $X2=3.36 $Y2=1.54
r43 16 17 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.36 $Y=1.625
+ $X2=3.36 $Y2=2.295
r44 14 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=2.38
+ $X2=3.36 $Y2=2.38
r45 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.235 $Y=2.38
+ $X2=2.645 $Y2=2.38
r46 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.52 $Y=2.295
+ $X2=2.645 $Y2=2.38
r47 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.52 $Y=2.295
+ $X2=2.52 $Y2=1.96
r48 3 29 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.485 $X2=4.2 $Y2=1.62
r49 3 22 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.485 $X2=4.2 $Y2=2.3
r50 2 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=2.3
r51 2 25 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=1.62
r52 1 12 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.375
+ $Y=1.485 $X2=2.52 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%A_27_47# 1 2 3 4 5 16 18 20 24 25 26 27 30
+ 32 36 42
r80 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.2 $Y=0.725 $X2=4.2
+ $Y2=0.39
r81 33 42 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=0.815
+ $X2=3.36 $Y2=0.815
r82 32 34 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.035 $Y=0.815
+ $X2=4.2 $Y2=0.725
r83 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.035 $Y=0.815
+ $X2=3.525 $Y2=0.815
r84 28 42 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.36 $Y=0.725 $X2=3.36
+ $Y2=0.815
r85 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.36 $Y=0.725
+ $X2=3.36 $Y2=0.39
r86 26 42 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=0.815
+ $X2=3.36 $Y2=0.815
r87 26 27 31.7323 $w=1.78e-07 $l=5.15e-07 $layer=LI1_cond $X=3.195 $Y=0.815
+ $X2=2.68 $Y2=0.815
r88 25 27 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.595 $Y=0.725
+ $X2=2.68 $Y2=0.815
r89 24 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.475
+ $X2=2.595 $Y2=0.39
r90 24 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.595 $Y=0.475
+ $X2=2.595 $Y2=0.725
r91 21 39 4.53113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.365 $Y=0.39
+ $X2=0.227 $Y2=0.39
r92 21 23 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.365 $Y=0.39
+ $X2=1.12 $Y2=0.39
r93 20 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=0.39
+ $X2=2.595 $Y2=0.39
r94 20 23 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=2.51 $Y=0.39
+ $X2=1.12 $Y2=0.39
r95 16 39 2.79091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.227 $Y=0.475
+ $X2=0.227 $Y2=0.39
r96 16 18 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=0.227 $Y=0.475
+ $X2=0.227 $Y2=0.73
r97 5 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.065
+ $Y=0.235 $X2=4.2 $Y2=0.39
r98 4 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.225
+ $Y=0.235 $X2=3.36 $Y2=0.39
r99 3 41 91 $w=1.7e-07 $l=7.63577e-07 $layer=licon1_NDIFF $count=2 $X=1.825
+ $Y=0.235 $X2=2.515 $Y2=0.39
r100 2 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r101 1 39 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
r102 1 18 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_2%VGND 1 2 9 13 16 17 19 20 21 34 35
r55 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r56 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r57 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r58 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r59 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r60 24 28 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r61 21 29 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r62 21 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r63 19 31 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.45
+ $Y2=0
r64 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.78
+ $Y2=0
r65 18 34 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.865 $Y=0 $X2=4.37
+ $Y2=0
r66 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=0 $X2=3.78
+ $Y2=0
r67 16 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.855 $Y=0 $X2=2.53
+ $Y2=0
r68 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0 $X2=2.94
+ $Y2=0
r69 15 31 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=3.45
+ $Y2=0
r70 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.94
+ $Y2=0
r71 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0
r72 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0.39
r73 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085 $X2=2.94
+ $Y2=0
r74 7 9 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.39
r75 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.235 $X2=3.78 $Y2=0.39
r76 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.235 $X2=2.94 $Y2=0.39
.ends


* NGSPICE file created from sky130_fd_sc_hd__buf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
M1000 VPWR a_27_47# X VPB phighvt w=1e+06u l=150000u
+  ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u
M1001 VPWR A a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1002 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=3.6625e+11p pd=3.78e+06u as=1.755e+11p ps=1.84e+06u
M1004 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1005 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


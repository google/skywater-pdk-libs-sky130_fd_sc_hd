* File: sky130_fd_sc_hd__a32oi_1.pex.spice
* Created: Tue Sep  1 18:55:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A32OI_1%B2 1 3 6 8 14
c26 6 0 1.78086e-19 $X=0.47 $Y=1.985
r27 11 14 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r29 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r31 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%B1 3 6 10 11 13 16
c44 16 0 1.95172e-19 $X=0.915 $Y=0.995
c45 13 0 1.78086e-19 $X=1.16 $Y=1.53
r46 13 18 12.8421 $w=1.88e-07 $l=2.2e-07 $layer=LI1_cond $X=1.16 $Y=1.52
+ $X2=0.94 $Y2=1.52
r47 11 17 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=0.915 $Y2=1.325
r48 11 16 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=0.915 $Y2=0.995
r49 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r50 8 18 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.94 $Y=1.425 $X2=0.94
+ $Y2=1.52
r51 8 10 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.94 $Y=1.425
+ $X2=0.94 $Y2=1.16
r52 6 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.985
+ $X2=0.89 $Y2=1.325
r53 3 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.85 $Y=0.56 $X2=0.85
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%A1 3 6 9 11 12 15 18
c45 18 0 3.14664e-20 $X=1.42 $Y=0.995
c46 15 0 1.95172e-19 $X=1.62 $Y=0.51
r47 15 23 11.3385 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.555 $Y=0.51
+ $X2=1.555 $Y2=0.765
r48 12 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.16
+ $X2=1.42 $Y2=1.325
r49 12 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.16
+ $X2=1.42 $Y2=0.995
r50 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.16 $X2=1.42 $Y2=1.16
r51 9 11 0.384081 $w=1.9e-07 $l=1.23693e-07 $layer=LI1_cond $X=1.5 $Y=1.075
+ $X2=1.42 $Y2=1.165
r52 9 23 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=1.5 $Y=1.075 $X2=1.5
+ $Y2=0.765
r53 6 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.47 $Y=1.985
+ $X2=1.47 $Y2=1.325
r54 3 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.47 $Y=0.56 $X2=1.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%A2 3 6 7 8 10 11 12 13 18
c40 11 0 3.14664e-20 $X=2.08 $Y=0.51
r41 20 28 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=0.995
+ $X2=2.065 $Y2=1.16
r42 19 28 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=1.16
+ $X2=2.065 $Y2=1.16
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.9
+ $Y=1.16 $X2=1.9 $Y2=1.16
r44 13 28 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.08 $Y=1.16
+ $X2=2.065 $Y2=1.16
r45 12 20 8.04091 $w=1.98e-07 $l=1.45e-07 $layer=LI1_cond $X=2.065 $Y=0.85
+ $X2=2.065 $Y2=0.995
r46 11 12 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=2.065 $Y=0.51
+ $X2=2.065 $Y2=0.85
r47 9 18 25.55 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=1.9 $Y=1.275 $X2=1.9
+ $Y2=1.16
r48 9 10 36.4065 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.9 $Y=1.275 $X2=1.9
+ $Y2=1.41
r49 7 18 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=1.9 $Y=1.095 $X2=1.9
+ $Y2=1.16
r50 7 8 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.9 $Y=1.095 $X2=1.9
+ $Y2=0.96
r51 6 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.89 $Y=1.985
+ $X2=1.89 $Y2=1.41
r52 3 8 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.84 $Y=0.56 $X2=1.84
+ $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%A3 3 6 7 10 12 13 17
r23 10 13 57.4123 $w=4.4e-07 $l=2.5e-07 $layer=POLY_cond $X=2.465 $Y=1.16
+ $X2=2.465 $Y2=1.41
r24 10 12 51.0924 $w=4.4e-07 $l=2e-07 $layer=POLY_cond $X=2.465 $Y=1.16
+ $X2=2.465 $Y2=0.96
r25 7 17 2.23053 $w=3.08e-07 $l=6e-08 $layer=LI1_cond $X=2.51 $Y=1.17 $X2=2.57
+ $Y2=1.17
r26 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.16 $X2=2.51 $Y2=1.16
r27 6 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.32 $Y=1.985
+ $X2=2.32 $Y2=1.41
r28 3 12 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.32 $Y=0.56 $X2=2.32
+ $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%A_27_297# 1 2 3 10 12 14 16 17 18 29
r38 19 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.87
+ $X2=1.22 $Y2=1.87
r39 18 29 3.40825 $w=1.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.015 $Y=1.87
+ $X2=2.1 $Y2=1.85
r40 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.015 $Y=1.87
+ $X2=1.345 $Y2=1.87
r41 17 27 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=2.255
+ $X2=1.22 $Y2=2.36
r42 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.955
+ $X2=1.22 $Y2=1.87
r43 16 17 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=1.22 $Y=1.955 $X2=1.22
+ $Y2=2.255
r44 15 23 3.8266 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=2.36
+ $X2=0.215 $Y2=2.36
r45 14 27 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=2.36
+ $X2=1.22 $Y2=2.36
r46 14 15 39.6104 $w=2.08e-07 $l=7.5e-07 $layer=LI1_cond $X=1.095 $Y=2.36
+ $X2=0.345 $Y2=2.36
r47 10 23 3.09071 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=0.215 $Y=2.255
+ $X2=0.215 $Y2=2.36
r48 10 12 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=2.255
+ $X2=0.215 $Y2=2
r49 3 29 300 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=1.485 $X2=2.1 $Y2=1.91
r50 2 27 600 $w=1.7e-07 $l=9.51131e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.26 $Y2=2.3
r51 2 25 600 $w=1.7e-07 $l=5.11664e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.26 $Y2=1.87
r52 1 23 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r53 1 12 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%Y 1 2 7 8 11 14
r38 14 19 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=0.68 $Y=1.935 $X2=0.6
+ $Y2=1.935
r39 14 19 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.6 $Y=1.785 $X2=0.6
+ $Y2=1.935
r40 13 14 44.6803 $w=2.58e-07 $l=9.8e-07 $layer=LI1_cond $X=0.6 $Y=0.805 $X2=0.6
+ $Y2=1.785
r41 9 11 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=1.04 $Y=0.635
+ $X2=1.04 $Y2=0.53
r42 8 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=0.72
+ $X2=0.6 $Y2=0.805
r43 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.915 $Y=0.72
+ $X2=1.04 $Y2=0.635
r44 7 8 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.915 $Y=0.72
+ $X2=0.685 $Y2=0.72
r45 2 14 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
r46 1 11 182 $w=1.7e-07 $l=3.64349e-07 $layer=licon1_NDIFF $count=1 $X=0.925
+ $Y=0.235 $X2=1.08 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%VPWR 1 2 9 13 17 19 24 31 32 35 38
r41 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r42 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r43 32 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 29 38 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.525 $Y2=2.72
r46 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.695 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 28 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 28 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 25 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.68 $Y2=2.72
r51 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 24 38 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.525 $Y2=2.72
r53 24 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 19 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.68 $Y2=2.72
r55 19 21 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 17 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 17 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 13 16 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=2.525 $Y=1.66
+ $X2=2.525 $Y2=2.34
r59 11 38 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=2.635
+ $X2=2.525 $Y2=2.72
r60 11 16 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.525 $Y=2.635
+ $X2=2.525 $Y2=2.34
r61 7 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.635
+ $X2=1.68 $Y2=2.72
r62 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.68 $Y=2.635
+ $X2=1.68 $Y2=2.3
r63 2 16 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.485 $X2=2.53 $Y2=2.34
r64 2 13 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.485 $X2=2.53 $Y2=1.66
r65 1 9 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.68 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_1%VGND 1 2 7 9 13 15 17 27 28 34
r42 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r43 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r44 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r45 25 34 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.525
+ $Y2=0
r46 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.99
+ $Y2=0
r47 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r48 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r49 21 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r50 20 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r51 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 18 31 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r53 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r54 17 34 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.525
+ $Y2=0
r55 17 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.07
+ $Y2=0
r56 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r57 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 11 34 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0
r59 11 13 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0.38
r60 7 31 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r61 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r62 2 13 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.395
+ $Y=0.235 $X2=2.53 $Y2=0.38
r63 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__nand2_1.pex.spice
* Created: Tue Sep  1 19:15:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND2_1%B 1 3 6 8 14
r23 11 14 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.265 $Y=1.16
+ $X2=0.49 $Y2=1.16
r24 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.265
+ $Y=1.16 $X2=0.265 $Y2=1.16
r25 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r26 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r27 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r28 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_1%A 1 3 6 8 13
r23 10 13 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.105 $Y2=1.16
r24 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.16 $X2=1.105 $Y2=1.16
r25 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r26 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325 $X2=0.91
+ $Y2=1.985
r27 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r28 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995 $X2=0.91
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_1%VPWR 1 2 7 9 13 15 19 21 31
r22 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r23 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r25 22 27 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r26 22 24 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.69 $Y2=2.72
r27 21 30 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.207 $Y2=2.72
r28 21 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r29 19 25 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.69 $Y2=2.72
r30 19 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r31 15 18 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.165 $Y=1.66
+ $X2=1.165 $Y2=2.34
r32 13 30 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=1.165 $Y=2.635
+ $X2=1.207 $Y2=2.72
r33 13 18 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.165 $Y=2.635
+ $X2=1.165 $Y2=2.34
r34 9 12 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.225 $Y=1.66
+ $X2=0.225 $Y2=2.34
r35 7 27 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.182 $Y2=2.72
r36 7 12 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=2.635
+ $X2=0.225 $Y2=2.34
r37 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.34
r38 2 15 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.66
r39 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=2.34
r40 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_1%Y 1 2 7 9 15 17 31
c23 7 0 1.13229e-19 $X=0.7 $Y=1.65
r24 15 31 8.25864 $w=6.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.685 $Y=0.57
+ $X2=1.12 $Y2=0.57
r25 15 22 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=0.685 $Y=0.57
+ $X2=0.685 $Y2=0.885
r26 15 17 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.685 $Y=0.91
+ $X2=0.685 $Y2=1.19
r27 15 22 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.685 $Y=0.91
+ $X2=0.685 $Y2=0.885
r28 14 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.685 $Y=1.485
+ $X2=0.685 $Y2=1.19
r29 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.7 $Y=1.66 $X2=0.7
+ $Y2=2.34
r30 7 14 7.25185 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=1.65 $X2=0.7
+ $Y2=1.485
r31 7 9 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.7 $Y=1.65 $X2=0.7
+ $Y2=1.66
r32 2 11 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2.34
r33 2 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.66
r34 1 31 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_1%VGND 1 4 6 8 12 13 21
r16 16 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r17 13 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.23
+ $Y2=0
r18 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r19 10 16 4.61546 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r20 10 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=1.15
+ $Y2=0
r21 8 21 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r22 4 16 2.98373 $w=3.1e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.197 $Y2=0
r23 4 6 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r24 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends


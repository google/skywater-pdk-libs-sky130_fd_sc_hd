* File: sky130_fd_sc_hd__mux4_2.spice.SKY130_FD_SC_HD__MUX4_2.pxi
* Created: Thu Aug 27 14:28:23 2020
* 
x_PM_SKY130_FD_SC_HD__MUX4_2%S0 N_S0_M1025_g N_S0_M1016_g N_S0_c_175_n
+ N_S0_M1023_g N_S0_c_176_n N_S0_M1002_g N_S0_M1015_g N_S0_c_179_n N_S0_c_180_n
+ N_S0_M1018_g S0 S0 N_S0_c_193_n N_S0_c_194_n N_S0_c_195_n N_S0_c_196_n
+ N_S0_c_182_n N_S0_c_198_n N_S0_c_199_n N_S0_c_183_n N_S0_c_184_n
+ PM_SKY130_FD_SC_HD__MUX4_2%S0
x_PM_SKY130_FD_SC_HD__MUX4_2%A2 N_A2_M1013_g N_A2_M1000_g N_A2_c_378_n
+ N_A2_c_385_n A2 A2 N_A2_c_381_n N_A2_c_382_n PM_SKY130_FD_SC_HD__MUX4_2%A2
x_PM_SKY130_FD_SC_HD__MUX4_2%A_27_47# N_A_27_47#_M1025_s N_A_27_47#_M1016_s
+ N_A_27_47#_c_442_n N_A_27_47#_M1004_g N_A_27_47#_M1017_g N_A_27_47#_M1022_g
+ N_A_27_47#_c_443_n N_A_27_47#_M1005_g N_A_27_47#_c_667_p N_A_27_47#_c_602_p
+ N_A_27_47#_c_444_n N_A_27_47#_c_455_n N_A_27_47#_c_483_n N_A_27_47#_c_445_n
+ N_A_27_47#_c_446_n N_A_27_47#_c_447_n N_A_27_47#_c_448_n N_A_27_47#_c_456_n
+ N_A_27_47#_c_457_n N_A_27_47#_c_458_n N_A_27_47#_c_459_n N_A_27_47#_c_460_n
+ N_A_27_47#_c_461_n N_A_27_47#_c_449_n N_A_27_47#_c_450_n N_A_27_47#_c_451_n
+ PM_SKY130_FD_SC_HD__MUX4_2%A_27_47#
x_PM_SKY130_FD_SC_HD__MUX4_2%A3 N_A3_M1007_g N_A3_c_684_n N_A3_c_690_n
+ N_A3_M1003_g N_A3_c_691_n A3 A3 N_A3_c_687_n N_A3_c_688_n
+ PM_SKY130_FD_SC_HD__MUX4_2%A3
x_PM_SKY130_FD_SC_HD__MUX4_2%S1 N_S1_c_743_n N_S1_M1026_g N_S1_c_745_n
+ N_S1_M1014_g N_S1_c_750_n N_S1_c_751_n N_S1_c_746_n N_S1_c_747_n N_S1_M1019_g
+ N_S1_M1008_g S1 S1 PM_SKY130_FD_SC_HD__MUX4_2%S1
x_PM_SKY130_FD_SC_HD__MUX4_2%A_600_345# N_A_600_345#_M1014_d
+ N_A_600_345#_M1026_d N_A_600_345#_M1020_g N_A_600_345#_c_829_n
+ N_A_600_345#_M1012_g N_A_600_345#_c_831_n N_A_600_345#_c_832_n
+ N_A_600_345#_c_833_n N_A_600_345#_c_834_n N_A_600_345#_c_835_n
+ PM_SKY130_FD_SC_HD__MUX4_2%A_600_345#
x_PM_SKY130_FD_SC_HD__MUX4_2%A1 N_A1_M1001_g N_A1_M1027_g A1 A1 N_A1_c_900_n
+ PM_SKY130_FD_SC_HD__MUX4_2%A1
x_PM_SKY130_FD_SC_HD__MUX4_2%A0 N_A0_M1024_g N_A0_M1021_g N_A0_c_939_n
+ N_A0_c_940_n A0 A0 PM_SKY130_FD_SC_HD__MUX4_2%A0
x_PM_SKY130_FD_SC_HD__MUX4_2%A_788_316# N_A_788_316#_M1019_d
+ N_A_788_316#_M1020_d N_A_788_316#_c_987_n N_A_788_316#_M1009_g
+ N_A_788_316#_M1006_g N_A_788_316#_c_988_n N_A_788_316#_M1010_g
+ N_A_788_316#_M1011_g N_A_788_316#_c_989_n N_A_788_316#_c_995_n
+ N_A_788_316#_c_996_n N_A_788_316#_c_997_n N_A_788_316#_c_998_n
+ N_A_788_316#_c_999_n N_A_788_316#_c_990_n N_A_788_316#_c_1001_n
+ N_A_788_316#_c_1002_n N_A_788_316#_c_1003_n N_A_788_316#_c_1018_n
+ N_A_788_316#_c_991_n N_A_788_316#_c_1019_n
+ PM_SKY130_FD_SC_HD__MUX4_2%A_788_316#
x_PM_SKY130_FD_SC_HD__MUX4_2%VPWR N_VPWR_M1016_d N_VPWR_M1003_d N_VPWR_M1001_s
+ N_VPWR_M1021_d N_VPWR_M1011_d N_VPWR_c_1136_n N_VPWR_c_1137_n N_VPWR_c_1138_n
+ N_VPWR_c_1139_n N_VPWR_c_1140_n N_VPWR_c_1141_n N_VPWR_c_1142_n
+ N_VPWR_c_1143_n N_VPWR_c_1144_n N_VPWR_c_1145_n VPWR N_VPWR_c_1146_n
+ N_VPWR_c_1147_n N_VPWR_c_1148_n N_VPWR_c_1149_n N_VPWR_c_1150_n
+ N_VPWR_c_1135_n PM_SKY130_FD_SC_HD__MUX4_2%VPWR
x_PM_SKY130_FD_SC_HD__MUX4_2%A_288_47# N_A_288_47#_M1004_d N_A_288_47#_M1019_s
+ N_A_288_47#_M1023_d N_A_288_47#_M1020_s N_A_288_47#_c_1279_n
+ N_A_288_47#_c_1280_n N_A_288_47#_c_1267_n N_A_288_47#_c_1271_n
+ N_A_288_47#_c_1283_n N_A_288_47#_c_1272_n N_A_288_47#_c_1273_n
+ N_A_288_47#_c_1268_n N_A_288_47#_c_1269_n N_A_288_47#_c_1270_n
+ N_A_288_47#_c_1276_n N_A_288_47#_c_1316_n N_A_288_47#_c_1277_n
+ PM_SKY130_FD_SC_HD__MUX4_2%A_288_47#
x_PM_SKY130_FD_SC_HD__MUX4_2%A_872_316# N_A_872_316#_M1012_d
+ N_A_872_316#_M1015_d N_A_872_316#_M1008_d N_A_872_316#_M1022_d
+ N_A_872_316#_c_1405_n N_A_872_316#_c_1408_n N_A_872_316#_c_1406_n
+ N_A_872_316#_c_1410_n N_A_872_316#_c_1482_p N_A_872_316#_c_1417_n
+ N_A_872_316#_c_1455_n N_A_872_316#_c_1418_n N_A_872_316#_c_1456_n
+ N_A_872_316#_c_1411_n PM_SKY130_FD_SC_HD__MUX4_2%A_872_316#
x_PM_SKY130_FD_SC_HD__MUX4_2%X N_X_M1009_s N_X_M1006_s N_X_c_1505_n N_X_c_1503_n
+ X X X X PM_SKY130_FD_SC_HD__MUX4_2%X
x_PM_SKY130_FD_SC_HD__MUX4_2%VGND N_VGND_M1025_d N_VGND_M1007_d N_VGND_M1027_s
+ N_VGND_M1024_d N_VGND_M1010_d N_VGND_c_1534_n N_VGND_c_1535_n N_VGND_c_1536_n
+ N_VGND_c_1537_n N_VGND_c_1538_n N_VGND_c_1539_n VGND N_VGND_c_1540_n
+ N_VGND_c_1541_n N_VGND_c_1542_n N_VGND_c_1543_n N_VGND_c_1544_n
+ N_VGND_c_1545_n N_VGND_c_1546_n N_VGND_c_1547_n N_VGND_c_1548_n
+ N_VGND_c_1549_n PM_SKY130_FD_SC_HD__MUX4_2%VGND
cc_1 VNB N_S0_M1025_g 0.0351649f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_S0_c_175_n 0.00818586f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.615
cc_3 VNB N_S0_c_176_n 0.0148947f $X=-0.19 $Y=-0.24 $X2=1.835 $Y2=1.32
cc_4 VNB N_S0_M1002_g 0.0435516f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=0.415
cc_5 VNB N_S0_M1015_g 0.0457451f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=0.415
cc_6 VNB N_S0_c_179_n 0.0107197f $X=-0.19 $Y=-0.24 $X2=6.245 $Y2=1.32
cc_7 VNB N_S0_c_180_n 0.00197903f $X=-0.19 $Y=-0.24 $X2=5.855 $Y2=1.32
cc_8 VNB S0 0.00322235f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_9 VNB N_S0_c_182_n 0.00218622f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.53
cc_10 VNB N_S0_c_183_n 0.043471f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_11 VNB N_S0_c_184_n 0.0110759f $X=-0.19 $Y=-0.24 $X2=6.38 $Y2=1.32
cc_12 VNB N_A2_c_378_n 0.0128209f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.275
cc_13 VNB A2 0.00268106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB A2 0.00423678f $X=-0.19 $Y=-0.24 $X2=1.835 $Y2=1.32
cc_15 VNB N_A2_c_381_n 0.0274502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_382_n 0.0166423f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=0.415
cc_17 VNB N_A_27_47#_c_442_n 0.0180022f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_18 VNB N_A_27_47#_c_443_n 0.0180623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_444_n 0.00400149f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_20 VNB N_A_27_47#_c_445_n 0.00884926f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.53
cc_21 VNB N_A_27_47#_c_446_n 0.0309921f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.53
cc_22 VNB N_A_27_47#_c_447_n 0.0030285f $X=-0.19 $Y=-0.24 $X2=6.21 $Y2=1.53
cc_23 VNB N_A_27_47#_c_448_n 0.00540154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_449_n 0.00905904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_450_n 0.032928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_451_n 0.00415242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A3_c_684_n 0.0112092f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_28 VNB A3 0.00653171f $X=-0.19 $Y=-0.24 $X2=1.835 $Y2=1.32
cc_29 VNB A3 0.00177632f $X=-0.19 $Y=-0.24 $X2=1.44 $Y2=1.32
cc_30 VNB N_A3_c_687_n 0.0241632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A3_c_688_n 0.0172648f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=0.415
cc_32 VNB N_S1_c_743_n 0.0288831f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_33 VNB N_S1_M1026_g 0.00924061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_S1_c_745_n 0.0184815f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_35 VNB N_S1_c_746_n 0.0513215f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.275
cc_36 VNB N_S1_c_747_n 0.0179541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB S1 0.00677138f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=1.245
cc_38 VNB N_A_600_345#_c_829_n 0.0321009f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.275
cc_39 VNB N_A_600_345#_M1012_g 0.0381718f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=1.245
cc_40 VNB N_A_600_345#_c_831_n 0.0234246f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=0.415
cc_41 VNB N_A_600_345#_c_832_n 0.00740591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_600_345#_c_833_n 0.00626684f $X=-0.19 $Y=-0.24 $X2=5.78 $Y2=0.415
cc_43 VNB N_A_600_345#_c_834_n 0.00114392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_600_345#_c_835_n 0.00367345f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_45 VNB N_A1_M1027_g 0.0386874f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_46 VNB A1 0.0121957f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.615
cc_47 VNB N_A1_c_900_n 0.0307838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A0_M1024_g 0.0291922f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_49 VNB N_A0_c_939_n 0.0139105f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.615
cc_50 VNB N_A0_c_940_n 0.0257079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB A0 0.00260222f $X=-0.19 $Y=-0.24 $X2=1.835 $Y2=1.32
cc_52 VNB N_A_788_316#_c_987_n 0.0166938f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_53 VNB N_A_788_316#_c_988_n 0.0215f $X=-0.19 $Y=-0.24 $X2=1.44 $Y2=1.32
cc_54 VNB N_A_788_316#_c_989_n 0.00865735f $X=-0.19 $Y=-0.24 $X2=6.245 $Y2=1.32
cc_55 VNB N_A_788_316#_c_990_n 0.00267682f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.53
cc_56 VNB N_A_788_316#_c_991_n 0.0427465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_1135_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_288_47#_c_1267_n 0.0043778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_288_47#_c_1268_n 0.00668781f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.53
cc_60 VNB N_A_288_47#_c_1269_n 0.00364533f $X=-0.19 $Y=-0.24 $X2=6.065 $Y2=1.53
cc_61 VNB N_A_288_47#_c_1270_n 7.8042e-19 $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.53
cc_62 VNB N_A_872_316#_c_1405_n 0.0132662f $X=-0.19 $Y=-0.24 $X2=1.44 $Y2=1.32
cc_63 VNB N_A_872_316#_c_1406_n 0.0123594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_X_c_1503_n 0.00108687f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.275
cc_65 VNB N_VGND_c_1534_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1535_n 0.00290102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1536_n 0.010332f $X=-0.19 $Y=-0.24 $X2=6.32 $Y2=2.275
cc_68 VNB N_VGND_c_1537_n 0.00229342f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_69 VNB N_VGND_c_1538_n 0.00997672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1539_n 0.033359f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=1.53
cc_71 VNB N_VGND_c_1540_n 0.0153519f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.53
cc_72 VNB N_VGND_c_1541_n 0.0418082f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.53
cc_73 VNB N_VGND_c_1542_n 0.0541513f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_74 VNB N_VGND_c_1543_n 0.0497635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1544_n 0.0171843f $X=-0.19 $Y=-0.24 $X2=6.38 $Y2=1.41
cc_76 VNB N_VGND_c_1545_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_77 VNB N_VGND_c_1546_n 0.00516502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1547_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1548_n 0.00356594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1549_n 0.40003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VPB N_S0_M1016_g 0.0433005f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_82 VPB N_S0_c_175_n 0.0227389f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.615
cc_83 VPB N_S0_M1023_g 0.0330551f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=2.275
cc_84 VPB N_S0_c_176_n 0.0167376f $X=-0.19 $Y=1.305 $X2=1.835 $Y2=1.32
cc_85 VPB N_S0_c_179_n 0.01241f $X=-0.19 $Y=1.305 $X2=6.245 $Y2=1.32
cc_86 VPB N_S0_c_180_n 0.00449122f $X=-0.19 $Y=1.305 $X2=5.855 $Y2=1.32
cc_87 VPB N_S0_M1018_g 0.0376059f $X=-0.19 $Y=1.305 $X2=6.32 $Y2=2.275
cc_88 VPB S0 0.0154537f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_89 VPB N_S0_c_193_n 0.00677823f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.53
cc_90 VPB N_S0_c_194_n 0.0143774f $X=-0.19 $Y=1.305 $X2=0.375 $Y2=1.53
cc_91 VPB N_S0_c_195_n 0.043526f $X=-0.19 $Y=1.305 $X2=6.065 $Y2=1.53
cc_92 VPB N_S0_c_196_n 0.00423102f $X=-0.19 $Y=1.305 $X2=1.295 $Y2=1.53
cc_93 VPB N_S0_c_182_n 0.00302522f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.53
cc_94 VPB N_S0_c_198_n 0.00246888f $X=-0.19 $Y=1.305 $X2=6.21 $Y2=1.53
cc_95 VPB N_S0_c_199_n 0.00362396f $X=-0.19 $Y=1.305 $X2=6.21 $Y2=1.53
cc_96 VPB N_S0_c_183_n 0.0111047f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_97 VPB N_S0_c_184_n 0.0215929f $X=-0.19 $Y=1.305 $X2=6.38 $Y2=1.32
cc_98 VPB N_A2_M1000_g 0.0170662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A2_c_378_n 0.0174405f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=2.275
cc_100 VPB N_A2_c_385_n 0.0024879f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=2.275
cc_101 VPB N_A_27_47#_M1017_g 0.02251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_47#_M1022_g 0.0226804f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=0.415
cc_103 VPB N_A_27_47#_c_444_n 0.00369148f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_104 VPB N_A_27_47#_c_455_n 0.00645667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_47#_c_456_n 0.00858126f $X=-0.19 $Y=1.305 $X2=1.305 $Y2=1.32
cc_106 VPB N_A_27_47#_c_457_n 0.0027247f $X=-0.19 $Y=1.305 $X2=1.305 $Y2=1.45
cc_107 VPB N_A_27_47#_c_458_n 0.00188091f $X=-0.19 $Y=1.305 $X2=6.38 $Y2=1.41
cc_108 VPB N_A_27_47#_c_459_n 0.0277359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_27_47#_c_460_n 0.00526335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_27_47#_c_461_n 0.0275765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_27_47#_c_449_n 0.00473799f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_27_47#_c_451_n 0.00201397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A3_c_684_n 0.0117778f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_114 VPB N_A3_c_690_n 0.0237103f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_115 VPB N_A3_c_691_n 0.0181615f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=2.275
cc_116 VPB A3 9.23002e-19 $X=-0.19 $Y=1.305 $X2=1.44 $Y2=1.32
cc_117 VPB N_S1_M1026_g 0.0332464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_S1_c_750_n 0.096695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_S1_c_751_n 0.00958866f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.615
cc_120 VPB N_S1_M1008_g 0.0364991f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=0.415
cc_121 VPB S1 0.00178367f $X=-0.19 $Y=1.305 $X2=5.78 $Y2=1.245
cc_122 VPB N_A_600_345#_M1020_g 0.0238152f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.615
cc_123 VPB N_A_600_345#_c_831_n 0.0207153f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=0.415
cc_124 VPB N_A_600_345#_c_832_n 0.00224568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_600_345#_c_834_n 0.0131964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A1_M1001_g 0.0458456f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_127 VPB A1 0.0035535f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.615
cc_128 VPB N_A1_c_900_n 0.0163508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A0_M1021_g 0.0377501f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_130 VPB N_A0_c_939_n 0.00286793f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.615
cc_131 VPB N_A0_c_940_n 0.00429793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_788_316#_M1006_g 0.0185888f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_788_316#_M1011_g 0.0252934f $X=-0.19 $Y=1.305 $X2=5.78 $Y2=1.245
cc_134 VPB N_A_788_316#_c_989_n 0.00438187f $X=-0.19 $Y=1.305 $X2=6.245 $Y2=1.32
cc_135 VPB N_A_788_316#_c_995_n 0.00187498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_788_316#_c_996_n 0.00313433f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_137 VPB N_A_788_316#_c_997_n 0.00173284f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_138 VPB N_A_788_316#_c_998_n 0.00185715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_788_316#_c_999_n 0.00258066f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.53
cc_140 VPB N_A_788_316#_c_990_n 3.66738e-19 $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.53
cc_141 VPB N_A_788_316#_c_1001_n 0.00232217f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_788_316#_c_1002_n 0.00114749f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.53
cc_143 VPB N_A_788_316#_c_1003_n 0.00329434f $X=-0.19 $Y=1.305 $X2=6.21 $Y2=1.53
cc_144 VPB N_A_788_316#_c_991_n 0.005583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_1136_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_1137_n 0.00835502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_1138_n 0.013457f $X=-0.19 $Y=1.305 $X2=6.32 $Y2=2.275
cc_148 VPB N_VPWR_c_1139_n 0.00468459f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_149 VPB N_VPWR_c_1140_n 0.0100141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_1141_n 0.0427673f $X=-0.19 $Y=1.305 $X2=0.375 $Y2=1.53
cc_151 VPB N_VPWR_c_1142_n 0.0489906f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.53
cc_152 VPB N_VPWR_c_1143_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_1144_n 0.0519215f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.53
cc_154 VPB N_VPWR_c_1145_n 0.00324402f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.53
cc_155 VPB N_VPWR_c_1146_n 0.0153943f $X=-0.19 $Y=1.305 $X2=6.21 $Y2=1.53
cc_156 VPB N_VPWR_c_1147_n 0.0543338f $X=-0.19 $Y=1.305 $X2=6.38 $Y2=1.32
cc_157 VPB N_VPWR_c_1148_n 0.0200388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1149_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_1150_n 0.0066101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1135_n 0.0496551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_288_47#_c_1271_n 0.00997171f $X=-0.19 $Y=1.305 $X2=5.855 $Y2=1.32
cc_162 VPB N_A_288_47#_c_1272_n 0.00977075f $X=-0.19 $Y=1.305 $X2=6.32 $Y2=2.275
cc_163 VPB N_A_288_47#_c_1273_n 4.38232e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_288_47#_c_1268_n 0.00277353f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.53
cc_165 VPB N_A_288_47#_c_1269_n 0.00136736f $X=-0.19 $Y=1.305 $X2=6.065 $Y2=1.53
cc_166 VPB N_A_288_47#_c_1276_n 3.67896e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_288_47#_c_1277_n 0.00406359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_872_316#_c_1405_n 0.00645389f $X=-0.19 $Y=1.305 $X2=1.44 $Y2=1.32
cc_169 VPB N_A_872_316#_c_1408_n 0.0111242f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=1.245
cc_170 VPB N_A_872_316#_c_1406_n 0.00454851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_872_316#_c_1410_n 0.00168598f $X=-0.19 $Y=1.305 $X2=5.78
+ $Y2=0.415
cc_172 VPB N_A_872_316#_c_1411_n 0.00105233f $X=-0.19 $Y=1.305 $X2=6.065
+ $Y2=1.53
cc_173 VPB N_X_c_1503_n 8.99923e-19 $X=-0.19 $Y=1.305 $X2=1.365 $Y2=2.275
cc_174 N_S0_M1016_g N_A2_M1000_g 0.0254984f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_175 N_S0_c_175_n N_A2_c_378_n 0.0230379f $X=1.365 $Y=1.615 $X2=0 $Y2=0
cc_176 N_S0_M1023_g N_A2_c_378_n 0.00220051f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_177 N_S0_c_193_n N_A2_c_378_n 0.00592757f $X=1.005 $Y=1.53 $X2=0 $Y2=0
cc_178 N_S0_c_196_n N_A2_c_378_n 9.9583e-19 $X=1.295 $Y=1.53 $X2=0 $Y2=0
cc_179 N_S0_c_182_n N_A2_c_378_n 0.00193624f $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_180 N_S0_c_183_n N_A2_c_378_n 0.0139922f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_181 N_S0_M1016_g N_A2_c_385_n 0.0139922f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_182 N_S0_M1023_g N_A2_c_385_n 0.0367403f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_183 N_S0_M1025_g A2 3.07188e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_184 N_S0_c_175_n A2 0.00133318f $X=1.365 $Y=1.615 $X2=0 $Y2=0
cc_185 N_S0_c_193_n A2 0.00572305f $X=1.005 $Y=1.53 $X2=0 $Y2=0
cc_186 N_S0_c_196_n A2 0.0054611f $X=1.295 $Y=1.53 $X2=0 $Y2=0
cc_187 N_S0_c_182_n A2 0.00784362f $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_188 N_S0_M1025_g N_A2_c_381_n 0.0169506f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_189 N_S0_c_193_n N_A2_c_381_n 0.00146091f $X=1.005 $Y=1.53 $X2=0 $Y2=0
cc_190 N_S0_c_196_n N_A2_c_381_n 0.00118428f $X=1.295 $Y=1.53 $X2=0 $Y2=0
cc_191 N_S0_c_182_n N_A2_c_381_n 9.40361e-19 $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_192 N_S0_M1025_g N_A2_c_382_n 0.0142496f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_193 N_S0_M1002_g N_A_27_47#_c_442_n 0.0133998f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_194 N_S0_M1023_g N_A_27_47#_M1017_g 0.0201836f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_195 N_S0_M1018_g N_A_27_47#_M1022_g 0.0187022f $X=6.32 $Y=2.275 $X2=0 $Y2=0
cc_196 N_S0_M1015_g N_A_27_47#_c_443_n 0.0184915f $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_197 N_S0_M1025_g N_A_27_47#_c_444_n 0.00866746f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_198 N_S0_M1016_g N_A_27_47#_c_444_n 0.00916433f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_199 S0 N_A_27_47#_c_444_n 0.0525763f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_200 N_S0_c_193_n N_A_27_47#_c_444_n 0.0235359f $X=1.005 $Y=1.53 $X2=0 $Y2=0
cc_201 N_S0_c_194_n N_A_27_47#_c_444_n 0.00267828f $X=0.375 $Y=1.53 $X2=0 $Y2=0
cc_202 N_S0_c_196_n N_A_27_47#_c_444_n 0.00228258f $X=1.295 $Y=1.53 $X2=0 $Y2=0
cc_203 N_S0_c_182_n N_A_27_47#_c_444_n 0.0102687f $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_204 N_S0_c_183_n N_A_27_47#_c_444_n 0.00804141f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_205 N_S0_c_175_n N_A_27_47#_c_455_n 8.45937e-19 $X=1.365 $Y=1.615 $X2=0 $Y2=0
cc_206 N_S0_M1023_g N_A_27_47#_c_455_n 0.0106339f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_207 N_S0_c_176_n N_A_27_47#_c_455_n 0.00281568f $X=1.835 $Y=1.32 $X2=0 $Y2=0
cc_208 N_S0_c_193_n N_A_27_47#_c_455_n 0.014054f $X=1.005 $Y=1.53 $X2=0 $Y2=0
cc_209 N_S0_c_195_n N_A_27_47#_c_455_n 0.00431952f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_210 N_S0_c_196_n N_A_27_47#_c_455_n 0.00821549f $X=1.295 $Y=1.53 $X2=0 $Y2=0
cc_211 N_S0_c_182_n N_A_27_47#_c_455_n 0.024961f $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_212 N_S0_M1016_g N_A_27_47#_c_483_n 0.0183543f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_213 S0 N_A_27_47#_c_483_n 0.0123932f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_214 N_S0_c_193_n N_A_27_47#_c_483_n 0.00399372f $X=1.005 $Y=1.53 $X2=0 $Y2=0
cc_215 N_S0_c_194_n N_A_27_47#_c_483_n 0.00325766f $X=0.375 $Y=1.53 $X2=0 $Y2=0
cc_216 N_S0_c_183_n N_A_27_47#_c_483_n 0.00160965f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_217 N_S0_M1025_g N_A_27_47#_c_445_n 0.0139414f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_218 S0 N_A_27_47#_c_445_n 0.0127362f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_219 N_S0_c_194_n N_A_27_47#_c_445_n 0.00210605f $X=0.375 $Y=1.53 $X2=0 $Y2=0
cc_220 N_S0_c_183_n N_A_27_47#_c_445_n 0.00363508f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_221 N_S0_c_175_n N_A_27_47#_c_446_n 0.023246f $X=1.365 $Y=1.615 $X2=0 $Y2=0
cc_222 N_S0_M1002_g N_A_27_47#_c_446_n 0.0193792f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_223 N_S0_c_195_n N_A_27_47#_c_446_n 2.34296e-19 $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_224 N_S0_c_182_n N_A_27_47#_c_446_n 7.00375e-19 $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_225 N_S0_c_175_n N_A_27_47#_c_447_n 0.00107346f $X=1.365 $Y=1.615 $X2=0 $Y2=0
cc_226 N_S0_c_176_n N_A_27_47#_c_447_n 4.97671e-19 $X=1.835 $Y=1.32 $X2=0 $Y2=0
cc_227 N_S0_M1002_g N_A_27_47#_c_447_n 0.00191472f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_228 N_S0_c_195_n N_A_27_47#_c_447_n 0.00565103f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_229 N_S0_M1015_g N_A_27_47#_c_448_n 0.0126611f $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_230 N_S0_c_179_n N_A_27_47#_c_448_n 0.00529488f $X=6.245 $Y=1.32 $X2=0 $Y2=0
cc_231 N_S0_c_195_n N_A_27_47#_c_448_n 0.00494576f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_232 N_S0_c_198_n N_A_27_47#_c_448_n 0.00305817f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_233 N_S0_c_199_n N_A_27_47#_c_448_n 0.00943055f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_234 N_S0_c_195_n N_A_27_47#_c_456_n 0.301643f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_235 N_S0_M1023_g N_A_27_47#_c_457_n 0.0010293f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_236 N_S0_c_195_n N_A_27_47#_c_457_n 0.0259379f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_237 N_S0_c_195_n N_A_27_47#_c_458_n 0.0255939f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_238 N_S0_c_175_n N_A_27_47#_c_459_n 0.0163856f $X=1.365 $Y=1.615 $X2=0 $Y2=0
cc_239 N_S0_c_176_n N_A_27_47#_c_459_n 0.0206876f $X=1.835 $Y=1.32 $X2=0 $Y2=0
cc_240 N_S0_c_195_n N_A_27_47#_c_459_n 3.65383e-19 $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_241 N_S0_M1023_g N_A_27_47#_c_460_n 0.00425396f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_242 N_S0_c_176_n N_A_27_47#_c_460_n 0.00300332f $X=1.835 $Y=1.32 $X2=0 $Y2=0
cc_243 N_S0_c_195_n N_A_27_47#_c_460_n 0.0103825f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_244 N_S0_c_196_n N_A_27_47#_c_460_n 0.00138334f $X=1.295 $Y=1.53 $X2=0 $Y2=0
cc_245 N_S0_c_180_n N_A_27_47#_c_461_n 0.0215228f $X=5.855 $Y=1.32 $X2=0 $Y2=0
cc_246 N_S0_M1018_g N_A_27_47#_c_461_n 0.0168768f $X=6.32 $Y=2.275 $X2=0 $Y2=0
cc_247 N_S0_c_195_n N_A_27_47#_c_461_n 5.96199e-19 $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_248 N_S0_c_198_n N_A_27_47#_c_461_n 6.73758e-19 $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_249 N_S0_c_199_n N_A_27_47#_c_461_n 2.32403e-19 $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_250 N_S0_M1015_g N_A_27_47#_c_449_n 0.00815578f $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_251 N_S0_c_179_n N_A_27_47#_c_449_n 0.0061637f $X=6.245 $Y=1.32 $X2=0 $Y2=0
cc_252 N_S0_c_180_n N_A_27_47#_c_449_n 0.00445788f $X=5.855 $Y=1.32 $X2=0 $Y2=0
cc_253 N_S0_M1018_g N_A_27_47#_c_449_n 0.00197425f $X=6.32 $Y=2.275 $X2=0 $Y2=0
cc_254 N_S0_c_195_n N_A_27_47#_c_449_n 0.0165427f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_255 N_S0_c_198_n N_A_27_47#_c_449_n 0.00278449f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_256 N_S0_c_199_n N_A_27_47#_c_449_n 0.028941f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_257 N_S0_c_184_n N_A_27_47#_c_449_n 0.00105544f $X=6.38 $Y=1.32 $X2=0 $Y2=0
cc_258 N_S0_M1015_g N_A_27_47#_c_450_n 0.0213388f $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_259 N_S0_c_179_n N_A_27_47#_c_450_n 0.0224415f $X=6.245 $Y=1.32 $X2=0 $Y2=0
cc_260 N_S0_c_199_n N_A_27_47#_c_450_n 0.0014931f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_261 N_S0_c_175_n N_A_27_47#_c_451_n 0.00407077f $X=1.365 $Y=1.615 $X2=0 $Y2=0
cc_262 N_S0_c_176_n N_A_27_47#_c_451_n 0.0117963f $X=1.835 $Y=1.32 $X2=0 $Y2=0
cc_263 N_S0_M1002_g N_A_27_47#_c_451_n 0.00433144f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_264 N_S0_c_195_n N_A_27_47#_c_451_n 0.00800201f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_265 N_S0_c_196_n N_A_27_47#_c_451_n 2.65465e-19 $X=1.295 $Y=1.53 $X2=0 $Y2=0
cc_266 N_S0_c_182_n N_A_27_47#_c_451_n 0.0226549f $X=1.15 $Y=1.53 $X2=0 $Y2=0
cc_267 N_S0_M1002_g N_A3_c_684_n 0.00975299f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_268 N_S0_c_195_n N_A3_c_684_n 0.00281616f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_269 N_S0_c_195_n N_A3_c_691_n 0.00588092f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_270 N_S0_M1002_g A3 8.90548e-19 $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_271 N_S0_c_195_n A3 0.00539843f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_272 N_S0_M1002_g A3 2.79419e-19 $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_273 N_S0_c_195_n A3 0.0104635f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_274 N_S0_M1002_g N_A3_c_687_n 0.0143597f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_275 N_S0_c_195_n N_A3_c_687_n 9.68438e-19 $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_276 N_S0_M1002_g N_A3_c_688_n 0.0238303f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_277 N_S0_c_195_n N_S1_c_743_n 7.7475e-19 $X=6.065 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_278 N_S0_c_195_n N_S1_M1026_g 0.00682163f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_279 N_S0_c_195_n N_S1_c_746_n 0.00336531f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_280 N_S0_c_195_n N_S1_M1008_g 0.00625641f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_281 N_S0_c_195_n S1 0.0121766f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_282 N_S0_c_195_n N_A_600_345#_M1020_g 0.00412283f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_283 N_S0_c_195_n N_A_600_345#_c_829_n 0.00309622f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_284 N_S0_c_195_n N_A_600_345#_c_831_n 0.00452009f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_285 N_S0_c_195_n N_A_600_345#_c_834_n 0.0266831f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_286 N_S0_c_195_n N_A1_M1001_g 0.00948456f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_287 N_S0_M1015_g N_A1_M1027_g 0.0172309f $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_288 N_S0_c_195_n A1 0.0107577f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_289 N_S0_c_180_n N_A1_c_900_n 0.0172309f $X=5.855 $Y=1.32 $X2=0 $Y2=0
cc_290 N_S0_c_195_n N_A1_c_900_n 0.00151751f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_291 N_S0_M1018_g N_A0_M1021_g 0.0345762f $X=6.32 $Y=2.275 $X2=0 $Y2=0
cc_292 N_S0_c_199_n N_A0_M1021_g 9.18038e-19 $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_293 N_S0_c_184_n N_A0_M1021_g 0.0136507f $X=6.38 $Y=1.32 $X2=0 $Y2=0
cc_294 N_S0_M1015_g N_A0_c_939_n 2.01922e-19 $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_295 N_S0_c_199_n N_A0_c_939_n 0.00629593f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_296 N_S0_c_184_n N_A0_c_939_n 5.65638e-19 $X=6.38 $Y=1.32 $X2=0 $Y2=0
cc_297 N_S0_c_184_n N_A0_c_940_n 0.00525853f $X=6.38 $Y=1.32 $X2=0 $Y2=0
cc_298 N_S0_c_195_n N_A_788_316#_M1020_d 6.16189e-19 $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_299 N_S0_c_195_n N_A_788_316#_c_989_n 0.0139892f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_300 N_S0_M1018_g N_A_788_316#_c_995_n 0.00848933f $X=6.32 $Y=2.275 $X2=0
+ $Y2=0
cc_301 N_S0_M1018_g N_A_788_316#_c_997_n 7.58543e-19 $X=6.32 $Y=2.275 $X2=0
+ $Y2=0
cc_302 N_S0_c_198_n N_A_788_316#_c_997_n 9.4687e-19 $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_303 N_S0_c_199_n N_A_788_316#_c_997_n 0.00987457f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_304 N_S0_c_184_n N_A_788_316#_c_997_n 5.56235e-19 $X=6.38 $Y=1.32 $X2=0 $Y2=0
cc_305 N_S0_c_199_n N_A_788_316#_c_998_n 0.00454895f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_306 N_S0_M1018_g N_A_788_316#_c_1001_n 0.00380986f $X=6.32 $Y=2.275 $X2=0
+ $Y2=0
cc_307 N_S0_c_195_n N_A_788_316#_c_1001_n 0.00774624f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_308 N_S0_c_198_n N_A_788_316#_c_1001_n 0.0150323f $X=6.21 $Y=1.53 $X2=0 $Y2=0
cc_309 N_S0_c_199_n N_A_788_316#_c_1001_n 0.00544375f $X=6.21 $Y=1.53 $X2=0
+ $Y2=0
cc_310 N_S0_c_184_n N_A_788_316#_c_1001_n 9.57678e-19 $X=6.38 $Y=1.32 $X2=0
+ $Y2=0
cc_311 N_S0_M1018_g N_A_788_316#_c_1018_n 0.00100458f $X=6.32 $Y=2.275 $X2=0
+ $Y2=0
cc_312 N_S0_M1018_g N_A_788_316#_c_1019_n 0.00151791f $X=6.32 $Y=2.275 $X2=0
+ $Y2=0
cc_313 N_S0_M1016_g N_VPWR_c_1136_n 0.01126f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_314 N_S0_M1023_g N_VPWR_c_1136_n 0.00200626f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_315 N_S0_M1023_g N_VPWR_c_1142_n 0.00546481f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_316 N_S0_M1018_g N_VPWR_c_1144_n 0.00545391f $X=6.32 $Y=2.275 $X2=0 $Y2=0
cc_317 N_S0_M1016_g N_VPWR_c_1146_n 0.0033925f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_318 N_S0_M1016_g N_VPWR_c_1135_n 0.004976f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_319 N_S0_M1023_g N_VPWR_c_1135_n 0.00623554f $X=1.365 $Y=2.275 $X2=0 $Y2=0
cc_320 N_S0_M1018_g N_VPWR_c_1135_n 0.00557212f $X=6.32 $Y=2.275 $X2=0 $Y2=0
cc_321 N_S0_c_195_n N_A_288_47#_M1020_s 6.67976e-19 $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_322 N_S0_M1023_g N_A_288_47#_c_1279_n 0.00426873f $X=1.365 $Y=2.275 $X2=0
+ $Y2=0
cc_323 N_S0_M1002_g N_A_288_47#_c_1280_n 0.0106572f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_324 N_S0_M1002_g N_A_288_47#_c_1267_n 0.0163104f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_325 N_S0_c_195_n N_A_288_47#_c_1271_n 0.0139277f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_326 N_S0_c_195_n N_A_288_47#_c_1283_n 5.93677e-19 $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_327 N_S0_c_176_n N_A_288_47#_c_1268_n 0.00510606f $X=1.835 $Y=1.32 $X2=0
+ $Y2=0
cc_328 N_S0_M1002_g N_A_288_47#_c_1268_n 4.69181e-19 $X=1.91 $Y=0.415 $X2=0
+ $Y2=0
cc_329 N_S0_c_195_n N_A_288_47#_c_1268_n 0.0104059f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_330 N_S0_c_195_n N_A_288_47#_c_1269_n 0.0127493f $X=6.065 $Y=1.53 $X2=0 $Y2=0
cc_331 N_S0_c_195_n N_A_872_316#_M1008_d 2.14086e-19 $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_332 N_S0_c_195_n N_A_872_316#_c_1405_n 0.0203392f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_333 N_S0_c_195_n N_A_872_316#_c_1408_n 0.0198601f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_334 N_S0_M1015_g N_A_872_316#_c_1406_n 0.00711633f $X=5.78 $Y=0.415 $X2=0
+ $Y2=0
cc_335 N_S0_c_195_n N_A_872_316#_c_1406_n 0.0155282f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_336 N_S0_M1015_g N_A_872_316#_c_1417_n 0.0110411f $X=5.78 $Y=0.415 $X2=0
+ $Y2=0
cc_337 N_S0_M1018_g N_A_872_316#_c_1418_n 0.00246628f $X=6.32 $Y=2.275 $X2=0
+ $Y2=0
cc_338 N_S0_c_195_n N_A_872_316#_c_1418_n 9.00069e-19 $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_339 N_S0_c_198_n N_A_872_316#_c_1418_n 0.00117806f $X=6.21 $Y=1.53 $X2=0
+ $Y2=0
cc_340 N_S0_c_199_n N_A_872_316#_c_1418_n 0.00270797f $X=6.21 $Y=1.53 $X2=0
+ $Y2=0
cc_341 N_S0_c_195_n N_A_872_316#_c_1411_n 0.00369858f $X=6.065 $Y=1.53 $X2=0
+ $Y2=0
cc_342 N_S0_M1025_g N_VGND_c_1534_n 0.0112612f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_343 N_S0_M1002_g N_VGND_c_1535_n 0.00171495f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_344 N_S0_M1025_g N_VGND_c_1540_n 0.00339367f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_345 N_S0_M1002_g N_VGND_c_1541_n 0.00379702f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_346 N_S0_M1015_g N_VGND_c_1543_n 0.00366111f $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_347 N_S0_M1025_g N_VGND_c_1549_n 0.00497794f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_348 N_S0_M1002_g N_VGND_c_1549_n 0.00583199f $X=1.91 $Y=0.415 $X2=0 $Y2=0
cc_349 N_S0_M1015_g N_VGND_c_1549_n 0.00589952f $X=5.78 $Y=0.415 $X2=0 $Y2=0
cc_350 A2 N_A_27_47#_c_442_n 0.00301706f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_351 N_A2_c_382_n N_A_27_47#_c_442_n 0.0221667f $X=0.92 $Y=0.765 $X2=0 $Y2=0
cc_352 N_A2_M1000_g N_A_27_47#_c_444_n 0.00145462f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_353 N_A2_c_378_n N_A_27_47#_c_444_n 0.0087804f $X=0.887 $Y=1.675 $X2=0 $Y2=0
cc_354 A2 N_A_27_47#_c_444_n 0.0221499f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_355 N_A2_c_381_n N_A_27_47#_c_444_n 0.0017807f $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_356 N_A2_M1000_g N_A_27_47#_c_455_n 0.0120011f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_357 N_A2_c_385_n N_A_27_47#_c_455_n 2.31416e-19 $X=0.887 $Y=1.715 $X2=0 $Y2=0
cc_358 N_A2_c_381_n N_A_27_47#_c_455_n 0.00150087f $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_359 N_A2_M1000_g N_A_27_47#_c_483_n 0.00338175f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_360 A2 N_A_27_47#_c_445_n 0.00594711f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_361 A2 N_A_27_47#_c_445_n 0.00317992f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_362 N_A2_c_381_n N_A_27_47#_c_445_n 2.83902e-19 $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_363 N_A2_c_382_n N_A_27_47#_c_445_n 0.0011592f $X=0.92 $Y=0.765 $X2=0 $Y2=0
cc_364 A2 N_A_27_47#_c_446_n 0.0020763f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_365 N_A2_c_381_n N_A_27_47#_c_446_n 0.0144246f $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_366 A2 N_A_27_47#_c_447_n 0.00453132f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_367 A2 N_A_27_47#_c_447_n 0.0217226f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_368 N_A2_c_381_n N_A_27_47#_c_447_n 2.07055e-19 $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_369 N_A2_c_378_n N_A_27_47#_c_451_n 0.00344585f $X=0.887 $Y=1.675 $X2=0 $Y2=0
cc_370 A2 N_A_27_47#_c_451_n 0.00304052f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_371 N_A2_c_381_n N_A_27_47#_c_451_n 2.60449e-19 $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_372 N_A2_M1000_g N_VPWR_c_1136_n 0.00980825f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_373 N_A2_M1000_g N_VPWR_c_1142_n 0.0046653f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_374 N_A2_M1000_g N_VPWR_c_1135_n 0.00440885f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_375 N_A2_M1000_g N_A_288_47#_c_1279_n 7.3574e-19 $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_376 A2 N_A_288_47#_c_1267_n 0.00346305f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_377 A2 N_VGND_c_1534_n 4.02658e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_378 N_A2_c_382_n N_VGND_c_1534_n 0.00982698f $X=0.92 $Y=0.765 $X2=0 $Y2=0
cc_379 A2 N_VGND_c_1541_n 0.00747058f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_380 N_A2_c_381_n N_VGND_c_1541_n 0.00106747f $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_381 N_A2_c_382_n N_VGND_c_1541_n 0.0046653f $X=0.92 $Y=0.765 $X2=0 $Y2=0
cc_382 A2 N_VGND_c_1549_n 0.00740674f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_383 A2 N_VGND_c_1549_n 0.00586186f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_384 N_A2_c_381_n N_VGND_c_1549_n 0.00131849f $X=0.92 $Y=0.93 $X2=0 $Y2=0
cc_385 N_A2_c_382_n N_VGND_c_1549_n 0.00440885f $X=0.92 $Y=0.765 $X2=0 $Y2=0
cc_386 A2 A_193_47# 0.00485061f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_387 N_A_27_47#_c_451_n N_A3_c_684_n 2.69784e-19 $X=1.73 $Y=1.575 $X2=0 $Y2=0
cc_388 N_A_27_47#_M1017_g N_A3_c_690_n 0.0138424f $X=1.785 $Y=2.275 $X2=0 $Y2=0
cc_389 N_A_27_47#_c_456_n N_A3_c_690_n 0.00580906f $X=5.605 $Y=1.87 $X2=0 $Y2=0
cc_390 N_A_27_47#_c_459_n N_A3_c_690_n 0.00498599f $X=1.815 $Y=1.74 $X2=0 $Y2=0
cc_391 N_A_27_47#_c_456_n N_A3_c_691_n 0.00220307f $X=5.605 $Y=1.87 $X2=0 $Y2=0
cc_392 N_A_27_47#_c_459_n N_A3_c_691_n 0.00134881f $X=1.815 $Y=1.74 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_456_n N_S1_M1026_g 0.00310138f $X=5.605 $Y=1.87 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_456_n N_S1_c_750_n 7.54852e-19 $X=5.605 $Y=1.87 $X2=0 $Y2=0
cc_395 N_A_27_47#_c_456_n N_S1_M1008_g 0.00272158f $X=5.605 $Y=1.87 $X2=0 $Y2=0
cc_396 N_A_27_47#_c_456_n N_A_600_345#_M1020_g 0.00263087f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_456_n N_A_600_345#_c_834_n 0.0185716f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_M1022_g N_A1_M1001_g 0.0154632f $X=5.9 $Y=2.275 $X2=0 $Y2=0
cc_399 N_A_27_47#_c_456_n N_A1_M1001_g 0.00637365f $X=5.605 $Y=1.87 $X2=0 $Y2=0
cc_400 N_A_27_47#_c_461_n N_A1_M1001_g 0.00734459f $X=5.87 $Y=1.74 $X2=0 $Y2=0
cc_401 N_A_27_47#_c_449_n N_A1_M1001_g 0.00100677f $X=5.87 $Y=1.74 $X2=0 $Y2=0
cc_402 N_A_27_47#_c_443_n N_A0_M1024_g 0.0317614f $X=6.33 $Y=0.705 $X2=0 $Y2=0
cc_403 N_A_27_47#_c_448_n N_A0_M1024_g 2.38614e-19 $X=6.2 $Y=0.87 $X2=0 $Y2=0
cc_404 N_A_27_47#_c_448_n N_A0_c_939_n 0.00248128f $X=6.2 $Y=0.87 $X2=0 $Y2=0
cc_405 N_A_27_47#_c_449_n N_A0_c_939_n 0.00143247f $X=5.87 $Y=1.74 $X2=0 $Y2=0
cc_406 N_A_27_47#_c_450_n N_A0_c_939_n 3.79122e-19 $X=6.33 $Y=0.87 $X2=0 $Y2=0
cc_407 N_A_27_47#_c_450_n N_A0_c_940_n 0.00142667f $X=6.33 $Y=0.87 $X2=0 $Y2=0
cc_408 N_A_27_47#_c_443_n A0 0.00936228f $X=6.33 $Y=0.705 $X2=0 $Y2=0
cc_409 N_A_27_47#_c_448_n A0 0.0178996f $X=6.2 $Y=0.87 $X2=0 $Y2=0
cc_410 N_A_27_47#_c_456_n N_A_788_316#_M1020_d 0.00139404f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_456_n N_A_788_316#_c_989_n 0.0146457f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_M1022_g N_A_788_316#_c_1001_n 0.00125658f $X=5.9 $Y=2.275
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_c_456_n N_A_788_316#_c_1001_n 0.0865979f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_458_n N_A_788_316#_c_1001_n 0.0265153f $X=5.75 $Y=1.87 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_461_n N_A_788_316#_c_1001_n 9.1661e-19 $X=5.87 $Y=1.74 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_449_n N_A_788_316#_c_1001_n 0.00140404f $X=5.87 $Y=1.74
+ $X2=0 $Y2=0
cc_417 N_A_27_47#_c_456_n N_A_788_316#_c_1002_n 0.0274654f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_418 N_A_27_47#_c_456_n N_A_788_316#_c_1003_n 0.00376868f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_c_455_n N_VPWR_M1016_d 0.00123431f $X=1.56 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_420 N_A_27_47#_c_483_n N_VPWR_M1016_d 0.00236204f $X=0.665 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_421 N_A_27_47#_c_456_n N_VPWR_M1003_d 0.00361504f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_456_n N_VPWR_M1001_s 0.00166679f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_c_455_n N_VPWR_c_1136_n 0.00562223f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_c_483_n N_VPWR_c_1136_n 0.00756186f $X=0.665 $Y=1.87 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_456_n N_VPWR_c_1137_n 0.0081452f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_c_456_n N_VPWR_c_1138_n 0.00382585f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_M1017_g N_VPWR_c_1142_n 0.00390868f $X=1.785 $Y=2.275 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_M1022_g N_VPWR_c_1144_n 0.00385416f $X=5.9 $Y=2.275 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_602_p N_VPWR_c_1146_n 0.00713694f $X=0.26 $Y=2.21 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_c_483_n N_VPWR_c_1146_n 0.00247476f $X=0.665 $Y=1.87 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_M1016_s N_VPWR_c_1135_n 0.00375328f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_M1017_g N_VPWR_c_1135_n 0.0059629f $X=1.785 $Y=2.275 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_M1022_g N_VPWR_c_1135_n 0.00539892f $X=5.9 $Y=2.275 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_602_p N_VPWR_c_1135_n 0.00608739f $X=0.26 $Y=2.21 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_c_455_n N_VPWR_c_1135_n 0.0199013f $X=1.56 $Y=1.87 $X2=0 $Y2=0
cc_436 N_A_27_47#_c_483_n N_VPWR_c_1135_n 0.00502272f $X=0.665 $Y=1.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_456_n N_VPWR_c_1135_n 0.0370753f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_457_n N_VPWR_c_1135_n 0.0160199f $X=1.755 $Y=1.87 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_c_455_n A_193_369# 0.00364525f $X=1.56 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_440 N_A_27_47#_c_456_n N_A_288_47#_M1020_s 0.00110497f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_M1017_g N_A_288_47#_c_1279_n 0.00945162f $X=1.785 $Y=2.275
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_455_n N_A_288_47#_c_1279_n 0.00793212f $X=1.56 $Y=1.87 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_456_n N_A_288_47#_c_1279_n 0.00239538f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_457_n N_A_288_47#_c_1279_n 0.00325767f $X=1.755 $Y=1.87
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_459_n N_A_288_47#_c_1279_n 0.00203367f $X=1.815 $Y=1.74
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_460_n N_A_288_47#_c_1279_n 0.019174f $X=1.815 $Y=1.74 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_446_n N_A_288_47#_c_1280_n 0.00341595f $X=1.49 $Y=0.87 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_447_n N_A_288_47#_c_1280_n 0.017832f $X=1.645 $Y=0.87 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_442_n N_A_288_47#_c_1267_n 4.32952e-19 $X=1.365 $Y=0.705
+ $X2=0 $Y2=0
cc_450 N_A_27_47#_c_446_n N_A_288_47#_c_1267_n 3.02268e-19 $X=1.49 $Y=0.87 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_447_n N_A_288_47#_c_1267_n 0.024855f $X=1.645 $Y=0.87 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_451_n N_A_288_47#_c_1267_n 0.0143036f $X=1.73 $Y=1.575 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_M1017_g N_A_288_47#_c_1271_n 0.00391048f $X=1.785 $Y=2.275
+ $X2=0 $Y2=0
cc_454 N_A_27_47#_c_456_n N_A_288_47#_c_1271_n 0.0132084f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_c_457_n N_A_288_47#_c_1271_n 0.00147315f $X=1.755 $Y=1.87
+ $X2=0 $Y2=0
cc_456 N_A_27_47#_c_459_n N_A_288_47#_c_1271_n 0.0023745f $X=1.815 $Y=1.74 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_460_n N_A_288_47#_c_1271_n 0.0274922f $X=1.815 $Y=1.74 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_451_n N_A_288_47#_c_1271_n 0.00661642f $X=1.73 $Y=1.575
+ $X2=0 $Y2=0
cc_459 N_A_27_47#_c_456_n N_A_288_47#_c_1283_n 0.00766148f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_460 N_A_27_47#_c_456_n N_A_288_47#_c_1272_n 0.0018441f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_461 N_A_27_47#_c_456_n N_A_288_47#_c_1273_n 0.00419026f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_462 N_A_27_47#_c_459_n N_A_288_47#_c_1268_n 0.00156489f $X=1.815 $Y=1.74
+ $X2=0 $Y2=0
cc_463 N_A_27_47#_c_451_n N_A_288_47#_c_1268_n 0.0121557f $X=1.73 $Y=1.575 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_456_n N_A_288_47#_c_1269_n 0.00302831f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_465 N_A_27_47#_c_456_n N_A_288_47#_c_1276_n 0.0865557f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_M1017_g N_A_288_47#_c_1316_n 0.00114372f $X=1.785 $Y=2.275
+ $X2=0 $Y2=0
cc_467 N_A_27_47#_c_456_n N_A_288_47#_c_1316_n 0.0263636f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_459_n N_A_288_47#_c_1316_n 2.73637e-19 $X=1.815 $Y=1.74
+ $X2=0 $Y2=0
cc_469 N_A_27_47#_c_456_n N_A_288_47#_c_1277_n 0.0275563f $X=5.605 $Y=1.87 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_456_n A_372_413# 0.00325861f $X=5.605 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_471 N_A_27_47#_c_456_n N_A_872_316#_M1008_d 0.00209072f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_472 N_A_27_47#_c_456_n N_A_872_316#_c_1405_n 0.0108836f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_473 N_A_27_47#_c_456_n N_A_872_316#_c_1408_n 0.0143232f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_474 N_A_27_47#_c_448_n N_A_872_316#_c_1406_n 0.0274865f $X=6.2 $Y=0.87 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_449_n N_A_872_316#_c_1406_n 0.0406896f $X=5.87 $Y=1.74 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_M1022_g N_A_872_316#_c_1410_n 0.00337169f $X=5.9 $Y=2.275
+ $X2=0 $Y2=0
cc_477 N_A_27_47#_c_456_n N_A_872_316#_c_1410_n 0.0140427f $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_478 N_A_27_47#_c_458_n N_A_872_316#_c_1410_n 0.00275409f $X=5.75 $Y=1.87
+ $X2=0 $Y2=0
cc_479 N_A_27_47#_c_461_n N_A_872_316#_c_1410_n 4.04648e-19 $X=5.87 $Y=1.74
+ $X2=0 $Y2=0
cc_480 N_A_27_47#_c_449_n N_A_872_316#_c_1410_n 0.0172732f $X=5.87 $Y=1.74 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_448_n N_A_872_316#_c_1417_n 0.0259764f $X=6.2 $Y=0.87 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_450_n N_A_872_316#_c_1417_n 0.00325712f $X=6.33 $Y=0.87
+ $X2=0 $Y2=0
cc_483 N_A_27_47#_M1022_g N_A_872_316#_c_1418_n 0.00887377f $X=5.9 $Y=2.275
+ $X2=0 $Y2=0
cc_484 N_A_27_47#_c_456_n N_A_872_316#_c_1418_n 7.78043e-19 $X=5.605 $Y=1.87
+ $X2=0 $Y2=0
cc_485 N_A_27_47#_c_458_n N_A_872_316#_c_1418_n 7.97005e-19 $X=5.75 $Y=1.87
+ $X2=0 $Y2=0
cc_486 N_A_27_47#_c_461_n N_A_872_316#_c_1418_n 0.00193698f $X=5.87 $Y=1.74
+ $X2=0 $Y2=0
cc_487 N_A_27_47#_c_449_n N_A_872_316#_c_1418_n 0.0189711f $X=5.87 $Y=1.74 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_461_n N_A_872_316#_c_1411_n 5.13754e-19 $X=5.87 $Y=1.74
+ $X2=0 $Y2=0
cc_489 N_A_27_47#_c_449_n N_A_872_316#_c_1411_n 0.0142775f $X=5.87 $Y=1.74 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_c_456_n A_1060_369# 4.93895e-19 $X=5.605 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_491 N_A_27_47#_c_445_n N_VGND_M1025_d 8.65503e-19 $X=0.58 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_492 N_A_27_47#_c_442_n N_VGND_c_1534_n 0.00170649f $X=1.365 $Y=0.705 $X2=0
+ $Y2=0
cc_493 N_A_27_47#_c_445_n N_VGND_c_1534_n 0.0068368f $X=0.58 $Y=0.72 $X2=0 $Y2=0
cc_494 N_A_27_47#_c_667_p N_VGND_c_1540_n 0.00713381f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_445_n N_VGND_c_1540_n 0.0024638f $X=0.58 $Y=0.72 $X2=0 $Y2=0
cc_496 N_A_27_47#_c_442_n N_VGND_c_1541_n 0.0055032f $X=1.365 $Y=0.705 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_446_n N_VGND_c_1541_n 5.70717e-19 $X=1.49 $Y=0.87 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_c_447_n N_VGND_c_1541_n 9.49253e-19 $X=1.645 $Y=0.87 $X2=0
+ $Y2=0
cc_499 N_A_27_47#_c_443_n N_VGND_c_1543_n 0.00555329f $X=6.33 $Y=0.705 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_448_n N_VGND_c_1543_n 9.49253e-19 $X=6.2 $Y=0.87 $X2=0 $Y2=0
cc_501 N_A_27_47#_c_450_n N_VGND_c_1543_n 6.11083e-19 $X=6.33 $Y=0.87 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_M1025_s N_VGND_c_1549_n 0.00355099f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_503 N_A_27_47#_c_442_n N_VGND_c_1549_n 0.0101784f $X=1.365 $Y=0.705 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_c_443_n N_VGND_c_1549_n 0.0103474f $X=6.33 $Y=0.705 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_c_667_p N_VGND_c_1549_n 0.00618063f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_c_445_n N_VGND_c_1549_n 0.00495052f $X=0.58 $Y=0.72 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_446_n N_VGND_c_1549_n 7.31425e-19 $X=1.49 $Y=0.87 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_447_n N_VGND_c_1549_n 0.00203708f $X=1.645 $Y=0.87 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_c_448_n N_VGND_c_1549_n 0.00295441f $X=6.2 $Y=0.87 $X2=0 $Y2=0
cc_510 N_A_27_47#_c_450_n N_VGND_c_1549_n 8.53329e-19 $X=6.33 $Y=0.87 $X2=0
+ $Y2=0
cc_511 A3 N_S1_c_743_n 0.00214806f $X=2.445 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_512 N_A3_c_687_n N_S1_c_743_n 0.0207417f $X=2.405 $Y=0.93 $X2=-0.19 $Y2=-0.24
cc_513 N_A3_c_688_n N_S1_c_743_n 0.00103795f $X=2.405 $Y=0.765 $X2=-0.19
+ $Y2=-0.24
cc_514 N_A3_c_684_n N_S1_M1026_g 0.0126585f $X=2.39 $Y=1.5 $X2=0 $Y2=0
cc_515 N_A3_c_691_n N_S1_M1026_g 0.0187074f $X=2.505 $Y=1.575 $X2=0 $Y2=0
cc_516 A3 N_S1_M1026_g 6.79827e-19 $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_517 N_A3_c_688_n N_S1_c_745_n 0.0137149f $X=2.405 $Y=0.765 $X2=0 $Y2=0
cc_518 N_A3_c_690_n N_S1_c_751_n 0.0187074f $X=2.505 $Y=1.65 $X2=0 $Y2=0
cc_519 N_A3_c_684_n S1 5.90277e-19 $X=2.39 $Y=1.5 $X2=0 $Y2=0
cc_520 A3 S1 0.0478665f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_521 N_A3_c_687_n S1 3.38407e-19 $X=2.405 $Y=0.93 $X2=0 $Y2=0
cc_522 N_A3_c_690_n N_A_600_345#_c_834_n 0.00125935f $X=2.505 $Y=1.65 $X2=0
+ $Y2=0
cc_523 N_A3_c_690_n N_VPWR_c_1137_n 0.0064285f $X=2.505 $Y=1.65 $X2=0 $Y2=0
cc_524 N_A3_c_690_n N_VPWR_c_1142_n 0.00585385f $X=2.505 $Y=1.65 $X2=0 $Y2=0
cc_525 N_A3_c_690_n N_VPWR_c_1135_n 0.00587666f $X=2.505 $Y=1.65 $X2=0 $Y2=0
cc_526 N_A3_c_688_n N_A_288_47#_c_1280_n 0.00145818f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_527 N_A3_c_684_n N_A_288_47#_c_1267_n 9.61953e-19 $X=2.39 $Y=1.5 $X2=0 $Y2=0
cc_528 A3 N_A_288_47#_c_1267_n 0.0240227f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_529 A3 N_A_288_47#_c_1267_n 0.00948099f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_530 N_A3_c_687_n N_A_288_47#_c_1267_n 0.00133579f $X=2.405 $Y=0.93 $X2=0
+ $Y2=0
cc_531 N_A3_c_688_n N_A_288_47#_c_1267_n 0.00349406f $X=2.405 $Y=0.765 $X2=0
+ $Y2=0
cc_532 N_A3_c_684_n N_A_288_47#_c_1271_n 0.00798315f $X=2.39 $Y=1.5 $X2=0 $Y2=0
cc_533 N_A3_c_690_n N_A_288_47#_c_1271_n 0.0105472f $X=2.505 $Y=1.65 $X2=0 $Y2=0
cc_534 N_A3_c_684_n N_A_288_47#_c_1268_n 0.00307277f $X=2.39 $Y=1.5 $X2=0 $Y2=0
cc_535 A3 N_A_288_47#_c_1268_n 0.00647251f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_536 N_A3_c_690_n N_A_288_47#_c_1276_n 0.00410206f $X=2.505 $Y=1.65 $X2=0
+ $Y2=0
cc_537 N_A3_c_690_n N_A_288_47#_c_1316_n 4.9262e-19 $X=2.505 $Y=1.65 $X2=0 $Y2=0
cc_538 A3 N_VGND_c_1535_n 0.0115245f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_539 N_A3_c_687_n N_VGND_c_1535_n 3.61231e-19 $X=2.405 $Y=0.93 $X2=0 $Y2=0
cc_540 N_A3_c_688_n N_VGND_c_1535_n 0.00975119f $X=2.405 $Y=0.765 $X2=0 $Y2=0
cc_541 A3 N_VGND_c_1541_n 0.00314583f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_542 N_A3_c_688_n N_VGND_c_1541_n 0.00391931f $X=2.405 $Y=0.765 $X2=0 $Y2=0
cc_543 A3 N_VGND_c_1549_n 0.00579556f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_544 N_A3_c_688_n N_VGND_c_1549_n 0.00476517f $X=2.405 $Y=0.765 $X2=0 $Y2=0
cc_545 N_S1_c_750_n N_A_600_345#_M1020_g 0.00975169f $X=4.21 $Y=2.54 $X2=0 $Y2=0
cc_546 N_S1_M1008_g N_A_600_345#_M1020_g 0.0197432f $X=4.285 $Y=1.85 $X2=0 $Y2=0
cc_547 N_S1_M1008_g N_A_600_345#_c_829_n 0.0120884f $X=4.285 $Y=1.85 $X2=0 $Y2=0
cc_548 N_S1_c_747_n N_A_600_345#_M1012_g 0.0192711f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_549 N_S1_c_743_n N_A_600_345#_c_831_n 3.3029e-19 $X=2.925 $Y=1.095 $X2=0
+ $Y2=0
cc_550 N_S1_M1026_g N_A_600_345#_c_831_n 0.0156633f $X=2.925 $Y=2.045 $X2=0
+ $Y2=0
cc_551 N_S1_c_746_n N_A_600_345#_c_831_n 0.0490984f $X=3.805 $Y=0.805 $X2=0
+ $Y2=0
cc_552 S1 N_A_600_345#_c_831_n 0.00152957f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_553 N_S1_c_743_n N_A_600_345#_c_833_n 0.00109538f $X=2.925 $Y=1.095 $X2=0
+ $Y2=0
cc_554 N_S1_c_745_n N_A_600_345#_c_833_n 0.00538776f $X=2.93 $Y=0.73 $X2=0 $Y2=0
cc_555 N_S1_c_746_n N_A_600_345#_c_833_n 0.0116555f $X=3.805 $Y=0.805 $X2=0
+ $Y2=0
cc_556 N_S1_c_747_n N_A_600_345#_c_833_n 6.32935e-19 $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_557 S1 N_A_600_345#_c_833_n 0.0258653f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_558 N_S1_M1026_g N_A_600_345#_c_834_n 0.0179348f $X=2.925 $Y=2.045 $X2=0
+ $Y2=0
cc_559 N_S1_c_750_n N_A_600_345#_c_834_n 0.00578358f $X=4.21 $Y=2.54 $X2=0 $Y2=0
cc_560 N_S1_c_746_n N_A_600_345#_c_834_n 0.00300126f $X=3.805 $Y=0.805 $X2=0
+ $Y2=0
cc_561 S1 N_A_600_345#_c_834_n 0.0214342f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_562 N_S1_c_745_n N_A_600_345#_c_835_n 0.00233282f $X=2.93 $Y=0.73 $X2=0 $Y2=0
cc_563 N_S1_c_746_n N_A_600_345#_c_835_n 0.00530393f $X=3.805 $Y=0.805 $X2=0
+ $Y2=0
cc_564 N_S1_c_747_n N_A_600_345#_c_835_n 0.00108928f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_565 S1 N_A_600_345#_c_835_n 0.00330055f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_566 N_S1_c_747_n N_A_788_316#_c_989_n 0.00191245f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_567 N_S1_M1008_g N_A_788_316#_c_989_n 0.00238534f $X=4.285 $Y=1.85 $X2=0
+ $Y2=0
cc_568 N_S1_c_750_n N_A_788_316#_c_999_n 0.00293376f $X=4.21 $Y=2.54 $X2=0 $Y2=0
cc_569 N_S1_M1008_g N_A_788_316#_c_1002_n 0.00411296f $X=4.285 $Y=1.85 $X2=0
+ $Y2=0
cc_570 N_S1_M1008_g N_A_788_316#_c_1003_n 0.0125788f $X=4.285 $Y=1.85 $X2=0
+ $Y2=0
cc_571 N_S1_M1026_g N_VPWR_c_1137_n 0.00655497f $X=2.925 $Y=2.045 $X2=0 $Y2=0
cc_572 N_S1_M1008_g N_VPWR_c_1138_n 0.0110777f $X=4.285 $Y=1.85 $X2=0 $Y2=0
cc_573 N_S1_c_751_n N_VPWR_c_1147_n 0.0435688f $X=3 $Y=2.54 $X2=0 $Y2=0
cc_574 N_S1_c_750_n N_VPWR_c_1135_n 0.0304569f $X=4.21 $Y=2.54 $X2=0 $Y2=0
cc_575 N_S1_c_751_n N_VPWR_c_1135_n 0.00442783f $X=3 $Y=2.54 $X2=0 $Y2=0
cc_576 N_S1_M1026_g N_A_288_47#_c_1272_n 0.0024883f $X=2.925 $Y=2.045 $X2=0
+ $Y2=0
cc_577 N_S1_c_750_n N_A_288_47#_c_1272_n 0.0101272f $X=4.21 $Y=2.54 $X2=0 $Y2=0
cc_578 N_S1_M1008_g N_A_288_47#_c_1272_n 2.99929e-19 $X=4.285 $Y=1.85 $X2=0
+ $Y2=0
cc_579 N_S1_M1026_g N_A_288_47#_c_1273_n 0.00265256f $X=2.925 $Y=2.045 $X2=0
+ $Y2=0
cc_580 N_S1_c_746_n N_A_288_47#_c_1269_n 0.00890714f $X=3.805 $Y=0.805 $X2=0
+ $Y2=0
cc_581 N_S1_c_747_n N_A_288_47#_c_1269_n 0.00142837f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_582 N_S1_c_746_n N_A_288_47#_c_1270_n 0.00269638f $X=3.805 $Y=0.805 $X2=0
+ $Y2=0
cc_583 N_S1_c_747_n N_A_288_47#_c_1270_n 0.00362535f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_584 N_S1_M1026_g N_A_288_47#_c_1276_n 0.0049068f $X=2.925 $Y=2.045 $X2=0
+ $Y2=0
cc_585 N_S1_c_750_n N_A_288_47#_c_1276_n 0.00260084f $X=4.21 $Y=2.54 $X2=0 $Y2=0
cc_586 N_S1_M1026_g N_A_288_47#_c_1277_n 0.00136441f $X=2.925 $Y=2.045 $X2=0
+ $Y2=0
cc_587 N_S1_c_750_n N_A_288_47#_c_1277_n 0.00358607f $X=4.21 $Y=2.54 $X2=0 $Y2=0
cc_588 N_S1_M1008_g N_A_288_47#_c_1277_n 5.70583e-19 $X=4.285 $Y=1.85 $X2=0
+ $Y2=0
cc_589 N_S1_M1008_g N_A_872_316#_c_1405_n 0.0028409f $X=4.285 $Y=1.85 $X2=0
+ $Y2=0
cc_590 N_S1_c_743_n N_VGND_c_1535_n 0.00120134f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_591 N_S1_c_745_n N_VGND_c_1535_n 0.00710898f $X=2.93 $Y=0.73 $X2=0 $Y2=0
cc_592 N_S1_c_743_n N_VGND_c_1542_n 3.27123e-19 $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_593 N_S1_c_745_n N_VGND_c_1542_n 0.00426984f $X=2.93 $Y=0.73 $X2=0 $Y2=0
cc_594 N_S1_c_746_n N_VGND_c_1542_n 0.0030174f $X=3.805 $Y=0.805 $X2=0 $Y2=0
cc_595 N_S1_c_747_n N_VGND_c_1542_n 0.00565823f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_596 S1 N_VGND_c_1542_n 0.00312826f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_597 N_S1_c_745_n N_VGND_c_1549_n 0.00749741f $X=2.93 $Y=0.73 $X2=0 $Y2=0
cc_598 N_S1_c_746_n N_VGND_c_1549_n 0.00370828f $X=3.805 $Y=0.805 $X2=0 $Y2=0
cc_599 N_S1_c_747_n N_VGND_c_1549_n 0.0117171f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_600 S1 N_VGND_c_1549_n 0.00521238f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_601 N_A_600_345#_M1012_g N_A1_c_900_n 0.0030673f $X=4.305 $Y=0.445 $X2=0
+ $Y2=0
cc_602 N_A_600_345#_c_829_n N_A_788_316#_c_989_n 0.015488f $X=4.23 $Y=1.165
+ $X2=0 $Y2=0
cc_603 N_A_600_345#_M1012_g N_A_788_316#_c_989_n 0.00651443f $X=4.305 $Y=0.445
+ $X2=0 $Y2=0
cc_604 N_A_600_345#_c_832_n N_A_788_316#_c_989_n 0.007437f $X=3.865 $Y=1.225
+ $X2=0 $Y2=0
cc_605 N_A_600_345#_M1020_g N_A_788_316#_c_999_n 9.91098e-19 $X=3.865 $Y=1.85
+ $X2=0 $Y2=0
cc_606 N_A_600_345#_M1020_g N_VPWR_c_1135_n 4.46264e-19 $X=3.865 $Y=1.85 $X2=0
+ $Y2=0
cc_607 N_A_600_345#_M1020_g N_A_288_47#_c_1283_n 9.13114e-19 $X=3.865 $Y=1.85
+ $X2=0 $Y2=0
cc_608 N_A_600_345#_c_831_n N_A_288_47#_c_1283_n 0.00196696f $X=3.79 $Y=1.225
+ $X2=0 $Y2=0
cc_609 N_A_600_345#_c_834_n N_A_288_47#_c_1283_n 0.00717583f $X=3.395 $Y=1.225
+ $X2=0 $Y2=0
cc_610 N_A_600_345#_M1020_g N_A_288_47#_c_1272_n 0.00424598f $X=3.865 $Y=1.85
+ $X2=0 $Y2=0
cc_611 N_A_600_345#_c_834_n N_A_288_47#_c_1272_n 0.00300039f $X=3.395 $Y=1.225
+ $X2=0 $Y2=0
cc_612 N_A_600_345#_M1020_g N_A_288_47#_c_1273_n 0.0020343f $X=3.865 $Y=1.85
+ $X2=0 $Y2=0
cc_613 N_A_600_345#_M1020_g N_A_288_47#_c_1269_n 0.0114548f $X=3.865 $Y=1.85
+ $X2=0 $Y2=0
cc_614 N_A_600_345#_c_831_n N_A_288_47#_c_1269_n 0.0117196f $X=3.79 $Y=1.225
+ $X2=0 $Y2=0
cc_615 N_A_600_345#_c_832_n N_A_288_47#_c_1269_n 0.00405971f $X=3.865 $Y=1.225
+ $X2=0 $Y2=0
cc_616 N_A_600_345#_c_833_n N_A_288_47#_c_1269_n 0.021905f $X=3.33 $Y=1.06 $X2=0
+ $Y2=0
cc_617 N_A_600_345#_c_834_n N_A_288_47#_c_1269_n 0.0454283f $X=3.395 $Y=1.225
+ $X2=0 $Y2=0
cc_618 N_A_600_345#_c_833_n N_A_288_47#_c_1270_n 0.0159402f $X=3.33 $Y=1.06
+ $X2=0 $Y2=0
cc_619 N_A_600_345#_c_835_n N_A_288_47#_c_1270_n 0.00973816f $X=3.33 $Y=0.38
+ $X2=0 $Y2=0
cc_620 N_A_600_345#_M1026_d N_A_288_47#_c_1276_n 0.00287178f $X=3 $Y=1.725 $X2=0
+ $Y2=0
cc_621 N_A_600_345#_c_834_n N_A_288_47#_c_1276_n 0.00945466f $X=3.395 $Y=1.225
+ $X2=0 $Y2=0
cc_622 N_A_600_345#_M1012_g N_A_872_316#_c_1405_n 0.0130074f $X=4.305 $Y=0.445
+ $X2=0 $Y2=0
cc_623 N_A_600_345#_c_833_n N_VGND_c_1535_n 0.00289962f $X=3.33 $Y=1.06 $X2=0
+ $Y2=0
cc_624 N_A_600_345#_c_835_n N_VGND_c_1535_n 0.0115629f $X=3.33 $Y=0.38 $X2=0
+ $Y2=0
cc_625 N_A_600_345#_M1012_g N_VGND_c_1536_n 0.00319988f $X=4.305 $Y=0.445 $X2=0
+ $Y2=0
cc_626 N_A_600_345#_M1012_g N_VGND_c_1542_n 0.00585385f $X=4.305 $Y=0.445 $X2=0
+ $Y2=0
cc_627 N_A_600_345#_c_835_n N_VGND_c_1542_n 0.0205768f $X=3.33 $Y=0.38 $X2=0
+ $Y2=0
cc_628 N_A_600_345#_M1014_d N_VGND_c_1549_n 0.0021994f $X=3.005 $Y=0.235 $X2=0
+ $Y2=0
cc_629 N_A_600_345#_M1012_g N_VGND_c_1549_n 0.0121029f $X=4.305 $Y=0.445 $X2=0
+ $Y2=0
cc_630 N_A_600_345#_c_835_n N_VGND_c_1549_n 0.0154649f $X=3.33 $Y=0.38 $X2=0
+ $Y2=0
cc_631 N_A1_M1001_g N_A_788_316#_c_1001_n 0.00368747f $X=5.225 $Y=2.165 $X2=0
+ $Y2=0
cc_632 N_A1_M1001_g N_VPWR_c_1138_n 0.00654565f $X=5.225 $Y=2.165 $X2=0 $Y2=0
cc_633 N_A1_M1001_g N_VPWR_c_1144_n 0.00585385f $X=5.225 $Y=2.165 $X2=0 $Y2=0
cc_634 N_A1_M1001_g N_VPWR_c_1135_n 0.00724353f $X=5.225 $Y=2.165 $X2=0 $Y2=0
cc_635 N_A1_M1001_g N_A_872_316#_c_1405_n 0.00559084f $X=5.225 $Y=2.165 $X2=0
+ $Y2=0
cc_636 N_A1_M1027_g N_A_872_316#_c_1405_n 0.00319248f $X=5.245 $Y=0.445 $X2=0
+ $Y2=0
cc_637 A1 N_A_872_316#_c_1405_n 0.0522563f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_638 N_A1_c_900_n N_A_872_316#_c_1405_n 0.00121304f $X=5.245 $Y=1.23 $X2=0
+ $Y2=0
cc_639 N_A1_M1001_g N_A_872_316#_c_1408_n 0.0143119f $X=5.225 $Y=2.165 $X2=0
+ $Y2=0
cc_640 A1 N_A_872_316#_c_1408_n 0.0257056f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_641 N_A1_c_900_n N_A_872_316#_c_1408_n 0.0034176f $X=5.245 $Y=1.23 $X2=0
+ $Y2=0
cc_642 N_A1_M1001_g N_A_872_316#_c_1406_n 0.00624408f $X=5.225 $Y=2.165 $X2=0
+ $Y2=0
cc_643 N_A1_M1027_g N_A_872_316#_c_1406_n 0.0100135f $X=5.245 $Y=0.445 $X2=0
+ $Y2=0
cc_644 A1 N_A_872_316#_c_1406_n 0.0454653f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_645 N_A1_M1001_g N_A_872_316#_c_1410_n 0.00579011f $X=5.225 $Y=2.165 $X2=0
+ $Y2=0
cc_646 N_A1_M1001_g N_A_872_316#_c_1455_n 0.00141938f $X=5.225 $Y=2.165 $X2=0
+ $Y2=0
cc_647 N_A1_M1027_g N_A_872_316#_c_1456_n 9.53828e-19 $X=5.245 $Y=0.445 $X2=0
+ $Y2=0
cc_648 N_A1_M1027_g N_VGND_c_1536_n 0.00461751f $X=5.245 $Y=0.445 $X2=0 $Y2=0
cc_649 A1 N_VGND_c_1536_n 0.0281027f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_650 N_A1_c_900_n N_VGND_c_1536_n 8.19449e-19 $X=5.245 $Y=1.23 $X2=0 $Y2=0
cc_651 A1 N_VGND_c_1542_n 8.41908e-19 $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_652 N_A1_M1027_g N_VGND_c_1543_n 0.00585385f $X=5.245 $Y=0.445 $X2=0 $Y2=0
cc_653 N_A1_M1027_g N_VGND_c_1549_n 0.0122213f $X=5.245 $Y=0.445 $X2=0 $Y2=0
cc_654 A1 N_VGND_c_1549_n 0.00283021f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_655 N_A0_M1024_g N_A_788_316#_c_987_n 0.021383f $X=6.805 $Y=0.445 $X2=0 $Y2=0
cc_656 A0 N_A_788_316#_c_987_n 0.00118764f $X=6.585 $Y=0.425 $X2=0 $Y2=0
cc_657 N_A0_M1021_g N_A_788_316#_M1006_g 0.030867f $X=6.825 $Y=2.165 $X2=0 $Y2=0
cc_658 N_A0_M1021_g N_A_788_316#_c_995_n 0.011716f $X=6.825 $Y=2.165 $X2=0 $Y2=0
cc_659 N_A0_M1021_g N_A_788_316#_c_996_n 0.00624325f $X=6.825 $Y=2.165 $X2=0
+ $Y2=0
cc_660 N_A0_c_939_n N_A_788_316#_c_996_n 0.00731293f $X=6.69 $Y=0.995 $X2=0
+ $Y2=0
cc_661 N_A0_c_940_n N_A_788_316#_c_996_n 0.00219554f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_662 N_A0_M1021_g N_A_788_316#_c_997_n 0.00383803f $X=6.825 $Y=2.165 $X2=0
+ $Y2=0
cc_663 N_A0_c_939_n N_A_788_316#_c_997_n 0.01487f $X=6.69 $Y=0.995 $X2=0 $Y2=0
cc_664 N_A0_M1021_g N_A_788_316#_c_998_n 0.00168903f $X=6.825 $Y=2.165 $X2=0
+ $Y2=0
cc_665 N_A0_c_939_n N_A_788_316#_c_990_n 0.0260946f $X=6.69 $Y=0.995 $X2=0 $Y2=0
cc_666 N_A0_c_940_n N_A_788_316#_c_990_n 0.00197607f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_667 N_A0_M1021_g N_A_788_316#_c_1018_n 7.65852e-19 $X=6.825 $Y=2.165 $X2=0
+ $Y2=0
cc_668 N_A0_c_939_n N_A_788_316#_c_991_n 3.13104e-19 $X=6.69 $Y=0.995 $X2=0
+ $Y2=0
cc_669 N_A0_c_940_n N_A_788_316#_c_991_n 0.0202878f $X=6.86 $Y=1.16 $X2=0 $Y2=0
cc_670 N_A0_M1021_g N_A_788_316#_c_1019_n 0.00569174f $X=6.825 $Y=2.165 $X2=0
+ $Y2=0
cc_671 N_A0_M1021_g N_VPWR_c_1139_n 0.00989024f $X=6.825 $Y=2.165 $X2=0 $Y2=0
cc_672 N_A0_M1021_g N_VPWR_c_1144_n 0.00462191f $X=6.825 $Y=2.165 $X2=0 $Y2=0
cc_673 N_A0_M1021_g N_VPWR_c_1135_n 0.00751757f $X=6.825 $Y=2.165 $X2=0 $Y2=0
cc_674 N_A0_M1021_g N_A_872_316#_c_1418_n 2.89316e-19 $X=6.825 $Y=2.165 $X2=0
+ $Y2=0
cc_675 N_A0_M1024_g N_VGND_c_1537_n 0.00886296f $X=6.805 $Y=0.445 $X2=0 $Y2=0
cc_676 A0 N_VGND_c_1537_n 0.0332811f $X=6.585 $Y=0.425 $X2=0 $Y2=0
cc_677 N_A0_M1024_g N_VGND_c_1543_n 0.00430438f $X=6.805 $Y=0.445 $X2=0 $Y2=0
cc_678 A0 N_VGND_c_1543_n 0.0109051f $X=6.585 $Y=0.425 $X2=0 $Y2=0
cc_679 N_A0_M1024_g N_VGND_c_1549_n 0.00705731f $X=6.805 $Y=0.445 $X2=0 $Y2=0
cc_680 A0 N_VGND_c_1549_n 0.0105489f $X=6.585 $Y=0.425 $X2=0 $Y2=0
cc_681 A0 A_1281_47# 0.0052103f $X=6.585 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_682 N_A_788_316#_c_1001_n N_VPWR_M1001_s 5.58164e-19 $X=6.525 $Y=2.21 $X2=0
+ $Y2=0
cc_683 N_A_788_316#_c_996_n N_VPWR_M1021_d 0.00805037f $X=7.115 $Y=1.58 $X2=0
+ $Y2=0
cc_684 N_A_788_316#_c_989_n N_VPWR_c_1138_n 0.00185641f $X=4.095 $Y=0.51 $X2=0
+ $Y2=0
cc_685 N_A_788_316#_c_1001_n N_VPWR_c_1138_n 0.0179356f $X=6.525 $Y=2.21 $X2=0
+ $Y2=0
cc_686 N_A_788_316#_c_1002_n N_VPWR_c_1138_n 0.00275185f $X=4.515 $Y=2.21 $X2=0
+ $Y2=0
cc_687 N_A_788_316#_c_1003_n N_VPWR_c_1138_n 0.00868777f $X=4.37 $Y=2.21 $X2=0
+ $Y2=0
cc_688 N_A_788_316#_M1006_g N_VPWR_c_1139_n 0.00278284f $X=7.31 $Y=1.985 $X2=0
+ $Y2=0
cc_689 N_A_788_316#_c_995_n N_VPWR_c_1139_n 0.0201657f $X=6.76 $Y=2.125 $X2=0
+ $Y2=0
cc_690 N_A_788_316#_c_996_n N_VPWR_c_1139_n 0.0133801f $X=7.115 $Y=1.58 $X2=0
+ $Y2=0
cc_691 N_A_788_316#_c_1018_n N_VPWR_c_1139_n 0.00268915f $X=6.67 $Y=2.21 $X2=0
+ $Y2=0
cc_692 N_A_788_316#_c_1019_n N_VPWR_c_1139_n 0.0113595f $X=6.76 $Y=2.21 $X2=0
+ $Y2=0
cc_693 N_A_788_316#_M1011_g N_VPWR_c_1141_n 0.0243935f $X=7.73 $Y=1.985 $X2=0
+ $Y2=0
cc_694 N_A_788_316#_c_1001_n N_VPWR_c_1144_n 0.00322607f $X=6.525 $Y=2.21 $X2=0
+ $Y2=0
cc_695 N_A_788_316#_c_1018_n N_VPWR_c_1144_n 8.0313e-19 $X=6.67 $Y=2.21 $X2=0
+ $Y2=0
cc_696 N_A_788_316#_c_1019_n N_VPWR_c_1144_n 0.0101875f $X=6.76 $Y=2.21 $X2=0
+ $Y2=0
cc_697 N_A_788_316#_c_999_n N_VPWR_c_1147_n 0.00647892f $X=4.18 $Y=2.21 $X2=0
+ $Y2=0
cc_698 N_A_788_316#_c_1001_n N_VPWR_c_1147_n 0.00125241f $X=6.525 $Y=2.21 $X2=0
+ $Y2=0
cc_699 N_A_788_316#_c_1002_n N_VPWR_c_1147_n 7.76522e-19 $X=4.515 $Y=2.21 $X2=0
+ $Y2=0
cc_700 N_A_788_316#_c_1003_n N_VPWR_c_1147_n 0.0111567f $X=4.37 $Y=2.21 $X2=0
+ $Y2=0
cc_701 N_A_788_316#_M1006_g N_VPWR_c_1148_n 0.00541763f $X=7.31 $Y=1.985 $X2=0
+ $Y2=0
cc_702 N_A_788_316#_M1011_g N_VPWR_c_1148_n 0.00421428f $X=7.73 $Y=1.985 $X2=0
+ $Y2=0
cc_703 N_A_788_316#_M1006_g N_VPWR_c_1135_n 0.00968077f $X=7.31 $Y=1.985 $X2=0
+ $Y2=0
cc_704 N_A_788_316#_M1011_g N_VPWR_c_1135_n 0.00780481f $X=7.73 $Y=1.985 $X2=0
+ $Y2=0
cc_705 N_A_788_316#_c_999_n N_VPWR_c_1135_n 0.00286413f $X=4.18 $Y=2.21 $X2=0
+ $Y2=0
cc_706 N_A_788_316#_c_1001_n N_VPWR_c_1135_n 0.17108f $X=6.525 $Y=2.21 $X2=0
+ $Y2=0
cc_707 N_A_788_316#_c_1002_n N_VPWR_c_1135_n 0.0297601f $X=4.515 $Y=2.21 $X2=0
+ $Y2=0
cc_708 N_A_788_316#_c_1003_n N_VPWR_c_1135_n 0.00197276f $X=4.37 $Y=2.21 $X2=0
+ $Y2=0
cc_709 N_A_788_316#_c_1018_n N_VPWR_c_1135_n 0.0297101f $X=6.67 $Y=2.21 $X2=0
+ $Y2=0
cc_710 N_A_788_316#_c_1019_n N_VPWR_c_1135_n 0.00215271f $X=6.76 $Y=2.21 $X2=0
+ $Y2=0
cc_711 N_A_788_316#_c_999_n N_A_288_47#_c_1272_n 0.0131455f $X=4.18 $Y=2.21
+ $X2=0 $Y2=0
cc_712 N_A_788_316#_c_1002_n N_A_288_47#_c_1272_n 7.53591e-19 $X=4.515 $Y=2.21
+ $X2=0 $Y2=0
cc_713 N_A_788_316#_c_989_n N_A_288_47#_c_1270_n 0.0987982f $X=4.095 $Y=0.51
+ $X2=0 $Y2=0
cc_714 N_A_788_316#_c_999_n N_A_288_47#_c_1277_n 8.20074e-19 $X=4.18 $Y=2.21
+ $X2=0 $Y2=0
cc_715 N_A_788_316#_c_1002_n N_A_872_316#_M1008_d 0.00107375f $X=4.515 $Y=2.21
+ $X2=0 $Y2=0
cc_716 N_A_788_316#_c_1001_n N_A_872_316#_M1022_d 0.00299297f $X=6.525 $Y=2.21
+ $X2=0 $Y2=0
cc_717 N_A_788_316#_c_989_n N_A_872_316#_c_1405_n 0.0611274f $X=4.095 $Y=0.51
+ $X2=0 $Y2=0
cc_718 N_A_788_316#_c_1001_n N_A_872_316#_c_1405_n 4.40444e-19 $X=6.525 $Y=2.21
+ $X2=0 $Y2=0
cc_719 N_A_788_316#_c_1002_n N_A_872_316#_c_1405_n 3.97141e-19 $X=4.515 $Y=2.21
+ $X2=0 $Y2=0
cc_720 N_A_788_316#_c_1003_n N_A_872_316#_c_1405_n 0.00600827f $X=4.37 $Y=2.21
+ $X2=0 $Y2=0
cc_721 N_A_788_316#_c_1001_n N_A_872_316#_c_1410_n 0.00351097f $X=6.525 $Y=2.21
+ $X2=0 $Y2=0
cc_722 N_A_788_316#_c_1001_n N_A_872_316#_c_1455_n 0.00522075f $X=6.525 $Y=2.21
+ $X2=0 $Y2=0
cc_723 N_A_788_316#_c_1001_n N_A_872_316#_c_1418_n 0.0249706f $X=6.525 $Y=2.21
+ $X2=0 $Y2=0
cc_724 N_A_788_316#_c_1018_n N_A_872_316#_c_1418_n 0.00153799f $X=6.67 $Y=2.21
+ $X2=0 $Y2=0
cc_725 N_A_788_316#_c_1019_n N_A_872_316#_c_1418_n 0.0062331f $X=6.76 $Y=2.21
+ $X2=0 $Y2=0
cc_726 N_A_788_316#_c_1001_n A_1060_369# 0.00249485f $X=6.525 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_727 N_A_788_316#_c_995_n A_1279_413# 0.00367035f $X=6.76 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_728 N_A_788_316#_c_1001_n A_1279_413# 0.00278888f $X=6.525 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_729 N_A_788_316#_c_1018_n A_1279_413# 0.00833367f $X=6.67 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_730 N_A_788_316#_c_1019_n A_1279_413# 0.00590254f $X=6.76 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_731 N_A_788_316#_M1006_g N_X_c_1505_n 0.00297963f $X=7.31 $Y=1.985 $X2=0
+ $Y2=0
cc_732 N_A_788_316#_M1011_g N_X_c_1505_n 0.0038203f $X=7.73 $Y=1.985 $X2=0 $Y2=0
cc_733 N_A_788_316#_c_996_n N_X_c_1505_n 0.0137876f $X=7.115 $Y=1.58 $X2=0 $Y2=0
cc_734 N_A_788_316#_c_991_n N_X_c_1505_n 0.00399972f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_735 N_A_788_316#_c_987_n N_X_c_1503_n 0.00379229f $X=7.31 $Y=0.995 $X2=0
+ $Y2=0
cc_736 N_A_788_316#_M1006_g N_X_c_1503_n 7.75191e-19 $X=7.31 $Y=1.985 $X2=0
+ $Y2=0
cc_737 N_A_788_316#_c_988_n N_X_c_1503_n 0.00933041f $X=7.73 $Y=0.995 $X2=0
+ $Y2=0
cc_738 N_A_788_316#_M1011_g N_X_c_1503_n 0.00938036f $X=7.73 $Y=1.985 $X2=0
+ $Y2=0
cc_739 N_A_788_316#_c_998_n N_X_c_1503_n 0.00546874f $X=7.2 $Y=1.495 $X2=0 $Y2=0
cc_740 N_A_788_316#_c_990_n N_X_c_1503_n 0.0234288f $X=7.34 $Y=1.16 $X2=0 $Y2=0
cc_741 N_A_788_316#_c_991_n N_X_c_1503_n 0.0217592f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_742 N_A_788_316#_c_988_n X 0.00932983f $X=7.73 $Y=0.995 $X2=0 $Y2=0
cc_743 N_A_788_316#_c_991_n X 0.00340328f $X=7.73 $Y=1.16 $X2=0 $Y2=0
cc_744 N_A_788_316#_M1011_g X 0.00359498f $X=7.73 $Y=1.985 $X2=0 $Y2=0
cc_745 N_A_788_316#_c_995_n X 0.00454339f $X=6.76 $Y=2.125 $X2=0 $Y2=0
cc_746 N_A_788_316#_M1006_g X 0.00459943f $X=7.31 $Y=1.985 $X2=0 $Y2=0
cc_747 N_A_788_316#_M1011_g X 0.00770132f $X=7.73 $Y=1.985 $X2=0 $Y2=0
cc_748 N_A_788_316#_M1006_g X 0.00290299f $X=7.31 $Y=1.985 $X2=0 $Y2=0
cc_749 N_A_788_316#_M1011_g X 0.00333096f $X=7.73 $Y=1.985 $X2=0 $Y2=0
cc_750 N_A_788_316#_c_990_n X 0.00153049f $X=7.34 $Y=1.16 $X2=0 $Y2=0
cc_751 N_A_788_316#_c_987_n N_VGND_c_1537_n 0.0132977f $X=7.31 $Y=0.995 $X2=0
+ $Y2=0
cc_752 N_A_788_316#_c_988_n N_VGND_c_1537_n 8.10162e-19 $X=7.73 $Y=0.995 $X2=0
+ $Y2=0
cc_753 N_A_788_316#_c_990_n N_VGND_c_1537_n 0.00961319f $X=7.34 $Y=1.16 $X2=0
+ $Y2=0
cc_754 N_A_788_316#_c_988_n N_VGND_c_1539_n 0.016039f $X=7.73 $Y=0.995 $X2=0
+ $Y2=0
cc_755 N_A_788_316#_c_989_n N_VGND_c_1542_n 0.0077748f $X=4.095 $Y=0.51 $X2=0
+ $Y2=0
cc_756 N_A_788_316#_c_987_n N_VGND_c_1544_n 0.0046653f $X=7.31 $Y=0.995 $X2=0
+ $Y2=0
cc_757 N_A_788_316#_c_988_n N_VGND_c_1544_n 0.00421428f $X=7.73 $Y=0.995 $X2=0
+ $Y2=0
cc_758 N_A_788_316#_M1019_d N_VGND_c_1549_n 0.0052901f $X=3.955 $Y=0.235 $X2=0
+ $Y2=0
cc_759 N_A_788_316#_c_987_n N_VGND_c_1549_n 0.00789179f $X=7.31 $Y=0.995 $X2=0
+ $Y2=0
cc_760 N_A_788_316#_c_988_n N_VGND_c_1549_n 0.00780481f $X=7.73 $Y=0.995 $X2=0
+ $Y2=0
cc_761 N_A_788_316#_c_989_n N_VGND_c_1549_n 0.00690003f $X=4.095 $Y=0.51 $X2=0
+ $Y2=0
cc_762 N_VPWR_c_1135_n A_193_369# 0.00441963f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_763 N_VPWR_c_1135_n N_A_288_47#_M1023_d 0.00192946f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_764 N_VPWR_c_1136_n N_A_288_47#_c_1279_n 0.00115476f $X=0.68 $Y=2.34 $X2=0
+ $Y2=0
cc_765 N_VPWR_c_1142_n N_A_288_47#_c_1279_n 0.0180901f $X=2.595 $Y=2.72 $X2=0
+ $Y2=0
cc_766 N_VPWR_c_1135_n N_A_288_47#_c_1279_n 0.00858407f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_767 N_VPWR_c_1137_n N_A_288_47#_c_1271_n 0.00423173f $X=2.715 $Y=2.22 $X2=0
+ $Y2=0
cc_768 N_VPWR_c_1142_n N_A_288_47#_c_1271_n 0.00582929f $X=2.595 $Y=2.72 $X2=0
+ $Y2=0
cc_769 N_VPWR_c_1135_n N_A_288_47#_c_1271_n 8.66284e-19 $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_770 N_VPWR_c_1137_n N_A_288_47#_c_1272_n 0.00289411f $X=2.715 $Y=2.22 $X2=0
+ $Y2=0
cc_771 N_VPWR_c_1147_n N_A_288_47#_c_1272_n 0.0172466f $X=4.755 $Y=2.72 $X2=0
+ $Y2=0
cc_772 N_VPWR_c_1135_n N_A_288_47#_c_1272_n 0.00412848f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_773 N_VPWR_M1003_d N_A_288_47#_c_1276_n 5.30843e-19 $X=2.58 $Y=1.725 $X2=0
+ $Y2=0
cc_774 N_VPWR_c_1137_n N_A_288_47#_c_1276_n 0.014737f $X=2.715 $Y=2.22 $X2=0
+ $Y2=0
cc_775 N_VPWR_c_1142_n N_A_288_47#_c_1276_n 0.00180834f $X=2.595 $Y=2.72 $X2=0
+ $Y2=0
cc_776 N_VPWR_c_1147_n N_A_288_47#_c_1276_n 0.00243737f $X=4.755 $Y=2.72 $X2=0
+ $Y2=0
cc_777 N_VPWR_c_1135_n N_A_288_47#_c_1276_n 0.093852f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_778 N_VPWR_c_1137_n N_A_288_47#_c_1316_n 0.00163392f $X=2.715 $Y=2.22 $X2=0
+ $Y2=0
cc_779 N_VPWR_c_1142_n N_A_288_47#_c_1316_n 8.27583e-19 $X=2.595 $Y=2.72 $X2=0
+ $Y2=0
cc_780 N_VPWR_c_1135_n N_A_288_47#_c_1316_n 0.0298306f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_781 N_VPWR_c_1137_n N_A_288_47#_c_1277_n 0.00250319f $X=2.715 $Y=2.22 $X2=0
+ $Y2=0
cc_782 N_VPWR_c_1147_n N_A_288_47#_c_1277_n 8.27838e-19 $X=4.755 $Y=2.72 $X2=0
+ $Y2=0
cc_783 N_VPWR_c_1135_n N_A_288_47#_c_1277_n 0.0296902f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_784 N_VPWR_c_1135_n A_372_413# 0.00300836f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_785 N_VPWR_c_1135_n N_A_872_316#_M1022_d 0.00130544f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_786 N_VPWR_c_1138_n N_A_872_316#_c_1408_n 0.0125871f $X=5.015 $Y=2.24 $X2=0
+ $Y2=0
cc_787 N_VPWR_c_1138_n N_A_872_316#_c_1410_n 3.9298e-19 $X=5.015 $Y=2.24 $X2=0
+ $Y2=0
cc_788 N_VPWR_c_1138_n N_A_872_316#_c_1455_n 0.00347614f $X=5.015 $Y=2.24 $X2=0
+ $Y2=0
cc_789 N_VPWR_c_1144_n N_A_872_316#_c_1455_n 0.00567337f $X=7.015 $Y=2.72 $X2=0
+ $Y2=0
cc_790 N_VPWR_c_1135_n N_A_872_316#_c_1455_n 0.00186252f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_791 N_VPWR_c_1144_n N_A_872_316#_c_1418_n 0.0233641f $X=7.015 $Y=2.72 $X2=0
+ $Y2=0
cc_792 N_VPWR_c_1135_n N_A_872_316#_c_1418_n 0.00706654f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_793 N_VPWR_c_1135_n A_1060_369# 0.00267305f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_794 N_VPWR_c_1135_n A_1279_413# 0.00221859f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_795 N_VPWR_c_1135_n N_X_M1006_s 0.00215535f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_796 N_VPWR_c_1141_n N_X_c_1505_n 0.0735075f $X=8.02 $Y=1.66 $X2=0 $Y2=0
cc_797 N_VPWR_c_1148_n X 0.0228774f $X=7.935 $Y=2.72 $X2=0 $Y2=0
cc_798 N_VPWR_c_1135_n X 0.0148499f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_799 N_VPWR_c_1141_n N_VGND_c_1539_n 0.0086927f $X=8.02 $Y=1.66 $X2=0 $Y2=0
cc_800 N_A_288_47#_c_1279_n A_372_413# 0.0041168f $X=2.07 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_801 N_A_288_47#_c_1271_n A_372_413# 0.0134763f $X=2.155 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_802 N_A_288_47#_c_1276_n A_372_413# 0.00266219f $X=3.305 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_803 N_A_288_47#_c_1316_n A_372_413# 0.00398835f $X=2.215 $Y=2.21 $X2=-0.19
+ $Y2=-0.24
cc_804 N_A_288_47#_c_1280_n N_VGND_c_1535_n 0.00748073f $X=1.9 $Y=0.45 $X2=0
+ $Y2=0
cc_805 N_A_288_47#_c_1267_n N_VGND_c_1535_n 3.77264e-19 $X=1.985 $Y=1.235 $X2=0
+ $Y2=0
cc_806 N_A_288_47#_c_1280_n N_VGND_c_1541_n 0.0202971f $X=1.9 $Y=0.45 $X2=0
+ $Y2=0
cc_807 N_A_288_47#_c_1270_n N_VGND_c_1542_n 0.00895969f $X=3.67 $Y=0.51 $X2=0
+ $Y2=0
cc_808 N_A_288_47#_M1004_d N_VGND_c_1549_n 0.00348335f $X=1.44 $Y=0.235 $X2=0
+ $Y2=0
cc_809 N_A_288_47#_M1019_s N_VGND_c_1549_n 0.00264447f $X=3.545 $Y=0.235 $X2=0
+ $Y2=0
cc_810 N_A_288_47#_c_1280_n N_VGND_c_1549_n 0.0203474f $X=1.9 $Y=0.45 $X2=0
+ $Y2=0
cc_811 N_A_288_47#_c_1270_n N_VGND_c_1549_n 0.00841871f $X=3.67 $Y=0.51 $X2=0
+ $Y2=0
cc_812 N_A_288_47#_c_1280_n A_397_47# 0.00244815f $X=1.9 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_813 N_A_288_47#_c_1267_n A_397_47# 0.00145797f $X=1.985 $Y=1.235 $X2=-0.19
+ $Y2=-0.24
cc_814 N_A_872_316#_c_1410_n A_1060_369# 0.00496775f $X=5.41 $Y=2.155 $X2=-0.19
+ $Y2=-0.24
cc_815 N_A_872_316#_c_1455_n A_1060_369# 0.00306462f $X=5.495 $Y=2.24 $X2=-0.19
+ $Y2=-0.24
cc_816 N_A_872_316#_c_1418_n A_1060_369# 0.00812168f $X=6.11 $Y=2.24 $X2=-0.19
+ $Y2=-0.24
cc_817 N_A_872_316#_c_1456_n N_VGND_c_1536_n 0.0207476f $X=4.515 $Y=0.42 $X2=0
+ $Y2=0
cc_818 N_A_872_316#_c_1456_n N_VGND_c_1542_n 0.0127262f $X=4.515 $Y=0.42 $X2=0
+ $Y2=0
cc_819 N_A_872_316#_c_1482_p N_VGND_c_1543_n 0.0080925f $X=5.495 $Y=0.38 $X2=0
+ $Y2=0
cc_820 N_A_872_316#_c_1417_n N_VGND_c_1543_n 0.0333963f $X=6.055 $Y=0.38 $X2=0
+ $Y2=0
cc_821 N_A_872_316#_M1012_d N_VGND_c_1549_n 0.00403727f $X=4.38 $Y=0.235 $X2=0
+ $Y2=0
cc_822 N_A_872_316#_M1015_d N_VGND_c_1549_n 0.00340843f $X=5.855 $Y=0.235 $X2=0
+ $Y2=0
cc_823 N_A_872_316#_c_1482_p N_VGND_c_1549_n 0.00641762f $X=5.495 $Y=0.38 $X2=0
+ $Y2=0
cc_824 N_A_872_316#_c_1417_n N_VGND_c_1549_n 0.0256442f $X=6.055 $Y=0.38 $X2=0
+ $Y2=0
cc_825 N_A_872_316#_c_1456_n N_VGND_c_1549_n 0.00779458f $X=4.515 $Y=0.42 $X2=0
+ $Y2=0
cc_826 N_A_872_316#_c_1406_n A_1064_47# 0.00347944f $X=5.41 $Y=1.565 $X2=-0.19
+ $Y2=-0.24
cc_827 N_A_872_316#_c_1482_p A_1064_47# 0.00236827f $X=5.495 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_828 N_A_872_316#_c_1417_n A_1064_47# 0.00762432f $X=6.055 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_829 N_X_c_1503_n N_VGND_c_1537_n 0.00173729f $X=7.61 $Y=1.495 $X2=0 $Y2=0
cc_830 X N_VGND_c_1539_n 0.0469672f $X=7.505 $Y=0.425 $X2=0 $Y2=0
cc_831 X N_VGND_c_1544_n 0.019081f $X=7.505 $Y=0.425 $X2=0 $Y2=0
cc_832 N_X_M1009_s N_VGND_c_1549_n 0.00389051f $X=7.385 $Y=0.235 $X2=0 $Y2=0
cc_833 X N_VGND_c_1549_n 0.0119356f $X=7.505 $Y=0.425 $X2=0 $Y2=0
cc_834 N_VGND_c_1549_n A_193_47# 0.00497208f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_835 N_VGND_c_1549_n A_397_47# 0.0089813f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_836 N_VGND_c_1549_n A_1064_47# 0.00329874f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_837 N_VGND_c_1549_n A_1281_47# 0.00726162f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a31o_4.spice.SKY130_FD_SC_HD__A31O_4.pxi
* Created: Thu Aug 27 14:04:49 2020
* 
x_PM_SKY130_FD_SC_HD__A31O_4%A3 N_A3_M1021_g N_A3_M1005_g N_A3_M1023_g
+ N_A3_M1012_g N_A3_c_108_n N_A3_c_100_n N_A3_c_101_n A3 A3 N_A3_c_102_n
+ N_A3_c_103_n N_A3_c_104_n N_A3_c_105_n PM_SKY130_FD_SC_HD__A31O_4%A3
x_PM_SKY130_FD_SC_HD__A31O_4%A2 N_A2_c_191_n N_A2_M1008_g N_A2_M1003_g
+ N_A2_c_192_n N_A2_M1018_g N_A2_M1014_g N_A2_c_193_n N_A2_c_194_n N_A2_c_215_n
+ N_A2_c_195_n N_A2_c_196_n A2 A2 N_A2_c_198_n N_A2_c_199_n N_A2_c_253_p
+ PM_SKY130_FD_SC_HD__A31O_4%A2
x_PM_SKY130_FD_SC_HD__A31O_4%A1 N_A1_M1011_g N_A1_M1002_g N_A1_M1010_g
+ N_A1_M1020_g A1 N_A1_c_283_n PM_SKY130_FD_SC_HD__A31O_4%A1
x_PM_SKY130_FD_SC_HD__A31O_4%B1 N_B1_c_324_n N_B1_M1004_g N_B1_M1000_g
+ N_B1_c_325_n N_B1_M1022_g N_B1_M1006_g N_B1_c_326_n B1 B1 N_B1_c_328_n
+ N_B1_c_329_n PM_SKY130_FD_SC_HD__A31O_4%B1
x_PM_SKY130_FD_SC_HD__A31O_4%A_277_47# N_A_277_47#_M1011_s N_A_277_47#_M1004_d
+ N_A_277_47#_M1000_d N_A_277_47#_c_388_n N_A_277_47#_M1013_g
+ N_A_277_47#_M1001_g N_A_277_47#_c_389_n N_A_277_47#_M1015_g
+ N_A_277_47#_M1007_g N_A_277_47#_c_390_n N_A_277_47#_M1016_g
+ N_A_277_47#_M1009_g N_A_277_47#_c_391_n N_A_277_47#_M1017_g
+ N_A_277_47#_M1019_g N_A_277_47#_c_416_n N_A_277_47#_c_404_n
+ N_A_277_47#_c_407_n N_A_277_47#_c_392_n N_A_277_47#_c_412_n
+ N_A_277_47#_c_400_n N_A_277_47#_c_393_n N_A_277_47#_c_487_p
+ N_A_277_47#_c_394_n N_A_277_47#_c_413_n N_A_277_47#_c_450_n
+ N_A_277_47#_c_403_n PM_SKY130_FD_SC_HD__A31O_4%A_277_47#
x_PM_SKY130_FD_SC_HD__A31O_4%A_27_297# N_A_27_297#_M1005_d N_A_27_297#_M1003_d
+ N_A_27_297#_M1020_s N_A_27_297#_M1012_d N_A_27_297#_M1006_s
+ N_A_27_297#_c_544_n N_A_27_297#_c_547_n N_A_27_297#_c_548_n
+ N_A_27_297#_c_551_n N_A_27_297#_c_560_n N_A_27_297#_c_580_p
+ N_A_27_297#_c_567_n N_A_27_297#_c_552_n N_A_27_297#_c_554_n
+ N_A_27_297#_c_555_n PM_SKY130_FD_SC_HD__A31O_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A31O_4%VPWR N_VPWR_M1005_s N_VPWR_M1002_d N_VPWR_M1014_s
+ N_VPWR_M1001_s N_VPWR_M1007_s N_VPWR_M1019_s N_VPWR_c_596_n N_VPWR_c_597_n
+ N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n
+ N_VPWR_c_603_n N_VPWR_c_604_n N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n
+ N_VPWR_c_608_n N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n VPWR
+ N_VPWR_c_612_n N_VPWR_c_613_n N_VPWR_c_595_n N_VPWR_c_615_n
+ PM_SKY130_FD_SC_HD__A31O_4%VPWR
x_PM_SKY130_FD_SC_HD__A31O_4%X N_X_M1013_s N_X_M1016_s N_X_M1001_d N_X_M1009_d
+ N_X_c_711_n N_X_c_715_n N_X_c_718_n X X X X N_X_c_707_n X
+ PM_SKY130_FD_SC_HD__A31O_4%X
x_PM_SKY130_FD_SC_HD__A31O_4%VGND N_VGND_M1021_d N_VGND_M1023_d N_VGND_M1022_s
+ N_VGND_M1015_d N_VGND_M1017_d N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n
+ N_VGND_c_761_n N_VGND_c_762_n N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n
+ N_VGND_c_766_n N_VGND_c_767_n N_VGND_c_768_n VGND N_VGND_c_769_n
+ N_VGND_c_770_n N_VGND_c_771_n N_VGND_c_772_n PM_SKY130_FD_SC_HD__A31O_4%VGND
cc_1 VNB N_A3_c_100_n 0.00394903f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.16
cc_2 VNB N_A3_c_101_n 0.0198644f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.16
cc_3 VNB N_A3_c_102_n 0.031696f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_4 VNB N_A3_c_103_n 0.0101544f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_5 VNB N_A3_c_104_n 0.0216903f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=0.995
cc_6 VNB N_A3_c_105_n 0.0173116f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=0.995
cc_7 VNB N_A2_c_191_n 0.0151526f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_A2_c_192_n 0.0163642f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=0.995
cc_9 VNB N_A2_c_193_n 0.00183228f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.53
cc_10 VNB N_A2_c_194_n 0.00799885f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.445
cc_11 VNB N_A2_c_195_n 0.00408923f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.16
cc_12 VNB N_A2_c_196_n 0.0212658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB A2 0.00173313f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_14 VNB N_A2_c_198_n 0.0203822f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.325
cc_15 VNB N_A2_c_199_n 0.00382732f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.16
cc_16 VNB N_A1_M1011_g 0.0174436f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_17 VNB N_A1_M1002_g 4.44034e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_M1010_g 0.0174371f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=1.325
cc_19 VNB N_A1_M1020_g 4.44034e-19 $X=-0.19 $Y=-0.24 $X2=2.525 $Y2=1.53
cc_20 VNB N_A1_c_283_n 0.0296083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B1_c_324_n 0.0163199f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_22 VNB N_B1_c_325_n 0.0193103f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=0.995
cc_23 VNB N_B1_c_326_n 0.027613f $X=-0.19 $Y=-0.24 $X2=2.525 $Y2=1.53
cc_24 VNB B1 0.00341511f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.16
cc_25 VNB N_B1_c_328_n 0.0321487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B1_c_329_n 0.0029435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_277_47#_c_388_n 0.0196354f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=0.56
cc_28 VNB N_A_277_47#_c_389_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.445
cc_29 VNB N_A_277_47#_c_390_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_277_47#_c_391_n 0.018648f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.16
cc_31 VNB N_A_277_47#_c_392_n 9.28168e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_277_47#_c_393_n 0.00801713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_277_47#_c_394_n 0.0798337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_595_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB X 0.00295327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_707_n 0.0103056f $X=-0.19 $Y=-0.24 $X2=0.337 $Y2=1.19
cc_37 VNB X 0.0231598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_758_n 0.0110531f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.53
cc_39 VNB N_VGND_c_759_n 0.00680105f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.16
cc_40 VNB N_VGND_c_760_n 0.00265724f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_41 VNB N_VGND_c_761_n 3.27478e-19 $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_42 VNB N_VGND_c_762_n 0.0126456f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.325
cc_43 VNB N_VGND_c_763_n 0.0627995f $X=-0.19 $Y=-0.24 $X2=2.69 $Y2=1.325
cc_44 VNB N_VGND_c_764_n 0.00435829f $X=-0.19 $Y=-0.24 $X2=0.337 $Y2=1.16
cc_45 VNB N_VGND_c_765_n 0.0184104f $X=-0.19 $Y=-0.24 $X2=0.337 $Y2=1.19
cc_46 VNB N_VGND_c_766_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_767_n 0.011903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_768_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_769_n 0.0203086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_770_n 0.0119952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_771_n 0.319183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_772_n 0.0164282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_A3_M1005_g 0.0228245f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_54 VPB N_A3_M1012_g 0.0185778f $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.985
cc_55 VPB N_A3_c_108_n 0.0205416f $X=-0.19 $Y=1.305 $X2=2.525 $Y2=1.53
cc_56 VPB N_A3_c_100_n 0.00262354f $X=-0.19 $Y=1.305 $X2=2.69 $Y2=1.16
cc_57 VPB N_A3_c_101_n 0.00446581f $X=-0.19 $Y=1.305 $X2=2.69 $Y2=1.16
cc_58 VPB N_A3_c_102_n 0.00644551f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_59 VPB N_A3_c_103_n 0.00681416f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_60 VPB N_A2_M1003_g 0.018381f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_A2_M1014_g 0.0190115f $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.985
cc_62 VPB N_A2_c_196_n 0.00406366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A2_c_198_n 0.00411157f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.325
cc_64 VPB N_A1_M1002_g 0.0192155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A1_M1020_g 0.0192155f $X=-0.19 $Y=1.305 $X2=2.525 $Y2=1.53
cc_66 VPB N_B1_M1000_g 0.0187402f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_B1_M1006_g 0.0230839f $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.985
cc_68 VPB N_B1_c_326_n 0.00469308f $X=-0.19 $Y=1.305 $X2=2.525 $Y2=1.53
cc_69 VPB N_A_277_47#_M1001_g 0.0209439f $X=-0.19 $Y=1.305 $X2=2.525 $Y2=1.53
cc_70 VPB N_A_277_47#_M1007_g 0.0182696f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_71 VPB N_A_277_47#_M1009_g 0.0182793f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=0.995
cc_72 VPB N_A_277_47#_M1019_g 0.021532f $X=-0.19 $Y=1.305 $X2=0.337 $Y2=1.19
cc_73 VPB N_A_277_47#_c_392_n 0.00121211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_277_47#_c_400_n 0.0199067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_277_47#_c_393_n 0.00365242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_277_47#_c_394_n 0.0190404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_277_47#_c_403_n 0.00151257f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_596_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_597_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_598_n 0.00271082f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=0.995
cc_81 VPB N_VPWR_c_599_n 0.00694843f $X=-0.19 $Y=1.305 $X2=2.69 $Y2=1.325
cc_82 VPB N_VPWR_c_600_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_601_n 0.00272466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_602_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_603_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_604_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_605_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_606_n 0.0401329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_607_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_608_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_609_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_610_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_611_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_612_n 0.0159043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_613_n 0.0128037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_595_n 0.0567464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_615_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB X 0.00915601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 N_A3_c_104_n N_A2_c_191_n 0.0420887f $X=0.385 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_100 N_A3_M1005_g N_A2_M1003_g 0.0429906f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A3_c_108_n N_A2_M1003_g 0.0104551f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_102 N_A3_c_103_n N_A2_M1003_g 8.27705e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A3_c_105_n N_A2_c_192_n 0.0309828f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A3_M1012_g N_A2_M1014_g 0.0335848f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A3_c_108_n N_A2_M1014_g 0.0106172f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_106 N_A3_c_100_n N_A2_M1014_g 0.00245189f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A3_c_102_n N_A2_c_193_n 5.05982e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A3_c_104_n N_A2_c_193_n 0.00164339f $X=0.385 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A3_c_108_n N_A2_c_194_n 0.0179673f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_110 N_A3_c_104_n N_A2_c_215_n 5.81733e-19 $X=0.385 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A3_c_108_n N_A2_c_195_n 0.0214436f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_112 N_A3_c_102_n N_A2_c_195_n 0.00100418f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A3_c_103_n N_A2_c_195_n 0.0120224f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A3_c_108_n N_A2_c_196_n 0.00289889f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_115 N_A3_c_102_n N_A2_c_196_n 0.0213019f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A3_c_103_n N_A2_c_196_n 7.27926e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A3_c_105_n A2 9.10852e-19 $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A3_c_108_n N_A2_c_198_n 0.00285374f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_119 N_A3_c_100_n N_A2_c_198_n 0.0017953f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A3_c_101_n N_A2_c_198_n 0.0158737f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A3_c_108_n N_A2_c_199_n 0.0235556f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_122 N_A3_c_100_n N_A2_c_199_n 0.0142658f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A3_c_101_n N_A2_c_199_n 6.7729e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A3_c_108_n N_A1_M1002_g 0.0117787f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_125 N_A3_c_108_n N_A1_M1020_g 0.0115361f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_126 N_A3_c_108_n A1 0.0250371f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_127 N_A3_c_108_n N_A1_c_283_n 0.00198252f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_128 N_A3_c_105_n N_B1_c_324_n 0.0207775f $X=2.69 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_129 N_A3_M1012_g N_B1_M1000_g 0.0202313f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A3_c_108_n N_B1_M1000_g 0.00149396f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_131 N_A3_c_100_n N_B1_c_326_n 0.00289249f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A3_c_101_n N_B1_c_326_n 0.0223158f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A3_c_100_n N_A_277_47#_c_404_n 0.0190485f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A3_c_101_n N_A_277_47#_c_404_n 0.0027274f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A3_c_105_n N_A_277_47#_c_404_n 0.01126f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A3_c_105_n N_A_277_47#_c_407_n 4.61731e-19 $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A3_c_108_n N_A_277_47#_c_392_n 5.11068e-19 $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_138 N_A3_c_100_n N_A_277_47#_c_392_n 0.0184215f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A3_c_101_n N_A_277_47#_c_392_n 6.86012e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A3_c_105_n N_A_277_47#_c_392_n 5.98576e-19 $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A3_M1012_g N_A_277_47#_c_412_n 6.98201e-19 $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A3_c_108_n N_A_277_47#_c_413_n 0.005232f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_143 N_A3_c_108_n N_A_277_47#_c_403_n 0.00906828f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_144 N_A3_c_103_n N_A_27_297#_M1005_d 0.00869141f $X=0.36 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_145 N_A3_c_108_n N_A_27_297#_M1003_d 0.00165831f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_146 N_A3_c_108_n N_A_27_297#_M1020_s 0.00165831f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_147 N_A3_c_108_n N_A_27_297#_M1012_d 0.00244577f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_148 N_A3_M1005_g N_A_27_297#_c_544_n 0.00930137f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A3_c_108_n N_A_27_297#_c_544_n 0.0228196f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_150 N_A3_c_103_n N_A_27_297#_c_544_n 0.00960524f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A3_c_108_n N_A_27_297#_c_547_n 0.0315971f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_152 N_A3_M1012_g N_A_27_297#_c_548_n 0.00989364f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A3_c_108_n N_A_27_297#_c_548_n 0.041192f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_154 N_A3_c_101_n N_A_27_297#_c_548_n 3.3535e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A3_c_108_n N_A_27_297#_c_551_n 0.00354737f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_156 N_A3_c_102_n N_A_27_297#_c_552_n 4.91121e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A3_c_103_n N_A_27_297#_c_552_n 0.0144494f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A3_c_108_n N_A_27_297#_c_554_n 0.0126919f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_159 N_A3_c_108_n N_A_27_297#_c_555_n 0.0126919f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_160 N_A3_c_108_n N_VPWR_M1005_s 0.00166235f $X=2.525 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A3_c_108_n N_VPWR_M1002_d 0.00166235f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_162 N_A3_c_108_n N_VPWR_M1014_s 0.00230172f $X=2.525 $Y=1.53 $X2=0 $Y2=0
cc_163 N_A3_M1005_g N_VPWR_c_596_n 0.0106557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A3_M1012_g N_VPWR_c_598_n 0.00348971f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A3_M1012_g N_VPWR_c_606_n 0.00585385f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A3_M1005_g N_VPWR_c_612_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A3_M1005_g N_VPWR_c_595_n 0.00515525f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A3_M1012_g N_VPWR_c_595_n 0.00632196f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A3_c_102_n N_VGND_c_759_n 0.00305311f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A3_c_103_n N_VGND_c_759_n 0.0149476f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A3_c_104_n N_VGND_c_759_n 0.004898f $X=0.385 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A3_c_105_n N_VGND_c_760_n 0.00802411f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A3_c_104_n N_VGND_c_763_n 0.00585385f $X=0.385 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A3_c_105_n N_VGND_c_763_n 0.00419163f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A3_c_104_n N_VGND_c_771_n 0.0115954f $X=0.385 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A3_c_105_n N_VGND_c_771_n 0.00502958f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A2_c_191_n N_A1_M1011_g 0.0440811f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A2_c_193_n N_A1_M1011_g 0.00215578f $X=0.89 $Y=1.075 $X2=0 $Y2=0
cc_179 N_A2_c_194_n N_A1_M1011_g 0.0132056f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_180 N_A2_c_196_n N_A1_M1011_g 0.0221481f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A2_M1003_g N_A1_M1002_g 0.0284553f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A2_c_192_n N_A1_M1010_g 0.0433403f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_c_194_n N_A1_M1010_g 0.0115242f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_184 A2 N_A1_M1010_g 0.0034855f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_185 N_A2_c_198_n N_A1_M1010_g 0.021619f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_M1014_g N_A1_M1020_g 0.0284553f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A2_c_194_n A1 0.0250368f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_188 N_A2_c_195_n A1 0.00882575f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A2_c_196_n A1 3.26244e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A2_c_198_n A1 2.05292e-19 $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A2_c_199_n A1 0.0109198f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A2_c_194_n N_A1_c_283_n 0.00205431f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_193 N_A2_c_195_n N_A1_c_283_n 0.00130712f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A2_c_199_n N_A1_c_283_n 0.00145631f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A2_c_194_n N_A_277_47#_M1011_s 0.00162389f $X=1.985 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A2_c_191_n N_A_277_47#_c_416_n 8.22884e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_192_n N_A_277_47#_c_416_n 0.0104605f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_194_n N_A_277_47#_c_416_n 0.0311938f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_199 N_A2_c_198_n N_A_277_47#_c_416_n 0.00109245f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A2_c_199_n N_A_277_47#_c_416_n 0.00349402f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A2_c_253_p N_A_277_47#_c_416_n 0.00903247f $X=2.077 $Y=0.905 $X2=0
+ $Y2=0
cc_202 N_A2_c_192_n N_A_277_47#_c_413_n 0.00498236f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A2_c_253_p N_A_277_47#_c_413_n 0.0101484f $X=2.077 $Y=0.905 $X2=0 $Y2=0
cc_204 N_A2_M1003_g N_A_27_297#_c_544_n 0.00932032f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A2_M1014_g N_A_27_297#_c_548_n 0.00965817f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A2_M1003_g N_VPWR_c_596_n 0.00889341f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A2_M1003_g N_VPWR_c_597_n 5.47116e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A2_M1014_g N_VPWR_c_597_n 5.47116e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A2_M1014_g N_VPWR_c_598_n 0.00893525f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A2_M1003_g N_VPWR_c_602_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A2_M1014_g N_VPWR_c_604_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A2_M1003_g N_VPWR_c_595_n 0.00422825f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A2_M1014_g N_VPWR_c_595_n 0.00422825f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A2_c_215_n N_VGND_c_759_n 7.99711e-19 $X=0.975 $Y=0.82 $X2=0 $Y2=0
cc_215 N_A2_c_192_n N_VGND_c_760_n 0.00164507f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A2_c_191_n N_VGND_c_763_n 0.00439071f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A2_c_192_n N_VGND_c_763_n 0.00385416f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A2_c_194_n N_VGND_c_763_n 0.00457298f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_219 N_A2_c_215_n N_VGND_c_763_n 0.00227506f $X=0.975 $Y=0.82 $X2=0 $Y2=0
cc_220 N_A2_c_191_n N_VGND_c_771_n 0.0061773f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A2_c_192_n N_VGND_c_771_n 0.00558582f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_194_n N_VGND_c_771_n 0.0103392f $X=1.985 $Y=0.82 $X2=0 $Y2=0
cc_223 N_A2_c_215_n N_VGND_c_771_n 0.00391846f $X=0.975 $Y=0.82 $X2=0 $Y2=0
cc_224 N_A2_c_194_n A_193_47# 0.00302426f $X=1.985 $Y=0.82 $X2=-0.19 $Y2=-0.24
cc_225 N_A2_c_194_n A_361_47# 0.00126997f $X=1.985 $Y=0.82 $X2=-0.19 $Y2=-0.24
cc_226 N_A2_c_253_p A_361_47# 3.39504e-19 $X=2.077 $Y=0.905 $X2=-0.19 $Y2=-0.24
cc_227 N_A1_M1011_g N_A_277_47#_c_416_n 0.00417689f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A1_M1010_g N_A_277_47#_c_416_n 0.00847015f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A1_M1002_g N_A_27_297#_c_547_n 0.00936448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A1_M1020_g N_A_27_297#_c_547_n 0.00936448f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_M1002_g N_VPWR_c_596_n 5.47116e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A1_M1002_g N_VPWR_c_597_n 0.00894861f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_M1020_g N_VPWR_c_597_n 0.00894861f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A1_M1020_g N_VPWR_c_598_n 5.47116e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A1_M1002_g N_VPWR_c_602_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A1_M1020_g N_VPWR_c_604_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A1_M1002_g N_VPWR_c_595_n 0.00422825f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A1_M1020_g N_VPWR_c_595_n 0.00422825f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A1_M1011_g N_VGND_c_763_n 0.00428448f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_240 N_A1_M1010_g N_VGND_c_763_n 0.00385416f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_241 N_A1_M1011_g N_VGND_c_771_n 0.00600354f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_242 N_A1_M1010_g N_VGND_c_771_n 0.00541157f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_243 B1 N_A_277_47#_c_388_n 0.00628191f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_244 N_B1_c_324_n N_A_277_47#_c_404_n 0.0123226f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_245 N_B1_c_324_n N_A_277_47#_c_407_n 0.00609246f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B1_c_325_n N_A_277_47#_c_407_n 0.00968387f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B1_c_324_n N_A_277_47#_c_392_n 0.00306393f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B1_M1000_g N_A_277_47#_c_392_n 0.00269003f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B1_c_325_n N_A_277_47#_c_392_n 0.00116425f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B1_M1006_g N_A_277_47#_c_392_n 0.00291926f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B1_c_326_n N_A_277_47#_c_392_n 0.0197363f $X=3.605 $Y=1.16 $X2=0 $Y2=0
cc_252 B1 N_A_277_47#_c_392_n 0.00724458f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_253 N_B1_c_329_n N_A_277_47#_c_392_n 0.0121165f $X=3.922 $Y=1.18 $X2=0 $Y2=0
cc_254 N_B1_M1000_g N_A_277_47#_c_412_n 0.00706389f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B1_M1006_g N_A_277_47#_c_412_n 0.0114396f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_256 N_B1_M1006_g N_A_277_47#_c_400_n 0.0135958f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_257 N_B1_c_328_n N_A_277_47#_c_400_n 0.00651143f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B1_c_329_n N_A_277_47#_c_400_n 0.0333911f $X=3.922 $Y=1.18 $X2=0 $Y2=0
cc_259 N_B1_M1006_g N_A_277_47#_c_393_n 3.20984e-19 $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_260 N_B1_c_326_n N_A_277_47#_c_393_n 0.00356099f $X=3.605 $Y=1.16 $X2=0 $Y2=0
cc_261 B1 N_A_277_47#_c_393_n 0.00556902f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_262 N_B1_c_328_n N_A_277_47#_c_393_n 9.20525e-19 $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B1_c_329_n N_A_277_47#_c_393_n 0.0154251f $X=3.922 $Y=1.18 $X2=0 $Y2=0
cc_264 B1 N_A_277_47#_c_394_n 2.92178e-19 $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_265 N_B1_c_328_n N_A_277_47#_c_394_n 0.00632652f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_266 N_B1_c_329_n N_A_277_47#_c_394_n 6.55257e-19 $X=3.922 $Y=1.18 $X2=0 $Y2=0
cc_267 N_B1_c_324_n N_A_277_47#_c_450_n 4.64231e-19 $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B1_c_325_n N_A_277_47#_c_450_n 0.00382839f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B1_c_326_n N_A_277_47#_c_450_n 5.69051e-19 $X=3.605 $Y=1.16 $X2=0 $Y2=0
cc_270 B1 N_A_277_47#_c_450_n 0.0053915f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_271 N_B1_M1000_g N_A_277_47#_c_403_n 0.0027147f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B1_M1006_g N_A_277_47#_c_403_n 0.00161189f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B1_c_326_n N_A_277_47#_c_403_n 6.27456e-19 $X=3.605 $Y=1.16 $X2=0 $Y2=0
cc_274 N_B1_M1000_g N_A_27_297#_c_560_n 0.0112555f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B1_M1006_g N_A_27_297#_c_560_n 0.00938455f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B1_M1006_g N_VPWR_c_599_n 0.00235209f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B1_M1000_g N_VPWR_c_606_n 0.00357877f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B1_M1006_g N_VPWR_c_606_n 0.00357877f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B1_M1000_g N_VPWR_c_595_n 0.00539297f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B1_M1006_g N_VPWR_c_595_n 0.00655123f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_281 B1 X 0.00283121f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_282 B1 N_VGND_M1022_s 0.00718281f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_283 N_B1_c_324_n N_VGND_c_760_n 0.00292297f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B1_c_324_n N_VGND_c_769_n 0.00422176f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B1_c_325_n N_VGND_c_769_n 0.00542953f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B1_c_324_n N_VGND_c_771_n 0.00583754f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B1_c_325_n N_VGND_c_771_n 0.01108f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_288 B1 N_VGND_c_771_n 8.53685e-19 $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_289 N_B1_c_325_n N_VGND_c_772_n 0.0124359f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_290 B1 N_VGND_c_772_n 0.0167504f $X=3.83 $Y=0.765 $X2=0 $Y2=0
cc_291 N_B1_c_328_n N_VGND_c_772_n 0.00189644f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B1_c_329_n N_VGND_c_772_n 0.00275659f $X=3.922 $Y=1.18 $X2=0 $Y2=0
cc_293 N_A_277_47#_c_400_n N_A_27_297#_M1006_s 0.00390196f $X=4.225 $Y=1.54
+ $X2=0 $Y2=0
cc_294 N_A_277_47#_M1000_d N_A_27_297#_c_560_n 0.00316374f $X=3.185 $Y=1.485
+ $X2=0 $Y2=0
cc_295 N_A_277_47#_M1001_g N_A_27_297#_c_560_n 5.09561e-19 $X=4.47 $Y=1.985
+ $X2=0 $Y2=0
cc_296 N_A_277_47#_c_412_n N_A_27_297#_c_560_n 0.015159f $X=3.32 $Y=1.63 $X2=0
+ $Y2=0
cc_297 N_A_277_47#_c_400_n N_A_27_297#_c_560_n 0.00256303f $X=4.225 $Y=1.54
+ $X2=0 $Y2=0
cc_298 N_A_277_47#_M1001_g N_A_27_297#_c_567_n 0.00622395f $X=4.47 $Y=1.985
+ $X2=0 $Y2=0
cc_299 N_A_277_47#_c_400_n N_A_27_297#_c_567_n 0.0131641f $X=4.225 $Y=1.54 $X2=0
+ $Y2=0
cc_300 N_A_277_47#_c_400_n N_VPWR_M1001_s 0.00259685f $X=4.225 $Y=1.54 $X2=0
+ $Y2=0
cc_301 N_A_277_47#_c_393_n N_VPWR_M1001_s 0.00324062f $X=4.395 $Y=1.16 $X2=0
+ $Y2=0
cc_302 N_A_277_47#_M1001_g N_VPWR_c_599_n 0.0117895f $X=4.47 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_277_47#_M1007_g N_VPWR_c_599_n 5.47116e-19 $X=4.89 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_A_277_47#_c_400_n N_VPWR_c_599_n 0.00484144f $X=4.225 $Y=1.54 $X2=0
+ $Y2=0
cc_305 N_A_277_47#_c_393_n N_VPWR_c_599_n 0.0044907f $X=4.395 $Y=1.16 $X2=0
+ $Y2=0
cc_306 N_A_277_47#_M1001_g N_VPWR_c_600_n 5.47116e-19 $X=4.47 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_A_277_47#_M1007_g N_VPWR_c_600_n 0.00894861f $X=4.89 $Y=1.985 $X2=0
+ $Y2=0
cc_308 N_A_277_47#_M1009_g N_VPWR_c_600_n 0.00894861f $X=5.31 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_277_47#_M1019_g N_VPWR_c_600_n 5.47116e-19 $X=5.73 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_A_277_47#_M1009_g N_VPWR_c_601_n 5.47116e-19 $X=5.31 $Y=1.985 $X2=0
+ $Y2=0
cc_311 N_A_277_47#_M1019_g N_VPWR_c_601_n 0.0107417f $X=5.73 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A_277_47#_M1001_g N_VPWR_c_608_n 0.0046653f $X=4.47 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A_277_47#_M1007_g N_VPWR_c_608_n 0.0046653f $X=4.89 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_277_47#_M1009_g N_VPWR_c_610_n 0.0046653f $X=5.31 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_277_47#_M1019_g N_VPWR_c_610_n 0.0046653f $X=5.73 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A_277_47#_M1000_d N_VPWR_c_595_n 0.00216833f $X=3.185 $Y=1.485 $X2=0
+ $Y2=0
cc_317 N_A_277_47#_M1001_g N_VPWR_c_595_n 0.00761484f $X=4.47 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A_277_47#_M1007_g N_VPWR_c_595_n 0.00420105f $X=4.89 $Y=1.985 $X2=0
+ $Y2=0
cc_319 N_A_277_47#_M1009_g N_VPWR_c_595_n 0.00420105f $X=5.31 $Y=1.985 $X2=0
+ $Y2=0
cc_320 N_A_277_47#_M1019_g N_VPWR_c_595_n 0.00420105f $X=5.73 $Y=1.985 $X2=0
+ $Y2=0
cc_321 N_A_277_47#_M1007_g N_X_c_711_n 0.0108499f $X=4.89 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_277_47#_M1009_g N_X_c_711_n 0.0108499f $X=5.31 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_277_47#_c_487_p N_X_c_711_n 0.0184321f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A_277_47#_c_394_n N_X_c_711_n 0.00162506f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_277_47#_M1001_g N_X_c_715_n 0.00820753f $X=4.47 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_277_47#_c_487_p N_X_c_715_n 0.00734001f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_277_47#_c_394_n N_X_c_715_n 0.00173288f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_277_47#_c_487_p N_X_c_718_n 0.00619755f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_277_47#_c_394_n N_X_c_718_n 0.00173288f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_277_47#_c_388_n X 0.00727387f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_277_47#_c_389_n X 0.00952437f $X=4.89 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_277_47#_c_390_n X 0.00952437f $X=5.31 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_277_47#_c_391_n X 0.0113488f $X=5.73 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_277_47#_c_487_p X 0.0897744f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_277_47#_c_394_n X 0.0107215f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_277_47#_M1019_g X 0.0126743f $X=5.73 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_277_47#_c_487_p X 0.00904517f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A_277_47#_c_394_n X 0.0035519f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A_277_47#_c_391_n X 0.00493062f $X=5.73 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_277_47#_M1019_g X 0.0133915f $X=5.73 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A_277_47#_c_487_p X 0.0240872f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_342 N_A_277_47#_c_394_n X 0.00911658f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_277_47#_c_404_n N_VGND_M1023_d 0.00785605f $X=3.155 $Y=0.785 $X2=0
+ $Y2=0
cc_344 N_A_277_47#_c_404_n N_VGND_c_760_n 0.0170458f $X=3.155 $Y=0.785 $X2=0
+ $Y2=0
cc_345 N_A_277_47#_c_388_n N_VGND_c_761_n 0.00127119f $X=4.47 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_277_47#_c_389_n N_VGND_c_761_n 0.00936721f $X=4.89 $Y=0.995 $X2=0
+ $Y2=0
cc_347 N_A_277_47#_c_390_n N_VGND_c_761_n 0.00845732f $X=5.31 $Y=0.995 $X2=0
+ $Y2=0
cc_348 N_A_277_47#_c_391_n N_VGND_c_761_n 0.00116151f $X=5.73 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_277_47#_c_390_n N_VGND_c_762_n 0.00116151f $X=5.31 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_277_47#_c_391_n N_VGND_c_762_n 0.00955881f $X=5.73 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_277_47#_c_416_n N_VGND_c_763_n 0.028758f $X=2.35 $Y=0.48 $X2=0 $Y2=0
cc_352 N_A_277_47#_c_404_n N_VGND_c_763_n 0.00233045f $X=3.155 $Y=0.785 $X2=0
+ $Y2=0
cc_353 N_A_277_47#_c_413_n N_VGND_c_763_n 0.00567506f $X=2.435 $Y=0.48 $X2=0
+ $Y2=0
cc_354 N_A_277_47#_c_388_n N_VGND_c_765_n 0.00543421f $X=4.47 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A_277_47#_c_389_n N_VGND_c_765_n 0.00341689f $X=4.89 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_277_47#_c_390_n N_VGND_c_767_n 0.00341689f $X=5.31 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_277_47#_c_391_n N_VGND_c_767_n 0.00341689f $X=5.73 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A_277_47#_c_404_n N_VGND_c_769_n 0.00209524f $X=3.155 $Y=0.785 $X2=0
+ $Y2=0
cc_359 N_A_277_47#_c_407_n N_VGND_c_769_n 0.0149873f $X=3.32 $Y=0.38 $X2=0 $Y2=0
cc_360 N_A_277_47#_M1011_s N_VGND_c_771_n 0.0023595f $X=1.385 $Y=0.235 $X2=0
+ $Y2=0
cc_361 N_A_277_47#_M1004_d N_VGND_c_771_n 0.00217524f $X=3.185 $Y=0.235 $X2=0
+ $Y2=0
cc_362 N_A_277_47#_c_388_n N_VGND_c_771_n 0.0108857f $X=4.47 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_277_47#_c_389_n N_VGND_c_771_n 0.0040262f $X=4.89 $Y=0.995 $X2=0
+ $Y2=0
cc_364 N_A_277_47#_c_390_n N_VGND_c_771_n 0.0040262f $X=5.31 $Y=0.995 $X2=0
+ $Y2=0
cc_365 N_A_277_47#_c_391_n N_VGND_c_771_n 0.0040262f $X=5.73 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A_277_47#_c_416_n N_VGND_c_771_n 0.0321646f $X=2.35 $Y=0.48 $X2=0 $Y2=0
cc_367 N_A_277_47#_c_404_n N_VGND_c_771_n 0.00921236f $X=3.155 $Y=0.785 $X2=0
+ $Y2=0
cc_368 N_A_277_47#_c_407_n N_VGND_c_771_n 0.0119254f $X=3.32 $Y=0.38 $X2=0 $Y2=0
cc_369 N_A_277_47#_c_413_n N_VGND_c_771_n 0.00590183f $X=2.435 $Y=0.48 $X2=0
+ $Y2=0
cc_370 N_A_277_47#_c_388_n N_VGND_c_772_n 0.012965f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A_277_47#_c_407_n N_VGND_c_772_n 0.0161879f $X=3.32 $Y=0.38 $X2=0 $Y2=0
cc_372 N_A_277_47#_c_393_n N_VGND_c_772_n 0.00177637f $X=4.395 $Y=1.16 $X2=0
+ $Y2=0
cc_373 N_A_277_47#_c_416_n A_361_47# 0.00355608f $X=2.35 $Y=0.48 $X2=-0.19
+ $Y2=-0.24
cc_374 N_A_277_47#_c_416_n A_445_47# 0.00313334f $X=2.35 $Y=0.48 $X2=-0.19
+ $Y2=-0.24
cc_375 N_A_277_47#_c_413_n A_445_47# 0.00911237f $X=2.435 $Y=0.48 $X2=-0.19
+ $Y2=-0.24
cc_376 N_A_27_297#_c_544_n N_VPWR_M1005_s 0.00325599f $X=1.015 $Y=1.87 $X2=0.47
+ $Y2=0.995
cc_377 N_A_27_297#_c_547_n N_VPWR_M1002_d 0.00317853f $X=1.855 $Y=1.87 $X2=0.47
+ $Y2=0.56
cc_378 N_A_27_297#_c_548_n N_VPWR_M1014_s 0.00452059f $X=2.815 $Y=1.87 $X2=0.47
+ $Y2=0.56
cc_379 N_A_27_297#_c_544_n N_VPWR_c_596_n 0.0165384f $X=1.015 $Y=1.87 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_c_547_n N_VPWR_c_597_n 0.0165384f $X=1.855 $Y=1.87 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_c_548_n N_VPWR_c_598_n 0.0191766f $X=2.815 $Y=1.87 $X2=0.385
+ $Y2=0.995
cc_382 N_A_27_297#_c_560_n N_VPWR_c_599_n 0.010563f $X=3.655 $Y=2.38 $X2=2.69
+ $Y2=1.325
cc_383 N_A_27_297#_c_567_n N_VPWR_c_599_n 0.00949729f $X=3.74 $Y=1.96 $X2=2.69
+ $Y2=1.325
cc_384 N_A_27_297#_c_554_n N_VPWR_c_602_n 0.0113958f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_385 N_A_27_297#_c_555_n N_VPWR_c_604_n 0.0113958f $X=1.94 $Y=1.95 $X2=0 $Y2=0
cc_386 N_A_27_297#_c_560_n N_VPWR_c_606_n 0.0475374f $X=3.655 $Y=2.38 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_c_580_p N_VPWR_c_606_n 0.0117106f $X=2.985 $Y=2.38 $X2=0
+ $Y2=0
cc_388 N_A_27_297#_c_552_n N_VPWR_c_612_n 0.0116048f $X=0.26 $Y=1.95 $X2=0 $Y2=0
cc_389 N_A_27_297#_M1005_d N_VPWR_c_595_n 0.00378138f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_M1003_d N_VPWR_c_595_n 0.00268171f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_391 N_A_27_297#_M1020_s N_VPWR_c_595_n 0.00268171f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_392 N_A_27_297#_M1012_d N_VPWR_c_595_n 0.00324087f $X=2.705 $Y=1.485 $X2=0
+ $Y2=0
cc_393 N_A_27_297#_M1006_s N_VPWR_c_595_n 0.00348186f $X=3.605 $Y=1.485 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_544_n N_VPWR_c_595_n 0.0117708f $X=1.015 $Y=1.87 $X2=0
+ $Y2=0
cc_395 N_A_27_297#_c_547_n N_VPWR_c_595_n 0.0117708f $X=1.855 $Y=1.87 $X2=0
+ $Y2=0
cc_396 N_A_27_297#_c_548_n N_VPWR_c_595_n 0.0159311f $X=2.815 $Y=1.87 $X2=0
+ $Y2=0
cc_397 N_A_27_297#_c_560_n N_VPWR_c_595_n 0.0299868f $X=3.655 $Y=2.38 $X2=0
+ $Y2=0
cc_398 N_A_27_297#_c_580_p N_VPWR_c_595_n 0.00654177f $X=2.985 $Y=2.38 $X2=0
+ $Y2=0
cc_399 N_A_27_297#_c_552_n N_VPWR_c_595_n 0.00646998f $X=0.26 $Y=1.95 $X2=0
+ $Y2=0
cc_400 N_A_27_297#_c_554_n N_VPWR_c_595_n 0.00646998f $X=1.1 $Y=1.95 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_555_n N_VPWR_c_595_n 0.00646998f $X=1.94 $Y=1.95 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_595_n N_X_M1001_d 0.00268098f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_c_595_n N_X_M1009_d 0.00268171f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_M1007_s N_X_c_711_n 0.004065f $X=4.965 $Y=1.485 $X2=0 $Y2=0
cc_405 N_VPWR_c_600_n N_X_c_711_n 0.0165384f $X=5.1 $Y=2.21 $X2=0 $Y2=0
cc_406 N_VPWR_c_595_n N_X_c_711_n 0.0117708f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_407 N_VPWR_c_608_n N_X_c_715_n 0.0113958f $X=4.935 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_595_n N_X_c_715_n 0.00853629f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_610_n N_X_c_718_n 0.0113958f $X=5.775 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_595_n N_X_c_718_n 0.00646998f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_M1019_s X 0.0243091f $X=5.805 $Y=1.485 $X2=0 $Y2=0
cc_412 N_VPWR_c_601_n X 0.0212316f $X=5.94 $Y=2.21 $X2=0 $Y2=0
cc_413 N_VPWR_c_595_n X 0.0142995f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_M1019_s X 0.0181031f $X=5.805 $Y=1.485 $X2=0 $Y2=0
cc_415 X N_VGND_M1015_d 0.00305768f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_416 X N_VGND_M1017_d 0.00703534f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_417 X N_VGND_c_761_n 0.0160613f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_418 X N_VGND_c_762_n 0.0207342f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_419 X N_VGND_c_765_n 0.00615083f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_420 X N_VGND_c_767_n 0.00739173f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_421 X N_VGND_c_770_n 3.32968e-19 $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_422 N_X_c_707_n N_VGND_c_770_n 0.00331351f $X=6.21 $Y=0.825 $X2=0 $Y2=0
cc_423 N_X_M1013_s N_VGND_c_771_n 0.00323135f $X=4.545 $Y=0.235 $X2=0 $Y2=0
cc_424 N_X_M1016_s N_VGND_c_771_n 0.00323135f $X=5.385 $Y=0.235 $X2=0 $Y2=0
cc_425 X N_VGND_c_771_n 0.0276551f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_426 N_X_c_707_n N_VGND_c_771_n 0.00504033f $X=6.21 $Y=0.825 $X2=0 $Y2=0
cc_427 N_VGND_c_771_n A_109_47# 0.0112452f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_428 N_VGND_c_771_n A_193_47# 0.00355046f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_429 N_VGND_c_771_n A_361_47# 0.0023595f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_430 N_VGND_c_771_n A_445_47# 0.00300108f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__dlymetal6s2s_1.pex.spice
* Created: Tue Sep  1 19:06:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A 3 7 9 10 15 17
c31 17 0 1.57226e-19 $X=0.645 $Y=1.16
r32 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.42 $Y=1.16
+ $X2=0.645 $Y2=1.16
r33 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=1.16 $X2=0.42 $Y2=1.16
r34 9 10 8.38488 $w=4.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.327 $Y=1.19
+ $X2=0.327 $Y2=1.53
r35 9 15 0.739842 $w=4.83e-07 $l=3e-08 $layer=LI1_cond $X=0.327 $Y=1.19
+ $X2=0.327 $Y2=1.16
r36 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=1.325
+ $X2=0.645 $Y2=1.16
r37 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.645 $Y=1.325
+ $X2=0.645 $Y2=2.275
r38 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=0.995
+ $X2=0.645 $Y2=1.16
r39 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.645 $Y=0.995
+ $X2=0.645 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_62_47# 1 2 9 12 14 16 21 23 27 33
+ 34 35 38
c59 33 0 1.1704e-19 $X=1.065 $Y=1.16
c60 16 0 1.57226e-19 $X=0.74 $Y=1.955
r61 34 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.16
+ $X2=1.065 $Y2=1.325
r62 34 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.16
+ $X2=1.065 $Y2=0.995
r63 33 36 5.05753 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.16
+ $X2=0.945 $Y2=1.325
r64 33 35 5.05753 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.16
+ $X2=0.945 $Y2=0.995
r65 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.065
+ $Y=1.16 $X2=1.065 $Y2=1.16
r66 27 30 8.47774 $w=4.33e-07 $l=3.2e-07 $layer=LI1_cond $X=0.302 $Y=1.955
+ $X2=0.302 $Y2=2.275
r67 23 25 7.81542 $w=4.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.302 $Y=0.445
+ $X2=0.302 $Y2=0.74
r68 21 36 18.7487 $w=3.33e-07 $l=5.45e-07 $layer=LI1_cond $X=0.907 $Y=1.87
+ $X2=0.907 $Y2=1.325
r69 18 35 5.84822 $w=3.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.907 $Y=0.825
+ $X2=0.907 $Y2=0.995
r70 17 27 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.52 $Y=1.955
+ $X2=0.302 $Y2=1.955
r71 16 21 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=0.74 $Y=1.955
+ $X2=0.907 $Y2=1.87
r72 16 17 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.74 $Y=1.955
+ $X2=0.52 $Y2=1.955
r73 15 25 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.52 $Y=0.74
+ $X2=0.302 $Y2=0.74
r74 14 18 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=0.74 $Y=0.74
+ $X2=0.907 $Y2=0.825
r75 14 15 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.74 $Y=0.74
+ $X2=0.52 $Y2=0.74
r76 12 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.12 $Y=1.985
+ $X2=1.12 $Y2=1.325
r77 9 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.12 $Y=0.56 $X2=1.12
+ $Y2=0.995
r78 2 30 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.31
+ $Y=2.065 $X2=0.435 $Y2=2.275
r79 1 23 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.235 $X2=0.435 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%X 1 2 9 13 15 16 17 18 19 20 21 22 35
+ 37
r49 32 35 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.015 $Y=1.16
+ $X2=2.24 $Y2=1.16
r50 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=1.16 $X2=2.015 $Y2=1.16
r51 20 41 6.77908 $w=4.23e-07 $l=2.5e-07 $layer=LI1_cond $X=1.457 $Y=2.21
+ $X2=1.457 $Y2=1.96
r52 19 41 2.44047 $w=4.23e-07 $l=9e-08 $layer=LI1_cond $X=1.457 $Y=1.87
+ $X2=1.457 $Y2=1.96
r53 19 37 5.28768 $w=4.23e-07 $l=1.95e-07 $layer=LI1_cond $X=1.457 $Y=1.87
+ $X2=1.457 $Y2=1.675
r54 18 37 4.06575 $w=6.19e-07 $l=2.76141e-07 $layer=LI1_cond $X=1.67 $Y=1.53
+ $X2=1.457 $Y2=1.675
r55 18 22 8.51824 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=1.67 $Y=1.53
+ $X2=2.045 $Y2=1.53
r56 17 18 6.70113 $w=6.19e-07 $l=3.4e-07 $layer=LI1_cond $X=1.67 $Y=1.19
+ $X2=1.67 $Y2=1.53
r57 17 21 8.51824 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=1.67 $Y=1.19
+ $X2=2.045 $Y2=1.19
r58 17 33 0.591276 $w=6.19e-07 $l=3e-08 $layer=LI1_cond $X=1.67 $Y=1.19 $X2=1.67
+ $Y2=1.16
r59 16 33 6.10985 $w=6.19e-07 $l=3.1e-07 $layer=LI1_cond $X=1.67 $Y=0.85
+ $X2=1.67 $Y2=1.16
r60 15 16 6.70113 $w=6.19e-07 $l=3.4e-07 $layer=LI1_cond $X=1.67 $Y=0.51
+ $X2=1.67 $Y2=0.85
r61 15 46 1.37964 $w=6.19e-07 $l=7e-08 $layer=LI1_cond $X=1.67 $Y=0.51 $X2=1.67
+ $Y2=0.44
r62 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=1.325
+ $X2=2.24 $Y2=1.16
r63 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.24 $Y=1.325
+ $X2=2.24 $Y2=2.275
r64 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=0.995
+ $X2=2.24 $Y2=1.16
r65 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.24 $Y=0.995 $X2=2.24
+ $Y2=0.445
r66 2 41 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.195
+ $Y=1.485 $X2=1.33 $Y2=1.96
r67 1 46 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.235 $X2=1.33 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_381_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c67 26 0 1.27733e-19 $X=2.495 $Y=1.325
r68 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.16
+ $X2=2.66 $Y2=1.325
r69 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.16
+ $X2=2.66 $Y2=0.995
r70 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.16 $X2=2.66 $Y2=1.16
r71 28 30 13.2746 $w=3.86e-07 $l=4.2e-07 $layer=LI1_cond $X=2.532 $Y=0.74
+ $X2=2.532 $Y2=1.16
r72 26 30 5.34605 $w=3.86e-07 $l=1.82565e-07 $layer=LI1_cond $X=2.495 $Y=1.325
+ $X2=2.532 $Y2=1.16
r73 26 27 17.122 $w=3.48e-07 $l=5.2e-07 $layer=LI1_cond $X=2.495 $Y=1.325
+ $X2=2.495 $Y2=1.845
r74 24 27 7.55928 $w=1.95e-07 $l=2.18174e-07 $layer=LI1_cond $X=2.32 $Y=1.942
+ $X2=2.495 $Y2=1.845
r75 24 25 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=2.32 $Y=1.942
+ $X2=2.115 $Y2=1.942
r76 22 28 5.5624 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.32 $Y=0.74
+ $X2=2.532 $Y2=0.74
r77 22 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.32 $Y=0.74
+ $X2=2.115 $Y2=0.74
r78 18 23 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.987 $Y=0.655
+ $X2=2.115 $Y2=0.74
r79 18 20 9.71668 $w=2.53e-07 $l=2.15e-07 $layer=LI1_cond $X=1.987 $Y=0.655
+ $X2=1.987 $Y2=0.44
r80 14 25 7.07654 $w=1.95e-07 $l=1.80466e-07 $layer=LI1_cond $X=1.977 $Y=2.04
+ $X2=2.115 $Y2=1.942
r81 14 16 9.84815 $w=2.73e-07 $l=2.35e-07 $layer=LI1_cond $X=1.977 $Y=2.04
+ $X2=1.977 $Y2=2.275
r82 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.715 $Y=1.985
+ $X2=2.715 $Y2=1.325
r83 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.715 $Y=0.56
+ $X2=2.715 $Y2=0.995
r84 2 16 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.065 $X2=2.03 $Y2=2.275
r85 1 20 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.03 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_558_47# 1 2 9 13 17 19 21 24 25 31
r55 28 31 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.43 $Y=1.16
+ $X2=3.655 $Y2=1.16
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.16 $X2=3.43 $Y2=1.16
r57 24 27 10.8173 $w=6.69e-07 $l=2.72276e-07 $layer=LI1_cond $X=3 $Y=0.995
+ $X2=3.202 $Y2=1.16
r58 24 25 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3 $Y=0.995 $X2=3
+ $Y2=0.825
r59 19 27 14.5453 $w=6.69e-07 $l=6.23558e-07 $layer=LI1_cond $X=2.962 $Y=1.675
+ $X2=3.202 $Y2=1.16
r60 19 21 13.406 $w=2.43e-07 $l=2.85e-07 $layer=LI1_cond $X=2.962 $Y=1.675
+ $X2=2.962 $Y2=1.96
r61 15 25 6.82988 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=2.962 $Y=0.703
+ $X2=2.962 $Y2=0.825
r62 15 17 12.3711 $w=2.43e-07 $l=2.63e-07 $layer=LI1_cond $X=2.962 $Y=0.703
+ $X2=2.962 $Y2=0.44
r63 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.325
+ $X2=3.655 $Y2=1.16
r64 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.655 $Y=1.325
+ $X2=3.655 $Y2=2.275
r65 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=0.995
+ $X2=3.655 $Y2=1.16
r66 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.655 $Y=0.995
+ $X2=3.655 $Y2=0.445
r67 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=1.485 $X2=2.925 $Y2=1.96
r68 1 17 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.235 $X2=2.925 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_664_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c66 26 0 1.27733e-19 $X=3.91 $Y=1.325
r67 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.16
+ $X2=4.075 $Y2=1.325
r68 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.16
+ $X2=4.075 $Y2=0.995
r69 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.075
+ $Y=1.16 $X2=4.075 $Y2=1.16
r70 28 30 13.2746 $w=3.86e-07 $l=4.2e-07 $layer=LI1_cond $X=3.947 $Y=0.74
+ $X2=3.947 $Y2=1.16
r71 26 30 5.34605 $w=3.86e-07 $l=1.82565e-07 $layer=LI1_cond $X=3.91 $Y=1.325
+ $X2=3.947 $Y2=1.16
r72 26 27 17.122 $w=3.48e-07 $l=5.2e-07 $layer=LI1_cond $X=3.91 $Y=1.325
+ $X2=3.91 $Y2=1.845
r73 24 27 7.55928 $w=1.95e-07 $l=2.18174e-07 $layer=LI1_cond $X=3.735 $Y=1.942
+ $X2=3.91 $Y2=1.845
r74 24 25 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.735 $Y=1.942
+ $X2=3.53 $Y2=1.942
r75 22 28 5.5624 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.735 $Y=0.74
+ $X2=3.947 $Y2=0.74
r76 22 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.735 $Y=0.74
+ $X2=3.53 $Y2=0.74
r77 18 25 6.9753 $w=1.95e-07 $l=1.70082e-07 $layer=LI1_cond $X=3.402 $Y=2.04
+ $X2=3.53 $Y2=1.942
r78 18 20 10.6206 $w=2.53e-07 $l=2.35e-07 $layer=LI1_cond $X=3.402 $Y=2.04
+ $X2=3.402 $Y2=2.275
r79 14 23 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=3.402 $Y=0.655
+ $X2=3.53 $Y2=0.74
r80 14 16 9.71668 $w=2.53e-07 $l=2.15e-07 $layer=LI1_cond $X=3.402 $Y=0.655
+ $X2=3.402 $Y2=0.44
r81 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.13 $Y=1.985
+ $X2=4.13 $Y2=1.325
r82 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.56 $X2=4.13
+ $Y2=0.995
r83 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=2.065 $X2=3.445 $Y2=2.275
r84 1 16 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.235 $X2=3.445 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%VPWR 1 2 3 14 18 22 24 26 34 41 42 45
+ 48 51 56
r62 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 46 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r68 39 51 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=3.892 $Y2=2.72
r69 39 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=4.37 $Y2=2.72
r70 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 38 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r73 35 48 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.67 $Y=2.72
+ $X2=2.477 $Y2=2.72
r74 35 37 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.67 $Y=2.72
+ $X2=3.45 $Y2=2.72
r75 34 51 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.7 $Y=2.72
+ $X2=3.892 $Y2=2.72
r76 34 37 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.45
+ $Y2=2.72
r77 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r78 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r79 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 30 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r82 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 27 45 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=0.882 $Y2=2.72
r84 27 29 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 26 48 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.477 $Y2=2.72
r86 26 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 24 56 0.00711354 $w=4.8e-07 $l=2.5e-08 $layer=MET1_cond $X=0.205 $Y=2.72
+ $X2=0.23 $Y2=2.72
r88 20 51 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.892 $Y2=2.72
r89 20 22 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.892 $Y2=2.36
r90 16 48 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.477 $Y=2.635
+ $X2=2.477 $Y2=2.72
r91 16 18 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=2.477 $Y=2.635
+ $X2=2.477 $Y2=2.36
r92 12 45 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.882 $Y=2.635
+ $X2=0.882 $Y2=2.72
r93 12 14 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=0.882 $Y=2.635
+ $X2=0.882 $Y2=2.36
r94 3 22 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=2.065 $X2=3.895 $Y2=2.36
r95 2 18 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.065 $X2=2.48 $Y2=2.36
r96 1 14 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=2.065 $X2=0.885 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%A_841_47# 1 2 9 11 13 17 18
r17 17 18 40.1671 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=4.422 $Y=0.825
+ $X2=4.422 $Y2=1.495
r18 11 18 6.73749 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=4.385 $Y=1.625
+ $X2=4.385 $Y2=1.495
r19 11 13 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=4.385 $Y=1.625
+ $X2=4.385 $Y2=1.96
r20 7 17 6.73749 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=4.385 $Y=0.695
+ $X2=4.385 $Y2=0.825
r21 7 9 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=4.385 $Y=0.695
+ $X2=4.385 $Y2=0.44
r22 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.205
+ $Y=1.485 $X2=4.34 $Y2=1.96
r23 1 9 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.235 $X2=4.34 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S2S_1%VGND 1 2 3 14 18 22 24 26 34 41 42 45
+ 48 51 56
r65 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r66 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r67 46 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r68 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r69 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r70 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r71 39 51 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=3.892
+ $Y2=0
r72 39 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.37
+ $Y2=0
r73 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r74 38 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r75 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r76 35 48 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.477
+ $Y2=0
r77 35 37 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=3.45
+ $Y2=0
r78 34 51 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.892
+ $Y2=0
r79 34 37 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.45
+ $Y2=0
r80 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r81 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r82 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r83 30 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r84 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r85 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r86 27 45 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.882
+ $Y2=0
r87 27 29 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.15
+ $Y2=0
r88 26 48 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.477
+ $Y2=0
r89 26 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.07
+ $Y2=0
r90 24 56 0.00711354 $w=4.8e-07 $l=2.5e-08 $layer=MET1_cond $X=0.205 $Y=0
+ $X2=0.23 $Y2=0
r91 20 51 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.892 $Y2=0
r92 20 22 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.892 $Y2=0.38
r93 16 48 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.477 $Y=0.085
+ $X2=2.477 $Y2=0
r94 16 18 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=2.477 $Y=0.085
+ $X2=2.477 $Y2=0.38
r95 12 45 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.882 $Y=0.085
+ $X2=0.882 $Y2=0
r96 12 14 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.882 $Y=0.085
+ $X2=0.882 $Y2=0.38
r97 3 22 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.89 $Y2=0.38
r98 2 18 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.235 $X2=2.475 $Y2=0.38
r99 1 14 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.72
+ $Y=0.235 $X2=0.88 $Y2=0.38
.ends


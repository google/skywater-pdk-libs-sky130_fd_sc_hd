* File: sky130_fd_sc_hd__inv_6.spice.pex
* Created: Thu Aug 27 14:22:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__INV_6%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 44 45 46 51 64
c109 27 0 5.55636e-20 $X=1.9 $Y=1.985
r110 62 64 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=2.45 $Y=1.16
+ $X2=2.74 $Y2=1.16
r111 60 62 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.32 $Y=1.16
+ $X2=2.45 $Y2=1.16
r112 59 60 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.9 $Y=1.16
+ $X2=2.32 $Y2=1.16
r113 58 59 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.48 $Y=1.16
+ $X2=1.9 $Y2=1.16
r114 57 58 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.06 $Y=1.16
+ $X2=1.48 $Y2=1.16
r115 56 57 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.64 $Y=1.16
+ $X2=1.06 $Y2=1.16
r116 51 56 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.64 $Y2=1.16
r117 51 53 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.27 $Y2=1.16
r118 46 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.45
+ $Y=1.16 $X2=2.45 $Y2=1.16
r119 45 46 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=2.03 $Y=1.2 $X2=2.45
+ $Y2=1.2
r120 44 45 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.57 $Y=1.2 $X2=2.03
+ $Y2=1.2
r121 43 44 61.7709 $w=2.48e-07 $l=1.34e-06 $layer=LI1_cond $X=0.23 $Y=1.2
+ $X2=1.57 $Y2=1.2
r122 43 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r123 39 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.325
+ $X2=2.74 $Y2=1.16
r124 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.74 $Y=1.325
+ $X2=2.74 $Y2=1.985
r125 36 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=0.995
+ $X2=2.74 $Y2=1.16
r126 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.74 $Y=0.995
+ $X2=2.74 $Y2=0.56
r127 32 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.325
+ $X2=2.32 $Y2=1.16
r128 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.32 $Y=1.325
+ $X2=2.32 $Y2=1.985
r129 29 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=0.995
+ $X2=2.32 $Y2=1.16
r130 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.32 $Y=0.995
+ $X2=2.32 $Y2=0.56
r131 25 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=1.325
+ $X2=1.9 $Y2=1.16
r132 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.9 $Y=1.325
+ $X2=1.9 $Y2=1.985
r133 22 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=1.16
r134 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=0.56
r135 18 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=1.325
+ $X2=1.48 $Y2=1.16
r136 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.48 $Y=1.325
+ $X2=1.48 $Y2=1.985
r137 15 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.16
r138 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=0.56
r139 11 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.325
+ $X2=1.06 $Y2=1.16
r140 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.06 $Y=1.325
+ $X2=1.06 $Y2=1.985
r141 8 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=0.995
+ $X2=1.06 $Y2=1.16
r142 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.06 $Y=0.995
+ $X2=1.06 $Y2=0.56
r143 4 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.325
+ $X2=0.64 $Y2=1.16
r144 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.64 $Y=1.325
+ $X2=0.64 $Y2=1.985
r145 1 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=0.995
+ $X2=0.64 $Y2=1.16
r146 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.64 $Y=0.995
+ $X2=0.64 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__INV_6%VPWR 1 2 3 4 13 15 21 23 27 29 31 33 34 35 41
+ 50 54
r51 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 45 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 45 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 42 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.11 $Y2=2.72
r57 42 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 41 53 3.40825 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.042 $Y2=2.72
r59 41 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 40 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 37 47 4.38764 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r63 37 39 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 35 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 35 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r66 33 39 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.27 $Y2=2.72
r68 29 53 3.40825 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=2.95 $Y=2.635
+ $X2=3.042 $Y2=2.72
r69 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.95 $Y=2.635
+ $X2=2.95 $Y2=2.34
r70 25 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=2.635
+ $X2=2.11 $Y2=2.72
r71 25 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.11 $Y=2.635
+ $X2=2.11 $Y2=2
r72 24 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=2.72
+ $X2=1.27 $Y2=2.72
r73 23 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.11 $Y2=2.72
r74 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.355 $Y2=2.72
r75 19 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.635
+ $X2=1.27 $Y2=2.72
r76 19 21 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.27 $Y=2.635
+ $X2=1.27 $Y2=2
r77 15 18 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.277 $Y=1.66
+ $X2=0.277 $Y2=2.34
r78 13 47 3.08989 $w=2.95e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.277 $Y=2.635
+ $X2=0.212 $Y2=2.72
r79 13 18 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.277 $Y=2.635
+ $X2=0.277 $Y2=2.34
r80 4 31 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.485 $X2=2.95 $Y2=2.34
r81 3 27 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.975
+ $Y=1.485 $X2=2.11 $Y2=2
r82 2 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.485 $X2=1.27 $Y2=2
r83 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r84 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__INV_6%Y 1 2 3 4 5 6 19 21 25 27 28 29 33 37 39 45 49
+ 54 55 56 57 58 64 65 77
c99 65 0 5.55636e-20 $X=2.96 $Y=1.495
r100 76 77 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=1.59
+ $X2=2.365 $Y2=1.59
r101 58 65 0.583732 $w=1.88e-07 $l=1e-08 $layer=LI1_cond $X=2.95 $Y=1.59
+ $X2=2.96 $Y2=1.59
r102 58 76 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=2.95 $Y=1.59
+ $X2=2.53 $Y2=1.59
r103 58 65 0.823174 $w=3.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.96 $Y=1.47
+ $X2=2.96 $Y2=1.495
r104 57 58 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.96 $Y=1.19
+ $X2=2.96 $Y2=1.47
r105 56 64 0.616162 $w=1.78e-07 $l=1e-08 $layer=LI1_cond $X=2.95 $Y=0.815
+ $X2=2.96 $Y2=0.815
r106 56 70 25.8788 $w=1.78e-07 $l=4.2e-07 $layer=LI1_cond $X=2.95 $Y=0.815
+ $X2=2.53 $Y2=0.815
r107 56 57 8.89028 $w=3.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.96 $Y=0.92
+ $X2=2.96 $Y2=1.19
r108 56 64 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=2.96 $Y=0.92
+ $X2=2.96 $Y2=0.905
r109 47 70 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.53 $Y=0.725 $X2=2.53
+ $Y2=0.815
r110 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.53 $Y=0.725
+ $X2=2.53 $Y2=0.42
r111 45 76 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=2.53 $Y=2.34
+ $X2=2.53 $Y2=1.685
r112 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=1.58
+ $X2=1.69 $Y2=1.58
r113 42 77 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.855 $Y=1.58
+ $X2=2.365 $Y2=1.58
r114 40 55 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=0.815
+ $X2=1.69 $Y2=0.815
r115 39 70 5.23737 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=0.815
+ $X2=2.53 $Y2=0.815
r116 39 40 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.445 $Y=0.815
+ $X2=1.775 $Y2=0.815
r117 35 55 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=0.725 $X2=1.69
+ $Y2=0.815
r118 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.69 $Y=0.725
+ $X2=1.69 $Y2=0.42
r119 31 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=1.665
+ $X2=1.69 $Y2=1.58
r120 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.69 $Y=1.665
+ $X2=1.69 $Y2=2.34
r121 30 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=1.58
+ $X2=0.85 $Y2=1.58
r122 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=1.58
+ $X2=1.69 $Y2=1.58
r123 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.525 $Y=1.58
+ $X2=1.015 $Y2=1.58
r124 27 55 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.815
+ $X2=1.69 $Y2=0.815
r125 27 28 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=1.605 $Y=0.815
+ $X2=0.935 $Y2=0.815
r126 23 28 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.85 $Y=0.725
+ $X2=0.935 $Y2=0.815
r127 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.85 $Y=0.725
+ $X2=0.85 $Y2=0.42
r128 19 52 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=1.665
+ $X2=0.85 $Y2=1.58
r129 19 21 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.85 $Y=1.665
+ $X2=0.85 $Y2=2.34
r130 6 76 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.485 $X2=2.53 $Y2=1.66
r131 6 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.485 $X2=2.53 $Y2=2.34
r132 5 54 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.485 $X2=1.69 $Y2=1.66
r133 5 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.485 $X2=1.69 $Y2=2.34
r134 4 52 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.485 $X2=0.85 $Y2=1.66
r135 4 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.485 $X2=0.85 $Y2=2.34
r136 3 49 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.53 $Y2=0.42
r137 2 37 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.42
r138 1 25 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.715
+ $Y=0.235 $X2=0.85 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__INV_6%VGND 1 2 3 4 13 15 19 21 25 27 29 31 32 33 39
+ 48 52
r56 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r57 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r58 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r59 43 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r60 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r61 40 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.11
+ $Y2=0
r62 40 42 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.53
+ $Y2=0
r63 39 51 3.93418 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=3.002
+ $Y2=0
r64 39 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=2.53
+ $Y2=0
r65 38 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r66 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r67 35 45 4.1239 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r68 35 37 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=1.15
+ $Y2=0
r69 33 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r70 33 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 31 37 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.15
+ $Y2=0
r72 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.27
+ $Y2=0
r73 27 51 3.20898 $w=2.5e-07 $l=1.27609e-07 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=3.002 $Y2=0
r74 27 29 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=2.91 $Y=0.085 $X2=2.91
+ $Y2=0.385
r75 23 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0
r76 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.38
r77 22 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.27
+ $Y2=0
r78 21 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.11
+ $Y2=0
r79 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.355
+ $Y2=0
r80 17 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=0.085
+ $X2=1.27 $Y2=0
r81 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.27 $Y=0.085
+ $X2=1.27 $Y2=0.38
r82 13 45 3.12417 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.197 $Y2=0
r83 13 15 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.262 $Y2=0.38
r84 4 29 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.235 $X2=2.95 $Y2=0.385
r85 3 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.38
r86 2 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.135
+ $Y=0.235 $X2=1.27 $Y2=0.38
r87 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends


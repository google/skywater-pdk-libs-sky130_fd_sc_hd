* File: sky130_fd_sc_hd__o22ai_1.spice.pex
* Created: Thu Aug 27 14:37:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O22AI_1%B1 1 3 6 8 14
r32 11 14 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r34 8 12 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.205 $Y=0.85
+ $X2=0.205 $Y2=1.16
r35 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r36 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r37 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_1%B2 3 7 10 11 13 16
c46 13 0 3.05135e-20 $X=1.15 $Y=1.53
c47 11 0 2.81177e-21 $X=0.92 $Y=1.16
c48 3 0 2.57224e-19 $X=0.845 $Y=1.985
r49 13 18 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.15 $Y=1.54
+ $X2=0.92 $Y2=1.54
r50 11 17 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.912 $Y=1.16
+ $X2=0.912 $Y2=1.325
r51 11 16 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.912 $Y=1.16
+ $X2=0.912 $Y2=0.995
r52 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.92
+ $Y=1.16 $X2=0.92 $Y2=1.16
r53 8 18 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.92 $Y=1.415
+ $X2=0.92 $Y2=1.54
r54 8 10 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.92 $Y=1.415
+ $X2=0.92 $Y2=1.16
r55 7 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.56
+ $X2=0.905 $Y2=0.995
r56 3 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.845 $Y=1.985
+ $X2=0.845 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_1%A2 3 6 9 12 14 19 21 24
c52 19 0 1.36372e-19 $X=1.625 $Y=1.615
c53 9 0 1.20852e-19 $X=1.495 $Y=1.445
r54 19 21 15.555 $w=2e-07 $l=2.55e-07 $layer=LI1_cond $X=1.625 $Y=1.615
+ $X2=1.625 $Y2=1.87
r55 16 19 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.495 $Y=1.53
+ $X2=1.625 $Y2=1.53
r56 12 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.16 $X2=1.4
+ $Y2=1.325
r57 12 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.16 $X2=1.4
+ $Y2=0.995
r58 11 14 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.4 $Y=1.16
+ $X2=1.495 $Y2=1.16
r59 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=1.16 $X2=1.4 $Y2=1.16
r60 9 16 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.495 $Y=1.445
+ $X2=1.495 $Y2=1.53
r61 8 14 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.495 $Y=1.245
+ $X2=1.495 $Y2=1.16
r62 8 9 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=1.495 $Y=1.245 $X2=1.495
+ $Y2=1.445
r63 6 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.46 $Y=1.985
+ $X2=1.46 $Y2=1.325
r64 3 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.56 $X2=1.41
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_1%A1 3 7 8 11 13
c27 8 0 2.81177e-21 $X=2.07 $Y=1.19
r28 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.16
+ $X2=1.91 $Y2=1.325
r29 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.16
+ $X2=1.91 $Y2=0.995
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r31 8 12 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.07 $Y=1.175
+ $X2=1.92 $Y2=1.175
r32 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.56 $X2=1.83
+ $Y2=0.995
r33 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.82 $Y=1.985
+ $X2=1.82 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_1%VPWR 1 2 7 9 11 13 17 19 32
c31 13 0 3.05135e-20 $X=2.03 $Y=1.64
r32 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r33 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r35 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r36 22 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r37 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 20 28 3.66972 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r39 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 19 31 4.71668 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=2.097 $Y2=2.72
r41 19 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 17 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r44 13 16 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.055 $Y=1.64
+ $X2=2.055 $Y2=2.32
r45 11 31 2.96544 $w=3.2e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.097 $Y2=2.72
r46 11 16 11.3444 $w=3.18e-07 $l=3.15e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2.32
r47 7 28 3.24547 $w=2.1e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.172 $Y2=2.72
r48 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.34
r49 2 16 400 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.485 $X2=2.03 $Y2=2.32
r50 2 13 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.485 $X2=2.03 $Y2=1.64
r51 1 9 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_1%Y 1 2 8 12 14
r31 14 18 2.51957 $w=4.6e-07 $l=9.5e-08 $layer=LI1_cond $X=1.15 $Y=2.15
+ $X2=1.055 $Y2=2.15
r32 9 12 6.16162 $w=1.78e-07 $l=1e-07 $layer=LI1_cond $X=0.58 $Y=0.735 $X2=0.68
+ $Y2=0.735
r33 8 18 12.5978 $w=4.6e-07 $l=6.12577e-07 $layer=LI1_cond $X=0.58 $Y=1.835
+ $X2=1.055 $Y2=2.15
r34 7 9 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.58 $Y=0.825 $X2=0.58
+ $Y2=0.735
r35 7 8 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.58 $Y=0.825
+ $X2=0.58 $Y2=1.835
r36 2 18 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.92
+ $Y=1.485 $X2=1.055 $Y2=1.96
r37 1 12 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_1%A_27_47# 1 2 3 10 14 15 16 20
r42 18 20 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=2.045 $Y=0.695
+ $X2=2.045 $Y2=0.39
r43 17 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0.78
+ $X2=1.18 $Y2=0.78
r44 16 18 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.875 $Y=0.78
+ $X2=2.045 $Y2=0.695
r45 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.875 $Y=0.78
+ $X2=1.345 $Y2=0.78
r46 15 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.695 $X2=1.18
+ $Y2=0.78
r47 14 23 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.18 $Y=0.475 $X2=1.18
+ $Y2=0.385
r48 14 15 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.18 $Y=0.475
+ $X2=1.18 $Y2=0.695
r49 10 23 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0.385
+ $X2=1.18 $Y2=0.385
r50 10 12 46.5202 $w=1.78e-07 $l=7.55e-07 $layer=LI1_cond $X=1.015 $Y=0.385
+ $X2=0.26 $Y2=0.385
r51 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.39
r52 2 25 182 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.18 $Y2=0.73
r53 2 23 182 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.18 $Y2=0.39
r54 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O22AI_1%VGND 1 6 8 10 17 18 21
r30 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r31 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r32 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r33 15 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.62
+ $Y2=0
r34 15 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=2.07
+ $Y2=0
r35 10 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.62
+ $Y2=0
r36 10 12 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=1.535 $Y=0 $X2=0.23
+ $Y2=0
r37 8 22 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r38 8 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r39 4 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085 $X2=1.62
+ $Y2=0
r40 4 6 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.36
r41 1 6 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__dlclkp_2.spice
* Created: Thu Aug 27 14:16:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlclkp_2.pex.spice"
.subckt sky130_fd_sc_hd__dlclkp_2  VNB VPB CLK GATE VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* GATE	GATE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_CLK_M1018_g N_A_27_47#_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_193_47#_M1012_d N_A_27_47#_M1012_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_397_119# N_GATE_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.117125 AS=0.1302 PD=1.085 PS=1.46 NRD=63.96 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1003 N_A_477_413#_M1003_d N_A_27_47#_M1003_g A_397_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.123615 AS=0.117125 PD=1.13037 PS=1.085 NRD=81.42 NRS=63.96 M=1
+ R=2.8 SA=75000.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 A_652_47# N_A_193_47#_M1005_g N_A_477_413#_M1003_d VNB NSHORT L=0.15
+ W=0.39 AD=0.0646389 AS=0.114785 PD=0.717407 PS=1.04963 NRD=34.068 NRS=3.072
+ M=1 R=2.6 SA=75000.9 SB=75001.2 A=0.0585 P=1.08 MULT=1
MM1021 N_VGND_M1021_d N_A_643_307#_M1021_g A_652_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0901822 AS=0.0696111 PD=0.808598 PS=0.772593 NRD=30 NRS=31.632 M=1 R=2.8
+ SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_643_307#_M1017_d N_A_477_413#_M1017_g N_VGND_M1021_d VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.139568 PD=1.82 PS=1.2514 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 A_1041_47# N_A_643_307#_M1006_g N_A_957_369#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_CLK_M1001_g A_1041_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0769738 AS=0.0441 PD=0.769346 PS=0.63 NRD=15.708 NRS=14.28 M=1 R=2.8
+ SA=75000.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1001_d N_A_957_369#_M1007_g N_GCLK_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.119126 AS=0.08775 PD=1.19065 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_957_369#_M1009_g N_GCLK_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.195 AS=0.08775 PD=1.9 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_CLK_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 A_381_369# N_GATE_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.116891 AS=0.1664 PD=1.17132 PS=1.8 NRD=39.2818 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 N_A_477_413#_M1004_d N_A_193_47#_M1004_g A_381_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0987 AS=0.0767094 PD=0.89 PS=0.768679 NRD=56.2829 NRS=59.8683 M=1
+ R=2.8 SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1020 A_601_413# N_A_27_47#_M1020_g N_A_477_413#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0987 PD=0.63 PS=0.89 NRD=23.443 NRS=32.8202 M=1 R=2.8
+ SA=75001.3 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_643_307#_M1002_g A_601_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A_477_413#_M1019_g N_A_643_307#_M1019_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.183659 AS=0.26 PD=1.62195 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_957_369#_M1010_d N_A_643_307#_M1010_g N_VPWR_M1019_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2016 AS=0.117541 PD=1.27 PS=1.03805 NRD=76.9482 NRS=16.9223
+ M=1 R=4.26667 SA=75000.7 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_CLK_M1016_g N_A_957_369#_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.117541 AS=0.2016 PD=1.03805 PS=1.27 NRD=16.9223 NRS=30.7714 M=1
+ R=4.26667 SA=75001.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1016_d N_A_957_369#_M1008_g N_GCLK_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.183659 AS=0.135 PD=1.62195 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.3
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A_957_369#_M1014_g N_GCLK_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.3 AS=0.135 PD=2.6 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75001.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=11.6029 P=17.87
c_146 VPB 0 1.42073e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__dlclkp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a2111o_1.pxi.spice
* Created: Thu Aug 27 13:58:30 2020
* 
x_PM_SKY130_FD_SC_HD__A2111O_1%A_85_193# N_A_85_193#_M1011_d N_A_85_193#_M1009_d
+ N_A_85_193#_M1006_s N_A_85_193#_M1000_g N_A_85_193#_c_61_n N_A_85_193#_M1001_g
+ N_A_85_193#_c_62_n N_A_85_193#_c_77_p N_A_85_193#_c_105_p N_A_85_193#_c_66_n
+ N_A_85_193#_c_67_n N_A_85_193#_c_83_p N_A_85_193#_c_91_p N_A_85_193#_c_98_p
+ N_A_85_193#_c_68_n N_A_85_193#_c_79_p N_A_85_193#_c_63_n
+ PM_SKY130_FD_SC_HD__A2111O_1%A_85_193#
x_PM_SKY130_FD_SC_HD__A2111O_1%D1 N_D1_M1011_g N_D1_M1006_g D1 D1 D1 D1
+ N_D1_c_144_n N_D1_c_145_n N_D1_c_146_n PM_SKY130_FD_SC_HD__A2111O_1%D1
x_PM_SKY130_FD_SC_HD__A2111O_1%C1 N_C1_M1004_g N_C1_M1002_g C1 C1 C1 C1
+ N_C1_c_188_n N_C1_c_189_n N_C1_c_192_n PM_SKY130_FD_SC_HD__A2111O_1%C1
x_PM_SKY130_FD_SC_HD__A2111O_1%B1 N_B1_M1009_g N_B1_M1003_g B1 B1 B1 B1
+ N_B1_c_221_n N_B1_c_222_n PM_SKY130_FD_SC_HD__A2111O_1%B1
x_PM_SKY130_FD_SC_HD__A2111O_1%A1 N_A1_c_257_n N_A1_M1010_g N_A1_c_258_n
+ N_A1_M1007_g A1 A1 PM_SKY130_FD_SC_HD__A2111O_1%A1
x_PM_SKY130_FD_SC_HD__A2111O_1%A2 N_A2_M1008_g N_A2_M1005_g A2 N_A2_c_298_n
+ N_A2_c_299_n PM_SKY130_FD_SC_HD__A2111O_1%A2
x_PM_SKY130_FD_SC_HD__A2111O_1%X N_X_M1001_s N_X_M1000_s X X X X X X N_X_c_321_n
+ X PM_SKY130_FD_SC_HD__A2111O_1%X
x_PM_SKY130_FD_SC_HD__A2111O_1%VPWR N_VPWR_M1000_d N_VPWR_M1010_d N_VPWR_c_338_n
+ N_VPWR_c_339_n VPWR N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n
+ N_VPWR_c_337_n N_VPWR_c_344_n N_VPWR_c_345_n PM_SKY130_FD_SC_HD__A2111O_1%VPWR
x_PM_SKY130_FD_SC_HD__A2111O_1%A_516_297# N_A_516_297#_M1003_d
+ N_A_516_297#_M1005_d N_A_516_297#_c_392_n N_A_516_297#_c_397_n
+ N_A_516_297#_c_394_n N_A_516_297#_c_412_n
+ PM_SKY130_FD_SC_HD__A2111O_1%A_516_297#
x_PM_SKY130_FD_SC_HD__A2111O_1%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_M1008_d
+ N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n
+ VGND N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n N_VGND_c_422_n
+ PM_SKY130_FD_SC_HD__A2111O_1%VGND
cc_1 VNB N_A_85_193#_c_61_n 0.0202635f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.96
cc_2 VNB N_A_85_193#_c_62_n 0.00151605f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.16
cc_3 VNB N_A_85_193#_c_63_n 0.0487262f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.15
cc_4 VNB D1 2.31601e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_D1_c_144_n 0.0260437f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=0.825
cc_6 VNB N_D1_c_145_n 0.0205404f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.16
cc_7 VNB N_D1_c_146_n 0.0047979f $X=-0.19 $Y=-0.24 $X2=2.6 $Y2=0.74
cc_8 VNB C1 0.00187364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C1_c_188_n 0.0227383f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_10 VNB N_C1_c_189_n 0.0176571f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.465
cc_11 VNB B1 0.00240734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_221_n 0.0261653f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=0.825
cc_13 VNB N_B1_c_222_n 0.0171614f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.16
cc_14 VNB N_A1_c_257_n 0.0276709f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=0.235
cc_15 VNB N_A1_c_258_n 0.0160695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB A1 0.0056504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB A2 0.0176892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_298_n 0.0331962f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.985
cc_19 VNB N_A2_c_299_n 0.0196332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_321_n 0.0178526f $X=-0.19 $Y=-0.24 $X2=1.585 $Y2=0.737
cc_21 VNB N_VPWR_c_337_n 0.17485f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.74
cc_22 VNB N_VGND_c_414_n 0.00569825f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.96
cc_23 VNB N_VGND_c_415_n 0.0127185f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_24 VNB N_VGND_c_416_n 0.00512327f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.465
cc_25 VNB N_VGND_c_417_n 0.0195573f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.16
cc_26 VNB N_VGND_c_418_n 0.00660388f $X=-0.19 $Y=-0.24 $X2=1.585 $Y2=0.737
cc_27 VNB N_VGND_c_419_n 0.0332781f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.39
cc_28 VNB N_VGND_c_420_n 0.0192517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_421_n 0.0205586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_422_n 0.222331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_A_85_193#_M1000_g 0.0246597f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_32 VPB N_A_85_193#_c_62_n 0.00232925f $X=-0.19 $Y=1.305 $X2=0.805 $Y2=1.16
cc_33 VPB N_A_85_193#_c_66_n 0.0115687f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.555
cc_34 VPB N_A_85_193#_c_67_n 0.00184063f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.555
cc_35 VPB N_A_85_193#_c_68_n 0.00296658f $X=-0.19 $Y=1.305 $X2=1.26 $Y2=1.63
cc_36 VPB N_A_85_193#_c_63_n 0.0149584f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.15
cc_37 VPB N_D1_M1006_g 0.0220508f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB D1 0.00344192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_D1_c_144_n 0.0109921f $X=-0.19 $Y=1.305 $X2=0.805 $Y2=0.825
cc_40 VPB C1 0.00177625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_C1_c_188_n 0.00879047f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_42 VPB N_C1_c_192_n 0.0155573f $X=-0.19 $Y=1.305 $X2=0.805 $Y2=1.16
cc_43 VPB N_B1_M1003_g 0.0201943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB B1 0.00320115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_B1_c_221_n 0.0085622f $X=-0.19 $Y=1.305 $X2=0.805 $Y2=0.825
cc_46 VPB N_A1_c_257_n 0.00628024f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=0.235
cc_47 VPB N_A1_M1010_g 0.0214578f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.485
cc_48 VPB A1 7.79524e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A2_M1005_g 0.0263149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A2_c_298_n 0.00674233f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_51 VPB N_X_c_321_n 0.00615372f $X=-0.19 $Y=1.305 $X2=1.585 $Y2=0.737
cc_52 VPB X 0.001239f $X=-0.19 $Y=1.305 $X2=1.26 $Y2=1.63
cc_53 VPB N_VPWR_c_338_n 0.0105686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_339_n 0.00496891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_340_n 0.0167189f $X=-0.19 $Y=1.305 $X2=0.805 $Y2=0.825
cc_56 VPB N_VPWR_c_341_n 0.0645247f $X=-0.19 $Y=1.305 $X2=1.585 $Y2=0.737
cc_57 VPB N_VPWR_c_342_n 0.0187397f $X=-0.19 $Y=1.305 $X2=2.6 $Y2=0.74
cc_58 VPB N_VPWR_c_337_n 0.057548f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.74
cc_59 VPB N_VPWR_c_344_n 0.00519718f $X=-0.19 $Y=1.305 $X2=2.72 $Y2=0.5
cc_60 VPB N_VPWR_c_345_n 0.00410958f $X=-0.19 $Y=1.305 $X2=1.26 $Y2=1.63
cc_61 N_A_85_193#_c_62_n N_D1_M1006_g 6.70019e-19 $X=0.805 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_85_193#_c_68_n N_D1_M1006_g 0.00724652f $X=1.26 $Y=1.63 $X2=0 $Y2=0
cc_63 N_A_85_193#_c_63_n N_D1_M1006_g 2.58508e-19 $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_64 N_A_85_193#_c_62_n D1 0.00532604f $X=0.805 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_85_193#_c_68_n D1 0.00879837f $X=1.26 $Y=1.63 $X2=0 $Y2=0
cc_66 N_A_85_193#_c_63_n D1 2.34781e-19 $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_67 N_A_85_193#_c_62_n N_D1_c_144_n 7.61856e-19 $X=0.805 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_85_193#_c_77_p N_D1_c_144_n 0.00306862f $X=1.585 $Y=0.737 $X2=0 $Y2=0
cc_69 N_A_85_193#_c_68_n N_D1_c_144_n 6.0605e-19 $X=1.26 $Y=1.63 $X2=0 $Y2=0
cc_70 N_A_85_193#_c_79_p N_D1_c_144_n 0.00146276f $X=1.75 $Y=0.737 $X2=0 $Y2=0
cc_71 N_A_85_193#_c_63_n N_D1_c_144_n 0.0113874f $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_72 N_A_85_193#_c_62_n N_D1_c_145_n 0.00338101f $X=0.805 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_85_193#_c_77_p N_D1_c_145_n 0.0110498f $X=1.585 $Y=0.737 $X2=0 $Y2=0
cc_74 N_A_85_193#_c_83_p N_D1_c_145_n 0.0107959f $X=1.75 $Y=0.39 $X2=0 $Y2=0
cc_75 N_A_85_193#_c_79_p N_D1_c_145_n 7.79452e-19 $X=1.75 $Y=0.737 $X2=0 $Y2=0
cc_76 N_A_85_193#_c_63_n N_D1_c_145_n 9.64409e-19 $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_77 N_A_85_193#_c_62_n N_D1_c_146_n 0.0104307f $X=0.805 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_85_193#_c_77_p N_D1_c_146_n 0.0152717f $X=1.585 $Y=0.737 $X2=0 $Y2=0
cc_79 N_A_85_193#_c_68_n N_D1_c_146_n 0.00456073f $X=1.26 $Y=1.63 $X2=0 $Y2=0
cc_80 N_A_85_193#_c_79_p N_D1_c_146_n 0.00673709f $X=1.75 $Y=0.737 $X2=0 $Y2=0
cc_81 N_A_85_193#_c_63_n N_D1_c_146_n 0.00196086f $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_82 N_A_85_193#_c_91_p C1 0.0170217f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A_85_193#_c_91_p N_C1_c_188_n 0.0034197f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A_85_193#_c_91_p N_C1_c_189_n 0.0106001f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A_85_193#_c_91_p B1 0.0188074f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_85_193#_c_91_p N_B1_c_221_n 0.0055091f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A_85_193#_c_91_p N_B1_c_222_n 0.0121263f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_85_193#_c_91_p N_A1_c_258_n 5.58779e-19 $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A_85_193#_c_98_p N_A1_c_258_n 0.00149039f $X=2.72 $Y=0.5 $X2=0 $Y2=0
cc_90 N_A_85_193#_M1009_d A1 0.00727297f $X=2.58 $Y=0.235 $X2=0 $Y2=0
cc_91 N_A_85_193#_c_91_p A1 0.0144642f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_85_193#_c_98_p A1 0.0287026f $X=2.72 $Y=0.5 $X2=0 $Y2=0
cc_93 N_A_85_193#_M1000_g N_X_c_321_n 0.00376139f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_85_193#_c_61_n N_X_c_321_n 0.00199737f $X=0.54 $Y=0.96 $X2=0 $Y2=0
cc_95 N_A_85_193#_c_62_n N_X_c_321_n 0.0379601f $X=0.805 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_85_193#_c_105_p N_X_c_321_n 0.0121826f $X=0.915 $Y=0.737 $X2=0 $Y2=0
cc_97 N_A_85_193#_c_63_n N_X_c_321_n 0.0159921f $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_98 N_A_85_193#_M1000_g X 0.00473458f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_85_193#_c_67_n X 0.0101403f $X=0.915 $Y=1.555 $X2=0 $Y2=0
cc_100 N_A_85_193#_c_67_n N_VPWR_M1000_d 0.00415129f $X=0.915 $Y=1.555 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_85_193#_M1000_g N_VPWR_c_338_n 0.0130927f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_85_193#_c_67_n N_VPWR_c_338_n 0.0181331f $X=0.915 $Y=1.555 $X2=0
+ $Y2=0
cc_103 N_A_85_193#_c_68_n N_VPWR_c_338_n 0.039861f $X=1.26 $Y=1.63 $X2=0 $Y2=0
cc_104 N_A_85_193#_c_63_n N_VPWR_c_338_n 0.00385044f $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_105 N_A_85_193#_M1000_g N_VPWR_c_340_n 0.00544582f $X=0.5 $Y=1.985 $X2=0
+ $Y2=0
cc_106 N_A_85_193#_c_68_n N_VPWR_c_341_n 0.0141722f $X=1.26 $Y=1.63 $X2=0 $Y2=0
cc_107 N_A_85_193#_M1006_s N_VPWR_c_337_n 0.00905805f $X=1.135 $Y=1.485 $X2=0
+ $Y2=0
cc_108 N_A_85_193#_M1000_g N_VPWR_c_337_n 0.0101021f $X=0.5 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_85_193#_c_68_n N_VPWR_c_337_n 0.00799167f $X=1.26 $Y=1.63 $X2=0 $Y2=0
cc_110 N_A_85_193#_c_62_n N_VGND_M1001_d 0.00152166f $X=0.805 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_85_193#_c_77_p N_VGND_M1001_d 0.0170098f $X=1.585 $Y=0.737 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_85_193#_c_105_p N_VGND_M1001_d 0.00566905f $X=0.915 $Y=0.737
+ $X2=-0.19 $Y2=-0.24
cc_113 N_A_85_193#_c_91_p N_VGND_M1004_d 0.00922042f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_85_193#_c_91_p N_VGND_c_414_n 0.0188848f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_85_193#_c_77_p N_VGND_c_417_n 0.00407811f $X=1.585 $Y=0.737 $X2=0
+ $Y2=0
cc_116 N_A_85_193#_c_83_p N_VGND_c_417_n 0.01843f $X=1.75 $Y=0.39 $X2=0 $Y2=0
cc_117 N_A_85_193#_c_91_p N_VGND_c_417_n 0.00251419f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_85_193#_c_91_p N_VGND_c_419_n 0.00251419f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A_85_193#_c_98_p N_VGND_c_419_n 0.0124668f $X=2.72 $Y=0.5 $X2=0 $Y2=0
cc_120 N_A_85_193#_c_61_n N_VGND_c_420_n 0.00585385f $X=0.54 $Y=0.96 $X2=0 $Y2=0
cc_121 N_A_85_193#_c_61_n N_VGND_c_421_n 0.00507064f $X=0.54 $Y=0.96 $X2=0 $Y2=0
cc_122 N_A_85_193#_c_77_p N_VGND_c_421_n 0.0286599f $X=1.585 $Y=0.737 $X2=0
+ $Y2=0
cc_123 N_A_85_193#_c_105_p N_VGND_c_421_n 0.0176019f $X=0.915 $Y=0.737 $X2=0
+ $Y2=0
cc_124 N_A_85_193#_c_83_p N_VGND_c_421_n 0.0119188f $X=1.75 $Y=0.39 $X2=0 $Y2=0
cc_125 N_A_85_193#_c_63_n N_VGND_c_421_n 0.0022468f $X=0.54 $Y=1.15 $X2=0 $Y2=0
cc_126 N_A_85_193#_M1011_d N_VGND_c_422_n 0.00243471f $X=1.61 $Y=0.235 $X2=0
+ $Y2=0
cc_127 N_A_85_193#_M1009_d N_VGND_c_422_n 0.0109769f $X=2.58 $Y=0.235 $X2=0
+ $Y2=0
cc_128 N_A_85_193#_c_61_n N_VGND_c_422_n 0.0128004f $X=0.54 $Y=0.96 $X2=0 $Y2=0
cc_129 N_A_85_193#_c_77_p N_VGND_c_422_n 0.00883577f $X=1.585 $Y=0.737 $X2=0
+ $Y2=0
cc_130 N_A_85_193#_c_105_p N_VGND_c_422_n 0.00111289f $X=0.915 $Y=0.737 $X2=0
+ $Y2=0
cc_131 N_A_85_193#_c_83_p N_VGND_c_422_n 0.0123586f $X=1.75 $Y=0.39 $X2=0 $Y2=0
cc_132 N_A_85_193#_c_91_p N_VGND_c_422_n 0.00933929f $X=2.6 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_85_193#_c_98_p N_VGND_c_422_n 0.00776141f $X=2.72 $Y=0.5 $X2=0 $Y2=0
cc_134 D1 C1 0.0155871f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_135 N_D1_c_144_n C1 0.00201874f $X=1.53 $Y=1.16 $X2=0 $Y2=0
cc_136 N_D1_c_146_n C1 0.0203079f $X=1.617 $Y=1.17 $X2=0 $Y2=0
cc_137 D1 N_C1_c_188_n 0.00133746f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_138 N_D1_c_144_n N_C1_c_188_n 0.0427505f $X=1.53 $Y=1.16 $X2=0 $Y2=0
cc_139 N_D1_c_146_n N_C1_c_188_n 7.9158e-19 $X=1.617 $Y=1.17 $X2=0 $Y2=0
cc_140 N_D1_c_145_n N_C1_c_189_n 0.0108956f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_141 N_D1_M1006_g N_C1_c_192_n 0.0427505f $X=1.595 $Y=1.985 $X2=0 $Y2=0
cc_142 N_D1_M1006_g N_VPWR_c_338_n 0.00309092f $X=1.595 $Y=1.985 $X2=0 $Y2=0
cc_143 N_D1_M1006_g N_VPWR_c_341_n 0.00357668f $X=1.595 $Y=1.985 $X2=0 $Y2=0
cc_144 D1 N_VPWR_c_341_n 0.0121075f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_145 N_D1_M1006_g N_VPWR_c_337_n 0.0066169f $X=1.595 $Y=1.985 $X2=0 $Y2=0
cc_146 D1 N_VPWR_c_337_n 0.00713192f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_147 N_D1_c_145_n N_VGND_c_417_n 0.00417376f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_148 N_D1_c_145_n N_VGND_c_421_n 0.00961048f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_149 N_D1_c_145_n N_VGND_c_422_n 0.00725697f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_150 C1 N_B1_M1003_g 0.00383306f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_151 N_C1_c_192_n N_B1_M1003_g 0.0406955f $X=2.07 $Y=1.38 $X2=0 $Y2=0
cc_152 C1 B1 0.070615f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_153 N_C1_c_188_n B1 0.0030349f $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_154 N_C1_c_192_n B1 9.59884e-19 $X=2.07 $Y=1.38 $X2=0 $Y2=0
cc_155 C1 N_B1_c_221_n 3.90035e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_156 N_C1_c_188_n N_B1_c_221_n 0.023893f $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_157 N_C1_c_189_n N_B1_c_222_n 0.0191988f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_158 C1 N_VPWR_c_341_n 0.0197479f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_159 N_C1_c_192_n N_VPWR_c_341_n 0.00357668f $X=2.07 $Y=1.38 $X2=0 $Y2=0
cc_160 C1 N_VPWR_c_337_n 0.0119459f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_161 N_C1_c_192_n N_VPWR_c_337_n 0.00548133f $X=2.07 $Y=1.38 $X2=0 $Y2=0
cc_162 C1 A_414_297# 0.00957729f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_163 N_C1_c_189_n N_VGND_c_414_n 0.00323586f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_164 N_C1_c_189_n N_VGND_c_417_n 0.00428022f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_165 N_C1_c_189_n N_VGND_c_422_n 0.00598352f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_166 B1 N_A1_c_257_n 3.54494e-19 $X=2.445 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_167 N_B1_c_221_n N_A1_c_257_n 0.0222681f $X=2.595 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_168 N_B1_M1003_g N_A1_M1010_g 0.0148559f $X=2.505 $Y=1.985 $X2=0 $Y2=0
cc_169 B1 N_A1_M1010_g 0.00459244f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_170 N_B1_c_222_n N_A1_c_258_n 0.0107816f $X=2.595 $Y=0.96 $X2=0 $Y2=0
cc_171 B1 A1 0.0212799f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_172 N_B1_c_221_n A1 0.00260566f $X=2.595 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B1_c_222_n A1 0.00311983f $X=2.595 $Y=0.96 $X2=0 $Y2=0
cc_174 N_B1_M1003_g N_VPWR_c_341_n 0.00357668f $X=2.505 $Y=1.985 $X2=0 $Y2=0
cc_175 B1 N_VPWR_c_341_n 0.0162318f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_176 N_B1_M1003_g N_VPWR_c_337_n 0.00611252f $X=2.505 $Y=1.985 $X2=0 $Y2=0
cc_177 B1 N_VPWR_c_337_n 0.0100203f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_178 B1 N_A_516_297#_M1003_d 0.0100165f $X=2.445 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_179 N_B1_M1003_g N_A_516_297#_c_392_n 0.00261795f $X=2.505 $Y=1.985 $X2=0
+ $Y2=0
cc_180 B1 N_A_516_297#_c_392_n 0.0596742f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_181 N_B1_M1003_g N_A_516_297#_c_394_n 6.44406e-19 $X=2.505 $Y=1.985 $X2=0
+ $Y2=0
cc_182 B1 N_A_516_297#_c_394_n 0.0137128f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_183 N_B1_c_222_n N_VGND_c_414_n 0.00329221f $X=2.595 $Y=0.96 $X2=0 $Y2=0
cc_184 N_B1_c_222_n N_VGND_c_419_n 0.00427293f $X=2.595 $Y=0.96 $X2=0 $Y2=0
cc_185 N_B1_c_222_n N_VGND_c_422_n 0.00648099f $X=2.595 $Y=0.96 $X2=0 $Y2=0
cc_186 N_A1_c_257_n N_A2_M1005_g 0.0299153f $X=3.215 $Y=1.33 $X2=0 $Y2=0
cc_187 N_A1_c_257_n A2 0.00176546f $X=3.215 $Y=1.33 $X2=0 $Y2=0
cc_188 A1 A2 0.0180848f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_189 N_A1_c_257_n N_A2_c_298_n 0.0197022f $X=3.215 $Y=1.33 $X2=0 $Y2=0
cc_190 A1 N_A2_c_298_n 5.34593e-19 $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A1_c_258_n N_A2_c_299_n 0.0409425f $X=3.225 $Y=0.965 $X2=0 $Y2=0
cc_192 A1 N_A2_c_299_n 0.0011504f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_193 N_A1_M1010_g N_VPWR_c_339_n 0.0028339f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A1_M1010_g N_VPWR_c_341_n 0.0057934f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A1_M1010_g N_VPWR_c_337_n 0.0110254f $X=3.215 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A1_M1010_g N_A_516_297#_c_392_n 0.0104547f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A1_M1010_g N_A_516_297#_c_397_n 0.0125122f $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_198 A1 N_A_516_297#_c_397_n 0.0154521f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A1_c_257_n N_A_516_297#_c_394_n 0.00376783f $X=3.215 $Y=1.33 $X2=0
+ $Y2=0
cc_200 N_A1_M1010_g N_A_516_297#_c_394_n 8.92169e-19 $X=3.215 $Y=1.985 $X2=0
+ $Y2=0
cc_201 A1 N_A_516_297#_c_394_n 0.0183287f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A1_c_258_n N_VGND_c_419_n 0.00363877f $X=3.225 $Y=0.965 $X2=0 $Y2=0
cc_203 A1 N_VGND_c_419_n 0.0277971f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_204 N_A1_c_258_n N_VGND_c_422_n 0.00588464f $X=3.225 $Y=0.965 $X2=0 $Y2=0
cc_205 A1 N_VGND_c_422_n 0.0203098f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_206 A1 A_660_47# 0.00507531f $X=2.905 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_207 N_A2_M1005_g N_VPWR_c_339_n 0.00291728f $X=3.635 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A2_M1005_g N_VPWR_c_342_n 0.00585385f $X=3.635 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A2_M1005_g N_VPWR_c_337_n 0.011589f $X=3.635 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A2_M1005_g N_A_516_297#_c_392_n 6.18506e-19 $X=3.635 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A2_M1005_g N_A_516_297#_c_397_n 0.0164998f $X=3.635 $Y=1.985 $X2=0
+ $Y2=0
cc_212 A2 N_A_516_297#_c_397_n 0.0286794f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_213 N_A2_c_298_n N_A_516_297#_c_397_n 0.00407812f $X=3.71 $Y=1.16 $X2=0 $Y2=0
cc_214 A2 N_VGND_c_416_n 0.0125224f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_215 N_A2_c_298_n N_VGND_c_416_n 0.00412826f $X=3.71 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A2_c_299_n N_VGND_c_416_n 0.00751723f $X=3.725 $Y=0.965 $X2=0 $Y2=0
cc_217 N_A2_c_299_n N_VGND_c_419_n 0.00585385f $X=3.725 $Y=0.965 $X2=0 $Y2=0
cc_218 N_A2_c_299_n N_VGND_c_422_n 0.011606f $X=3.725 $Y=0.965 $X2=0 $Y2=0
cc_219 X N_VPWR_c_340_n 0.0165311f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_220 N_X_M1000_s N_VPWR_c_337_n 0.00354753f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_221 X N_VPWR_c_337_n 0.00972063f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_222 N_X_c_321_n N_VGND_c_420_n 0.0211142f $X=0.3 $Y=0.4 $X2=0 $Y2=0
cc_223 N_X_M1001_s N_VGND_c_422_n 0.00265902f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_224 N_X_c_321_n N_VGND_c_422_n 0.0126319f $X=0.3 $Y=0.4 $X2=0 $Y2=0
cc_225 N_VPWR_c_337_n A_334_297# 0.00797857f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_226 N_VPWR_c_337_n A_414_297# 0.00920902f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_227 N_VPWR_c_337_n N_A_516_297#_M1003_d 0.0108501f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_228 N_VPWR_c_337_n N_A_516_297#_M1005_d 0.00311237f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_341_n N_A_516_297#_c_392_n 0.0173544f $X=3.325 $Y=2.72 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_337_n N_A_516_297#_c_392_n 0.0108549f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_231 N_VPWR_M1010_d N_A_516_297#_c_397_n 0.00489584f $X=3.29 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_339_n N_A_516_297#_c_397_n 0.0126919f $X=3.425 $Y=2.005 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_342_n N_A_516_297#_c_412_n 0.0167113f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_337_n N_A_516_297#_c_412_n 0.010297f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VGND_c_422_n A_660_47# 0.00258177f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

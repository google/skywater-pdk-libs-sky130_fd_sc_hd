* File: sky130_fd_sc_hd__and2_4.spice.pex
* Created: Thu Aug 27 14:07:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND2_4%A 3 6 8 11 12 13
r27 11 14 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.16
+ $X2=0.382 $Y2=1.325
r28 11 13 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.382 $Y=1.16
+ $X2=0.382 $Y2=0.995
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.16 $X2=0.35 $Y2=1.16
r30 8 12 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.53 $X2=0.28
+ $Y2=1.16
r31 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r32 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_4%B 3 6 8 11 12 13
c38 11 0 1.91186e-19 $X=0.895 $Y=1.16
r39 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.16
+ $X2=0.895 $Y2=1.325
r40 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.16
+ $X2=0.895 $Y2=0.995
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=1.16 $X2=0.895 $Y2=1.16
r42 8 12 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.895 $Y2=1.16
r43 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.985
+ $X2=0.905 $Y2=1.325
r44 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.835 $Y=0.56
+ $X2=0.835 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_4%A_27_47# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 37 39 40 43 45 46 48 50 56 59 66
c108 48 0 1.91186e-19 $X=1.255 $Y=1.02
r109 63 64 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.84 $Y=1.16
+ $X2=2.27 $Y2=1.16
r110 57 66 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.52 $Y=1.16 $X2=2.7
+ $Y2=1.16
r111 57 64 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.52 $Y=1.16
+ $X2=2.27 $Y2=1.16
r112 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.16 $X2=2.52 $Y2=1.16
r113 54 63 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.5 $Y=1.16
+ $X2=1.84 $Y2=1.16
r114 54 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.5 $Y=1.16 $X2=1.41
+ $Y2=1.16
r115 53 56 35.0893 $w=3.33e-07 $l=1.02e-06 $layer=LI1_cond $X=1.5 $Y=1.187
+ $X2=2.52 $Y2=1.187
r116 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.5
+ $Y=1.16 $X2=1.5 $Y2=1.16
r117 51 59 0.271299 $w=3.35e-07 $l=1.05e-07 $layer=LI1_cond $X=1.36 $Y=1.187
+ $X2=1.255 $Y2=1.187
r118 51 53 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.36 $Y=1.187
+ $X2=1.5 $Y2=1.187
r119 49 59 7.47207 $w=2.1e-07 $l=1.68e-07 $layer=LI1_cond $X=1.255 $Y=1.355
+ $X2=1.255 $Y2=1.187
r120 49 50 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=1.255 $Y=1.355
+ $X2=1.255 $Y2=1.58
r121 48 59 7.47207 $w=2.1e-07 $l=1.67e-07 $layer=LI1_cond $X=1.255 $Y=1.02
+ $X2=1.255 $Y2=1.187
r122 47 48 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.255 $Y=0.805
+ $X2=1.255 $Y2=1.02
r123 45 50 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.255 $Y2=1.58
r124 45 46 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=0.785 $Y2=1.665
r125 41 46 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.695 $Y=1.75
+ $X2=0.785 $Y2=1.665
r126 41 43 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.695 $Y=1.75
+ $X2=0.695 $Y2=1.96
r127 39 47 6.83868 $w=1.9e-07 $l=1.44914e-07 $layer=LI1_cond $X=1.15 $Y=0.71
+ $X2=1.255 $Y2=0.805
r128 39 40 42.3206 $w=1.88e-07 $l=7.25e-07 $layer=LI1_cond $X=1.15 $Y=0.71
+ $X2=0.425 $Y2=0.71
r129 35 40 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.425 $Y2=0.71
r130 35 37 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.26 $Y2=0.38
r131 31 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.16
r132 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.985
r133 28 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=1.16
r134 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=0.56
r135 24 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.325
+ $X2=2.27 $Y2=1.16
r136 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.27 $Y=1.325
+ $X2=2.27 $Y2=1.985
r137 21 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.27 $Y2=1.16
r138 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.27 $Y2=0.56
r139 17 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.16
r140 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.985
r141 14 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=0.995
+ $X2=1.84 $Y2=1.16
r142 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.84 $Y=0.995
+ $X2=1.84 $Y2=0.56
r143 10 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r144 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.985
r145 7 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r146 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r147 2 43 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.96
r148 1 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_4%VPWR 1 2 3 4 13 15 19 23 25 27 29 31 36 41 50
+ 53 57
r55 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 45 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 45 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 42 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=2.72
+ $X2=2.055 $Y2=2.72
r62 42 44 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.22 $Y=2.72
+ $X2=2.53 $Y2=2.72
r63 41 56 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.75 $Y=2.72
+ $X2=2.985 $Y2=2.72
r64 41 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.75 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 40 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 40 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=2.72
+ $X2=1.155 $Y2=2.72
r69 37 39 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.32 $Y=2.72
+ $X2=1.61 $Y2=2.72
r70 36 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=2.72
+ $X2=2.055 $Y2=2.72
r71 36 39 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.89 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 35 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r73 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r74 32 47 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r75 32 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 31 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=2.72
+ $X2=1.155 $Y2=2.72
r77 31 34 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=0.69
+ $Y2=2.72
r78 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 29 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 25 56 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.915 $Y=2.635
+ $X2=2.985 $Y2=2.72
r81 25 27 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.915 $Y=2.635
+ $X2=2.915 $Y2=2.02
r82 21 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2.72
r83 21 23 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2.02
r84 17 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.635
+ $X2=1.155 $Y2=2.72
r85 17 19 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.155 $Y=2.635
+ $X2=1.155 $Y2=2.02
r86 13 47 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r87 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2
r88 4 27 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=2.775
+ $Y=1.485 $X2=2.915 $Y2=2.02
r89 3 23 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=1.915
+ $Y=1.485 $X2=2.055 $Y2=2.02
r90 2 19 300 $w=1.7e-07 $l=6.1632e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.155 $Y2=2.02
r91 1 15 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_4%X 1 2 3 4 15 17 19 20 23 27 29 31 36 38 40 42
+ 45 47
r56 45 47 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=0.845
+ $X2=2.995 $Y2=0.85
r57 42 45 3.11269 $w=2.8e-07 $l=1.15e-07 $layer=LI1_cond $X=2.995 $Y=0.73
+ $X2=2.995 $Y2=0.845
r58 42 47 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=2.995 $Y=0.89
+ $X2=2.995 $Y2=0.85
r59 41 42 26.5473 $w=2.78e-07 $l=6.45e-07 $layer=LI1_cond $X=2.995 $Y=1.535
+ $X2=2.995 $Y2=0.89
r60 34 36 4.38803 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.625 $Y=0.68
+ $X2=1.72 $Y2=0.68
r61 32 40 4.43576 $w=2.27e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=1.65
+ $X2=2.485 $Y2=1.65
r62 31 41 6.90206 $w=2.3e-07 $l=1.88944e-07 $layer=LI1_cond $X=2.855 $Y=1.65
+ $X2=2.995 $Y2=1.535
r63 31 32 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.855 $Y=1.65
+ $X2=2.58 $Y2=1.65
r64 30 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=0.73
+ $X2=2.485 $Y2=0.73
r65 29 42 3.78936 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=2.855 $Y=0.73
+ $X2=2.995 $Y2=0.73
r66 29 30 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.855 $Y=0.73
+ $X2=2.58 $Y2=0.73
r67 25 40 1.99853 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.485 $Y=1.765
+ $X2=2.485 $Y2=1.65
r68 25 27 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.485 $Y=1.765
+ $X2=2.485 $Y2=1.96
r69 21 38 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.485 $Y=0.615
+ $X2=2.485 $Y2=0.73
r70 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.485 $Y=0.615
+ $X2=2.485 $Y2=0.42
r71 19 40 4.43576 $w=2.27e-07 $l=9.64883e-08 $layer=LI1_cond $X=2.39 $Y=1.647
+ $X2=2.485 $Y2=1.65
r72 19 20 34.3172 $w=2.23e-07 $l=6.7e-07 $layer=LI1_cond $X=2.39 $Y=1.647
+ $X2=1.72 $Y2=1.647
r73 17 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.39 $Y=0.73
+ $X2=2.485 $Y2=0.73
r74 17 36 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.39 $Y=0.73
+ $X2=1.72 $Y2=0.73
r75 13 20 6.87974 $w=2.25e-07 $l=1.5331e-07 $layer=LI1_cond $X=1.625 $Y=1.76
+ $X2=1.72 $Y2=1.647
r76 13 15 11.6746 $w=1.88e-07 $l=2e-07 $layer=LI1_cond $X=1.625 $Y=1.76
+ $X2=1.625 $Y2=1.96
r77 4 40 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.485 $X2=2.485 $Y2=1.62
r78 4 27 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=2.345
+ $Y=1.485 $X2=2.485 $Y2=1.96
r79 3 15 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.485 $X2=1.625 $Y2=1.96
r80 2 38 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.235 $X2=2.485 $Y2=0.76
r81 2 23 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.235 $X2=2.485 $Y2=0.42
r82 1 34 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.625 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__AND2_4%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r60 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r61 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r62 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r63 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r64 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r65 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r66 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.055
+ $Y2=0
r67 35 37 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.53
+ $Y2=0
r68 34 46 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.985
+ $Y2=0
r69 34 37 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.53
+ $Y2=0
r70 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r71 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r72 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r73 30 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r74 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.61
+ $Y2=0
r75 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.055
+ $Y2=0
r76 29 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.61
+ $Y2=0
r77 27 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r78 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r79 24 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r80 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.69
+ $Y2=0
r81 22 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r82 18 46 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.985 $Y2=0
r83 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.36
r84 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r85 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.36
r86 10 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r87 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r88 3 20 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.235 $X2=2.915 $Y2=0.36
r89 2 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.235 $X2=2.055 $Y2=0.36
r90 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.12 $Y2=0.36
.ends


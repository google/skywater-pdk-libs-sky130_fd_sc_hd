* File: sky130_fd_sc_hd__nor4bb_1.spice
* Created: Thu Aug 27 14:33:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor4bb_1.spice.pex"
.subckt sky130_fd_sc_hd__nor4bb_1  VNB VPB C_N D_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_C_N_M1002_g N_A_27_410#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.1092 PD=0.71 PS=1.36 NRD=4.284 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_205_93#_M1008_d N_D_N_M1008_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0609 PD=1.36 PS=0.71 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_205_93#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_27_410#_M1005_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=4.608 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_C_N_M1010_g N_A_27_410#_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.122612 AS=0.1092 PD=1.32 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_205_93#_M1011_d N_D_N_M1011_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1085 AS=0.122612 PD=1.36 PS=1.32 NRD=0 NRS=111.128 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_393_297# N_A_205_93#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.2559 PD=1.27 PS=2.52 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 A_477_297# N_A_27_410#_M1004_g A_393_297# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1001 A_573_297# N_B_M1001_g A_477_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.165 PD=1.27 PS=1.33 NRD=15.7403 NRS=21.6503 M=1 R=6.66667 SA=75001.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_573_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75001.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_38 VNB 0 1.59638e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__nor4bb_1.spice.SKY130_FD_SC_HD__NOR4BB_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__dlygate4sd3_1.spice.pex
* Created: Thu Aug 27 14:18:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A 3 7 9 11 18
c31 18 0 7.47284e-20 $X=0.49 $Y=1.16
r32 18 21 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.16
+ $X2=0.505 $Y2=1.325
r33 18 20 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.16
+ $X2=0.505 $Y2=0.995
r34 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r35 11 19 4.27171 $w=5.58e-07 $l=2e-07 $layer=LI1_cond $X=0.69 $Y=1.335 $X2=0.49
+ $Y2=1.335
r36 9 19 5.55322 $w=5.58e-07 $l=2.6e-07 $layer=LI1_cond $X=0.23 $Y=1.335
+ $X2=0.49 $Y2=1.335
r37 7 21 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.58 $Y=2.275
+ $X2=0.58 $Y2=1.325
r38 3 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.58 $Y=0.445
+ $X2=0.58 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_49_47# 1 2 9 13 15 16 17 18 22 25 29
c58 17 0 7.47284e-20 $X=0.945 $Y=1.895
r59 23 29 119.312 $w=5e-07 $l=1.115e-06 $layer=POLY_cond $X=1.175 $Y=1.16
+ $X2=1.175 $Y2=2.275
r60 23 25 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.175 $Y=1.16
+ $X2=1.175 $Y2=0.445
r61 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.16 $X2=1.06 $Y2=1.16
r62 20 22 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=1.05 $Y=1.785
+ $X2=1.05 $Y2=1.16
r63 19 22 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.05 $Y=0.885
+ $X2=1.05 $Y2=1.16
r64 17 20 6.82129 $w=2.2e-07 $l=1.53786e-07 $layer=LI1_cond $X=0.945 $Y=1.895
+ $X2=1.05 $Y2=1.785
r65 17 18 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=0.945 $Y=1.895
+ $X2=0.485 $Y2=1.895
r66 15 19 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.945 $Y=0.8
+ $X2=1.05 $Y2=0.885
r67 15 16 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.945 $Y=0.8
+ $X2=0.485 $Y2=0.8
r68 11 18 6.96441 $w=2.2e-07 $l=1.90208e-07 $layer=LI1_cond $X=0.342 $Y=2.005
+ $X2=0.485 $Y2=1.895
r69 11 13 8.2895 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=0.342 $Y=2.005
+ $X2=0.342 $Y2=2.21
r70 7 16 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.342 $Y=0.715
+ $X2=0.485 $Y2=0.8
r71 7 9 8.2895 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=0.342 $Y=0.715
+ $X2=0.342 $Y2=0.51
r72 2 13 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=2.065 $X2=0.37 $Y2=2.21
r73 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_285_47# 1 2 7 9 13 17 21 25 28
c58 25 0 1.28874e-19 $X=2.08 $Y=1.16
c59 7 0 7.47284e-20 $X=2.465 $Y=0.995
r60 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.16 $X2=2.08 $Y2=1.16
r61 23 28 0.164012 $w=5.6e-07 $l=2e-07 $layer=LI1_cond $X=1.725 $Y=1.335
+ $X2=1.525 $Y2=1.335
r62 23 25 7.58228 $w=5.58e-07 $l=3.55e-07 $layer=LI1_cond $X=1.725 $Y=1.335
+ $X2=2.08 $Y2=1.335
r63 19 28 6.76825 $w=4e-07 $l=2.8e-07 $layer=LI1_cond $X=1.525 $Y=1.615
+ $X2=1.525 $Y2=1.335
r64 19 21 17.1426 $w=3.98e-07 $l=5.95e-07 $layer=LI1_cond $X=1.525 $Y=1.615
+ $X2=1.525 $Y2=2.21
r65 15 28 6.76825 $w=4e-07 $l=2.8e-07 $layer=LI1_cond $X=1.525 $Y=1.055
+ $X2=1.525 $Y2=1.335
r66 15 17 15.702 $w=3.98e-07 $l=5.45e-07 $layer=LI1_cond $X=1.525 $Y=1.055
+ $X2=1.525 $Y2=0.51
r67 7 26 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=2.465 $Y=1.16
+ $X2=2.08 $Y2=1.16
r68 7 13 101.656 $w=5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.465 $Y=1.325
+ $X2=2.465 $Y2=2.275
r69 7 9 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.465 $Y=0.995 $X2=2.465
+ $Y2=0.445
r70 2 21 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=2.065 $X2=1.56 $Y2=2.21
r71 1 17 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.235 $X2=1.56 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%A_391_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c68 31 0 1.28874e-19 $X=3.06 $Y=1.16
c69 24 0 7.47284e-20 $X=2.59 $Y=1.895
r70 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.16
+ $X2=3.06 $Y2=1.325
r71 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.16
+ $X2=3.06 $Y2=0.995
r72 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.16 $X2=3.06 $Y2=1.16
r73 28 30 8.67984 $w=5.06e-07 $l=3.6e-07 $layer=LI1_cond $X=2.867 $Y=0.8
+ $X2=2.867 $Y2=1.16
r74 26 30 4.15671 $w=5.06e-07 $l=1.89222e-07 $layer=LI1_cond $X=2.815 $Y=1.325
+ $X2=2.867 $Y2=1.16
r75 26 27 12.2266 $w=4.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.815 $Y=1.325
+ $X2=2.815 $Y2=1.785
r76 24 27 7.91732 $w=2.2e-07 $l=2.74545e-07 $layer=LI1_cond $X=2.59 $Y=1.895
+ $X2=2.815 $Y2=1.785
r77 24 25 20.6916 $w=2.18e-07 $l=3.95e-07 $layer=LI1_cond $X=2.59 $Y=1.895
+ $X2=2.195 $Y2=1.895
r78 22 28 7.23163 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=2.59 $Y=0.8
+ $X2=2.867 $Y2=0.8
r79 22 23 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.59 $Y=0.8
+ $X2=2.195 $Y2=0.8
r80 18 25 6.94494 $w=2.2e-07 $l=1.87083e-07 $layer=LI1_cond $X=2.055 $Y=2.005
+ $X2=2.195 $Y2=1.895
r81 18 20 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=2.055 $Y=2.005
+ $X2=2.055 $Y2=2.21
r82 14 23 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.055 $Y=0.715
+ $X2=2.195 $Y2=0.8
r83 14 16 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=2.055 $Y=0.715
+ $X2=2.055 $Y2=0.51
r84 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.115 $Y=1.985
+ $X2=3.115 $Y2=1.325
r85 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.115 $Y=0.56
+ $X2=3.115 $Y2=0.995
r86 2 20 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=2.065 $X2=2.08 $Y2=2.21
r87 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.08 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%VPWR 1 2 11 15 18 19 20 30 31 34
r42 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r45 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 25 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 24 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 22 34 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.79 $Y2=2.72
r51 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 18 27 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 18 19 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.715 $Y=2.72
+ $X2=2.877 $Y2=2.72
r55 17 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.04 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 17 19 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=3.04 $Y=2.72
+ $X2=2.877 $Y2=2.72
r57 13 19 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.877 $Y=2.635
+ $X2=2.877 $Y2=2.72
r58 13 15 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=2.877 $Y=2.635
+ $X2=2.877 $Y2=2.34
r59 9 34 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=2.635
+ $X2=0.79 $Y2=2.72
r60 9 11 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.79 $Y=2.635
+ $X2=0.79 $Y2=2.34
r61 2 15 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=2.065 $X2=2.875 $Y2=2.34
r62 1 11 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=2.065 $X2=0.79 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%X 1 2 7 8 9 10 11 12 24 43
r16 43 44 1.9254 $w=3.83e-07 $l=3.5e-08 $layer=LI1_cond $X=3.402 $Y=1.53
+ $X2=3.402 $Y2=1.495
r17 24 41 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.455 $Y=0.85
+ $X2=3.455 $Y2=0.825
r18 11 12 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=3.402 $Y=1.87
+ $X2=3.402 $Y2=2.21
r19 11 29 5.47785 $w=3.83e-07 $l=1.83e-07 $layer=LI1_cond $X=3.402 $Y=1.87
+ $X2=3.402 $Y2=1.687
r20 10 29 3.95123 $w=3.83e-07 $l=1.32e-07 $layer=LI1_cond $X=3.402 $Y=1.555
+ $X2=3.402 $Y2=1.687
r21 10 43 0.74834 $w=3.83e-07 $l=2.5e-08 $layer=LI1_cond $X=3.402 $Y=1.555
+ $X2=3.402 $Y2=1.53
r22 10 44 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.455 $Y=1.47
+ $X2=3.455 $Y2=1.495
r23 9 10 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=3.455 $Y=1.19
+ $X2=3.455 $Y2=1.47
r24 8 41 1.77574 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=3.402 $Y=0.795
+ $X2=3.402 $Y2=0.825
r25 8 9 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=3.455 $Y=0.88
+ $X2=3.455 $Y2=1.19
r26 8 24 1.23476 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=3.455 $Y=0.88 $X2=3.455
+ $Y2=0.85
r27 7 8 8.53107 $w=3.83e-07 $l=2.85e-07 $layer=LI1_cond $X=3.402 $Y=0.51
+ $X2=3.402 $Y2=0.795
r28 2 12 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.485 $X2=3.325 $Y2=2.21
r29 1 7 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.235 $X2=3.325 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLYGATE4SD3_1%VGND 1 2 11 15 18 19 20 30 31 34
r43 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r45 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r46 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r47 25 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r48 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r49 24 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r50 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r51 22 34 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.79
+ $Y2=0
r52 22 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.15
+ $Y2=0
r53 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r54 18 27 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.53
+ $Y2=0
r55 18 19 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.877
+ $Y2=0
r56 17 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.45
+ $Y2=0
r57 17 19 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.877
+ $Y2=0
r58 13 19 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.877 $Y=0.085
+ $X2=2.877 $Y2=0
r59 13 15 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=2.877 $Y=0.085
+ $X2=2.877 $Y2=0.38
r60 9 34 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r61 9 11 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.38
r62 2 15 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.875 $Y2=0.38
r63 1 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.655
+ $Y=0.235 $X2=0.79 $Y2=0.38
.ends


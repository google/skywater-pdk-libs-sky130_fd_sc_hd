* File: sky130_fd_sc_hd__o2bb2ai_1.pex.spice
* Created: Tue Sep  1 19:24:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%A1_N 1 3 6 8 14
c23 8 0 6.1502e-21 $X=0.23 $Y=1.19
r24 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.27 $Y=1.16
+ $X2=0.485 $Y2=1.16
r25 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r26 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.16
r27 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.985
r28 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.16
r29 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%A2_N 3 6 10 13 14 15 19
c40 15 0 6.1502e-21 $X=0.905 $Y=0.995
r41 14 19 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.905 $Y=1.16
+ $X2=0.715 $Y2=1.16
r42 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.16
+ $X2=0.905 $Y2=0.995
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.16 $X2=0.905 $Y2=1.16
r44 10 19 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.715 $Y2=1.16
r45 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r46 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r47 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.845 $Y=0.56
+ $X2=0.845 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%A_112_297# 1 2 7 9 12 14 15 18 20 21 24 29
+ 30 32 34
r60 32 35 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=1.16
+ $X2=1.32 $Y2=1.325
r61 32 34 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=1.16
+ $X2=1.32 $Y2=0.995
r62 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=1.16 $X2=1.385 $Y2=1.16
r63 30 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.255 $Y=0.825
+ $X2=1.255 $Y2=0.995
r64 29 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.255 $Y=1.495
+ $X2=1.255 $Y2=1.325
r65 22 30 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.17 $Y=0.655
+ $X2=1.17 $Y2=0.825
r66 22 24 8.98228 $w=3.38e-07 $l=2.65e-07 $layer=LI1_cond $X=1.17 $Y=0.655
+ $X2=1.17 $Y2=0.39
r67 20 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.17 $Y=1.58
+ $X2=1.255 $Y2=1.495
r68 20 21 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.17 $Y=1.58
+ $X2=0.82 $Y2=1.58
r69 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.695 $Y=1.665
+ $X2=0.82 $Y2=1.58
r70 16 18 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.695 $Y=1.665
+ $X2=0.695 $Y2=1.96
r71 14 33 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=1.385 $Y2=1.16
r72 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=1.895 $Y2=1.16
r73 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.325
+ $X2=1.895 $Y2=1.16
r74 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.895 $Y=1.325
+ $X2=1.895 $Y2=1.985
r75 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=1.16
r76 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=0.56
r77 2 18 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=1.485 $X2=0.695 $Y2=1.96
r78 1 24 91 $w=1.7e-07 $l=3.1305e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.235 $X2=1.165 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%B2 1 3 6 8 11 14
c41 11 0 1.58219e-19 $X=2.315 $Y=1.16
r42 13 14 14.7118 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.53 $Y=1.325
+ $X2=2.53 $Y2=1.53
r43 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.315
+ $Y=1.16 $X2=2.315 $Y2=1.16
r44 8 13 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.445 $Y=1.2
+ $X2=2.53 $Y2=1.325
r45 8 10 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.445 $Y=1.2 $X2=2.315
+ $Y2=1.2
r46 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.16
r47 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.985
r48 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%B1 1 3 6 8 13
c25 8 0 1.58219e-19 $X=2.99 $Y=1.19
r26 10 13 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=2.95 $Y2=1.16
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r28 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.325
+ $X2=2.735 $Y2=1.16
r29 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.735 $Y=1.325
+ $X2=2.735 $Y2=1.985
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.735 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.735 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%VPWR 1 2 3 10 12 18 20 22 26 28 33 42 46
r46 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 37 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r49 37 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r51 34 42 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=1.77 $Y=2.72 $X2=1.38
+ $Y2=2.72
r52 34 36 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.77 $Y=2.72
+ $X2=2.53 $Y2=2.72
r53 33 45 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.82 $Y=2.72 $X2=3.02
+ $Y2=2.72
r54 33 36 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.82 $Y=2.72
+ $X2=2.53 $Y2=2.72
r55 32 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 29 39 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.2
+ $Y2=2.72
r58 29 31 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.69
+ $Y2=2.72
r59 28 42 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=1.38
+ $Y2=2.72
r60 28 31 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=0.69
+ $Y2=2.72
r61 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 26 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 22 25 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.945 $Y=1.63
+ $X2=2.945 $Y2=2.31
r64 20 45 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=3.02 $Y2=2.72
r65 20 25 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.945 $Y=2.635
+ $X2=2.945 $Y2=2.31
r66 16 42 3.08259 $w=7.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=2.635
+ $X2=1.38 $Y2=2.72
r67 16 18 10.3507 $w=7.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.38 $Y=2.635
+ $X2=1.38 $Y2=1.96
r68 12 15 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.275 $Y=1.63
+ $X2=0.275 $Y2=2.31
r69 10 39 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.2 $Y2=2.72
r70 10 15 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.275 $Y2=2.31
r71 3 25 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=1.485 $X2=2.945 $Y2=2.31
r72 3 22 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=1.485 $X2=2.945 $Y2=1.63
r73 2 18 150 $w=1.7e-07 $l=8.29156e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=1.485 $X2=1.605 $Y2=1.96
r74 1 15 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.31
r75 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%Y 1 2 8 10 16 19
r34 19 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.105 $Y=1.87
+ $X2=2.105 $Y2=2.3
r35 16 19 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.105 $Y=1.665
+ $X2=2.105 $Y2=1.87
r36 13 16 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.725 $Y=1.58
+ $X2=2.105 $Y2=1.58
r37 10 12 9.71523 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=1.685 $Y=0.605
+ $X2=1.685 $Y2=0.79
r38 8 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=1.495
+ $X2=1.725 $Y2=1.58
r39 8 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.725 $Y=1.495
+ $X2=1.725 $Y2=0.79
r40 2 24 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.485 $X2=2.105 $Y2=2.3
r41 2 16 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.485 $X2=2.105 $Y2=1.62
r42 1 10 182 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.685 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%VGND 1 2 7 9 13 16 17 18 28 29
r43 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r44 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r46 23 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r47 22 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r48 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r49 20 32 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r50 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r51 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r52 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r53 16 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.44 $Y=0 $X2=2.07
+ $Y2=0
r54 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0 $X2=2.525
+ $Y2=0
r55 15 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.61 $Y=0 $X2=2.99
+ $Y2=0
r56 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0 $X2=2.525
+ $Y2=0
r57 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0
r58 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0.39
r59 7 32 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r60 7 9 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.39
r61 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.235 $X2=2.525 $Y2=0.39
r62 1 9 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O2BB2AI_1%A_394_47# 1 2 9 11 12 15
r30 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.945 $Y=0.725
+ $X2=2.945 $Y2=0.39
r31 11 13 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.78 $Y=0.815
+ $X2=2.945 $Y2=0.725
r32 11 12 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.78 $Y=0.815
+ $X2=2.27 $Y2=0.815
r33 7 12 7.31368 $w=1.8e-07 $l=1.84594e-07 $layer=LI1_cond $X=2.125 $Y=0.725
+ $X2=2.27 $Y2=0.815
r34 7 9 4.76873 $w=2.88e-07 $l=1.2e-07 $layer=LI1_cond $X=2.125 $Y=0.725
+ $X2=2.125 $Y2=0.605
r35 2 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.81
+ $Y=0.235 $X2=2.945 $Y2=0.39
r36 1 9 182 $w=1.7e-07 $l=4.32262e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.105 $Y2=0.605
.ends


* File: sky130_fd_sc_hd__and2b_2.pxi.spice
* Created: Tue Sep  1 18:57:14 2020
* 
x_PM_SKY130_FD_SC_HD__AND2B_2%A_N N_A_N_M1008_g N_A_N_M1005_g A_N N_A_N_c_58_n
+ A_N A_N PM_SKY130_FD_SC_HD__AND2B_2%A_N
x_PM_SKY130_FD_SC_HD__AND2B_2%A_27_413# N_A_27_413#_M1008_d N_A_27_413#_M1005_s
+ N_A_27_413#_M1000_g N_A_27_413#_M1003_g N_A_27_413#_c_95_n N_A_27_413#_c_96_n
+ N_A_27_413#_c_97_n N_A_27_413#_c_89_n N_A_27_413#_c_90_n N_A_27_413#_c_91_n
+ N_A_27_413#_c_92_n N_A_27_413#_c_93_n PM_SKY130_FD_SC_HD__AND2B_2%A_27_413#
x_PM_SKY130_FD_SC_HD__AND2B_2%B N_B_c_150_n N_B_M1006_g N_B_M1002_g B B
+ PM_SKY130_FD_SC_HD__AND2B_2%B
x_PM_SKY130_FD_SC_HD__AND2B_2%A_212_413# N_A_212_413#_M1003_s
+ N_A_212_413#_M1000_d N_A_212_413#_c_182_n N_A_212_413#_M1007_g
+ N_A_212_413#_M1001_g N_A_212_413#_c_183_n N_A_212_413#_M1009_g
+ N_A_212_413#_M1004_g N_A_212_413#_c_190_n N_A_212_413#_c_184_n
+ N_A_212_413#_c_185_n N_A_212_413#_c_186_n N_A_212_413#_c_206_n
+ N_A_212_413#_c_187_n PM_SKY130_FD_SC_HD__AND2B_2%A_212_413#
x_PM_SKY130_FD_SC_HD__AND2B_2%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_M1004_d
+ N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_262_n VPWR N_VPWR_c_263_n
+ N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_259_n
+ PM_SKY130_FD_SC_HD__AND2B_2%VPWR
x_PM_SKY130_FD_SC_HD__AND2B_2%X N_X_M1007_s N_X_M1001_s N_X_c_304_n X
+ N_X_c_303_n N_X_c_301_n N_X_c_315_n X X PM_SKY130_FD_SC_HD__AND2B_2%X
x_PM_SKY130_FD_SC_HD__AND2B_2%VGND N_VGND_M1008_s N_VGND_M1002_d N_VGND_M1009_d
+ N_VGND_c_325_n N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n
+ VGND N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n
+ PM_SKY130_FD_SC_HD__AND2B_2%VGND
cc_1 VNB N_A_N_M1008_g 0.0394803f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_A_N_c_58_n 0.0326513f $X=-0.19 $Y=-0.24 $X2=0.365 $Y2=1.16
cc_3 VNB A_N 0.0221698f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0.85
cc_4 VNB N_A_27_413#_M1000_g 0.0104956f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_5 VNB N_A_27_413#_M1003_g 0.02179f $X=-0.19 $Y=-0.24 $X2=0.365 $Y2=1.16
cc_6 VNB N_A_27_413#_c_89_n 0.0040409f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_7 VNB N_A_27_413#_c_90_n 0.00373597f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.53
cc_8 VNB N_A_27_413#_c_91_n 0.00458034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_413#_c_92_n 0.00788638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_413#_c_93_n 0.0513758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_c_150_n 0.0182419f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_12 VNB N_B_M1002_g 0.0372957f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_13 VNB N_A_212_413#_c_182_n 0.0158203f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_14 VNB N_A_212_413#_c_183_n 0.0207514f $X=-0.19 $Y=-0.24 $X2=0.372 $Y2=0.995
cc_15 VNB N_A_212_413#_c_184_n 0.00291494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_212_413#_c_185_n 0.0149587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_212_413#_c_186_n 0.0042882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_212_413#_c_187_n 0.0508429f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_259_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_301_n 7.86697e-19 $X=-0.19 $Y=-0.24 $X2=0.372 $Y2=1.325
cc_21 VNB N_VGND_c_325_n 0.0103099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_326_n 0.0180257f $X=-0.19 $Y=-0.24 $X2=0.365 $Y2=1.16
cc_23 VNB N_VGND_c_327_n 4.09712e-19 $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.85
cc_24 VNB N_VGND_c_328_n 0.0101057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_329_n 0.0250683f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.16
cc_26 VNB N_VGND_c_330_n 0.0387178f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.53
cc_27 VNB N_VGND_c_331_n 0.0153481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_332_n 0.00529996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_333_n 0.183316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_A_N_M1005_g 0.0640217f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_31 VPB N_A_N_c_58_n 0.00732313f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.16
cc_32 VPB A_N 0.0147197f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0.85
cc_33 VPB N_A_27_413#_M1000_g 0.05115f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_34 VPB N_A_27_413#_c_95_n 0.0021894f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0.85
cc_35 VPB N_A_27_413#_c_96_n 0.00886909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_413#_c_97_n 0.0109634f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.16
cc_37 VPB N_A_27_413#_c_90_n 0.00961334f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.53
cc_38 VPB N_B_c_150_n 0.0664143f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_39 VPB N_B_M1006_g 0.0257968f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_40 VPB B 0.00643373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_212_413#_M1001_g 0.021985f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.16
cc_42 VPB N_A_212_413#_M1004_g 0.0253035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_212_413#_c_190_n 0.00613575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_212_413#_c_185_n 0.00731252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_212_413#_c_186_n 0.00249332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_212_413#_c_187_n 0.00985248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_260_n 0.00227888f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.16
cc_48 VPB N_VPWR_c_261_n 0.0100799f $X=-0.19 $Y=1.305 $X2=0.372 $Y2=0.995
cc_49 VPB N_VPWR_c_262_n 0.0380806f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.85
cc_50 VPB N_VPWR_c_263_n 0.015299f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.16
cc_51 VPB N_VPWR_c_264_n 0.0189132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_265_n 0.00507571f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_266_n 0.018616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_267_n 0.0197068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_259_n 0.0444927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_X_c_301_n 0.00148119f $X=-0.19 $Y=1.305 $X2=0.372 $Y2=1.325
cc_57 N_A_N_c_58_n N_A_27_413#_M1000_g 0.0216609f $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_N_M1005_g N_A_27_413#_c_95_n 0.00239329f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_59 N_A_N_M1005_g N_A_27_413#_c_96_n 0.0188468f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_60 A_N N_A_27_413#_c_96_n 0.00847314f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_61 N_A_N_c_58_n N_A_27_413#_c_97_n 6.06494e-19 $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_62 A_N N_A_27_413#_c_97_n 0.0158932f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_63 N_A_N_M1008_g N_A_27_413#_c_89_n 0.00513589f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_64 A_N N_A_27_413#_c_89_n 0.00303884f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_65 N_A_N_c_58_n N_A_27_413#_c_90_n 0.00838026f $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_66 A_N N_A_27_413#_c_90_n 0.0366833f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_67 N_A_N_M1008_g N_A_27_413#_c_92_n 0.00295745f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_68 A_N N_A_27_413#_c_92_n 0.0269815f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_69 N_A_N_M1008_g N_A_27_413#_c_93_n 0.0216609f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_70 A_N N_A_27_413#_c_93_n 3.62695e-19 $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_71 N_A_N_M1005_g N_A_212_413#_c_190_n 7.69706e-19 $X=0.47 $Y=2.275 $X2=0
+ $Y2=0
cc_72 N_A_N_M1005_g N_VPWR_c_260_n 0.0101169f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_73 N_A_N_M1005_g N_VPWR_c_263_n 0.00347311f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_74 N_A_N_M1005_g N_VPWR_c_259_n 0.00511644f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_75 N_A_N_M1008_g N_VGND_c_326_n 0.0119738f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_N_c_58_n N_VGND_c_326_n 8.02374e-19 $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_77 A_N N_VGND_c_326_n 0.0209484f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_78 N_A_N_M1008_g N_VGND_c_330_n 0.0046653f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A_N_M1008_g N_VGND_c_333_n 0.00857541f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_80 A_N N_VGND_c_333_n 0.00196247f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_81 N_A_27_413#_M1000_g N_B_c_150_n 0.0398867f $X=0.985 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_82 N_A_27_413#_c_93_n N_B_c_150_n 0.00277424f $X=1.09 $Y=0.97 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_27_413#_M1000_g N_B_M1002_g 2.7762e-19 $X=0.985 $Y=2.275 $X2=0 $Y2=0
cc_84 N_A_27_413#_M1003_g N_B_M1002_g 0.0380868f $X=1.41 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_27_413#_c_93_n N_B_M1002_g 0.00320805f $X=1.09 $Y=0.97 $X2=0 $Y2=0
cc_86 N_A_27_413#_M1000_g N_A_212_413#_c_190_n 0.0172006f $X=0.985 $Y=2.275
+ $X2=0 $Y2=0
cc_87 N_A_27_413#_c_96_n N_A_212_413#_c_190_n 0.017661f $X=0.62 $Y=1.9 $X2=0
+ $Y2=0
cc_88 N_A_27_413#_c_90_n N_A_212_413#_c_190_n 0.0216612f $X=0.737 $Y=1.785 $X2=0
+ $Y2=0
cc_89 N_A_27_413#_M1003_g N_A_212_413#_c_184_n 0.00586327f $X=1.41 $Y=0.445
+ $X2=0 $Y2=0
cc_90 N_A_27_413#_c_91_n N_A_212_413#_c_184_n 0.00621632f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_91 N_A_27_413#_c_92_n N_A_212_413#_c_184_n 0.0103761f $X=1.09 $Y=0.97 $X2=0
+ $Y2=0
cc_92 N_A_27_413#_c_93_n N_A_212_413#_c_184_n 0.00420658f $X=1.09 $Y=0.97 $X2=0
+ $Y2=0
cc_93 N_A_27_413#_M1000_g N_A_212_413#_c_185_n 0.00635329f $X=0.985 $Y=2.275
+ $X2=0 $Y2=0
cc_94 N_A_27_413#_c_90_n N_A_212_413#_c_185_n 0.019776f $X=0.737 $Y=1.785 $X2=0
+ $Y2=0
cc_95 N_A_27_413#_c_92_n N_A_212_413#_c_185_n 0.0274557f $X=1.09 $Y=0.97 $X2=0
+ $Y2=0
cc_96 N_A_27_413#_c_93_n N_A_212_413#_c_185_n 0.0141397f $X=1.09 $Y=0.97 $X2=0
+ $Y2=0
cc_97 N_A_27_413#_M1003_g N_A_212_413#_c_206_n 0.00610483f $X=1.41 $Y=0.445
+ $X2=0 $Y2=0
cc_98 N_A_27_413#_c_91_n N_A_212_413#_c_206_n 0.0182853f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_99 N_A_27_413#_c_92_n N_A_212_413#_c_206_n 0.00405807f $X=1.09 $Y=0.97 $X2=0
+ $Y2=0
cc_100 N_A_27_413#_c_93_n N_A_212_413#_c_206_n 0.0062871f $X=1.09 $Y=0.97 $X2=0
+ $Y2=0
cc_101 N_A_27_413#_M1000_g N_VPWR_c_260_n 0.00465679f $X=0.985 $Y=2.275 $X2=0
+ $Y2=0
cc_102 N_A_27_413#_c_96_n N_VPWR_c_260_n 0.0252018f $X=0.62 $Y=1.9 $X2=0 $Y2=0
cc_103 N_A_27_413#_c_95_n N_VPWR_c_263_n 0.0102625f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_104 N_A_27_413#_c_96_n N_VPWR_c_263_n 0.0025049f $X=0.62 $Y=1.9 $X2=0 $Y2=0
cc_105 N_A_27_413#_M1000_g N_VPWR_c_266_n 0.00564994f $X=0.985 $Y=2.275 $X2=0
+ $Y2=0
cc_106 N_A_27_413#_M1005_s N_VPWR_c_259_n 0.00375546f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_107 N_A_27_413#_M1000_g N_VPWR_c_259_n 0.0105412f $X=0.985 $Y=2.275 $X2=0
+ $Y2=0
cc_108 N_A_27_413#_c_95_n N_VPWR_c_259_n 0.00640243f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_109 N_A_27_413#_c_96_n N_VPWR_c_259_n 0.00577167f $X=0.62 $Y=1.9 $X2=0 $Y2=0
cc_110 N_A_27_413#_M1003_g N_VGND_c_327_n 0.00183913f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_111 N_A_27_413#_M1003_g N_VGND_c_330_n 0.00388886f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_112 N_A_27_413#_c_91_n N_VGND_c_330_n 0.0139933f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_27_413#_M1008_d N_VGND_c_333_n 0.00388065f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_114 N_A_27_413#_M1003_g N_VGND_c_333_n 0.00681766f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_c_91_n N_VGND_c_333_n 0.00898141f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_116 N_A_27_413#_c_92_n N_VGND_c_333_n 0.00993011f $X=1.09 $Y=0.97 $X2=0 $Y2=0
cc_117 N_A_27_413#_c_93_n N_VGND_c_333_n 0.00515873f $X=1.09 $Y=0.97 $X2=0 $Y2=0
cc_118 N_B_M1002_g N_A_212_413#_c_182_n 0.0247788f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_119 N_B_c_150_n N_A_212_413#_M1001_g 0.0161917f $X=1.425 $Y=1.895 $X2=0 $Y2=0
cc_120 N_B_c_150_n N_A_212_413#_c_190_n 0.0107208f $X=1.425 $Y=1.895 $X2=0 $Y2=0
cc_121 B N_A_212_413#_c_190_n 0.025312f $X=2.095 $Y=1.87 $X2=0 $Y2=0
cc_122 N_B_M1002_g N_A_212_413#_c_184_n 0.00557851f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B_c_150_n N_A_212_413#_c_185_n 0.036453f $X=1.425 $Y=1.895 $X2=0 $Y2=0
cc_124 N_B_M1002_g N_A_212_413#_c_185_n 0.0154812f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_125 B N_A_212_413#_c_185_n 0.0317236f $X=2.095 $Y=1.87 $X2=0 $Y2=0
cc_126 B N_A_212_413#_c_186_n 0.0149134f $X=2.095 $Y=1.87 $X2=0 $Y2=0
cc_127 N_B_M1002_g N_A_212_413#_c_187_n 0.0220914f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_128 B N_A_212_413#_c_187_n 0.00172058f $X=2.095 $Y=1.87 $X2=0 $Y2=0
cc_129 B N_VPWR_M1006_d 0.00771626f $X=2.095 $Y=1.87 $X2=0 $Y2=0
cc_130 N_B_M1006_g N_VPWR_c_266_n 0.00585385f $X=1.425 $Y=2.275 $X2=0 $Y2=0
cc_131 N_B_c_150_n N_VPWR_c_267_n 0.00202247f $X=1.425 $Y=1.895 $X2=0 $Y2=0
cc_132 N_B_M1006_g N_VPWR_c_267_n 0.00363903f $X=1.425 $Y=2.275 $X2=0 $Y2=0
cc_133 B N_VPWR_c_267_n 0.0451162f $X=2.095 $Y=1.87 $X2=0 $Y2=0
cc_134 N_B_M1006_g N_VPWR_c_259_n 0.0119149f $X=1.425 $Y=2.275 $X2=0 $Y2=0
cc_135 B N_VPWR_c_259_n 0.00319716f $X=2.095 $Y=1.87 $X2=0 $Y2=0
cc_136 N_B_c_150_n N_X_c_303_n 5.1312e-19 $X=1.425 $Y=1.895 $X2=0 $Y2=0
cc_137 N_B_M1002_g N_VGND_c_327_n 0.0163118f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_138 N_B_M1002_g N_VGND_c_330_n 0.0046653f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_139 N_B_M1002_g N_VGND_c_333_n 0.00799591f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A_212_413#_c_190_n N_VPWR_c_260_n 0.0159244f $X=1.205 $Y=2.225 $X2=0
+ $Y2=0
cc_141 N_A_212_413#_M1004_g N_VPWR_c_262_n 0.00494189f $X=2.74 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_212_413#_M1001_g N_VPWR_c_264_n 0.0055908f $X=2.32 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_212_413#_M1004_g N_VPWR_c_264_n 0.00566002f $X=2.74 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_212_413#_c_190_n N_VPWR_c_266_n 0.0129171f $X=1.205 $Y=2.225 $X2=0
+ $Y2=0
cc_145 N_A_212_413#_M1001_g N_VPWR_c_267_n 0.00949595f $X=2.32 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_212_413#_M1000_d N_VPWR_c_259_n 0.00308576f $X=1.06 $Y=2.065 $X2=0
+ $Y2=0
cc_147 N_A_212_413#_M1001_g N_VPWR_c_259_n 0.0113689f $X=2.32 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_212_413#_M1004_g N_VPWR_c_259_n 0.0111778f $X=2.74 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_212_413#_c_190_n N_VPWR_c_259_n 0.0105781f $X=1.205 $Y=2.225 $X2=0
+ $Y2=0
cc_150 N_A_212_413#_c_183_n N_X_c_304_n 0.00516243f $X=2.74 $Y=0.985 $X2=0 $Y2=0
cc_151 N_A_212_413#_M1001_g N_X_c_303_n 0.00384387f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_212_413#_M1004_g N_X_c_303_n 0.00545323f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_212_413#_c_187_n N_X_c_303_n 8.13882e-19 $X=2.74 $Y=1.155 $X2=0 $Y2=0
cc_154 N_A_212_413#_c_182_n N_X_c_301_n 0.0040252f $X=2.32 $Y=0.985 $X2=0 $Y2=0
cc_155 N_A_212_413#_M1001_g N_X_c_301_n 0.0039659f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_212_413#_c_183_n N_X_c_301_n 0.00979203f $X=2.74 $Y=0.985 $X2=0 $Y2=0
cc_157 N_A_212_413#_M1004_g N_X_c_301_n 0.0119105f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_212_413#_c_185_n N_X_c_301_n 0.00483562f $X=1.905 $Y=1.135 $X2=0
+ $Y2=0
cc_159 N_A_212_413#_c_186_n N_X_c_301_n 0.0289559f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_212_413#_c_187_n N_X_c_301_n 0.0264604f $X=2.74 $Y=1.155 $X2=0 $Y2=0
cc_161 N_A_212_413#_c_183_n N_X_c_315_n 0.00315687f $X=2.74 $Y=0.985 $X2=0 $Y2=0
cc_162 N_A_212_413#_c_187_n N_X_c_315_n 8.20839e-19 $X=2.74 $Y=1.155 $X2=0 $Y2=0
cc_163 N_A_212_413#_M1001_g X 0.0135943f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_212_413#_M1004_g X 0.00671036f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_212_413#_c_182_n N_VGND_c_327_n 0.00907204f $X=2.32 $Y=0.985 $X2=0
+ $Y2=0
cc_166 N_A_212_413#_c_183_n N_VGND_c_327_n 6.65279e-19 $X=2.74 $Y=0.985 $X2=0
+ $Y2=0
cc_167 N_A_212_413#_c_185_n N_VGND_c_327_n 0.00129558f $X=1.905 $Y=1.135 $X2=0
+ $Y2=0
cc_168 N_A_212_413#_c_186_n N_VGND_c_327_n 0.0155077f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_169 N_A_212_413#_c_187_n N_VGND_c_327_n 6.3588e-19 $X=2.74 $Y=1.155 $X2=0
+ $Y2=0
cc_170 N_A_212_413#_c_183_n N_VGND_c_329_n 0.0054252f $X=2.74 $Y=0.985 $X2=0
+ $Y2=0
cc_171 N_A_212_413#_c_206_n N_VGND_c_330_n 0.0165109f $X=1.2 $Y=0.445 $X2=0
+ $Y2=0
cc_172 N_A_212_413#_c_182_n N_VGND_c_331_n 0.0046653f $X=2.32 $Y=0.985 $X2=0
+ $Y2=0
cc_173 N_A_212_413#_c_183_n N_VGND_c_331_n 0.00564131f $X=2.74 $Y=0.985 $X2=0
+ $Y2=0
cc_174 N_A_212_413#_M1003_s N_VGND_c_333_n 0.00239557f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_175 N_A_212_413#_c_182_n N_VGND_c_333_n 0.00796766f $X=2.32 $Y=0.985 $X2=0
+ $Y2=0
cc_176 N_A_212_413#_c_183_n N_VGND_c_333_n 0.0111716f $X=2.74 $Y=0.985 $X2=0
+ $Y2=0
cc_177 N_A_212_413#_c_206_n N_VGND_c_333_n 0.0136184f $X=1.2 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_259_n N_X_M1001_s 0.00227401f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_179 N_VPWR_c_264_n X 0.0105213f $X=2.865 $Y=2.72 $X2=0 $Y2=0
cc_180 N_VPWR_c_259_n X 0.0108709f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_181 N_X_c_304_n N_VGND_c_331_n 0.0140878f $X=2.562 $Y=0.658 $X2=0 $Y2=0
cc_182 N_X_M1007_s N_VGND_c_333_n 0.00393857f $X=2.395 $Y=0.235 $X2=0 $Y2=0
cc_183 N_X_c_304_n N_VGND_c_333_n 0.00889354f $X=2.562 $Y=0.658 $X2=0 $Y2=0
cc_184 N_VGND_c_333_n A_297_47# 0.0105263f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

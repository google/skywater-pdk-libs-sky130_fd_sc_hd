* File: sky130_fd_sc_hd__a22oi_1.spice.pex
* Created: Thu Aug 27 14:02:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A22OI_1%B2 3 6 8 9 13 15
c30 13 0 7.30641e-20 $X=0.41 $Y=1.16
c31 6 0 1.14647e-19 $X=0.47 $Y=1.985
r32 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=1.325
r33 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=0.995
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r35 9 14 0.797386 $w=4.48e-07 $l=3e-08 $layer=LI1_cond $X=0.35 $Y=1.19 $X2=0.35
+ $Y2=1.16
r36 8 14 8.23965 $w=4.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.35 $Y=0.85 $X2=0.35
+ $Y2=1.16
r37 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r38 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_1%B1 3 6 8 9 13 15
c41 8 0 7.30641e-20 $X=1.155 $Y=0.85
r42 14 17 10.2591 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=0.93 $Y=1.175
+ $X2=1.115 $Y2=1.175
r43 13 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=1.325
r44 13 15 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=0.995
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=1.16 $X2=0.93 $Y2=1.16
r46 9 17 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.115 $Y2=1.175
r47 8 17 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=1.115 $Y=0.85
+ $X2=1.115 $Y2=1.075
r48 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.985
+ $X2=0.89 $Y2=1.325
r49 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.85 $Y=0.56 $X2=0.85
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_1%A1 3 6 8 9 13 15 25
c35 25 0 1.81634e-19 $X=1.635 $Y=1.19
c36 8 0 6.4496e-20 $X=1.635 $Y=0.85
r37 17 21 0.416767 $w=2.1e-07 $l=1e-07 $layer=LI1_cond $X=1.595 $Y=1.075
+ $X2=1.595 $Y2=1.175
r38 13 16 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.712 $Y=1.16
+ $X2=1.712 $Y2=1.325
r39 13 15 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.712 $Y=1.16
+ $X2=1.712 $Y2=0.995
r40 13 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r41 9 25 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.635 $Y2=1.175
r42 9 21 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.595 $Y2=1.175
r43 8 17 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=1.595 $Y=0.85
+ $X2=1.595 $Y2=1.075
r44 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.985
+ $X2=1.83 $Y2=1.325
r45 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.56 $X2=1.83
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_1%A2 3 6 8 11 12 13
c33 11 0 2.4613e-19 $X=2.25 $Y=1.16
c34 6 0 1.71143e-19 $X=2.25 $Y=1.985
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.25 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r37 8 12 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.095 $Y=1.16
+ $X2=2.25 $Y2=1.16
r38 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.325
+ $X2=2.25 $Y2=1.16
r39 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.25 $Y=1.325 $X2=2.25
+ $Y2=1.985
r40 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.19 $Y=0.56 $X2=2.19
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_1%Y 1 2 3 4 13 14 16 19 25 28 29 30 32 36 37
+ 39 40 48 55
c91 55 0 1.71143e-19 $X=1.84 $Y=1.555
c92 36 0 1.14647e-19 $X=1.1 $Y=2.34
c93 32 0 1.81018e-19 $X=2.59 $Y=1.495
r94 40 55 10.2115 $w=2.18e-07 $l=1.83e-07 $layer=LI1_cond $X=1.657 $Y=1.555
+ $X2=1.84 $Y2=1.555
r95 40 48 2.20012 $w=2.18e-07 $l=4.2e-08 $layer=LI1_cond $X=1.657 $Y=1.555
+ $X2=1.615 $Y2=1.555
r96 40 48 2.64949 $w=1.78e-07 $l=4.3e-08 $layer=LI1_cond $X=1.572 $Y=1.535
+ $X2=1.615 $Y2=1.535
r97 40 45 70.6737 $w=1.78e-07 $l=1.147e-06 $layer=LI1_cond $X=1.572 $Y=1.535
+ $X2=0.425 $Y2=1.535
r98 39 45 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.535
+ $X2=0.425 $Y2=1.535
r99 36 37 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=2.36
+ $X2=0.935 $Y2=2.36
r100 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.59 $Y=0.825
+ $X2=2.59 $Y2=1.495
r101 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=0.74
+ $X2=2.59 $Y2=0.825
r102 29 30 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.505 $Y=0.74
+ $X2=2.125 $Y2=0.74
r103 28 30 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.035 $Y=0.655
+ $X2=2.125 $Y2=0.74
r104 27 28 9.24242 $w=1.78e-07 $l=1.5e-07 $layer=LI1_cond $X=2.035 $Y=0.505
+ $X2=2.035 $Y2=0.655
r105 25 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=1.58
+ $X2=2.59 $Y2=1.495
r106 25 55 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.505 $Y=1.58
+ $X2=1.84 $Y2=1.58
r107 21 24 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=1.06 $Y=0.38
+ $X2=1.62 $Y2=0.38
r108 19 27 7.0541 $w=2.5e-07 $l=1.63936e-07 $layer=LI1_cond $X=1.945 $Y=0.38
+ $X2=2.035 $Y2=0.505
r109 19 24 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.945 $Y=0.38
+ $X2=1.62 $Y2=0.38
r110 18 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.26 $Y2=2.38
r111 18 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.935 $Y2=2.38
r112 14 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=2.38
r113 14 16 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=1.66
r114 13 39 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.26 $Y=1.625 $X2=0.26
+ $Y2=1.535
r115 13 16 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.66
r116 4 36 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r117 3 34 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r118 3 16 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r119 2 24 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.42
r120 1 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.925
+ $Y=0.235 $X2=1.06 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_1%A_109_297# 1 2 7 9 14
r27 12 14 5.26246 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.68 $Y=1.96
+ $X2=0.825 $Y2=1.96
r28 9 10 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.955 $Y=1.935
+ $X2=1.475 $Y2=1.935
r29 7 10 19.463 $w=2.57e-07 $l=4.12492e-07 $layer=LI1_cond $X=1.065 $Y=1.94
+ $X2=1.475 $Y2=1.935
r30 7 14 9.53746 $w=2.88e-07 $l=2.4e-07 $layer=LI1_cond $X=1.065 $Y=1.94
+ $X2=0.825 $Y2=1.94
r31 2 9 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2
r32 1 12 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_1%VPWR 1 2 9 11 13 15 17 25 31 35
c40 2 0 1.81018e-19 $X=2.325 $Y=1.485
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r43 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r45 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 26 31 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=1.622 $Y2=2.72
r47 26 28 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=2.07 $Y2=2.72
r48 25 34 4.10655 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=2.72 $X2=2.56
+ $Y2=2.72
r49 25 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 24 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 19 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 17 31 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.622 $Y2=2.72
r54 17 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 15 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 15 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 11 34 3.14151 $w=2.65e-07 $l=1.14039e-07 $layer=LI1_cond $X=2.492 $Y=2.635
+ $X2=2.56 $Y2=2.72
r58 11 13 26.7454 $w=2.63e-07 $l=6.15e-07 $layer=LI1_cond $X=2.492 $Y=2.635
+ $X2=2.492 $Y2=2.02
r59 7 31 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.622 $Y=2.635
+ $X2=1.622 $Y2=2.72
r60 7 9 9.06588 $w=3.73e-07 $l=2.95e-07 $layer=LI1_cond $X=1.622 $Y=2.635
+ $X2=1.622 $Y2=2.34
r61 2 13 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.02
r62 1 9 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.485 $X2=1.62 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_1%VGND 1 2 7 9 11 13 15 17 30
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r34 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r35 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r36 21 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r37 20 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r38 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r39 18 26 5.92045 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.272
+ $Y2=0
r40 18 20 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.69
+ $Y2=0
r41 17 29 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.532
+ $Y2=0
r42 17 23 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.07
+ $Y2=0
r43 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r44 15 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r45 11 29 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=2.47 $Y=0.085
+ $X2=2.532 $Y2=0
r46 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.47 $Y=0.085
+ $X2=2.47 $Y2=0.4
r47 7 26 2.88432 $w=4.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.272 $Y2=0
r48 7 9 11.2963 $w=4.48e-07 $l=4.25e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.32 $Y2=0.51
r49 2 13 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.235 $X2=2.47 $Y2=0.4
r50 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends


* File: sky130_fd_sc_hd__a2bb2oi_2.spice.pex
* Created: Thu Aug 27 14:03:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%B1 3 6 8 10 13 17 18 20 21 23 29 31 41
c75 31 0 1.20878e-19 $X=0.545 $Y=0.995
r76 29 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.16
+ $X2=0.545 $Y2=1.325
r77 29 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.16
+ $X2=0.545 $Y2=0.995
r78 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.545
+ $Y=1.16 $X2=0.545 $Y2=1.16
r79 23 41 7.2872 $w=5.38e-07 $l=5.3e-08 $layer=LI1_cond $X=0.657 $Y=1.345
+ $X2=0.71 $Y2=1.345
r80 23 30 2.48076 $w=5.38e-07 $l=1.12e-07 $layer=LI1_cond $X=0.657 $Y=1.345
+ $X2=0.545 $Y2=1.345
r81 23 41 2.0877 $w=1.68e-07 $l=3.2e-08 $layer=LI1_cond $X=0.742 $Y=1.53
+ $X2=0.71 $Y2=1.53
r82 21 30 6.97712 $w=5.38e-07 $l=3.15e-07 $layer=LI1_cond $X=0.23 $Y=1.345
+ $X2=0.545 $Y2=1.345
r83 20 23 62.5005 $w=1.68e-07 $l=9.58e-07 $layer=LI1_cond $X=1.7 $Y=1.53
+ $X2=0.742 $Y2=1.53
r84 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=1.16 $X2=1.865 $Y2=1.16
r85 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.865 $Y=1.445
+ $X2=1.7 $Y2=1.53
r86 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.865 $Y=1.445
+ $X2=1.865 $Y2=1.16
r87 11 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.325
+ $X2=1.865 $Y2=1.16
r88 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.865 $Y=1.325
+ $X2=1.865 $Y2=1.985
r89 8 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=0.995
+ $X2=1.865 $Y2=1.16
r90 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.865 $Y=0.995
+ $X2=1.865 $Y2=0.56
r91 6 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.605 $Y=1.985
+ $X2=0.605 $Y2=1.325
r92 3 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.605 $Y=0.56
+ $X2=0.605 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%B2 1 3 6 8 10 13 15 22
c43 1 0 6.86556e-20 $X=1.025 $Y=0.995
r44 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.235 $Y=1.16
+ $X2=1.445 $Y2=1.16
r45 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.025 $Y=1.16
+ $X2=1.235 $Y2=1.16
r46 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.235
+ $Y=1.16 $X2=1.235 $Y2=1.16
r47 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.325
+ $X2=1.445 $Y2=1.16
r48 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.445 $Y=1.325
+ $X2=1.445 $Y2=1.985
r49 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.445 $Y2=1.16
r50 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.445 $Y2=0.56
r51 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=1.325
+ $X2=1.025 $Y2=1.16
r52 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.025 $Y=1.325
+ $X2=1.025 $Y2=1.985
r53 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%A_442_21# 1 2 3 10 12 15 17 19 22 24 26 30
+ 32 36 40 44 45 47
r106 48 50 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.285 $Y=1.16
+ $X2=2.705 $Y2=1.16
r107 45 50 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.915 $Y=1.16
+ $X2=2.705 $Y2=1.16
r108 44 46 21.0935 $w=2.14e-07 $l=3.7e-07 $layer=LI1_cond $X=2.975 $Y=1.16
+ $X2=2.975 $Y2=1.53
r109 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.16 $X2=2.915 $Y2=1.16
r110 42 44 19.6682 $w=2.14e-07 $l=3.45e-07 $layer=LI1_cond $X=2.975 $Y=0.815
+ $X2=2.975 $Y2=1.16
r111 38 40 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.695 $Y=1.615
+ $X2=4.695 $Y2=1.62
r112 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.695 $Y=0.725
+ $X2=4.695 $Y2=0.39
r113 33 47 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=0.815
+ $X2=3.855 $Y2=0.815
r114 32 34 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.53 $Y=0.815
+ $X2=4.695 $Y2=0.725
r115 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.53 $Y=0.815
+ $X2=4.02 $Y2=0.815
r116 28 47 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.855 $Y=0.725
+ $X2=3.855 $Y2=0.815
r117 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.855 $Y=0.725
+ $X2=3.855 $Y2=0.39
r118 27 46 2.08775 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.12 $Y=1.53
+ $X2=2.975 $Y2=1.53
r119 26 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.57 $Y=1.53
+ $X2=4.695 $Y2=1.615
r120 26 27 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=4.57 $Y=1.53
+ $X2=3.12 $Y2=1.53
r121 25 42 1.75188 $w=1.8e-07 $l=1.45e-07 $layer=LI1_cond $X=3.12 $Y=0.815
+ $X2=2.975 $Y2=0.815
r122 24 47 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=0.815
+ $X2=3.855 $Y2=0.815
r123 24 25 35.1212 $w=1.78e-07 $l=5.7e-07 $layer=LI1_cond $X=3.69 $Y=0.815
+ $X2=3.12 $Y2=0.815
r124 20 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.325
+ $X2=2.705 $Y2=1.16
r125 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.705 $Y=1.325
+ $X2=2.705 $Y2=1.985
r126 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.705 $Y2=1.16
r127 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.705 $Y2=0.56
r128 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.325
+ $X2=2.285 $Y2=1.16
r129 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.285 $Y=1.325
+ $X2=2.285 $Y2=1.985
r130 10 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=0.995
+ $X2=2.285 $Y2=1.16
r131 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.285 $Y=0.995
+ $X2=2.285 $Y2=0.56
r132 3 40 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.56
+ $Y=1.485 $X2=4.695 $Y2=1.62
r133 2 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.56
+ $Y=0.235 $X2=4.695 $Y2=0.39
r134 1 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.72
+ $Y=0.235 $X2=3.855 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%A1_N 1 3 6 8 10 13 15 22
r47 20 22 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.845 $Y=1.16
+ $X2=4.065 $Y2=1.16
r48 17 20 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=3.645 $Y=1.16
+ $X2=3.845 $Y2=1.16
r49 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.16 $X2=3.845 $Y2=1.16
r50 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.065 $Y=1.325
+ $X2=4.065 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.065 $Y=1.325
+ $X2=4.065 $Y2=1.985
r52 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.065 $Y=0.995
+ $X2=4.065 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.065 $Y=0.995
+ $X2=4.065 $Y2=0.56
r54 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.325
+ $X2=3.645 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.645 $Y=1.325
+ $X2=3.645 $Y2=1.985
r56 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=0.995
+ $X2=3.645 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.645 $Y=0.995
+ $X2=3.645 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%A2_N 1 3 6 8 10 13 15 22
r39 20 22 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=4.705 $Y=1.16
+ $X2=4.905 $Y2=1.16
r40 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.705
+ $Y=1.16 $X2=4.705 $Y2=1.16
r41 17 20 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=4.485 $Y=1.16
+ $X2=4.705 $Y2=1.16
r42 15 21 8.04091 $w=1.98e-07 $l=1.45e-07 $layer=LI1_cond $X=4.85 $Y=1.175
+ $X2=4.705 $Y2=1.175
r43 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.325
+ $X2=4.905 $Y2=1.16
r44 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.905 $Y=1.325
+ $X2=4.905 $Y2=1.985
r45 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=0.995
+ $X2=4.905 $Y2=1.16
r46 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.905 $Y=0.995
+ $X2=4.905 $Y2=0.56
r47 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.485 $Y=1.325
+ $X2=4.485 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.485 $Y=1.325
+ $X2=4.485 $Y2=1.985
r49 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.485 $Y=0.995
+ $X2=4.485 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.485 $Y=0.995
+ $X2=4.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%A_54_297# 1 2 3 4 15 17 18 21 23 29 30 33
+ 35
r43 31 33 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.915 $Y=2.295
+ $X2=2.915 $Y2=1.96
r44 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.79 $Y=2.38
+ $X2=2.915 $Y2=2.295
r45 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.79 $Y=2.38 $X2=2.2
+ $Y2=2.38
r46 26 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.075 $Y=2.295
+ $X2=2.2 $Y2=2.38
r47 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.075 $Y=2.295
+ $X2=2.075 $Y2=1.96
r48 25 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=1.955
+ $X2=2.075 $Y2=1.96
r49 24 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.36 $Y=1.87
+ $X2=1.235 $Y2=1.87
r50 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.95 $Y=1.87
+ $X2=2.075 $Y2=1.955
r51 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.95 $Y=1.87 $X2=1.36
+ $Y2=1.87
r52 19 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=1.955
+ $X2=1.235 $Y2=1.87
r53 19 21 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.235 $Y=1.955
+ $X2=1.235 $Y2=1.96
r54 17 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.11 $Y=1.87
+ $X2=1.235 $Y2=1.87
r55 17 18 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.11 $Y=1.87 $X2=0.52
+ $Y2=1.87
r56 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.395 $Y=1.955
+ $X2=0.52 $Y2=1.87
r57 13 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.395 $Y=1.955
+ $X2=0.395 $Y2=1.96
r58 4 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.78
+ $Y=1.485 $X2=2.915 $Y2=1.96
r59 3 28 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=1.485 $X2=2.075 $Y2=1.96
r60 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.1
+ $Y=1.485 $X2=1.235 $Y2=1.96
r61 1 15 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.27
+ $Y=1.485 $X2=0.395 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%VPWR 1 2 3 14 16 20 24 26 28 38 39 42 45
+ 48
r76 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r77 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r78 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r79 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 39 49 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=3.91 $Y2=2.72
r81 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r82 36 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.98 $Y=2.72
+ $X2=3.855 $Y2=2.72
r83 36 38 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.98 $Y=2.72
+ $X2=5.29 $Y2=2.72
r84 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r85 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r86 32 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r87 32 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r88 31 34 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r90 29 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.78 $Y=2.72
+ $X2=1.655 $Y2=2.72
r91 29 31 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.78 $Y=2.72
+ $X2=2.07 $Y2=2.72
r92 28 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.855 $Y2=2.72
r93 28 34 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.45 $Y2=2.72
r94 26 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 22 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=2.635
+ $X2=3.855 $Y2=2.72
r96 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.855 $Y=2.635
+ $X2=3.855 $Y2=2.3
r97 18 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=2.635
+ $X2=1.655 $Y2=2.72
r98 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.655 $Y=2.635
+ $X2=1.655 $Y2=2.3
r99 17 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.94 $Y=2.72
+ $X2=0.815 $Y2=2.72
r100 16 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.53 $Y=2.72
+ $X2=1.655 $Y2=2.72
r101 16 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.53 $Y=2.72
+ $X2=0.94 $Y2=2.72
r102 12 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.635
+ $X2=0.815 $Y2=2.72
r103 12 14 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=2.635
+ $X2=0.815 $Y2=2.3
r104 3 24 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.485 $X2=3.855 $Y2=2.3
r105 2 20 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.485 $X2=1.655 $Y2=2.3
r106 1 14 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.485 $X2=0.815 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%Y 1 2 3 10 14 21 23 24 25 33
c50 21 0 1.20878e-19 $X=1.4 $Y=0.775
r51 29 33 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=2.515 $Y=1.515
+ $X2=2.515 $Y2=1.53
r52 25 33 1.39088 $w=2.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.515 $Y=1.565
+ $X2=2.515 $Y2=1.53
r53 25 29 1.39088 $w=2.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.515 $Y=1.48
+ $X2=2.515 $Y2=1.515
r54 24 25 11.5244 $w=2.88e-07 $l=2.9e-07 $layer=LI1_cond $X=2.515 $Y=1.19
+ $X2=2.515 $Y2=1.48
r55 22 24 11.3257 $w=2.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.515 $Y=0.905
+ $X2=2.515 $Y2=1.19
r56 22 23 3.21907 $w=3.1e-07 $l=9.94987e-08 $layer=LI1_cond $X=2.515 $Y=0.905
+ $X2=2.495 $Y2=0.815
r57 19 21 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0.775
+ $X2=1.4 $Y2=0.775
r58 12 23 3.21907 $w=3.1e-07 $l=9e-08 $layer=LI1_cond $X=2.495 $Y=0.725
+ $X2=2.495 $Y2=0.815
r59 12 14 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=0.725
+ $X2=2.495 $Y2=0.39
r60 10 23 3.35592 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0.815
+ $X2=2.495 $Y2=0.815
r61 10 21 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=2.33 $Y=0.815 $X2=1.4
+ $Y2=0.815
r62 3 25 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=1.485 $X2=2.495 $Y2=1.62
r63 2 14 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.235 $X2=2.495 $Y2=0.39
r64 1 19 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.235 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%A_662_297# 1 2 3 12 14 16 17 18 20 23
r34 18 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=2.295
+ $X2=5.115 $Y2=2.38
r35 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.115 $Y=2.295
+ $X2=5.115 $Y2=1.62
r36 16 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.99 $Y=2.38
+ $X2=5.115 $Y2=2.38
r37 16 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.99 $Y=2.38 $X2=4.4
+ $Y2=2.38
r38 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.275 $Y=2.295
+ $X2=4.4 $Y2=2.38
r39 14 25 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=4.275 $Y=1.965
+ $X2=4.275 $Y2=1.875
r40 14 15 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=4.275 $Y=1.965
+ $X2=4.275 $Y2=2.295
r41 13 23 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.56 $Y=1.875
+ $X2=3.435 $Y2=1.875
r42 12 25 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.15 $Y=1.875
+ $X2=4.275 $Y2=1.875
r43 12 13 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=4.15 $Y=1.875
+ $X2=3.56 $Y2=1.875
r44 3 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.485 $X2=5.115 $Y2=2.3
r45 3 20 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.485 $X2=5.115 $Y2=1.62
r46 2 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.14
+ $Y=1.485 $X2=4.275 $Y2=1.96
r47 1 23 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=3.31
+ $Y=1.485 $X2=3.435 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%VGND 1 2 3 4 5 18 22 26 30 33 34 36 37 39
+ 40 41 47 64 65 68 73 76
r83 75 76 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.435 $Y=0.235
+ $X2=3.52 $Y2=0.235
r84 71 75 8.31648 $w=6.38e-07 $l=4.45e-07 $layer=LI1_cond $X=2.99 $Y=0.235
+ $X2=3.435 $Y2=0.235
r85 71 73 10.3234 $w=6.38e-07 $l=1.6e-07 $layer=LI1_cond $X=2.99 $Y=0.235
+ $X2=2.83 $Y2=0.235
r86 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r87 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r88 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r89 62 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r90 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r91 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r92 59 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r93 58 76 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=3.52
+ $Y2=0
r94 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r95 55 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r96 55 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r97 54 73 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.83
+ $Y2=0
r98 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r99 52 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.075
+ $Y2=0
r100 52 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.53
+ $Y2=0
r101 50 69 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r102 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r103 47 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0 $X2=2.075
+ $Y2=0
r104 47 49 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=1.99 $Y=0 $X2=0.69
+ $Y2=0
r105 41 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r106 41 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r107 39 61 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.03 $Y=0 $X2=4.83
+ $Y2=0
r108 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0 $X2=5.115
+ $Y2=0
r109 38 64 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.2 $Y=0 $X2=5.29
+ $Y2=0
r110 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.2 $Y=0 $X2=5.115
+ $Y2=0
r111 36 58 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=3.91
+ $Y2=0
r112 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.275
+ $Y2=0
r113 35 61 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.36 $Y=0 $X2=4.83
+ $Y2=0
r114 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.36 $Y=0 $X2=4.275
+ $Y2=0
r115 33 44 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.31 $Y=0 $X2=0.23
+ $Y2=0
r116 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=0 $X2=0.395
+ $Y2=0
r117 32 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.69
+ $Y2=0
r118 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.395
+ $Y2=0
r119 28 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0
r120 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0.39
r121 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.275 $Y=0.085
+ $X2=4.275 $Y2=0
r122 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.275 $Y=0.085
+ $X2=4.275 $Y2=0.39
r123 20 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0
r124 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0.39
r125 16 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.395 $Y=0.085
+ $X2=0.395 $Y2=0
r126 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.395 $Y=0.085
+ $X2=0.395 $Y2=0.39
r127 5 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.98
+ $Y=0.235 $X2=5.115 $Y2=0.39
r128 4 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.14
+ $Y=0.235 $X2=4.275 $Y2=0.39
r129 3 75 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=2.78
+ $Y=0.235 $X2=3.435 $Y2=0.39
r130 2 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.235 $X2=2.075 $Y2=0.39
r131 1 18 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.27
+ $Y=0.235 $X2=0.395 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_2%A_136_47# 1 2 7 9 13
c21 9 0 6.86556e-20 $X=0.815 $Y=0.73
r22 11 16 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=0.9 $Y=0.365
+ $X2=0.775 $Y2=0.365
r23 11 13 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=0.9 $Y=0.365
+ $X2=1.655 $Y2=0.365
r24 7 16 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.775 $Y=0.475
+ $X2=0.775 $Y2=0.365
r25 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.775 $Y=0.475
+ $X2=0.775 $Y2=0.73
r26 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.235 $X2=1.655 $Y2=0.39
r27 1 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.68
+ $Y=0.235 $X2=0.815 $Y2=0.39
r28 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.68
+ $Y=0.235 $X2=0.815 $Y2=0.73
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o41a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.650000 1.075000 7.735000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 1.075000 6.360000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.330000 1.075000 4.960000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.075000 4.040000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 1.075000 3.165000 1.275000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 1.685000 0.905000 ;
        RECT 0.085000 0.905000 0.345000 1.465000 ;
        RECT 0.085000 1.465000 1.685000 1.665000 ;
        RECT 0.515000 0.255000 0.845000 0.715000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 0.255000 1.685000 0.715000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.085000  0.085000 0.345000 0.545000 ;
        RECT 1.015000  0.085000 1.185000 0.545000 ;
        RECT 1.855000  0.085000 2.105000 0.885000 ;
        RECT 3.655000  0.085000 3.875000 0.545000 ;
        RECT 4.445000  0.085000 4.715000 0.545000 ;
        RECT 5.305000  0.085000 5.915000 0.545000 ;
        RECT 6.685000  0.085000 6.955000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.085000 1.835000 0.345000 2.635000 ;
        RECT 1.015000 1.835000 1.185000 2.635000 ;
        RECT 1.855000 1.465000 2.025000 2.635000 ;
        RECT 2.715000 1.835000 2.965000 2.635000 ;
        RECT 6.655000 1.785000 6.985000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 1.075000 2.665000 1.245000 ;
      RECT 0.515000 1.245000 2.545000 1.295000 ;
      RECT 2.195000 1.295000 2.545000 1.445000 ;
      RECT 2.195000 1.445000 3.825000 1.615000 ;
      RECT 2.195000 1.615000 2.545000 2.465000 ;
      RECT 2.295000 0.255000 3.485000 0.465000 ;
      RECT 2.295000 0.635000 3.045000 0.905000 ;
      RECT 2.295000 0.905000 2.665000 1.075000 ;
      RECT 3.135000 1.835000 3.405000 2.295000 ;
      RECT 3.135000 2.295000 4.325000 2.465000 ;
      RECT 3.235000 0.465000 3.485000 0.735000 ;
      RECT 3.235000 0.735000 7.595000 0.905000 ;
      RECT 3.575000 1.615000 3.825000 2.125000 ;
      RECT 3.995000 1.445000 5.165000 1.615000 ;
      RECT 3.995000 1.615000 4.325000 2.295000 ;
      RECT 4.075000 0.255000 4.245000 0.735000 ;
      RECT 4.495000 1.785000 4.665000 2.295000 ;
      RECT 4.495000 2.295000 6.145000 2.465000 ;
      RECT 4.835000 1.615000 5.165000 2.115000 ;
      RECT 4.915000 0.255000 5.085000 0.735000 ;
      RECT 5.395000 1.445000 7.595000 1.615000 ;
      RECT 5.395000 1.615000 5.645000 2.115000 ;
      RECT 5.815000 1.785000 6.145000 2.295000 ;
      RECT 6.240000 0.255000 6.410000 0.735000 ;
      RECT 6.315000 1.615000 6.485000 2.455000 ;
      RECT 7.265000 0.255000 7.595000 0.735000 ;
      RECT 7.265000 1.615000 7.595000 2.465000 ;
  END
END sky130_fd_sc_hd__o41a_4
END LIBRARY

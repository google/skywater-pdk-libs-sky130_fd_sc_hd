* File: sky130_fd_sc_hd__and4_4.spice.pex
* Created: Thu Aug 27 14:08:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4_4%A 1 3 6 8 9 16
r31 13 16 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r32 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r33 8 9 16.7716 $w=2.03e-07 $l=3.1e-07 $layer=LI1_cond $X=0.227 $Y=0.85
+ $X2=0.227 $Y2=1.16
r34 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r35 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r36 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_4%B 3 6 8 9 10 15 16 17
r37 16 25 4.90054 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.042 $Y=1.16
+ $X2=1.042 $Y2=0.995
r38 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.925 $Y2=1.325
r39 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.16
+ $X2=0.925 $Y2=0.995
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.16 $X2=0.925 $Y2=1.16
r41 10 16 0.853661 $w=4.03e-07 $l=3e-08 $layer=LI1_cond $X=1.042 $Y=1.19
+ $X2=1.042 $Y2=1.16
r42 9 25 4.70716 $w=3.53e-07 $l=1.45e-07 $layer=LI1_cond $X=1.067 $Y=0.85
+ $X2=1.067 $Y2=0.995
r43 8 9 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=1.067 $Y=0.51
+ $X2=1.067 $Y2=0.85
r44 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.985
+ $X2=0.89 $Y2=1.325
r45 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.865 $Y=0.56
+ $X2=0.865 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_4%C 3 6 8 9 10 15 17
r36 15 18 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.452 $Y=1.16
+ $X2=1.452 $Y2=1.325
r37 15 17 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.452 $Y=1.16
+ $X2=1.452 $Y2=0.995
r38 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.16 $X2=1.5 $Y2=1.16
r39 10 16 1.2131 $w=2.83e-07 $l=3e-08 $layer=LI1_cond $X=1.557 $Y=1.19 $X2=1.557
+ $Y2=1.16
r40 9 16 12.5353 $w=2.83e-07 $l=3.1e-07 $layer=LI1_cond $X=1.557 $Y=0.85
+ $X2=1.557 $Y2=1.16
r41 8 9 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.557 $Y=0.51
+ $X2=1.557 $Y2=0.85
r42 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.35 $Y=1.985
+ $X2=1.35 $Y2=1.325
r43 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.35 $Y=0.56 $X2=1.35
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_4%D 3 7 8 12 13 14
c43 12 0 1.11144e-19 $X=1.99 $Y=1.16
r44 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.16
+ $X2=1.99 $Y2=1.325
r45 12 14 55.0811 $w=2.7e-07 $l=1.95e-07 $layer=POLY_cond $X=1.99 $Y=1.16
+ $X2=1.99 $Y2=0.965
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.16 $X2=1.99 $Y2=1.16
r47 8 13 11.2615 $w=2.63e-07 $l=2.25e-07 $layer=LI1_cond $X=1.99 $Y=0.935
+ $X2=1.99 $Y2=1.16
r48 7 14 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=1.935 $Y=0.56
+ $X2=1.935 $Y2=0.965
r49 3 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.93 $Y=1.985
+ $X2=1.93 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_4%A_27_47# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 39 42 44 48 50 53 54 59 65 67 68 76
c132 53 0 2.21114e-19 $X=2.33 $Y=1.495
r133 73 74 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.83 $Y=1.16
+ $X2=3.25 $Y2=1.16
r134 63 65 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.26 $Y=0.42
+ $X2=0.585 $Y2=0.42
r135 60 76 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.42 $Y=1.16
+ $X2=3.67 $Y2=1.16
r136 60 74 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=3.42 $Y=1.16
+ $X2=3.25 $Y2=1.16
r137 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.16 $X2=3.42 $Y2=1.16
r138 57 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.74 $Y=1.16 $X2=2.83
+ $Y2=1.16
r139 57 70 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.74 $Y=1.16
+ $X2=2.41 $Y2=1.16
r140 56 59 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.74 $Y=1.19
+ $X2=3.42 $Y2=1.19
r141 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.16 $X2=2.74 $Y2=1.16
r142 54 69 19.2442 $w=2.3e-07 $l=3.6e-07 $layer=LI1_cond $X=2.69 $Y=1.19
+ $X2=2.33 $Y2=1.19
r143 54 56 2.50531 $w=2.28e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=1.19 $X2=2.74
+ $Y2=1.19
r144 52 69 1.89258 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.33 $Y=1.305
+ $X2=2.33 $Y2=1.19
r145 52 53 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.33 $Y=1.305
+ $X2=2.33 $Y2=1.495
r146 51 68 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.645 $Y=1.58
+ $X2=1.55 $Y2=1.58
r147 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.245 $Y=1.58
+ $X2=2.33 $Y2=1.495
r148 50 51 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.245 $Y=1.58
+ $X2=1.645 $Y2=1.58
r149 46 68 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.665
+ $X2=1.55 $Y2=1.58
r150 46 48 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.55 $Y=1.665
+ $X2=1.55 $Y2=1.96
r151 45 67 1.74598 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.765 $Y=1.58
+ $X2=0.632 $Y2=1.58
r152 44 68 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.55 $Y2=1.58
r153 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=0.765 $Y2=1.58
r154 40 67 4.70473 $w=1.9e-07 $l=9.80051e-08 $layer=LI1_cond $X=0.66 $Y=1.665
+ $X2=0.632 $Y2=1.58
r155 40 42 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.66 $Y=1.665
+ $X2=0.66 $Y2=1.96
r156 39 67 4.70473 $w=1.9e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.585 $Y=1.495
+ $X2=0.632 $Y2=1.58
r157 38 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0.585
+ $X2=0.585 $Y2=0.42
r158 38 39 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.585 $Y=0.585
+ $X2=0.585 $Y2=1.495
r159 34 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r160 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.985
r161 31 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=1.16
r162 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=0.56
r163 27 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.325
+ $X2=3.25 $Y2=1.16
r164 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.25 $Y=1.325
+ $X2=3.25 $Y2=1.985
r165 24 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=1.16
r166 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=0.56
r167 20 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.325
+ $X2=2.83 $Y2=1.16
r168 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.83 $Y=1.325
+ $X2=2.83 $Y2=1.985
r169 17 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=0.995
+ $X2=2.83 $Y2=1.16
r170 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.83 $Y=0.995
+ $X2=2.83 $Y2=0.56
r171 13 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.325
+ $X2=2.41 $Y2=1.16
r172 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.41 $Y=1.325
+ $X2=2.41 $Y2=1.985
r173 10 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=0.995
+ $X2=2.41 $Y2=1.16
r174 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.41 $Y=0.995
+ $X2=2.41 $Y2=0.56
r175 3 48 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.425
+ $Y=1.485 $X2=1.56 $Y2=1.96
r176 2 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
r177 1 63 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_4%VPWR 1 2 3 4 5 16 18 22 24 28 30 34 36 38 40
+ 42 47 56 59 62 66
c69 3 0 1.09969e-19 $X=2.005 $Y=1.485
r70 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r72 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r75 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 51 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r77 51 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r78 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r79 48 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=3.08 $Y2=2.72
r80 48 50 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 47 65 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.927 $Y2=2.72
r82 47 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 46 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r84 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r85 43 53 4.29151 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r86 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r87 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=1.12 $Y2=2.72
r88 42 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 40 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 40 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 36 65 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.927 $Y2=2.72
r92 36 38 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2
r93 32 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r94 32 34 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r95 31 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.19 $Y2=2.72
r96 30 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=2.72
+ $X2=3.08 $Y2=2.72
r97 30 31 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.955 $Y=2.72
+ $X2=2.355 $Y2=2.72
r98 26 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r99 26 28 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.02
r100 25 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.12 $Y2=2.72
r101 24 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.19 $Y2=2.72
r102 24 25 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.285 $Y2=2.72
r103 20 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r104 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.02
r105 16 53 3.06854 $w=2.8e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.192 $Y2=2.72
r106 16 18 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2
r107 5 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=2
r108 4 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.905
+ $Y=1.485 $X2=3.04 $Y2=2
r109 3 28 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=2.005
+ $Y=1.485 $X2=2.19 $Y2=2.02
r110 2 22 300 $w=1.7e-07 $l=6.07577e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.12 $Y2=2.02
r111 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_4%X 1 2 3 4 15 17 19 23 24 26 29 33 35 37 38 39
+ 40 41 47 50 57 60
c67 47 0 1.00756e-19 $X=3.925 $Y=0.81
r68 56 57 5.14764 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=1.615
+ $X2=3.375 $Y2=1.615
r69 48 60 0.954516 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=3.925 $Y=1.485
+ $X2=3.925 $Y2=1.615
r70 47 50 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.925 $Y=0.81
+ $X2=3.925 $Y2=0.85
r71 41 60 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.905 $Y=1.615
+ $X2=3.925 $Y2=1.615
r72 41 56 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=3.905 $Y=1.615
+ $X2=3.46 $Y2=1.615
r73 41 48 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=3.925 $Y=1.465
+ $X2=3.925 $Y2=1.485
r74 40 41 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=3.925 $Y=1.19
+ $X2=3.925 $Y2=1.465
r75 39 47 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.725
+ $X2=3.925 $Y2=0.81
r76 39 40 14.6591 $w=2.48e-07 $l=3.18e-07 $layer=LI1_cond $X=3.925 $Y=0.872
+ $X2=3.925 $Y2=1.19
r77 39 50 1.01415 $w=2.48e-07 $l=2.2e-08 $layer=LI1_cond $X=3.925 $Y=0.872
+ $X2=3.925 $Y2=0.85
r78 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.46 $Y2=0.725
r79 35 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.8 $Y=0.725
+ $X2=3.925 $Y2=0.725
r80 35 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.8 $Y=0.725
+ $X2=3.545 $Y2=0.725
r81 31 56 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.46 $Y=1.745
+ $X2=3.46 $Y2=1.615
r82 31 33 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.46 $Y=1.745
+ $X2=3.46 $Y2=1.96
r83 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=0.64 $X2=3.46
+ $Y2=0.725
r84 27 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.46 $Y=0.64
+ $X2=3.46 $Y2=0.42
r85 26 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.785 $Y=1.57
+ $X2=3.375 $Y2=1.57
r86 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=0.725
+ $X2=3.46 $Y2=0.725
r87 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.375 $Y=0.725
+ $X2=2.705 $Y2=0.725
r88 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.7 $Y=1.655
+ $X2=2.785 $Y2=1.57
r89 21 37 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.7 $Y=1.655 $X2=2.7
+ $Y2=1.795
r90 17 37 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.66 $Y=1.92
+ $X2=2.66 $Y2=1.795
r91 17 19 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=2.66 $Y=1.92 $X2=2.66
+ $Y2=1.96
r92 13 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.62 $Y=0.64
+ $X2=2.705 $Y2=0.725
r93 13 15 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.62 $Y=0.64
+ $X2=2.62 $Y2=0.42
r94 4 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=1.485 $X2=3.46 $Y2=1.96
r95 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.485 $X2=2.62 $Y2=1.96
r96 2 29 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.46 $Y2=0.42
r97 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4_4%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
c69 18 0 1.00756e-19 $X=3.88 $Y=0.085
r70 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r71 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r72 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r74 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r75 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r76 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.04
+ $Y2=0
r77 35 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.45
+ $Y2=0
r78 34 46 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.927
+ $Y2=0
r79 34 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.45
+ $Y2=0
r80 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r81 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r82 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r83 30 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.18
+ $Y2=0
r84 30 32 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.53
+ $Y2=0
r85 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=3.04
+ $Y2=0
r86 29 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.53
+ $Y2=0
r87 24 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.18
+ $Y2=0
r88 24 26 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=0.23 $Y2=0
r89 22 41 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r90 22 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r91 18 46 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.927 $Y2=0
r92 18 20 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.88 $Y=0.085 $X2=3.88
+ $Y2=0.385
r93 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0
r94 14 16 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.04 $Y=0.085 $X2=3.04
+ $Y2=0.385
r95 10 40 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r96 10 12 11.1527 $w=3.08e-07 $l=3e-07 $layer=LI1_cond $X=2.18 $Y=0.085 $X2=2.18
+ $Y2=0.385
r97 3 20 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.385
r98 2 16 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.235 $X2=3.04 $Y2=0.385
r99 1 12 182 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.235 $X2=2.19 $Y2=0.385
.ends


* File: sky130_fd_sc_hd__fa_2.spice.SKY130_FD_SC_HD__FA_2.pxi
* Created: Thu Aug 27 14:21:10 2020
* 
x_PM_SKY130_FD_SC_HD__FA_2%A_80_21# N_A_80_21#_M1026_d N_A_80_21#_M1013_d
+ N_A_80_21#_c_185_n N_A_80_21#_M1008_g N_A_80_21#_M1005_g N_A_80_21#_c_186_n
+ N_A_80_21#_M1014_g N_A_80_21#_M1019_g N_A_80_21#_M1027_g N_A_80_21#_M1020_g
+ N_A_80_21#_c_345_p N_A_80_21#_c_189_n N_A_80_21#_c_190_n N_A_80_21#_c_191_n
+ N_A_80_21#_c_355_p N_A_80_21#_c_204_n N_A_80_21#_c_205_n N_A_80_21#_c_231_p
+ N_A_80_21#_c_217_p N_A_80_21#_c_275_p N_A_80_21#_c_291_p N_A_80_21#_c_192_n
+ N_A_80_21#_c_193_n N_A_80_21#_c_194_n N_A_80_21#_c_195_n N_A_80_21#_c_196_n
+ N_A_80_21#_c_197_n N_A_80_21#_c_198_n N_A_80_21#_c_199_n
+ PM_SKY130_FD_SC_HD__FA_2%A_80_21#
x_PM_SKY130_FD_SC_HD__FA_2%A N_A_c_411_n N_A_M1002_g N_A_M1004_g N_A_M1029_g
+ N_A_M1030_g N_A_M1021_g N_A_M1012_g N_A_M1009_g N_A_M1022_g A N_A_c_418_n
+ N_A_c_419_n N_A_c_420_n N_A_c_421_n N_A_c_422_n N_A_c_423_n N_A_c_424_n
+ N_A_c_425_n N_A_c_426_n N_A_c_427_n N_A_c_428_n N_A_c_429_n N_A_c_430_n
+ PM_SKY130_FD_SC_HD__FA_2%A
x_PM_SKY130_FD_SC_HD__FA_2%B N_B_M1013_g N_B_M1026_g N_B_c_678_n N_B_M1028_g
+ N_B_c_687_n N_B_M1023_g N_B_c_679_n N_B_c_680_n N_B_c_688_n N_B_c_689_n
+ N_B_c_681_n N_B_M1017_g N_B_M1024_g N_B_M1006_g N_B_M1010_g N_B_c_683_n B
+ N_B_c_693_n N_B_c_694_n N_B_c_695_n N_B_c_763_n N_B_c_696_n N_B_c_697_n
+ N_B_c_698_n N_B_c_699_n N_B_c_700_n N_B_c_684_n N_B_c_702_n N_B_c_703_n
+ PM_SKY130_FD_SC_HD__FA_2%B
x_PM_SKY130_FD_SC_HD__FA_2%CIN N_CIN_M1025_g N_CIN_M1000_g N_CIN_M1015_g
+ N_CIN_M1016_g N_CIN_M1007_g N_CIN_M1003_g N_CIN_c_912_n N_CIN_c_913_n
+ N_CIN_c_914_n N_CIN_c_927_n N_CIN_c_928_n N_CIN_c_915_n N_CIN_c_916_n
+ N_CIN_c_917_n N_CIN_c_918_n N_CIN_c_931_n N_CIN_c_919_n N_CIN_c_920_n
+ N_CIN_c_933_n N_CIN_c_934_n CIN N_CIN_c_921_n N_CIN_c_936_n N_CIN_c_937_n
+ PM_SKY130_FD_SC_HD__FA_2%CIN
x_PM_SKY130_FD_SC_HD__FA_2%A_1086_47# N_A_1086_47#_M1027_d N_A_1086_47#_M1020_d
+ N_A_1086_47#_c_1138_n N_A_1086_47#_M1018_g N_A_1086_47#_M1001_g
+ N_A_1086_47#_M1011_g N_A_1086_47#_c_1139_n N_A_1086_47#_M1031_g
+ N_A_1086_47#_c_1185_n N_A_1086_47#_c_1151_n N_A_1086_47#_c_1164_n
+ N_A_1086_47#_c_1140_n N_A_1086_47#_c_1141_n N_A_1086_47#_c_1169_n
+ N_A_1086_47#_c_1172_n N_A_1086_47#_c_1142_n N_A_1086_47#_c_1143_n
+ N_A_1086_47#_c_1233_p N_A_1086_47#_c_1155_n N_A_1086_47#_c_1196_n
+ N_A_1086_47#_c_1149_n N_A_1086_47#_c_1144_n N_A_1086_47#_c_1145_n
+ PM_SKY130_FD_SC_HD__FA_2%A_1086_47#
x_PM_SKY130_FD_SC_HD__FA_2%VPWR N_VPWR_M1005_d N_VPWR_M1019_d N_VPWR_M1030_d
+ N_VPWR_M1024_s N_VPWR_M1016_d N_VPWR_M1022_d N_VPWR_M1011_d N_VPWR_c_1283_n
+ N_VPWR_c_1284_n N_VPWR_c_1285_n N_VPWR_c_1286_n N_VPWR_c_1287_n
+ N_VPWR_c_1288_n N_VPWR_c_1289_n N_VPWR_c_1290_n VPWR VPWR N_VPWR_c_1292_n
+ N_VPWR_c_1293_n N_VPWR_c_1294_n N_VPWR_c_1295_n N_VPWR_c_1296_n
+ N_VPWR_c_1297_n N_VPWR_c_1282_n N_VPWR_c_1299_n N_VPWR_c_1300_n
+ N_VPWR_c_1301_n N_VPWR_c_1302_n N_VPWR_c_1303_n N_VPWR_c_1304_n
+ PM_SKY130_FD_SC_HD__FA_2%VPWR
x_PM_SKY130_FD_SC_HD__FA_2%COUT N_COUT_M1008_s N_COUT_M1005_s N_COUT_c_1419_n
+ N_COUT_c_1422_n N_COUT_c_1423_n N_COUT_c_1433_n N_COUT_c_1420_n
+ N_COUT_c_1442_n COUT COUT N_COUT_c_1447_n COUT PM_SKY130_FD_SC_HD__FA_2%COUT
x_PM_SKY130_FD_SC_HD__FA_2%A_473_371# N_A_473_371#_M1000_d N_A_473_371#_M1023_d
+ N_A_473_371#_c_1477_n N_A_473_371#_c_1465_n N_A_473_371#_c_1471_n
+ N_A_473_371#_c_1466_n PM_SKY130_FD_SC_HD__FA_2%A_473_371#
x_PM_SKY130_FD_SC_HD__FA_2%A_829_369# N_A_829_369#_M1024_d N_A_829_369#_M1012_d
+ N_A_829_369#_c_1499_n N_A_829_369#_c_1488_n N_A_829_369#_c_1491_n
+ N_A_829_369#_c_1506_n PM_SKY130_FD_SC_HD__FA_2%A_829_369#
x_PM_SKY130_FD_SC_HD__FA_2%SUM N_SUM_M1018_d N_SUM_M1001_s N_SUM_c_1514_n
+ N_SUM_c_1517_n N_SUM_c_1518_n N_SUM_c_1515_n N_SUM_c_1537_n N_SUM_c_1541_n
+ N_SUM_c_1544_n SUM PM_SKY130_FD_SC_HD__FA_2%SUM
x_PM_SKY130_FD_SC_HD__FA_2%VGND N_VGND_M1008_d N_VGND_M1014_d N_VGND_M1029_d
+ N_VGND_M1017_s N_VGND_M1015_d N_VGND_M1009_d N_VGND_M1031_s N_VGND_c_1565_n
+ N_VGND_c_1566_n N_VGND_c_1567_n N_VGND_c_1568_n N_VGND_c_1569_n
+ N_VGND_c_1570_n N_VGND_c_1571_n N_VGND_c_1572_n N_VGND_c_1573_n VGND VGND
+ N_VGND_c_1575_n N_VGND_c_1576_n N_VGND_c_1577_n N_VGND_c_1578_n
+ N_VGND_c_1579_n N_VGND_c_1580_n N_VGND_c_1581_n N_VGND_c_1582_n
+ N_VGND_c_1583_n N_VGND_c_1584_n N_VGND_c_1585_n PM_SKY130_FD_SC_HD__FA_2%VGND
x_PM_SKY130_FD_SC_HD__FA_2%A_473_47# N_A_473_47#_M1025_d N_A_473_47#_M1028_d
+ N_A_473_47#_c_1740_n N_A_473_47#_c_1715_n N_A_473_47#_c_1716_n
+ N_A_473_47#_c_1732_n PM_SKY130_FD_SC_HD__FA_2%A_473_47#
x_PM_SKY130_FD_SC_HD__FA_2%A_829_47# N_A_829_47#_M1017_d N_A_829_47#_M1021_d
+ N_A_829_47#_c_1773_n N_A_829_47#_c_1750_n N_A_829_47#_c_1751_n
+ N_A_829_47#_c_1770_n PM_SKY130_FD_SC_HD__FA_2%A_829_47#
cc_1 VNB N_A_80_21#_c_185_n 0.0191332f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_186_n 0.0162873f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.995
cc_3 VNB N_A_80_21#_M1027_g 0.0230444f $X=-0.19 $Y=-0.24 $X2=5.355 $Y2=0.445
cc_4 VNB N_A_80_21#_M1020_g 0.00523751f $X=-0.19 $Y=-0.24 $X2=5.355 $Y2=2.165
cc_5 VNB N_A_80_21#_c_189_n 0.00158238f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.075
cc_6 VNB N_A_80_21#_c_190_n 3.11126e-19 $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.43
cc_7 VNB N_A_80_21#_c_191_n 0.00269814f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=0.74
cc_8 VNB N_A_80_21#_c_192_n 9.01538e-19 $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.16
cc_9 VNB N_A_80_21#_c_193_n 0.0123286f $X=-0.19 $Y=-0.24 $X2=5.625 $Y2=0.85
cc_10 VNB N_A_80_21#_c_194_n 0.00176616f $X=-0.19 $Y=-0.24 $X2=2.215 $Y2=0.85
cc_11 VNB N_A_80_21#_c_195_n 0.00665295f $X=-0.19 $Y=-0.24 $X2=2.07 $Y2=0.85
cc_12 VNB N_A_80_21#_c_196_n 0.00132437f $X=-0.19 $Y=-0.24 $X2=5.77 $Y2=0.85
cc_13 VNB N_A_80_21#_c_197_n 0.0320057f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.16
cc_14 VNB N_A_80_21#_c_198_n 0.0252305f $X=-0.19 $Y=-0.24 $X2=5.415 $Y2=1.04
cc_15 VNB N_A_80_21#_c_199_n 0.00649189f $X=-0.19 $Y=-0.24 $X2=5.415 $Y2=1.04
cc_16 VNB N_A_c_411_n 0.0224371f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=0.235
cc_17 VNB N_A_M1004_g 0.0287956f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_18 VNB N_A_M1029_g 0.0299029f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_19 VNB N_A_M1021_g 0.0198556f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.985
cc_20 VNB N_A_M1012_g 0.00424732f $X=-0.19 $Y=-0.24 $X2=5.355 $Y2=0.445
cc_21 VNB N_A_M1009_g 0.0288631f $X=-0.19 $Y=-0.24 $X2=5.355 $Y2=2.165
cc_22 VNB A 0.00864784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_c_418_n 0.0031034f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.075
cc_24 VNB N_A_c_419_n 0.00107886f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.245
cc_25 VNB N_A_c_420_n 0.00614383f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.43
cc_26 VNB N_A_c_421_n 8.64789e-19 $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=0.74
cc_27 VNB N_A_c_422_n 0.00558474f $X=-0.19 $Y=-0.24 $X2=1.075 $Y2=0.74
cc_28 VNB N_A_c_423_n 0.00124236f $X=-0.19 $Y=-0.24 $X2=1.305 $Y2=1.58
cc_29 VNB N_A_c_424_n 0.00253456f $X=-0.19 $Y=-0.24 $X2=2.072 $Y2=2.335
cc_30 VNB N_A_c_425_n 0.00170256f $X=-0.19 $Y=-0.24 $X2=2.072 $Y2=1.995
cc_31 VNB N_A_c_426_n 0.0224949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_c_427_n 0.0244928f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.16
cc_33 VNB N_A_c_428_n 0.00666652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_c_429_n 0.0203718f $X=-0.19 $Y=-0.24 $X2=5.415 $Y2=1.04
cc_35 VNB N_A_c_430_n 0.0122585f $X=-0.19 $Y=-0.24 $X2=5.415 $Y2=1.04
cc_36 VNB N_B_M1026_g 0.0419701f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_37 VNB N_B_c_678_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_38 VNB N_B_c_679_n 0.0530718f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.56
cc_39 VNB N_B_c_680_n 0.00947258f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.56
cc_40 VNB N_B_c_681_n 0.0171497f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.985
cc_41 VNB N_B_M1006_g 0.0415238f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_42 VNB N_B_c_683_n 0.00469281f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.075
cc_43 VNB N_B_c_684_n 0.0213523f $X=-0.19 $Y=-0.24 $X2=5.77 $Y2=0.85
cc_44 VNB N_CIN_M1025_g 0.0283499f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_CIN_M1003_g 0.0416782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_CIN_c_912_n 0.0134432f $X=-0.19 $Y=-0.24 $X2=5.355 $Y2=2.165
cc_47 VNB N_CIN_c_913_n 0.00664345f $X=-0.19 $Y=-0.24 $X2=5.355 $Y2=2.165
cc_48 VNB N_CIN_c_914_n 3.21027e-19 $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_49 VNB N_CIN_c_915_n 0.00215826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_CIN_c_916_n 0.0152367f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.825
cc_51 VNB N_CIN_c_917_n 0.00451859f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.075
cc_52 VNB N_CIN_c_918_n 5.41591e-19 $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.43
cc_53 VNB N_CIN_c_919_n 0.0190028f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.665
cc_54 VNB N_CIN_c_920_n 0.00303344f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.995
cc_55 VNB N_CIN_c_921_n 0.0187439f $X=-0.19 $Y=-0.24 $X2=2.07 $Y2=0.85
cc_56 VNB N_A_1086_47#_c_1138_n 0.017346f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_57 VNB N_A_1086_47#_c_1139_n 0.0202605f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.985
cc_58 VNB N_A_1086_47#_c_1140_n 0.00364909f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_59 VNB N_A_1086_47#_c_1141_n 0.0033791f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_60 VNB N_A_1086_47#_c_1142_n 0.00165814f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.245
cc_61 VNB N_A_1086_47#_c_1143_n 4.74296e-19 $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=0.74
cc_62 VNB N_A_1086_47#_c_1144_n 0.00104403f $X=-0.19 $Y=-0.24 $X2=2.07 $Y2=0.85
cc_63 VNB N_A_1086_47#_c_1145_n 0.0396472f $X=-0.19 $Y=-0.24 $X2=5.77 $Y2=0.85
cc_64 VNB N_VPWR_c_1282_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_COUT_c_1419_n 0.0212177f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_66 VNB N_COUT_c_1420_n 0.0103707f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.325
cc_67 VNB N_SUM_c_1514_n 0.00175733f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.325
cc_68 VNB N_SUM_c_1515_n 0.0105213f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=0.56
cc_69 VNB SUM 0.0202808f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_70 VNB N_VGND_c_1565_n 0.0022431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1566_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1567_n 0.0049662f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_73 VNB N_VGND_c_1568_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.245
cc_74 VNB N_VGND_c_1569_n 0.00280508f $X=-0.19 $Y=-0.24 $X2=1.305 $Y2=1.58
cc_75 VNB N_VGND_c_1570_n 0.0118239f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.665
cc_76 VNB N_VGND_c_1571_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.995
cc_77 VNB N_VGND_c_1572_n 0.0456861f $X=-0.19 $Y=-0.24 $X2=2.072 $Y2=2.335
cc_78 VNB N_VGND_c_1573_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=2.08 $Y2=2.335
cc_79 VNB VGND 0.0108394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1575_n 0.0173899f $X=-0.19 $Y=-0.24 $X2=5.625 $Y2=0.85
cc_81 VNB N_VGND_c_1576_n 0.0332962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1577_n 0.0159136f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.16
cc_83 VNB N_VGND_c_1578_n 0.0116974f $X=-0.19 $Y=-0.24 $X2=5.415 $Y2=0.875
cc_84 VNB N_VGND_c_1579_n 0.0202688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1580_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1581_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1582_n 0.00507318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1583_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1584_n 0.393053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1585_n 0.00417638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_473_47#_c_1715_n 0.00310751f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_92 VNB N_A_473_47#_c_1716_n 0.00259269f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_93 VNB N_A_829_47#_c_1750_n 0.00540238f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_94 VNB N_A_829_47#_c_1751_n 0.00218811f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_95 VPB N_A_80_21#_M1005_g 0.0220043f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_96 VPB N_A_80_21#_M1019_g 0.0184668f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_97 VPB N_A_80_21#_M1020_g 0.0378103f $X=-0.19 $Y=1.305 $X2=5.355 $Y2=2.165
cc_98 VPB N_A_80_21#_c_190_n 0.00216775f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.43
cc_99 VPB N_A_80_21#_c_204_n 0.00288707f $X=-0.19 $Y=1.305 $X2=1.305 $Y2=1.58
cc_100 VPB N_A_80_21#_c_205_n 0.00184251f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.91
cc_101 VPB N_A_80_21#_c_197_n 0.00400826f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.16
cc_102 VPB N_A_c_411_n 0.00442823f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=0.235
cc_103 VPB N_A_M1002_g 0.0367825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_M1030_g 0.0374744f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=0.56
cc_105 VPB N_A_M1012_g 0.0364185f $X=-0.19 $Y=1.305 $X2=5.355 $Y2=0.445
cc_106 VPB N_A_M1022_g 0.0396698f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_107 VPB A 0.00144132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_c_419_n 0.00245924f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.245
cc_109 VPB N_A_c_421_n 2.32744e-19 $X=-0.19 $Y=1.305 $X2=1.535 $Y2=0.74
cc_110 VPB N_A_c_423_n 5.14832e-19 $X=-0.19 $Y=1.305 $X2=1.305 $Y2=1.58
cc_111 VPB N_A_c_424_n 0.00178219f $X=-0.19 $Y=1.305 $X2=2.072 $Y2=2.335
cc_112 VPB N_A_c_425_n 7.64837e-19 $X=-0.19 $Y=1.305 $X2=2.072 $Y2=1.995
cc_113 VPB N_A_c_426_n 0.00700974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_c_429_n 0.00482402f $X=-0.19 $Y=1.305 $X2=5.415 $Y2=1.04
cc_115 VPB N_B_M1013_g 0.0200155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_B_M1026_g 0.0031866f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_117 VPB N_B_c_687_n 0.0199086f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_118 VPB N_B_c_688_n 0.0399721f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.325
cc_119 VPB N_B_c_689_n 0.00881125f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.985
cc_120 VPB N_B_M1006_g 0.00322479f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_121 VPB N_B_M1010_g 0.0205486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB B 0.00696233f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.245
cc_123 VPB N_B_c_693_n 0.00733903f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=0.74
cc_124 VPB N_B_c_694_n 0.0016476f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=0.74
cc_125 VPB N_B_c_695_n 0.0105272f $X=-0.19 $Y=1.305 $X2=1.305 $Y2=1.58
cc_126 VPB N_B_c_696_n 0.00168228f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.16
cc_127 VPB N_B_c_697_n 0.00813082f $X=-0.19 $Y=1.305 $X2=1.007 $Y2=1.58
cc_128 VPB N_B_c_698_n 0.0246507f $X=-0.19 $Y=1.305 $X2=5.625 $Y2=0.85
cc_129 VPB N_B_c_699_n 0.0389846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_B_c_700_n 0.00182223f $X=-0.19 $Y=1.305 $X2=5.77 $Y2=0.85
cc_131 VPB N_B_c_684_n 0.00173871f $X=-0.19 $Y=1.305 $X2=5.77 $Y2=0.85
cc_132 VPB N_B_c_702_n 0.0184685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_B_c_703_n 0.0243326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_CIN_M1000_g 0.0344566f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_135 VPB N_CIN_M1016_g 0.0188895f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=0.995
cc_136 VPB N_CIN_M1007_g 0.0179457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_CIN_M1003_g 0.00271333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_CIN_c_914_n 0.00267764f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_139 VPB N_CIN_c_927_n 0.00934831f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_140 VPB N_CIN_c_928_n 0.00271596f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_141 VPB N_CIN_c_915_n 0.0069689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_CIN_c_918_n 0.00124245f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.43
cc_143 VPB N_CIN_c_931_n 0.0171474f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=0.74
cc_144 VPB N_CIN_c_919_n 0.00639429f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.665
cc_145 VPB N_CIN_c_933_n 0.0233104f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.16
cc_146 VPB N_CIN_c_934_n 0.00366471f $X=-0.19 $Y=1.305 $X2=1.007 $Y2=1.58
cc_147 VPB N_CIN_c_921_n 0.00233543f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=0.85
cc_148 VPB N_CIN_c_936_n 0.0253827f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=0.85
cc_149 VPB N_CIN_c_937_n 0.00644752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_1086_47#_M1001_g 0.0182265f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_151 VPB N_A_1086_47#_M1011_g 0.0221267f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=0.56
cc_152 VPB N_A_1086_47#_c_1143_n 0.00157521f $X=-0.19 $Y=1.305 $X2=1.535
+ $Y2=0.74
cc_153 VPB N_A_1086_47#_c_1149_n 0.00199451f $X=-0.19 $Y=1.305 $X2=5.625
+ $Y2=0.85
cc_154 VPB N_A_1086_47#_c_1145_n 0.00771186f $X=-0.19 $Y=1.305 $X2=5.77 $Y2=0.85
cc_155 VPB N_VPWR_c_1283_n 0.00231272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_1284_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_1285_n 0.00765493f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_158 VPB N_VPWR_c_1286_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.245
cc_159 VPB N_VPWR_c_1287_n 0.0027527f $X=-0.19 $Y=1.305 $X2=1.305 $Y2=1.58
cc_160 VPB N_VPWR_c_1288_n 0.00412306f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.995
cc_161 VPB N_VPWR_c_1289_n 0.0159536f $X=-0.19 $Y=1.305 $X2=2.072 $Y2=2.335
cc_162 VPB N_VPWR_c_1290_n 0.00324402f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=2.335
cc_163 VPB VPWR 0.0111867f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1292_n 0.0180274f $X=-0.19 $Y=1.305 $X2=5.625 $Y2=0.85
cc_165 VPB N_VPWR_c_1293_n 0.0354897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1294_n 0.0153149f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=1.16
cc_167 VPB N_VPWR_c_1295_n 0.0116974f $X=-0.19 $Y=1.305 $X2=5.415 $Y2=0.875
cc_168 VPB N_VPWR_c_1296_n 0.0484432f $X=-0.19 $Y=1.305 $X2=5.415 $Y2=1.04
cc_169 VPB N_VPWR_c_1297_n 0.0115308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1282_n 0.0610372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1299_n 0.0051592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1300_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1301_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1302_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1303_n 0.00510002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1304_n 0.00416482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_COUT_c_1419_n 0.00548844f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_178 VPB N_COUT_c_1422_n 0.00218591f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_179 VPB N_COUT_c_1423_n 0.00963798f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.325
cc_180 VPB N_A_473_371#_c_1465_n 0.00158421f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.325
cc_181 VPB N_A_473_371#_c_1466_n 0.0032459f $X=-0.19 $Y=1.305 $X2=0.475
+ $Y2=1.985
cc_182 VPB N_SUM_c_1517_n 0.0172425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_SUM_c_1518_n 0.00156228f $X=-0.19 $Y=1.305 $X2=0.895 $Y2=0.995
cc_184 VPB SUM 0.00583754f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_185 N_A_80_21#_c_189_n N_A_c_411_n 4.68892e-19 $X=0.99 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_186 N_A_80_21#_c_190_n N_A_c_411_n 4.6773e-19 $X=0.99 $Y=1.43 $X2=-0.19
+ $Y2=-0.24
cc_187 N_A_80_21#_c_191_n N_A_c_411_n 0.0018936f $X=1.535 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_80_21#_c_204_n N_A_c_411_n 0.00189849f $X=1.305 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_80_21#_c_192_n N_A_c_411_n 0.00112398f $X=0.99 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_80_21#_c_197_n N_A_c_411_n 0.0185562f $X=0.895 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_191 N_A_80_21#_M1019_g N_A_M1002_g 0.0343293f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_80_21#_c_190_n N_A_M1002_g 0.00289362f $X=0.99 $Y=1.43 $X2=0 $Y2=0
cc_193 N_A_80_21#_c_204_n N_A_M1002_g 0.00742995f $X=1.305 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A_80_21#_c_205_n N_A_M1002_g 0.00710889f $X=1.39 $Y=1.91 $X2=0 $Y2=0
cc_195 N_A_80_21#_c_217_p N_A_M1002_g 0.00937325f $X=1.475 $Y=1.995 $X2=0 $Y2=0
cc_196 N_A_80_21#_c_186_n N_A_M1004_g 0.0229188f $X=0.895 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_80_21#_c_189_n N_A_M1004_g 0.00329971f $X=0.99 $Y=1.075 $X2=0 $Y2=0
cc_198 N_A_80_21#_c_191_n N_A_M1004_g 0.012185f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_80_21#_c_195_n N_A_M1004_g 0.00857598f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_200 N_A_80_21#_c_193_n N_A_M1029_g 0.00338905f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_201 N_A_80_21#_M1027_g N_A_M1021_g 0.0165256f $X=5.355 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A_80_21#_c_193_n N_A_M1021_g 0.00113591f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_203 N_A_80_21#_c_199_n N_A_M1021_g 7.05654e-19 $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_204 N_A_80_21#_M1020_g N_A_M1012_g 0.044851f $X=5.355 $Y=2.165 $X2=0 $Y2=0
cc_205 N_A_80_21#_c_189_n A 0.00621074f $X=0.99 $Y=1.075 $X2=0 $Y2=0
cc_206 N_A_80_21#_c_190_n A 0.00578614f $X=0.99 $Y=1.43 $X2=0 $Y2=0
cc_207 N_A_80_21#_c_191_n A 0.0211381f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_80_21#_c_204_n A 0.0180302f $X=1.305 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A_80_21#_c_231_p A 0.0027377f $X=1.9 $Y=1.995 $X2=0 $Y2=0
cc_210 N_A_80_21#_c_192_n A 0.0137902f $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_80_21#_c_195_n A 0.0175056f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_212 N_A_80_21#_c_197_n A 3.14871e-19 $X=0.895 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_80_21#_c_193_n N_A_c_418_n 0.0499403f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_214 N_A_80_21#_c_194_n N_A_c_418_n 0.0274258f $X=2.215 $Y=0.85 $X2=0 $Y2=0
cc_215 N_A_80_21#_c_195_n N_A_c_418_n 0.00511587f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_216 N_A_80_21#_c_190_n N_A_c_419_n 2.70135e-19 $X=0.99 $Y=1.43 $X2=0 $Y2=0
cc_217 N_A_80_21#_c_191_n N_A_c_419_n 4.27198e-19 $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A_80_21#_c_231_p N_A_c_419_n 0.00328892f $X=1.9 $Y=1.995 $X2=0 $Y2=0
cc_219 N_A_80_21#_c_192_n N_A_c_419_n 8.4171e-19 $X=0.99 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_80_21#_c_195_n N_A_c_419_n 0.00150462f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_221 N_A_80_21#_c_193_n N_A_c_420_n 0.124008f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_222 N_A_80_21#_c_193_n N_A_c_421_n 0.0266325f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_223 N_A_80_21#_M1020_g N_A_c_422_n 0.00200174f $X=5.355 $Y=2.165 $X2=0 $Y2=0
cc_224 N_A_80_21#_c_193_n N_A_c_422_n 0.0490684f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_225 N_A_80_21#_c_196_n N_A_c_422_n 0.0249445f $X=5.77 $Y=0.85 $X2=0 $Y2=0
cc_226 N_A_80_21#_c_198_n N_A_c_422_n 0.00198965f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_227 N_A_80_21#_c_199_n N_A_c_422_n 0.0168241f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_228 N_A_80_21#_M1020_g N_A_c_423_n 4.24426e-19 $X=5.355 $Y=2.165 $X2=0 $Y2=0
cc_229 N_A_80_21#_c_193_n N_A_c_423_n 0.0261862f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_230 N_A_80_21#_c_199_n N_A_c_423_n 3.07492e-19 $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_231 N_A_80_21#_c_193_n N_A_c_424_n 0.00306165f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_232 N_A_80_21#_c_199_n N_A_c_425_n 0.00133594f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_233 N_A_80_21#_c_193_n N_A_c_426_n 0.00187757f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_234 N_A_80_21#_c_193_n N_A_c_427_n 0.00347599f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_235 N_A_80_21#_c_198_n N_A_c_427_n 0.0196997f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_236 N_A_80_21#_c_199_n N_A_c_427_n 0.00115543f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_237 N_A_80_21#_c_193_n N_A_c_428_n 0.00253419f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_238 N_A_80_21#_c_198_n N_A_c_428_n 0.00311574f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_239 N_A_80_21#_c_199_n N_A_c_428_n 0.014709f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_240 N_A_80_21#_c_199_n N_A_c_430_n 0.0106157f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_241 N_A_80_21#_c_205_n N_B_M1013_g 0.00311481f $X=1.39 $Y=1.91 $X2=0 $Y2=0
cc_242 N_A_80_21#_c_231_p N_B_M1013_g 0.0101713f $X=1.9 $Y=1.995 $X2=0 $Y2=0
cc_243 N_A_80_21#_c_194_n N_B_M1026_g 0.00290518f $X=2.215 $Y=0.85 $X2=0 $Y2=0
cc_244 N_A_80_21#_c_195_n N_B_M1026_g 0.0246037f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_245 N_A_80_21#_c_193_n N_B_c_679_n 0.0124329f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_246 N_A_80_21#_c_193_n N_B_c_680_n 0.00188483f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_247 N_A_80_21#_c_199_n N_B_M1006_g 0.00137141f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_248 N_A_80_21#_c_193_n N_B_c_683_n 0.00336351f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_249 N_A_80_21#_c_190_n B 0.00181899f $X=0.99 $Y=1.43 $X2=0 $Y2=0
cc_250 N_A_80_21#_c_204_n B 0.0147872f $X=1.305 $Y=1.58 $X2=0 $Y2=0
cc_251 N_A_80_21#_c_205_n B 0.00194117f $X=1.39 $Y=1.91 $X2=0 $Y2=0
cc_252 N_A_80_21#_c_231_p B 0.0126623f $X=1.9 $Y=1.995 $X2=0 $Y2=0
cc_253 N_A_80_21#_c_275_p B 0.0140727f $X=2.072 $Y=2.08 $X2=0 $Y2=0
cc_254 N_A_80_21#_c_195_n B 0.0061929f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_255 N_A_80_21#_c_275_p N_B_c_693_n 6.81732e-19 $X=2.072 $Y=2.08 $X2=0 $Y2=0
cc_256 N_A_80_21#_c_204_n N_B_c_694_n 6.71852e-19 $X=1.305 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A_80_21#_c_275_p N_B_c_694_n 0.00362931f $X=2.072 $Y=2.08 $X2=0 $Y2=0
cc_258 N_A_80_21#_M1020_g N_B_c_695_n 0.00173774f $X=5.355 $Y=2.165 $X2=0 $Y2=0
cc_259 N_A_80_21#_c_198_n N_B_c_695_n 5.89663e-19 $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_260 N_A_80_21#_c_199_n N_B_c_695_n 0.00221477f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_261 N_A_80_21#_c_204_n N_B_c_698_n 5.79882e-19 $X=1.305 $Y=1.58 $X2=0 $Y2=0
cc_262 N_A_80_21#_c_231_p N_B_c_698_n 0.00127292f $X=1.9 $Y=1.995 $X2=0 $Y2=0
cc_263 N_A_80_21#_c_195_n N_B_c_698_n 9.62187e-19 $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_264 N_A_80_21#_c_193_n N_B_c_684_n 0.00135025f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_265 N_A_80_21#_c_193_n N_CIN_M1025_g 0.00462124f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_266 N_A_80_21#_c_194_n N_CIN_M1025_g 0.0024037f $X=2.215 $Y=0.85 $X2=0 $Y2=0
cc_267 N_A_80_21#_c_195_n N_CIN_M1025_g 0.00449075f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_268 N_A_80_21#_c_275_p N_CIN_M1000_g 0.00277646f $X=2.072 $Y=2.08 $X2=0 $Y2=0
cc_269 N_A_80_21#_c_291_p N_CIN_M1000_g 0.0042364f $X=2.08 $Y=2.335 $X2=0 $Y2=0
cc_270 N_A_80_21#_M1020_g N_CIN_M1007_g 0.0251353f $X=5.355 $Y=2.165 $X2=0 $Y2=0
cc_271 N_A_80_21#_M1027_g N_CIN_M1003_g 0.0126f $X=5.355 $Y=0.445 $X2=0 $Y2=0
cc_272 N_A_80_21#_M1020_g N_CIN_M1003_g 0.00538209f $X=5.355 $Y=2.165 $X2=0
+ $Y2=0
cc_273 N_A_80_21#_c_196_n N_CIN_M1003_g 0.00134755f $X=5.77 $Y=0.85 $X2=0 $Y2=0
cc_274 N_A_80_21#_c_198_n N_CIN_M1003_g 0.0160461f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_275 N_A_80_21#_c_199_n N_CIN_M1003_g 0.0149352f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_276 N_A_80_21#_c_193_n N_CIN_c_913_n 0.00117521f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_277 N_A_80_21#_c_193_n N_CIN_c_916_n 0.021158f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_278 N_A_80_21#_c_193_n N_CIN_c_917_n 0.00158362f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_279 N_A_80_21#_M1020_g N_CIN_c_931_n 0.0148758f $X=5.355 $Y=2.165 $X2=0 $Y2=0
cc_280 N_A_80_21#_c_198_n N_CIN_c_931_n 0.00169335f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_281 N_A_80_21#_c_199_n N_CIN_c_931_n 0.0114048f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_282 N_A_80_21#_c_275_p N_CIN_c_919_n 8.27068e-19 $X=2.072 $Y=2.08 $X2=0 $Y2=0
cc_283 N_A_80_21#_c_193_n N_CIN_c_919_n 9.52651e-19 $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_284 N_A_80_21#_c_194_n N_CIN_c_919_n 9.74524e-19 $X=2.215 $Y=0.85 $X2=0 $Y2=0
cc_285 N_A_80_21#_c_195_n N_CIN_c_919_n 2.46291e-19 $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_286 N_A_80_21#_c_275_p N_CIN_c_920_n 5.50643e-19 $X=2.072 $Y=2.08 $X2=0 $Y2=0
cc_287 N_A_80_21#_c_193_n N_CIN_c_920_n 0.00500146f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_288 N_A_80_21#_c_194_n N_CIN_c_920_n 0.0013906f $X=2.215 $Y=0.85 $X2=0 $Y2=0
cc_289 N_A_80_21#_c_195_n N_CIN_c_920_n 0.00266523f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_290 N_A_80_21#_c_193_n N_CIN_c_921_n 0.00174757f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_291 N_A_80_21#_M1020_g N_CIN_c_936_n 0.0153265f $X=5.355 $Y=2.165 $X2=0 $Y2=0
cc_292 N_A_80_21#_c_199_n N_CIN_c_936_n 7.33058e-19 $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_293 N_A_80_21#_M1020_g N_CIN_c_937_n 0.00668536f $X=5.355 $Y=2.165 $X2=0
+ $Y2=0
cc_294 N_A_80_21#_c_199_n N_CIN_c_937_n 0.0119833f $X=5.415 $Y=1.04 $X2=0 $Y2=0
cc_295 N_A_80_21#_c_196_n N_A_1086_47#_c_1151_n 0.00212136f $X=5.77 $Y=0.85
+ $X2=0 $Y2=0
cc_296 N_A_80_21#_c_199_n N_A_1086_47#_c_1151_n 0.00815626f $X=5.415 $Y=1.04
+ $X2=0 $Y2=0
cc_297 N_A_80_21#_c_196_n N_A_1086_47#_c_1141_n 0.00161347f $X=5.77 $Y=0.85
+ $X2=0 $Y2=0
cc_298 N_A_80_21#_c_199_n N_A_1086_47#_c_1141_n 0.00199818f $X=5.415 $Y=1.04
+ $X2=0 $Y2=0
cc_299 N_A_80_21#_c_193_n N_A_1086_47#_c_1155_n 4.08874e-19 $X=5.625 $Y=0.85
+ $X2=0 $Y2=0
cc_300 N_A_80_21#_c_196_n N_A_1086_47#_c_1155_n 0.00101125f $X=5.77 $Y=0.85
+ $X2=0 $Y2=0
cc_301 N_A_80_21#_c_199_n N_A_1086_47#_c_1155_n 0.0120345f $X=5.415 $Y=1.04
+ $X2=0 $Y2=0
cc_302 N_A_80_21#_c_190_n N_VPWR_M1019_d 0.00185736f $X=0.99 $Y=1.43 $X2=0 $Y2=0
cc_303 N_A_80_21#_c_204_n N_VPWR_M1019_d 0.00422101f $X=1.305 $Y=1.58 $X2=0
+ $Y2=0
cc_304 N_A_80_21#_M1019_g N_VPWR_c_1283_n 0.00176026f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_305 N_A_80_21#_c_190_n N_VPWR_c_1283_n 0.00271926f $X=0.99 $Y=1.43 $X2=0
+ $Y2=0
cc_306 N_A_80_21#_c_204_n N_VPWR_c_1283_n 0.0050401f $X=1.305 $Y=1.58 $X2=0
+ $Y2=0
cc_307 N_A_80_21#_M1020_g N_VPWR_c_1286_n 0.00114511f $X=5.355 $Y=2.165 $X2=0
+ $Y2=0
cc_308 N_A_80_21#_M1005_g N_VPWR_c_1292_n 0.00585385f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_309 N_A_80_21#_M1019_g N_VPWR_c_1292_n 0.00585385f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_A_80_21#_c_231_p N_VPWR_c_1293_n 0.00646093f $X=1.9 $Y=1.995 $X2=0
+ $Y2=0
cc_311 N_A_80_21#_c_217_p N_VPWR_c_1293_n 0.00265378f $X=1.475 $Y=1.995 $X2=0
+ $Y2=0
cc_312 N_A_80_21#_c_291_p N_VPWR_c_1293_n 0.0201907f $X=2.08 $Y=2.335 $X2=0
+ $Y2=0
cc_313 N_A_80_21#_M1020_g N_VPWR_c_1296_n 0.00585385f $X=5.355 $Y=2.165 $X2=0
+ $Y2=0
cc_314 N_A_80_21#_M1013_d N_VPWR_c_1282_n 0.00261911f $X=1.89 $Y=1.855 $X2=0
+ $Y2=0
cc_315 N_A_80_21#_M1005_g N_VPWR_c_1282_n 0.0114961f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A_80_21#_M1019_g N_VPWR_c_1282_n 0.0105934f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_317 N_A_80_21#_M1020_g N_VPWR_c_1282_n 0.0108663f $X=5.355 $Y=2.165 $X2=0
+ $Y2=0
cc_318 N_A_80_21#_c_231_p N_VPWR_c_1282_n 0.0111822f $X=1.9 $Y=1.995 $X2=0 $Y2=0
cc_319 N_A_80_21#_c_217_p N_VPWR_c_1282_n 0.00425201f $X=1.475 $Y=1.995 $X2=0
+ $Y2=0
cc_320 N_A_80_21#_c_291_p N_VPWR_c_1282_n 0.0129355f $X=2.08 $Y=2.335 $X2=0
+ $Y2=0
cc_321 N_A_80_21#_M1005_g N_VPWR_c_1304_n 0.00311917f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A_80_21#_c_185_n N_COUT_c_1419_n 0.0158983f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_80_21#_c_345_p N_COUT_c_1419_n 0.0136881f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_324 N_A_80_21#_c_189_n N_COUT_c_1419_n 0.0053138f $X=0.99 $Y=1.075 $X2=0
+ $Y2=0
cc_325 N_A_80_21#_c_190_n N_COUT_c_1419_n 0.00529562f $X=0.99 $Y=1.43 $X2=0
+ $Y2=0
cc_326 N_A_80_21#_M1005_g N_COUT_c_1422_n 0.0173022f $X=0.475 $Y=1.985 $X2=0
+ $Y2=0
cc_327 N_A_80_21#_M1019_g N_COUT_c_1422_n 0.00125156f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_328 N_A_80_21#_c_345_p N_COUT_c_1422_n 0.0153741f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_A_80_21#_c_190_n N_COUT_c_1422_n 0.0142073f $X=0.99 $Y=1.43 $X2=0 $Y2=0
cc_330 N_A_80_21#_c_197_n N_COUT_c_1422_n 0.00231083f $X=0.895 $Y=1.16 $X2=0
+ $Y2=0
cc_331 N_A_80_21#_c_185_n N_COUT_c_1433_n 0.00903078f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_A_80_21#_c_186_n N_COUT_c_1433_n 0.00380293f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A_80_21#_c_355_p N_COUT_c_1433_n 0.00524027f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_334 N_A_80_21#_c_185_n N_COUT_c_1420_n 0.0137294f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A_80_21#_c_186_n N_COUT_c_1420_n 0.00124912f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_A_80_21#_c_345_p N_COUT_c_1420_n 0.0106923f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_A_80_21#_c_189_n N_COUT_c_1420_n 0.00515875f $X=0.99 $Y=1.075 $X2=0
+ $Y2=0
cc_338 N_A_80_21#_c_355_p N_COUT_c_1420_n 0.00642327f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_339 N_A_80_21#_c_197_n N_COUT_c_1420_n 0.00123236f $X=0.895 $Y=1.16 $X2=0
+ $Y2=0
cc_340 N_A_80_21#_c_185_n N_COUT_c_1442_n 0.00226964f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A_80_21#_c_186_n N_COUT_c_1442_n 0.00306707f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_342 N_A_80_21#_c_345_p N_COUT_c_1442_n 0.00333874f $X=0.905 $Y=1.16 $X2=0
+ $Y2=0
cc_343 N_A_80_21#_c_197_n N_COUT_c_1442_n 7.11944e-19 $X=0.895 $Y=1.16 $X2=0
+ $Y2=0
cc_344 N_A_80_21#_c_345_p COUT 0.00151726f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A_80_21#_M1019_g N_COUT_c_1447_n 0.00176697f $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_A_80_21#_c_190_n N_COUT_c_1447_n 0.00545866f $X=0.99 $Y=1.43 $X2=0
+ $Y2=0
cc_347 N_A_80_21#_c_205_n N_COUT_c_1447_n 0.00309381f $X=1.39 $Y=1.91 $X2=0
+ $Y2=0
cc_348 N_A_80_21#_c_231_p A_289_371# 0.00634937f $X=1.9 $Y=1.995 $X2=-0.19
+ $Y2=-0.24
cc_349 N_A_80_21#_M1020_g N_A_829_369#_c_1488_n 0.0048174f $X=5.355 $Y=2.165
+ $X2=0 $Y2=0
cc_350 N_A_80_21#_c_189_n N_VGND_M1014_d 7.2386e-19 $X=0.99 $Y=1.075 $X2=0 $Y2=0
cc_351 N_A_80_21#_c_191_n N_VGND_M1014_d 0.00448661f $X=1.535 $Y=0.74 $X2=0
+ $Y2=0
cc_352 N_A_80_21#_c_355_p N_VGND_M1014_d 5.36799e-19 $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_353 N_A_80_21#_c_186_n N_VGND_c_1565_n 0.00285054f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_354 N_A_80_21#_c_191_n N_VGND_c_1565_n 0.016676f $X=1.535 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A_80_21#_c_355_p N_VGND_c_1565_n 0.00368134f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_356 N_A_80_21#_c_195_n N_VGND_c_1565_n 0.0161429f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_357 N_A_80_21#_c_193_n N_VGND_c_1566_n 0.00115864f $X=5.625 $Y=0.85 $X2=0
+ $Y2=0
cc_358 N_A_80_21#_c_193_n N_VGND_c_1567_n 0.00407154f $X=5.625 $Y=0.85 $X2=0
+ $Y2=0
cc_359 N_A_80_21#_M1027_g N_VGND_c_1568_n 0.00114511f $X=5.355 $Y=0.445 $X2=0
+ $Y2=0
cc_360 N_A_80_21#_c_193_n N_VGND_c_1568_n 0.00115864f $X=5.625 $Y=0.85 $X2=0
+ $Y2=0
cc_361 N_A_80_21#_M1027_g N_VGND_c_1572_n 0.00585385f $X=5.355 $Y=0.445 $X2=0
+ $Y2=0
cc_362 N_A_80_21#_c_185_n N_VGND_c_1575_n 0.00425388f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_80_21#_c_186_n N_VGND_c_1575_n 0.00474077f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_364 N_A_80_21#_c_355_p N_VGND_c_1575_n 0.0015722f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_365 N_A_80_21#_c_191_n N_VGND_c_1576_n 0.00299685f $X=1.535 $Y=0.74 $X2=0
+ $Y2=0
cc_366 N_A_80_21#_c_195_n N_VGND_c_1576_n 0.0394373f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_367 N_A_80_21#_M1026_d N_VGND_c_1584_n 0.00208923f $X=1.945 $Y=0.235 $X2=0
+ $Y2=0
cc_368 N_A_80_21#_c_185_n N_VGND_c_1584_n 0.00670042f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A_80_21#_c_186_n N_VGND_c_1584_n 0.00764688f $X=0.895 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_80_21#_M1027_g N_VGND_c_1584_n 0.00673586f $X=5.355 $Y=0.445 $X2=0
+ $Y2=0
cc_371 N_A_80_21#_c_191_n N_VGND_c_1584_n 0.00580564f $X=1.535 $Y=0.74 $X2=0
+ $Y2=0
cc_372 N_A_80_21#_c_355_p N_VGND_c_1584_n 0.00335468f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_373 N_A_80_21#_c_193_n N_VGND_c_1584_n 0.156698f $X=5.625 $Y=0.85 $X2=0 $Y2=0
cc_374 N_A_80_21#_c_194_n N_VGND_c_1584_n 0.0149056f $X=2.215 $Y=0.85 $X2=0
+ $Y2=0
cc_375 N_A_80_21#_c_195_n N_VGND_c_1584_n 0.018502f $X=2.07 $Y=0.85 $X2=0 $Y2=0
cc_376 N_A_80_21#_c_196_n N_VGND_c_1584_n 0.015806f $X=5.77 $Y=0.85 $X2=0 $Y2=0
cc_377 N_A_80_21#_c_199_n N_VGND_c_1584_n 0.00304902f $X=5.415 $Y=1.04 $X2=0
+ $Y2=0
cc_378 N_A_80_21#_c_185_n N_VGND_c_1585_n 0.00316354f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_80_21#_c_195_n A_294_47# 0.00723985f $X=2.07 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_380 N_A_80_21#_c_193_n N_A_473_47#_c_1715_n 0.0271275f $X=5.625 $Y=0.85 $X2=0
+ $Y2=0
cc_381 N_A_80_21#_c_193_n N_A_473_47#_c_1716_n 0.00797006f $X=5.625 $Y=0.85
+ $X2=0 $Y2=0
cc_382 N_A_80_21#_c_194_n N_A_473_47#_c_1716_n 0.00117968f $X=2.215 $Y=0.85
+ $X2=0 $Y2=0
cc_383 N_A_80_21#_c_195_n N_A_473_47#_c_1716_n 0.0081472f $X=2.07 $Y=0.85 $X2=0
+ $Y2=0
cc_384 N_A_80_21#_M1027_g N_A_829_47#_c_1750_n 0.00472067f $X=5.355 $Y=0.445
+ $X2=0 $Y2=0
cc_385 N_A_80_21#_c_193_n N_A_829_47#_c_1750_n 0.0286552f $X=5.625 $Y=0.85 $X2=0
+ $Y2=0
cc_386 N_A_80_21#_c_196_n N_A_829_47#_c_1750_n 0.00140299f $X=5.77 $Y=0.85 $X2=0
+ $Y2=0
cc_387 N_A_80_21#_c_199_n N_A_829_47#_c_1750_n 0.00128307f $X=5.415 $Y=1.04
+ $X2=0 $Y2=0
cc_388 N_A_80_21#_c_193_n N_A_829_47#_c_1751_n 0.00610599f $X=5.625 $Y=0.85
+ $X2=0 $Y2=0
cc_389 N_A_M1002_g N_B_M1013_g 0.0383136f $X=1.37 $Y=2.17 $X2=0 $Y2=0
cc_390 N_A_c_411_n N_B_M1026_g 0.00666585f $X=1.37 $Y=1.325 $X2=0 $Y2=0
cc_391 N_A_M1002_g N_B_M1026_g 0.00161938f $X=1.37 $Y=2.17 $X2=0 $Y2=0
cc_392 N_A_M1004_g N_B_M1026_g 0.0376795f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_393 A N_B_M1026_g 0.00577722f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_394 N_A_c_418_n N_B_M1026_g 0.0049792f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_395 N_A_c_419_n N_B_M1026_g 5.14482e-19 $X=1.755 $Y=1.19 $X2=0 $Y2=0
cc_396 N_A_M1029_g N_B_c_678_n 0.0218633f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_397 N_A_c_420_n N_B_c_680_n 5.6387e-19 $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_398 N_A_c_421_n N_B_c_680_n 3.21623e-19 $X=3.135 $Y=1.19 $X2=0 $Y2=0
cc_399 N_A_c_424_n N_B_c_680_n 4.12248e-19 $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_400 N_A_M1030_g N_B_c_689_n 0.0329021f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_401 N_A_M1009_g N_B_M1006_g 0.043667f $X=6.735 $Y=0.445 $X2=0 $Y2=0
cc_402 N_A_M1022_g N_B_M1006_g 0.00146789f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_403 N_A_c_425_n N_B_M1006_g 8.60102e-19 $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_404 N_A_c_430_n N_B_M1006_g 0.0135237f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_405 N_A_M1022_g N_B_M1010_g 0.0262997f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_406 N_A_M1002_g B 0.00114149f $X=1.37 $Y=2.17 $X2=0 $Y2=0
cc_407 A B 0.00723799f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_408 N_A_c_418_n B 0.00544203f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_409 N_A_c_419_n B 0.00310978f $X=1.755 $Y=1.19 $X2=0 $Y2=0
cc_410 N_A_M1030_g N_B_c_693_n 0.00360106f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_411 N_A_c_418_n N_B_c_693_n 0.0492111f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_412 N_A_c_420_n N_B_c_693_n 0.0518636f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_413 N_A_c_421_n N_B_c_693_n 0.0266263f $X=3.135 $Y=1.19 $X2=0 $Y2=0
cc_414 N_A_c_424_n N_B_c_693_n 0.00287761f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_415 N_A_c_426_n N_B_c_693_n 0.00189048f $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_416 N_A_c_418_n N_B_c_694_n 0.0274262f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_417 N_A_M1012_g N_B_c_695_n 0.00147663f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_418 N_A_c_420_n N_B_c_695_n 0.049641f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_419 N_A_c_422_n N_B_c_695_n 0.0886059f $X=6.085 $Y=1.19 $X2=0 $Y2=0
cc_420 N_A_c_423_n N_B_c_695_n 0.0275415f $X=4.995 $Y=1.19 $X2=0 $Y2=0
cc_421 N_A_c_425_n N_B_c_695_n 0.0266188f $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_422 N_A_c_428_n N_B_c_695_n 0.00168577f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_423 N_A_c_430_n N_B_c_695_n 0.00203106f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_424 N_A_c_420_n N_B_c_763_n 0.0274198f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_425 N_A_M1022_g N_B_c_696_n 0.00308106f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_426 N_A_c_429_n N_B_c_696_n 0.00186167f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A_c_430_n N_B_c_696_n 0.00780453f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_428 N_A_M1022_g N_B_c_697_n 0.0100188f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_429 N_A_c_425_n N_B_c_697_n 0.00127994f $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_430 N_A_c_429_n N_B_c_697_n 0.00165748f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_431 N_A_c_430_n N_B_c_697_n 0.0454517f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_432 N_A_M1002_g N_B_c_698_n 0.0189688f $X=1.37 $Y=2.17 $X2=0 $Y2=0
cc_433 A N_B_c_698_n 0.00201388f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_434 N_A_c_418_n N_B_c_698_n 0.00114706f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_435 N_A_c_419_n N_B_c_698_n 0.00226867f $X=1.755 $Y=1.19 $X2=0 $Y2=0
cc_436 N_A_c_420_n N_B_c_699_n 0.00153932f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_437 N_A_c_420_n N_B_c_700_n 0.00207379f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_438 N_A_c_420_n N_B_c_684_n 0.00138637f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_439 N_A_M1022_g N_B_c_703_n 0.0159725f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_440 N_A_c_425_n N_B_c_703_n 7.30893e-19 $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_441 N_A_c_430_n N_B_c_703_n 0.00296771f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_442 N_A_M1029_g N_CIN_M1025_g 0.0261054f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_443 N_A_c_426_n N_CIN_M1000_g 0.0412791f $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_444 N_A_M1012_g N_CIN_M1016_g 0.0298654f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_445 N_A_c_422_n N_CIN_M1003_g 0.00347129f $X=6.085 $Y=1.19 $X2=0 $Y2=0
cc_446 N_A_c_425_n N_CIN_M1003_g 0.00137964f $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_447 N_A_c_430_n N_CIN_M1003_g 0.0036571f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_448 N_A_M1021_g N_CIN_c_912_n 0.0141455f $X=4.91 $Y=0.445 $X2=0 $Y2=0
cc_449 N_A_M1021_g N_CIN_c_913_n 0.00744646f $X=4.91 $Y=0.445 $X2=0 $Y2=0
cc_450 N_A_c_427_n N_CIN_c_913_n 0.0209378f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_451 N_A_c_418_n N_CIN_c_914_n 6.22985e-19 $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_452 N_A_c_419_n N_CIN_c_914_n 9.00939e-19 $X=1.755 $Y=1.19 $X2=0 $Y2=0
cc_453 N_A_c_424_n N_CIN_c_914_n 0.00575336f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_454 N_A_c_426_n N_CIN_c_914_n 0.00450847f $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_455 N_A_M1030_g N_CIN_c_927_n 0.0111093f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_456 N_A_c_418_n N_CIN_c_927_n 0.00162254f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_457 N_A_c_420_n N_CIN_c_927_n 6.24857e-19 $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_458 N_A_c_421_n N_CIN_c_927_n 5.60263e-19 $X=3.135 $Y=1.19 $X2=0 $Y2=0
cc_459 N_A_c_424_n N_CIN_c_927_n 0.0202345f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_460 N_A_c_426_n N_CIN_c_927_n 0.00255109f $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_461 N_A_M1030_g N_CIN_c_915_n 0.00429073f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_462 N_A_c_420_n N_CIN_c_915_n 0.00318872f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_463 N_A_c_421_n N_CIN_c_915_n 0.00137624f $X=3.135 $Y=1.19 $X2=0 $Y2=0
cc_464 N_A_c_424_n N_CIN_c_915_n 0.00802988f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_465 N_A_c_426_n N_CIN_c_915_n 5.0579e-19 $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_466 N_A_c_420_n N_CIN_c_916_n 0.0373123f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_467 N_A_c_423_n N_CIN_c_916_n 0.00126698f $X=4.995 $Y=1.19 $X2=0 $Y2=0
cc_468 N_A_c_427_n N_CIN_c_916_n 2.96853e-19 $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_469 N_A_c_428_n N_CIN_c_916_n 0.0147988f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_470 N_A_M1029_g N_CIN_c_917_n 0.00195651f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_471 N_A_c_420_n N_CIN_c_917_n 0.00560548f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_472 N_A_c_421_n N_CIN_c_917_n 0.00142282f $X=3.135 $Y=1.19 $X2=0 $Y2=0
cc_473 N_A_c_424_n N_CIN_c_917_n 0.0168914f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_474 N_A_c_426_n N_CIN_c_917_n 0.0010498f $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_475 N_A_M1012_g N_CIN_c_918_n 7.9432e-19 $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_476 N_A_c_420_n N_CIN_c_918_n 0.00235868f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_477 N_A_c_423_n N_CIN_c_918_n 0.00166046f $X=4.995 $Y=1.19 $X2=0 $Y2=0
cc_478 N_A_c_428_n N_CIN_c_918_n 0.00105124f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_479 N_A_M1012_g N_CIN_c_931_n 0.0100247f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_480 N_A_c_420_n N_CIN_c_931_n 3.16966e-19 $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_481 N_A_c_422_n N_CIN_c_931_n 0.00292909f $X=6.085 $Y=1.19 $X2=0 $Y2=0
cc_482 N_A_c_423_n N_CIN_c_931_n 0.00113336f $X=4.995 $Y=1.19 $X2=0 $Y2=0
cc_483 N_A_c_427_n N_CIN_c_931_n 5.94361e-19 $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_484 N_A_c_428_n N_CIN_c_931_n 0.0170478f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_485 N_A_M1029_g N_CIN_c_919_n 0.0215001f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_486 N_A_c_424_n N_CIN_c_919_n 7.99315e-19 $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_487 A N_CIN_c_920_n 0.00559733f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_488 N_A_c_418_n N_CIN_c_920_n 0.0143043f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_489 N_A_c_419_n N_CIN_c_920_n 2.10722e-19 $X=1.755 $Y=1.19 $X2=0 $Y2=0
cc_490 N_A_c_424_n N_CIN_c_920_n 0.0106105f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_491 N_A_c_426_n N_CIN_c_920_n 8.25882e-19 $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_492 N_A_M1012_g N_CIN_c_933_n 0.0213309f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_493 N_A_c_420_n N_CIN_c_933_n 8.79356e-19 $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_494 N_A_M1012_g N_CIN_c_934_n 0.00147223f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_495 N_A_c_420_n N_CIN_c_934_n 0.00232417f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_496 N_A_M1012_g N_CIN_c_921_n 0.00733914f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_497 N_A_c_420_n N_CIN_c_921_n 0.00214774f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_498 N_A_c_423_n N_CIN_c_921_n 0.00137864f $X=4.995 $Y=1.19 $X2=0 $Y2=0
cc_499 N_A_c_428_n N_CIN_c_921_n 0.00203847f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_500 N_A_c_422_n N_CIN_c_937_n 0.00212697f $X=6.085 $Y=1.19 $X2=0 $Y2=0
cc_501 N_A_M1009_g N_A_1086_47#_c_1138_n 0.0239805f $X=6.735 $Y=0.445 $X2=0
+ $Y2=0
cc_502 N_A_M1022_g N_A_1086_47#_M1001_g 0.0316775f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_503 N_A_M1009_g N_A_1086_47#_c_1151_n 0.00349977f $X=6.735 $Y=0.445 $X2=0
+ $Y2=0
cc_504 N_A_c_422_n N_A_1086_47#_c_1151_n 0.00451776f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_505 N_A_c_425_n N_A_1086_47#_c_1151_n 0.00220053f $X=6.23 $Y=1.19 $X2=0 $Y2=0
cc_506 N_A_c_430_n N_A_1086_47#_c_1151_n 0.00641421f $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_507 N_A_M1009_g N_A_1086_47#_c_1164_n 0.00339087f $X=6.735 $Y=0.445 $X2=0
+ $Y2=0
cc_508 N_A_M1009_g N_A_1086_47#_c_1140_n 0.0118677f $X=6.735 $Y=0.445 $X2=0
+ $Y2=0
cc_509 N_A_c_429_n N_A_1086_47#_c_1140_n 0.00292686f $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_510 N_A_c_430_n N_A_1086_47#_c_1140_n 0.0297985f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_511 N_A_c_430_n N_A_1086_47#_c_1141_n 0.0146449f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_512 N_A_M1022_g N_A_1086_47#_c_1169_n 0.011406f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_513 N_A_c_429_n N_A_1086_47#_c_1169_n 7.79054e-19 $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_514 N_A_c_430_n N_A_1086_47#_c_1169_n 0.00240743f $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_515 N_A_M1022_g N_A_1086_47#_c_1172_n 0.00499834f $X=6.795 $Y=2.17 $X2=0
+ $Y2=0
cc_516 N_A_M1009_g N_A_1086_47#_c_1142_n 0.0021234f $X=6.735 $Y=0.445 $X2=0
+ $Y2=0
cc_517 N_A_c_429_n N_A_1086_47#_c_1142_n 2.15792e-19 $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_518 N_A_c_430_n N_A_1086_47#_c_1142_n 0.00663221f $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_519 N_A_M1022_g N_A_1086_47#_c_1143_n 0.00244048f $X=6.795 $Y=2.17 $X2=0
+ $Y2=0
cc_520 N_A_c_429_n N_A_1086_47#_c_1143_n 0.00108479f $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_521 N_A_c_430_n N_A_1086_47#_c_1143_n 0.00241069f $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_522 N_A_M1022_g N_A_1086_47#_c_1149_n 0.00113171f $X=6.795 $Y=2.17 $X2=0
+ $Y2=0
cc_523 N_A_c_429_n N_A_1086_47#_c_1144_n 5.97356e-19 $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_524 N_A_c_430_n N_A_1086_47#_c_1144_n 0.0159055f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_525 N_A_c_429_n N_A_1086_47#_c_1145_n 0.0195751f $X=6.795 $Y=1.16 $X2=0 $Y2=0
cc_526 N_A_c_430_n N_A_1086_47#_c_1145_n 0.00100447f $X=6.795 $Y=1.16 $X2=0
+ $Y2=0
cc_527 N_A_M1002_g N_VPWR_c_1283_n 0.00846964f $X=1.37 $Y=2.17 $X2=0 $Y2=0
cc_528 N_A_M1030_g N_VPWR_c_1284_n 0.00760687f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_529 N_A_M1012_g N_VPWR_c_1286_n 0.00761262f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_530 N_A_M1022_g N_VPWR_c_1287_n 0.00313672f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_531 N_A_M1002_g N_VPWR_c_1293_n 0.00382403f $X=1.37 $Y=2.17 $X2=0 $Y2=0
cc_532 N_A_M1030_g N_VPWR_c_1293_n 0.00337001f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_533 N_A_M1012_g N_VPWR_c_1296_n 0.00337001f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_534 N_A_M1022_g N_VPWR_c_1296_n 0.00422112f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_535 N_A_M1002_g N_VPWR_c_1282_n 0.00451477f $X=1.37 $Y=2.17 $X2=0 $Y2=0
cc_536 N_A_M1030_g N_VPWR_c_1282_n 0.00397658f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_537 N_A_M1012_g N_VPWR_c_1282_n 0.00403935f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_538 N_A_M1022_g N_VPWR_c_1282_n 0.00605013f $X=6.795 $Y=2.17 $X2=0 $Y2=0
cc_539 N_A_M1030_g N_A_473_371#_c_1465_n 0.0100291f $X=2.71 $Y=2.17 $X2=0 $Y2=0
cc_540 N_A_M1012_g N_A_829_369#_c_1488_n 0.0111197f $X=4.91 $Y=2.165 $X2=0 $Y2=0
cc_541 N_A_M1004_g N_VGND_c_1565_n 0.00801931f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_542 N_A_M1029_g N_VGND_c_1566_n 0.00760016f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_543 N_A_M1021_g N_VGND_c_1568_n 0.00760591f $X=4.91 $Y=0.445 $X2=0 $Y2=0
cc_544 N_A_M1009_g N_VGND_c_1569_n 0.00800495f $X=6.735 $Y=0.445 $X2=0 $Y2=0
cc_545 N_A_M1021_g N_VGND_c_1572_n 0.00337001f $X=4.91 $Y=0.445 $X2=0 $Y2=0
cc_546 N_A_M1009_g N_VGND_c_1572_n 0.00341689f $X=6.735 $Y=0.445 $X2=0 $Y2=0
cc_547 N_A_M1004_g N_VGND_c_1576_n 0.00341689f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_548 N_A_M1029_g N_VGND_c_1576_n 0.00337001f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_549 N_A_M1004_g N_VGND_c_1584_n 0.00418888f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_550 N_A_M1029_g N_VGND_c_1584_n 0.00377406f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_551 N_A_M1021_g N_VGND_c_1584_n 0.00383683f $X=4.91 $Y=0.445 $X2=0 $Y2=0
cc_552 N_A_M1009_g N_VGND_c_1584_n 0.00420045f $X=6.735 $Y=0.445 $X2=0 $Y2=0
cc_553 N_A_M1029_g N_A_473_47#_c_1715_n 0.0108136f $X=2.71 $Y=0.445 $X2=0 $Y2=0
cc_554 N_A_c_418_n N_A_473_47#_c_1715_n 0.00108134f $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_555 N_A_c_420_n N_A_473_47#_c_1715_n 0.00161385f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_556 N_A_c_421_n N_A_473_47#_c_1715_n 9.66928e-19 $X=3.135 $Y=1.19 $X2=0 $Y2=0
cc_557 N_A_c_424_n N_A_473_47#_c_1715_n 0.0169746f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_558 N_A_c_426_n N_A_473_47#_c_1715_n 0.00247695f $X=2.77 $Y=1.195 $X2=0 $Y2=0
cc_559 N_A_c_418_n N_A_473_47#_c_1716_n 5.45312e-19 $X=2.845 $Y=1.19 $X2=0 $Y2=0
cc_560 N_A_M1021_g N_A_829_47#_c_1750_n 0.00973522f $X=4.91 $Y=0.445 $X2=0 $Y2=0
cc_561 N_A_c_420_n N_A_829_47#_c_1750_n 0.00124068f $X=4.705 $Y=1.19 $X2=0 $Y2=0
cc_562 N_A_c_422_n N_A_829_47#_c_1750_n 7.16872e-19 $X=6.085 $Y=1.19 $X2=0 $Y2=0
cc_563 N_A_c_423_n N_A_829_47#_c_1750_n 4.03515e-19 $X=4.995 $Y=1.19 $X2=0 $Y2=0
cc_564 N_A_c_427_n N_A_829_47#_c_1750_n 0.00230741f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_565 N_A_c_428_n N_A_829_47#_c_1750_n 0.0230574f $X=4.915 $Y=1.04 $X2=0 $Y2=0
cc_566 N_B_M1026_g N_CIN_M1025_g 0.026095f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_567 N_B_M1013_g N_CIN_M1000_g 0.0123883f $X=1.815 $Y=2.17 $X2=0 $Y2=0
cc_568 N_B_M1026_g N_CIN_M1000_g 0.0165982f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_569 B N_CIN_M1000_g 0.00155132f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_570 N_B_c_693_n N_CIN_M1000_g 0.00426557f $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_571 N_B_c_694_n N_CIN_M1000_g 0.0024037f $X=2.215 $Y=1.53 $X2=0 $Y2=0
cc_572 N_B_c_699_n N_CIN_M1016_g 0.0268107f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_573 N_B_c_700_n N_CIN_M1016_g 3.15588e-19 $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_574 N_B_c_703_n N_CIN_M1007_g 0.0352431f $X=6.315 $Y=1.53 $X2=0 $Y2=0
cc_575 N_B_M1006_g N_CIN_M1003_g 0.0500916f $X=6.255 $Y=0.445 $X2=0 $Y2=0
cc_576 N_B_c_681_n N_CIN_c_912_n 0.00946436f $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_577 N_B_c_683_n N_CIN_c_913_n 0.00946436f $X=4.07 $Y=0.805 $X2=0 $Y2=0
cc_578 N_B_M1026_g N_CIN_c_914_n 8.26522e-19 $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_579 B N_CIN_c_914_n 0.00849277f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_580 N_B_c_693_n N_CIN_c_914_n 0.0085825f $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_581 N_B_c_694_n N_CIN_c_914_n 0.00173655f $X=2.215 $Y=1.53 $X2=0 $Y2=0
cc_582 N_B_c_680_n N_CIN_c_927_n 0.00203699f $X=3.205 $Y=0.805 $X2=0 $Y2=0
cc_583 N_B_c_688_n N_CIN_c_927_n 0.0111006f $X=3.77 $Y=1.695 $X2=0 $Y2=0
cc_584 N_B_c_689_n N_CIN_c_927_n 0.00751562f $X=3.205 $Y=1.695 $X2=0 $Y2=0
cc_585 N_B_c_693_n N_CIN_c_927_n 0.0266023f $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_586 N_B_c_763_n N_CIN_c_927_n 2.72288e-19 $X=4.075 $Y=1.53 $X2=0 $Y2=0
cc_587 N_B_c_699_n N_CIN_c_927_n 2.61162e-19 $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_588 N_B_c_700_n N_CIN_c_927_n 0.0100882f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_589 N_B_M1013_g N_CIN_c_928_n 2.1681e-19 $X=1.815 $Y=2.17 $X2=0 $Y2=0
cc_590 B N_CIN_c_928_n 0.00911713f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_591 N_B_c_693_n N_CIN_c_928_n 0.00591938f $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_592 N_B_c_694_n N_CIN_c_928_n 0.00122285f $X=2.215 $Y=1.53 $X2=0 $Y2=0
cc_593 N_B_c_693_n N_CIN_c_915_n 0.00984268f $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_594 N_B_c_763_n N_CIN_c_915_n 8.96072e-19 $X=4.075 $Y=1.53 $X2=0 $Y2=0
cc_595 N_B_c_699_n N_CIN_c_915_n 0.00315065f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_596 N_B_c_700_n N_CIN_c_915_n 0.00699272f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_597 N_B_c_684_n N_CIN_c_915_n 2.3672e-19 $X=3.957 $Y=1.355 $X2=0 $Y2=0
cc_598 N_B_c_679_n N_CIN_c_916_n 0.0147995f $X=3.995 $Y=0.805 $X2=0 $Y2=0
cc_599 N_B_c_688_n N_CIN_c_916_n 0.0061986f $X=3.77 $Y=1.695 $X2=0 $Y2=0
cc_600 N_B_c_693_n N_CIN_c_916_n 0.00184237f $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_601 N_B_c_695_n N_CIN_c_916_n 0.00209743f $X=6.545 $Y=1.53 $X2=0 $Y2=0
cc_602 N_B_c_763_n N_CIN_c_916_n 0.00103879f $X=4.075 $Y=1.53 $X2=0 $Y2=0
cc_603 N_B_c_699_n N_CIN_c_916_n 0.00231696f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_604 N_B_c_700_n N_CIN_c_916_n 0.0258113f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_605 N_B_c_684_n N_CIN_c_916_n 0.0188183f $X=3.957 $Y=1.355 $X2=0 $Y2=0
cc_606 N_B_c_679_n N_CIN_c_917_n 0.00347447f $X=3.995 $Y=0.805 $X2=0 $Y2=0
cc_607 N_B_c_695_n N_CIN_c_918_n 4.57159e-19 $X=6.545 $Y=1.53 $X2=0 $Y2=0
cc_608 N_B_c_763_n N_CIN_c_918_n 8.51268e-19 $X=4.075 $Y=1.53 $X2=0 $Y2=0
cc_609 N_B_c_684_n N_CIN_c_918_n 0.00397174f $X=3.957 $Y=1.355 $X2=0 $Y2=0
cc_610 N_B_c_695_n N_CIN_c_931_n 0.0425084f $X=6.545 $Y=1.53 $X2=0 $Y2=0
cc_611 N_B_M1026_g N_CIN_c_919_n 0.0214103f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_612 N_B_c_694_n N_CIN_c_919_n 9.74524e-19 $X=2.215 $Y=1.53 $X2=0 $Y2=0
cc_613 N_B_M1026_g N_CIN_c_920_n 0.0010142f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_614 B N_CIN_c_920_n 0.00197411f $X=1.985 $Y=1.445 $X2=0 $Y2=0
cc_615 N_B_c_693_n N_CIN_c_920_n 0.00216801f $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_616 N_B_c_694_n N_CIN_c_920_n 8.46704e-19 $X=2.215 $Y=1.53 $X2=0 $Y2=0
cc_617 N_B_c_699_n N_CIN_c_933_n 0.0216836f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_618 N_B_c_700_n N_CIN_c_933_n 3.87164e-19 $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_619 N_B_c_695_n N_CIN_c_934_n 0.0164483f $X=6.545 $Y=1.53 $X2=0 $Y2=0
cc_620 N_B_c_763_n N_CIN_c_934_n 0.00171886f $X=4.075 $Y=1.53 $X2=0 $Y2=0
cc_621 N_B_c_699_n N_CIN_c_934_n 0.00153667f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_622 N_B_c_700_n N_CIN_c_934_n 0.0135944f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_623 N_B_c_684_n N_CIN_c_921_n 0.0225963f $X=3.957 $Y=1.355 $X2=0 $Y2=0
cc_624 N_B_c_695_n N_CIN_c_936_n 0.00175799f $X=6.545 $Y=1.53 $X2=0 $Y2=0
cc_625 N_B_c_697_n N_CIN_c_936_n 0.00134146f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_626 N_B_c_703_n N_CIN_c_936_n 0.0500916f $X=6.315 $Y=1.53 $X2=0 $Y2=0
cc_627 N_B_M1006_g N_CIN_c_937_n 5.62374e-19 $X=6.255 $Y=0.445 $X2=0 $Y2=0
cc_628 N_B_M1010_g N_CIN_c_937_n 0.00428927f $X=6.255 $Y=2.17 $X2=0 $Y2=0
cc_629 N_B_c_695_n N_CIN_c_937_n 0.0141879f $X=6.545 $Y=1.53 $X2=0 $Y2=0
cc_630 N_B_c_697_n N_CIN_c_937_n 0.017102f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_631 N_B_c_703_n N_CIN_c_937_n 5.23813e-19 $X=6.315 $Y=1.53 $X2=0 $Y2=0
cc_632 N_B_c_697_n N_A_1086_47#_M1001_g 3.1636e-19 $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_633 N_B_M1010_g N_A_1086_47#_c_1185_n 0.0173719f $X=6.255 $Y=2.17 $X2=0 $Y2=0
cc_634 N_B_c_695_n N_A_1086_47#_c_1185_n 0.0120753f $X=6.545 $Y=1.53 $X2=0 $Y2=0
cc_635 N_B_c_697_n N_A_1086_47#_c_1185_n 0.011759f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_636 N_B_c_703_n N_A_1086_47#_c_1185_n 5.22774e-19 $X=6.315 $Y=1.53 $X2=0
+ $Y2=0
cc_637 N_B_M1006_g N_A_1086_47#_c_1151_n 0.0132015f $X=6.255 $Y=0.445 $X2=0
+ $Y2=0
cc_638 N_B_M1006_g N_A_1086_47#_c_1141_n 0.00438384f $X=6.255 $Y=0.445 $X2=0
+ $Y2=0
cc_639 N_B_c_696_n N_A_1086_47#_c_1169_n 8.48123e-19 $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_640 N_B_c_697_n N_A_1086_47#_c_1169_n 0.00776504f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_641 N_B_c_697_n N_A_1086_47#_c_1172_n 0.0071466f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_642 N_B_c_696_n N_A_1086_47#_c_1143_n 0.00138572f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_643 N_B_c_697_n N_A_1086_47#_c_1143_n 8.41183e-19 $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_644 N_B_M1010_g N_A_1086_47#_c_1196_n 0.00429324f $X=6.255 $Y=2.17 $X2=0
+ $Y2=0
cc_645 N_B_c_696_n N_A_1086_47#_c_1196_n 9.31973e-19 $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_646 N_B_c_697_n N_A_1086_47#_c_1196_n 0.0107388f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_647 N_B_c_696_n N_A_1086_47#_c_1149_n 0.00128946f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_648 N_B_c_697_n N_A_1086_47#_c_1149_n 0.0106926f $X=6.69 $Y=1.53 $X2=0 $Y2=0
cc_649 N_B_M1013_g N_VPWR_c_1283_n 0.00163718f $X=1.815 $Y=2.17 $X2=0 $Y2=0
cc_650 N_B_c_687_n N_VPWR_c_1284_n 0.00677587f $X=3.13 $Y=1.77 $X2=0 $Y2=0
cc_651 N_B_c_687_n N_VPWR_c_1285_n 0.00321545f $X=3.13 $Y=1.77 $X2=0 $Y2=0
cc_652 N_B_c_688_n N_VPWR_c_1285_n 0.00489764f $X=3.77 $Y=1.695 $X2=0 $Y2=0
cc_653 N_B_c_693_n N_VPWR_c_1285_n 5.45078e-19 $X=3.785 $Y=1.53 $X2=0 $Y2=0
cc_654 N_B_c_763_n N_VPWR_c_1285_n 0.00157163f $X=4.075 $Y=1.53 $X2=0 $Y2=0
cc_655 N_B_c_700_n N_VPWR_c_1285_n 0.0225991f $X=3.905 $Y=1.52 $X2=0 $Y2=0
cc_656 N_B_c_702_n N_VPWR_c_1285_n 0.0114275f $X=3.957 $Y=1.77 $X2=0 $Y2=0
cc_657 N_B_c_702_n N_VPWR_c_1286_n 5.31689e-19 $X=3.957 $Y=1.77 $X2=0 $Y2=0
cc_658 N_B_M1013_g N_VPWR_c_1293_n 0.00425831f $X=1.815 $Y=2.17 $X2=0 $Y2=0
cc_659 N_B_c_687_n N_VPWR_c_1294_n 0.00337001f $X=3.13 $Y=1.77 $X2=0 $Y2=0
cc_660 N_B_c_702_n N_VPWR_c_1295_n 0.0046653f $X=3.957 $Y=1.77 $X2=0 $Y2=0
cc_661 N_B_M1010_g N_VPWR_c_1296_n 0.00357877f $X=6.255 $Y=2.17 $X2=0 $Y2=0
cc_662 N_B_M1013_g N_VPWR_c_1282_n 0.00609368f $X=1.815 $Y=2.17 $X2=0 $Y2=0
cc_663 N_B_c_687_n N_VPWR_c_1282_n 0.0053254f $X=3.13 $Y=1.77 $X2=0 $Y2=0
cc_664 N_B_M1010_g N_VPWR_c_1282_n 0.00573192f $X=6.255 $Y=2.17 $X2=0 $Y2=0
cc_665 N_B_c_702_n N_VPWR_c_1282_n 0.00799591f $X=3.957 $Y=1.77 $X2=0 $Y2=0
cc_666 N_B_c_687_n N_A_473_371#_c_1465_n 0.0107429f $X=3.13 $Y=1.77 $X2=0 $Y2=0
cc_667 N_B_c_688_n N_A_473_371#_c_1465_n 0.00540826f $X=3.77 $Y=1.695 $X2=0
+ $Y2=0
cc_668 N_B_c_693_n N_A_473_371#_c_1465_n 0.00782028f $X=3.785 $Y=1.53 $X2=0
+ $Y2=0
cc_669 N_B_c_693_n N_A_473_371#_c_1471_n 0.00104195f $X=3.785 $Y=1.53 $X2=0
+ $Y2=0
cc_670 N_B_c_695_n N_A_829_369#_c_1488_n 0.00513411f $X=6.545 $Y=1.53 $X2=0
+ $Y2=0
cc_671 N_B_c_695_n N_A_829_369#_c_1491_n 0.00484515f $X=6.545 $Y=1.53 $X2=0
+ $Y2=0
cc_672 N_B_M1026_g N_VGND_c_1565_n 0.00121824f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_673 N_B_c_678_n N_VGND_c_1566_n 0.00676915f $X=3.13 $Y=0.73 $X2=0 $Y2=0
cc_674 N_B_c_678_n N_VGND_c_1567_n 0.00208038f $X=3.13 $Y=0.73 $X2=0 $Y2=0
cc_675 N_B_c_679_n N_VGND_c_1567_n 0.0045972f $X=3.995 $Y=0.805 $X2=0 $Y2=0
cc_676 N_B_c_681_n N_VGND_c_1567_n 0.00827538f $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_677 N_B_c_681_n N_VGND_c_1568_n 5.31689e-19 $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_678 N_B_M1006_g N_VGND_c_1569_n 0.00120942f $X=6.255 $Y=0.445 $X2=0 $Y2=0
cc_679 N_B_M1006_g N_VGND_c_1572_n 0.00357877f $X=6.255 $Y=0.445 $X2=0 $Y2=0
cc_680 N_B_M1026_g N_VGND_c_1576_n 0.00357668f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_681 N_B_c_678_n N_VGND_c_1577_n 0.00337001f $X=3.13 $Y=0.73 $X2=0 $Y2=0
cc_682 N_B_c_679_n N_VGND_c_1577_n 0.00469312f $X=3.995 $Y=0.805 $X2=0 $Y2=0
cc_683 N_B_c_681_n N_VGND_c_1578_n 0.0046653f $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_684 N_B_M1026_g N_VGND_c_1584_n 0.00544133f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_685 N_B_c_678_n N_VGND_c_1584_n 0.00512288f $X=3.13 $Y=0.73 $X2=0 $Y2=0
cc_686 N_B_c_679_n N_VGND_c_1584_n 0.00336079f $X=3.995 $Y=0.805 $X2=0 $Y2=0
cc_687 N_B_c_681_n N_VGND_c_1584_n 0.00446764f $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_688 N_B_M1006_g N_VGND_c_1584_n 0.00530375f $X=6.255 $Y=0.445 $X2=0 $Y2=0
cc_689 N_B_c_678_n N_A_473_47#_c_1715_n 0.00758462f $X=3.13 $Y=0.73 $X2=0 $Y2=0
cc_690 N_B_c_679_n N_A_473_47#_c_1715_n 0.00812182f $X=3.995 $Y=0.805 $X2=0
+ $Y2=0
cc_691 N_B_c_680_n N_A_473_47#_c_1715_n 0.00392189f $X=3.205 $Y=0.805 $X2=0
+ $Y2=0
cc_692 N_B_c_681_n N_A_473_47#_c_1715_n 0.00310565f $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_693 N_B_c_681_n N_A_473_47#_c_1732_n 0.00158481f $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_694 N_B_c_681_n N_A_829_47#_c_1751_n 0.00420459f $X=4.07 $Y=0.73 $X2=0 $Y2=0
cc_695 N_CIN_M1007_g N_A_1086_47#_c_1185_n 0.0125611f $X=5.78 $Y=2.165 $X2=0
+ $Y2=0
cc_696 N_CIN_c_931_n N_A_1086_47#_c_1185_n 0.0057196f $X=5.67 $Y=1.6 $X2=0 $Y2=0
cc_697 N_CIN_c_936_n N_A_1086_47#_c_1185_n 0.00187747f $X=5.835 $Y=1.52 $X2=0
+ $Y2=0
cc_698 N_CIN_c_937_n N_A_1086_47#_c_1185_n 0.011642f $X=5.835 $Y=1.52 $X2=0
+ $Y2=0
cc_699 N_CIN_M1003_g N_A_1086_47#_c_1151_n 0.00979993f $X=5.895 $Y=0.445 $X2=0
+ $Y2=0
cc_700 N_CIN_c_937_n N_A_1086_47#_c_1196_n 5.83799e-19 $X=5.835 $Y=1.52 $X2=0
+ $Y2=0
cc_701 N_CIN_M1000_g N_VPWR_c_1284_n 0.00119528f $X=2.29 $Y=2.17 $X2=0 $Y2=0
cc_702 N_CIN_M1016_g N_VPWR_c_1285_n 7.98505e-19 $X=4.49 $Y=2.165 $X2=0 $Y2=0
cc_703 N_CIN_M1016_g N_VPWR_c_1286_n 0.00640108f $X=4.49 $Y=2.165 $X2=0 $Y2=0
cc_704 N_CIN_M1000_g N_VPWR_c_1293_n 0.00541359f $X=2.29 $Y=2.17 $X2=0 $Y2=0
cc_705 N_CIN_M1016_g N_VPWR_c_1295_n 0.00337001f $X=4.49 $Y=2.165 $X2=0 $Y2=0
cc_706 N_CIN_M1007_g N_VPWR_c_1296_n 0.00357877f $X=5.78 $Y=2.165 $X2=0 $Y2=0
cc_707 N_CIN_M1000_g N_VPWR_c_1282_n 0.00988509f $X=2.29 $Y=2.17 $X2=0 $Y2=0
cc_708 N_CIN_M1016_g N_VPWR_c_1282_n 0.00397658f $X=4.49 $Y=2.165 $X2=0 $Y2=0
cc_709 N_CIN_M1007_g N_VPWR_c_1282_n 0.00542737f $X=5.78 $Y=2.165 $X2=0 $Y2=0
cc_710 N_CIN_c_927_n N_A_473_371#_c_1465_n 0.0442431f $X=3.245 $Y=1.655 $X2=0
+ $Y2=0
cc_711 N_CIN_c_927_n N_A_473_371#_c_1471_n 0.00577586f $X=3.245 $Y=1.655 $X2=0
+ $Y2=0
cc_712 N_CIN_c_928_n N_A_473_371#_c_1471_n 0.00557804f $X=2.495 $Y=1.655 $X2=0
+ $Y2=0
cc_713 N_CIN_M1016_g N_A_829_369#_c_1488_n 0.0110354f $X=4.49 $Y=2.165 $X2=0
+ $Y2=0
cc_714 N_CIN_c_931_n N_A_829_369#_c_1488_n 0.00893804f $X=5.67 $Y=1.6 $X2=0
+ $Y2=0
cc_715 N_CIN_c_933_n N_A_829_369#_c_1488_n 0.00113985f $X=4.49 $Y=1.52 $X2=0
+ $Y2=0
cc_716 N_CIN_c_934_n N_A_829_369#_c_1488_n 0.02703f $X=4.655 $Y=1.56 $X2=0 $Y2=0
cc_717 N_CIN_c_934_n N_A_829_369#_c_1491_n 0.00362847f $X=4.655 $Y=1.56 $X2=0
+ $Y2=0
cc_718 N_CIN_c_937_n A_1171_369# 0.00154519f $X=5.835 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_719 N_CIN_M1025_g N_VGND_c_1566_n 0.00118455f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_720 N_CIN_c_912_n N_VGND_c_1567_n 5.44952e-19 $X=4.492 $Y=0.73 $X2=0 $Y2=0
cc_721 N_CIN_c_916_n N_VGND_c_1567_n 0.00546777f $X=4.295 $Y=1.107 $X2=0 $Y2=0
cc_722 N_CIN_c_912_n N_VGND_c_1568_n 0.00639437f $X=4.492 $Y=0.73 $X2=0 $Y2=0
cc_723 N_CIN_M1003_g N_VGND_c_1572_n 0.00357877f $X=5.895 $Y=0.445 $X2=0 $Y2=0
cc_724 N_CIN_M1025_g N_VGND_c_1576_n 0.00585385f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_725 N_CIN_c_912_n N_VGND_c_1578_n 0.00337001f $X=4.492 $Y=0.73 $X2=0 $Y2=0
cc_726 N_CIN_M1025_g N_VGND_c_1584_n 0.00649423f $X=2.29 $Y=0.445 $X2=0 $Y2=0
cc_727 N_CIN_M1003_g N_VGND_c_1584_n 0.00532102f $X=5.895 $Y=0.445 $X2=0 $Y2=0
cc_728 N_CIN_c_912_n N_VGND_c_1584_n 0.00377406f $X=4.492 $Y=0.73 $X2=0 $Y2=0
cc_729 N_CIN_c_916_n N_A_473_47#_c_1715_n 5.77639e-19 $X=4.295 $Y=1.107 $X2=0
+ $Y2=0
cc_730 N_CIN_c_917_n N_A_473_47#_c_1715_n 0.0110711f $X=3.415 $Y=1.107 $X2=0
+ $Y2=0
cc_731 N_CIN_M1025_g N_A_473_47#_c_1716_n 0.00129924f $X=2.29 $Y=0.445 $X2=0
+ $Y2=0
cc_732 N_CIN_c_919_n N_A_473_47#_c_1716_n 2.17239e-19 $X=2.29 $Y=1.19 $X2=0
+ $Y2=0
cc_733 N_CIN_c_920_n N_A_473_47#_c_1716_n 0.00270907f $X=2.41 $Y=1.19 $X2=0
+ $Y2=0
cc_734 N_CIN_c_912_n N_A_829_47#_c_1750_n 0.00669222f $X=4.492 $Y=0.73 $X2=0
+ $Y2=0
cc_735 N_CIN_c_913_n N_A_829_47#_c_1750_n 0.00441497f $X=4.492 $Y=0.88 $X2=0
+ $Y2=0
cc_736 N_CIN_c_916_n N_A_829_47#_c_1750_n 0.00624534f $X=4.295 $Y=1.107 $X2=0
+ $Y2=0
cc_737 N_CIN_c_933_n N_A_829_47#_c_1750_n 9.85703e-19 $X=4.49 $Y=1.52 $X2=0
+ $Y2=0
cc_738 N_CIN_c_934_n N_A_829_47#_c_1750_n 0.00195538f $X=4.655 $Y=1.56 $X2=0
+ $Y2=0
cc_739 N_CIN_c_916_n N_A_829_47#_c_1751_n 0.0111405f $X=4.295 $Y=1.107 $X2=0
+ $Y2=0
cc_740 N_A_1086_47#_c_1169_n N_VPWR_M1022_d 0.00544362f $X=7.01 $Y=2.02 $X2=0
+ $Y2=0
cc_741 N_A_1086_47#_c_1172_n N_VPWR_M1022_d 0.00399486f $X=7.095 $Y=1.935 $X2=0
+ $Y2=0
cc_742 N_A_1086_47#_c_1149_n N_VPWR_M1022_d 0.001562f $X=7.215 $Y=1.555 $X2=0
+ $Y2=0
cc_743 N_A_1086_47#_M1001_g N_VPWR_c_1287_n 0.00671141f $X=7.27 $Y=1.985 $X2=0
+ $Y2=0
cc_744 N_A_1086_47#_M1011_g N_VPWR_c_1287_n 5.32661e-19 $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_745 N_A_1086_47#_c_1169_n N_VPWR_c_1287_n 0.0166961f $X=7.01 $Y=2.02 $X2=0
+ $Y2=0
cc_746 N_A_1086_47#_c_1149_n N_VPWR_c_1287_n 5.96676e-19 $X=7.215 $Y=1.555 $X2=0
+ $Y2=0
cc_747 N_A_1086_47#_M1011_g N_VPWR_c_1288_n 0.00307904f $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_748 N_A_1086_47#_M1001_g N_VPWR_c_1289_n 0.00486043f $X=7.27 $Y=1.985 $X2=0
+ $Y2=0
cc_749 N_A_1086_47#_M1011_g N_VPWR_c_1289_n 0.00557614f $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_750 N_A_1086_47#_c_1185_n N_VPWR_c_1296_n 0.0606537f $X=6.515 $Y=2.295 $X2=0
+ $Y2=0
cc_751 N_A_1086_47#_c_1169_n N_VPWR_c_1296_n 0.00312966f $X=7.01 $Y=2.02 $X2=0
+ $Y2=0
cc_752 N_A_1086_47#_c_1196_n N_VPWR_c_1296_n 0.0108964f $X=6.6 $Y=2.02 $X2=0
+ $Y2=0
cc_753 N_A_1086_47#_M1020_d N_VPWR_c_1282_n 0.00406702f $X=5.43 $Y=1.845 $X2=0
+ $Y2=0
cc_754 N_A_1086_47#_M1001_g N_VPWR_c_1282_n 0.00819893f $X=7.27 $Y=1.985 $X2=0
+ $Y2=0
cc_755 N_A_1086_47#_M1011_g N_VPWR_c_1282_n 0.0107219f $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_756 N_A_1086_47#_c_1185_n N_VPWR_c_1282_n 0.0375122f $X=6.515 $Y=2.295 $X2=0
+ $Y2=0
cc_757 N_A_1086_47#_c_1169_n N_VPWR_c_1282_n 0.00650684f $X=7.01 $Y=2.02 $X2=0
+ $Y2=0
cc_758 N_A_1086_47#_c_1196_n N_VPWR_c_1282_n 0.00642843f $X=6.6 $Y=2.02 $X2=0
+ $Y2=0
cc_759 N_A_1086_47#_c_1185_n A_1171_369# 0.00563231f $X=6.515 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_760 N_A_1086_47#_c_1185_n A_1266_371# 0.00398461f $X=6.515 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_761 N_A_1086_47#_c_1196_n A_1266_371# 0.0080653f $X=6.6 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_762 N_A_1086_47#_c_1138_n N_SUM_c_1514_n 0.00580287f $X=7.23 $Y=0.995 $X2=0
+ $Y2=0
cc_763 N_A_1086_47#_c_1139_n N_SUM_c_1514_n 0.00913962f $X=7.77 $Y=0.995 $X2=0
+ $Y2=0
cc_764 N_A_1086_47#_c_1140_n N_SUM_c_1514_n 0.0140032f $X=7.13 $Y=0.74 $X2=0
+ $Y2=0
cc_765 N_A_1086_47#_c_1142_n N_SUM_c_1514_n 0.00620674f $X=7.215 $Y=1.075 $X2=0
+ $Y2=0
cc_766 N_A_1086_47#_c_1233_p N_SUM_c_1514_n 0.0199585f $X=7.635 $Y=1.16 $X2=0
+ $Y2=0
cc_767 N_A_1086_47#_c_1145_n N_SUM_c_1514_n 0.00367134f $X=7.77 $Y=1.16 $X2=0
+ $Y2=0
cc_768 N_A_1086_47#_M1011_g N_SUM_c_1517_n 0.0124427f $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_769 N_A_1086_47#_c_1233_p N_SUM_c_1517_n 0.0106028f $X=7.635 $Y=1.16 $X2=0
+ $Y2=0
cc_770 N_A_1086_47#_c_1145_n N_SUM_c_1517_n 0.0025007f $X=7.77 $Y=1.16 $X2=0
+ $Y2=0
cc_771 N_A_1086_47#_M1001_g N_SUM_c_1518_n 0.0011776f $X=7.27 $Y=1.985 $X2=0
+ $Y2=0
cc_772 N_A_1086_47#_M1011_g N_SUM_c_1518_n 0.00206908f $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_773 N_A_1086_47#_c_1143_n N_SUM_c_1518_n 0.00436337f $X=7.215 $Y=1.47 $X2=0
+ $Y2=0
cc_774 N_A_1086_47#_c_1233_p N_SUM_c_1518_n 0.0134703f $X=7.635 $Y=1.16 $X2=0
+ $Y2=0
cc_775 N_A_1086_47#_c_1149_n N_SUM_c_1518_n 0.00923521f $X=7.215 $Y=1.555 $X2=0
+ $Y2=0
cc_776 N_A_1086_47#_c_1145_n N_SUM_c_1518_n 0.0012838f $X=7.77 $Y=1.16 $X2=0
+ $Y2=0
cc_777 N_A_1086_47#_c_1139_n N_SUM_c_1515_n 0.0104354f $X=7.77 $Y=0.995 $X2=0
+ $Y2=0
cc_778 N_A_1086_47#_c_1233_p N_SUM_c_1515_n 0.00504964f $X=7.635 $Y=1.16 $X2=0
+ $Y2=0
cc_779 N_A_1086_47#_c_1138_n N_SUM_c_1537_n 0.00299067f $X=7.23 $Y=0.995 $X2=0
+ $Y2=0
cc_780 N_A_1086_47#_c_1139_n N_SUM_c_1537_n 0.00276871f $X=7.77 $Y=0.995 $X2=0
+ $Y2=0
cc_781 N_A_1086_47#_c_1233_p N_SUM_c_1537_n 0.00214742f $X=7.635 $Y=1.16 $X2=0
+ $Y2=0
cc_782 N_A_1086_47#_c_1145_n N_SUM_c_1537_n 0.00153202f $X=7.77 $Y=1.16 $X2=0
+ $Y2=0
cc_783 N_A_1086_47#_M1011_g N_SUM_c_1541_n 0.00259906f $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_784 N_A_1086_47#_c_1233_p N_SUM_c_1541_n 0.00238329f $X=7.635 $Y=1.16 $X2=0
+ $Y2=0
cc_785 N_A_1086_47#_c_1145_n N_SUM_c_1541_n 7.88595e-19 $X=7.77 $Y=1.16 $X2=0
+ $Y2=0
cc_786 N_A_1086_47#_M1001_g N_SUM_c_1544_n 0.00136769f $X=7.27 $Y=1.985 $X2=0
+ $Y2=0
cc_787 N_A_1086_47#_M1011_g N_SUM_c_1544_n 0.00970798f $X=7.69 $Y=1.985 $X2=0
+ $Y2=0
cc_788 N_A_1086_47#_c_1149_n N_SUM_c_1544_n 0.00384346f $X=7.215 $Y=1.555 $X2=0
+ $Y2=0
cc_789 N_A_1086_47#_M1011_g SUM 0.00208251f $X=7.69 $Y=1.985 $X2=0 $Y2=0
cc_790 N_A_1086_47#_c_1139_n SUM 0.0123928f $X=7.77 $Y=0.995 $X2=0 $Y2=0
cc_791 N_A_1086_47#_c_1142_n SUM 0.00430679f $X=7.215 $Y=1.075 $X2=0 $Y2=0
cc_792 N_A_1086_47#_c_1143_n SUM 0.00431135f $X=7.215 $Y=1.47 $X2=0 $Y2=0
cc_793 N_A_1086_47#_c_1233_p SUM 0.0136853f $X=7.635 $Y=1.16 $X2=0 $Y2=0
cc_794 N_A_1086_47#_c_1140_n N_VGND_M1009_d 0.00651691f $X=7.13 $Y=0.74 $X2=0
+ $Y2=0
cc_795 N_A_1086_47#_c_1138_n N_VGND_c_1569_n 0.00409489f $X=7.23 $Y=0.995 $X2=0
+ $Y2=0
cc_796 N_A_1086_47#_c_1151_n N_VGND_c_1569_n 0.0124309f $X=6.38 $Y=0.38 $X2=0
+ $Y2=0
cc_797 N_A_1086_47#_c_1140_n N_VGND_c_1569_n 0.0179629f $X=7.13 $Y=0.74 $X2=0
+ $Y2=0
cc_798 N_A_1086_47#_c_1139_n N_VGND_c_1571_n 0.00438629f $X=7.77 $Y=0.995 $X2=0
+ $Y2=0
cc_799 N_A_1086_47#_c_1151_n N_VGND_c_1572_n 0.0115639f $X=6.38 $Y=0.38 $X2=0
+ $Y2=0
cc_800 N_A_1086_47#_c_1140_n N_VGND_c_1572_n 0.00378546f $X=7.13 $Y=0.74 $X2=0
+ $Y2=0
cc_801 N_A_1086_47#_c_1155_n N_VGND_c_1572_n 0.047666f $X=5.71 $Y=0.425 $X2=0
+ $Y2=0
cc_802 N_A_1086_47#_c_1138_n N_VGND_c_1579_n 0.00433127f $X=7.23 $Y=0.995 $X2=0
+ $Y2=0
cc_803 N_A_1086_47#_c_1139_n N_VGND_c_1579_n 0.00424416f $X=7.77 $Y=0.995 $X2=0
+ $Y2=0
cc_804 N_A_1086_47#_c_1140_n N_VGND_c_1579_n 0.00272228f $X=7.13 $Y=0.74 $X2=0
+ $Y2=0
cc_805 N_A_1086_47#_M1027_d N_VGND_c_1584_n 0.00285934f $X=5.43 $Y=0.235 $X2=0
+ $Y2=0
cc_806 N_A_1086_47#_c_1138_n N_VGND_c_1584_n 0.00645524f $X=7.23 $Y=0.995 $X2=0
+ $Y2=0
cc_807 N_A_1086_47#_c_1139_n N_VGND_c_1584_n 0.00701197f $X=7.77 $Y=0.995 $X2=0
+ $Y2=0
cc_808 N_A_1086_47#_c_1151_n N_VGND_c_1584_n 0.00651702f $X=6.38 $Y=0.38 $X2=0
+ $Y2=0
cc_809 N_A_1086_47#_c_1140_n N_VGND_c_1584_n 0.0122148f $X=7.13 $Y=0.74 $X2=0
+ $Y2=0
cc_810 N_A_1086_47#_c_1155_n N_VGND_c_1584_n 0.0226199f $X=5.71 $Y=0.425 $X2=0
+ $Y2=0
cc_811 N_A_1086_47#_c_1155_n N_A_829_47#_c_1770_n 0.0162015f $X=5.71 $Y=0.425
+ $X2=0 $Y2=0
cc_812 N_A_1086_47#_c_1151_n A_1194_47# 0.00288105f $X=6.38 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_813 N_A_1086_47#_c_1151_n A_1266_47# 0.00470231f $X=6.38 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_814 N_A_1086_47#_c_1164_n A_1266_47# 0.00165868f $X=6.465 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_815 N_VPWR_c_1282_n N_COUT_M1005_s 0.00320325f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_816 N_VPWR_M1005_d N_COUT_c_1423_n 0.00425861f $X=0.14 $Y=1.485 $X2=0 $Y2=0
cc_817 N_VPWR_c_1304_n N_COUT_c_1423_n 0.0124697f $X=0.265 $Y=1.96 $X2=0 $Y2=0
cc_818 N_VPWR_c_1292_n COUT 0.0128161f $X=0.98 $Y=2.72 $X2=0 $Y2=0
cc_819 N_VPWR_c_1282_n COUT 0.00939489f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_820 N_VPWR_c_1282_n A_289_371# 0.0034659f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_821 N_VPWR_c_1282_n N_A_473_371#_M1000_d 0.00409863f $X=8.05 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_822 N_VPWR_c_1282_n N_A_473_371#_M1023_d 0.00226128f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_823 N_VPWR_c_1293_n N_A_473_371#_c_1477_n 0.0111986f $X=2.755 $Y=2.72 $X2=0
+ $Y2=0
cc_824 N_VPWR_c_1282_n N_A_473_371#_c_1477_n 0.00642843f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_825 N_VPWR_M1030_d N_A_473_371#_c_1465_n 0.00319397f $X=2.785 $Y=1.855 $X2=0
+ $Y2=0
cc_826 N_VPWR_c_1284_n N_A_473_371#_c_1465_n 0.0158599f $X=2.92 $Y=2.36 $X2=0
+ $Y2=0
cc_827 N_VPWR_c_1285_n N_A_473_371#_c_1465_n 0.0131777f $X=3.86 $Y=2 $X2=0 $Y2=0
cc_828 N_VPWR_c_1293_n N_A_473_371#_c_1465_n 0.00255672f $X=2.755 $Y=2.72 $X2=0
+ $Y2=0
cc_829 N_VPWR_c_1294_n N_A_473_371#_c_1465_n 0.00255672f $X=3.695 $Y=2.72 $X2=0
+ $Y2=0
cc_830 N_VPWR_c_1282_n N_A_473_371#_c_1465_n 0.0101119f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_831 N_VPWR_c_1285_n N_A_473_371#_c_1466_n 0.0255946f $X=3.86 $Y=2 $X2=0 $Y2=0
cc_832 N_VPWR_c_1294_n N_A_473_371#_c_1466_n 0.0159201f $X=3.695 $Y=2.72 $X2=0
+ $Y2=0
cc_833 N_VPWR_c_1282_n N_A_473_371#_c_1466_n 0.00891562f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_834 N_VPWR_c_1282_n N_A_829_369#_M1024_d 0.00409863f $X=8.05 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_835 N_VPWR_c_1282_n N_A_829_369#_M1012_d 0.00516727f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_836 N_VPWR_c_1295_n N_A_829_369#_c_1499_n 0.0111986f $X=4.535 $Y=2.72 $X2=0
+ $Y2=0
cc_837 N_VPWR_c_1282_n N_A_829_369#_c_1499_n 0.00642843f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_838 N_VPWR_M1016_d N_A_829_369#_c_1488_n 0.00340913f $X=4.565 $Y=1.845 $X2=0
+ $Y2=0
cc_839 N_VPWR_c_1286_n N_A_829_369#_c_1488_n 0.0158599f $X=4.7 $Y=2.36 $X2=0
+ $Y2=0
cc_840 N_VPWR_c_1295_n N_A_829_369#_c_1488_n 0.00255672f $X=4.535 $Y=2.72 $X2=0
+ $Y2=0
cc_841 N_VPWR_c_1296_n N_A_829_369#_c_1488_n 0.00255672f $X=6.89 $Y=2.72 $X2=0
+ $Y2=0
cc_842 N_VPWR_c_1282_n N_A_829_369#_c_1488_n 0.0101119f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_843 N_VPWR_c_1296_n N_A_829_369#_c_1506_n 0.0114f $X=6.89 $Y=2.72 $X2=0 $Y2=0
cc_844 N_VPWR_c_1282_n N_A_829_369#_c_1506_n 0.00642843f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_845 N_VPWR_c_1282_n A_1171_369# 0.00261003f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_846 N_VPWR_c_1282_n A_1266_371# 0.00323344f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_847 N_VPWR_c_1282_n N_SUM_M1001_s 0.00414458f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_848 N_VPWR_M1011_d N_SUM_c_1517_n 0.0041678f $X=7.765 $Y=1.485 $X2=0 $Y2=0
cc_849 N_VPWR_c_1288_n N_SUM_c_1517_n 0.0113354f $X=7.9 $Y=1.96 $X2=0 $Y2=0
cc_850 N_VPWR_c_1289_n N_SUM_c_1541_n 0.01214f $X=7.815 $Y=2.72 $X2=0 $Y2=0
cc_851 N_VPWR_c_1282_n N_SUM_c_1541_n 0.00842369f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_852 N_COUT_c_1420_n N_VGND_M1008_d 0.00311706f $X=0.605 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_853 N_COUT_c_1420_n VGND 0.00139367f $X=0.605 $Y=0.82 $X2=0 $Y2=0
cc_854 N_COUT_c_1420_n N_VGND_c_1575_n 0.00194318f $X=0.605 $Y=0.82 $X2=0 $Y2=0
cc_855 N_COUT_c_1442_n N_VGND_c_1575_n 0.0127666f $X=0.685 $Y=0.4 $X2=0 $Y2=0
cc_856 N_COUT_M1008_s N_VGND_c_1584_n 0.00218954f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_857 N_COUT_c_1420_n N_VGND_c_1584_n 0.0069814f $X=0.605 $Y=0.82 $X2=0 $Y2=0
cc_858 N_COUT_c_1442_n N_VGND_c_1584_n 0.0114218f $X=0.685 $Y=0.4 $X2=0 $Y2=0
cc_859 N_COUT_c_1420_n N_VGND_c_1585_n 0.0127122f $X=0.605 $Y=0.82 $X2=0 $Y2=0
cc_860 N_SUM_c_1515_n N_VGND_M1031_s 0.00318975f $X=7.97 $Y=0.82 $X2=0 $Y2=0
cc_861 N_SUM_c_1515_n N_VGND_c_1570_n 0.00213959f $X=7.97 $Y=0.82 $X2=0 $Y2=0
cc_862 N_SUM_c_1515_n N_VGND_c_1571_n 0.0134519f $X=7.97 $Y=0.82 $X2=0 $Y2=0
cc_863 N_SUM_c_1515_n N_VGND_c_1579_n 0.00193763f $X=7.97 $Y=0.82 $X2=0 $Y2=0
cc_864 N_SUM_c_1537_n N_VGND_c_1579_n 0.0205316f $X=7.56 $Y=0.4 $X2=0 $Y2=0
cc_865 N_SUM_M1018_d N_VGND_c_1584_n 0.00628276f $X=7.305 $Y=0.235 $X2=0 $Y2=0
cc_866 N_SUM_c_1515_n N_VGND_c_1584_n 0.00816424f $X=7.97 $Y=0.82 $X2=0 $Y2=0
cc_867 N_SUM_c_1537_n N_VGND_c_1584_n 0.012337f $X=7.56 $Y=0.4 $X2=0 $Y2=0
cc_868 N_VGND_c_1584_n A_294_47# 0.00286569f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_869 N_VGND_c_1584_n N_A_473_47#_M1025_d 0.00227466f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_870 N_VGND_c_1584_n N_A_473_47#_M1028_d 0.00204709f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_871 N_VGND_c_1576_n N_A_473_47#_c_1740_n 0.0111986f $X=2.755 $Y=0 $X2=0 $Y2=0
cc_872 N_VGND_c_1584_n N_A_473_47#_c_1740_n 0.00304042f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_873 N_VGND_M1029_d N_A_473_47#_c_1715_n 0.00158918f $X=2.785 $Y=0.235 $X2=0
+ $Y2=0
cc_874 N_VGND_c_1566_n N_A_473_47#_c_1715_n 0.0147553f $X=2.92 $Y=0.36 $X2=0
+ $Y2=0
cc_875 N_VGND_c_1576_n N_A_473_47#_c_1715_n 0.00255672f $X=2.755 $Y=0 $X2=0
+ $Y2=0
cc_876 N_VGND_c_1577_n N_A_473_47#_c_1715_n 0.00255672f $X=3.695 $Y=0 $X2=0
+ $Y2=0
cc_877 N_VGND_c_1584_n N_A_473_47#_c_1715_n 0.00461038f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_878 N_VGND_c_1567_n N_A_473_47#_c_1732_n 0.0131643f $X=3.86 $Y=0.405 $X2=0
+ $Y2=0
cc_879 N_VGND_c_1577_n N_A_473_47#_c_1732_n 0.0114f $X=3.695 $Y=0 $X2=0 $Y2=0
cc_880 N_VGND_c_1584_n N_A_473_47#_c_1732_n 0.00304042f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_881 N_VGND_c_1584_n N_A_829_47#_M1017_d 0.00227466f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_882 N_VGND_c_1584_n N_A_829_47#_M1021_d 0.00263427f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_883 N_VGND_c_1578_n N_A_829_47#_c_1773_n 0.0111986f $X=4.535 $Y=0 $X2=0 $Y2=0
cc_884 N_VGND_c_1584_n N_A_829_47#_c_1773_n 0.00304042f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_885 N_VGND_M1015_d N_A_829_47#_c_1750_n 0.00158918f $X=4.565 $Y=0.235 $X2=0
+ $Y2=0
cc_886 N_VGND_c_1568_n N_A_829_47#_c_1750_n 0.0147553f $X=4.7 $Y=0.36 $X2=0
+ $Y2=0
cc_887 N_VGND_c_1572_n N_A_829_47#_c_1750_n 0.00255672f $X=6.78 $Y=0 $X2=0 $Y2=0
cc_888 N_VGND_c_1578_n N_A_829_47#_c_1750_n 0.00255672f $X=4.535 $Y=0 $X2=0
+ $Y2=0
cc_889 N_VGND_c_1584_n N_A_829_47#_c_1750_n 0.00461038f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_890 N_VGND_c_1572_n N_A_829_47#_c_1770_n 0.0114f $X=6.78 $Y=0 $X2=0 $Y2=0
cc_891 N_VGND_c_1584_n N_A_829_47#_c_1770_n 0.00304042f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_892 N_VGND_c_1584_n A_1194_47# 0.00168648f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_893 N_VGND_c_1584_n A_1266_47# 0.0030831f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24

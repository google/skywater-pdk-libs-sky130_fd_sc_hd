* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_467_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=1.3455e+12p pd=1.194e+07u as=1.4365e+12p ps=1.352e+07u
M1001 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=1.33e+12p ps=1.266e+07u
M1002 a_467_47# A4 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_889_297# A3 a_639_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=8.1e+11p ps=7.62e+06u
M1004 VPWR B1 a_79_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1005 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_639_297# A4 a_79_21# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_467_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_1083_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.04e+12p ps=8.08e+06u
M1009 VGND A3 a_467_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_79_21# A4 a_639_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1083_297# A2 a_889_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1 a_467_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.51e+11p ps=3.68e+06u
M1014 a_467_47# B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1015 a_79_21# B1 a_467_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_889_297# A2 a_1083_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1083_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_79_21# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_467_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_639_297# A3 a_889_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A4 a_467_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_467_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

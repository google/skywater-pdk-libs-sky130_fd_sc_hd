# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.265000 1.065000 ;
        RECT 0.085000 1.065000 0.575000 1.285000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.270000 1.075000 8.010000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 0.255000 2.335000 0.725000 ;
        RECT 2.005000 0.725000 8.655000 0.905000 ;
        RECT 2.845000 0.255000 3.175000 0.725000 ;
        RECT 3.685000 0.255000 4.015000 0.725000 ;
        RECT 4.525000 0.255000 4.855000 0.725000 ;
        RECT 5.365000 0.255000 5.695000 0.725000 ;
        RECT 5.405000 1.445000 8.655000 1.615000 ;
        RECT 5.405000 1.615000 5.655000 2.125000 ;
        RECT 6.205000 0.255000 6.535000 0.725000 ;
        RECT 6.245000 1.615000 6.495000 2.125000 ;
        RECT 7.045000 0.255000 7.375000 0.725000 ;
        RECT 7.085000 1.615000 7.335000 2.125000 ;
        RECT 7.885000 0.255000 8.215000 0.725000 ;
        RECT 7.925000 1.615000 8.175000 2.125000 ;
        RECT 8.180000 0.905000 8.655000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.740000 0.085000 ;
        RECT 0.435000  0.085000 0.655000 0.895000 ;
        RECT 1.325000  0.085000 1.835000 0.905000 ;
        RECT 2.505000  0.085000 2.675000 0.555000 ;
        RECT 3.345000  0.085000 3.515000 0.555000 ;
        RECT 4.185000  0.085000 4.355000 0.555000 ;
        RECT 5.025000  0.085000 5.195000 0.555000 ;
        RECT 5.865000  0.085000 6.035000 0.555000 ;
        RECT 6.705000  0.085000 6.875000 0.555000 ;
        RECT 7.545000  0.085000 7.715000 0.555000 ;
        RECT 8.385000  0.085000 8.655000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.740000 2.805000 ;
        RECT 0.195000 1.455000 0.415000 2.635000 ;
        RECT 1.085000 1.455000 1.330000 2.635000 ;
        RECT 2.045000 1.835000 2.295000 2.635000 ;
        RECT 2.885000 1.835000 3.135000 2.635000 ;
        RECT 3.725000 1.835000 3.975000 2.635000 ;
        RECT 4.565000 1.835000 4.815000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.585000 1.455000 0.915000 2.465000 ;
      RECT 0.745000 1.065000 1.155000 1.075000 ;
      RECT 0.745000 1.075000 5.000000 1.285000 ;
      RECT 0.745000 1.285000 0.915000 1.455000 ;
      RECT 0.825000 0.255000 1.155000 1.065000 ;
      RECT 1.555000 1.455000 5.235000 1.665000 ;
      RECT 1.555000 1.665000 1.875000 2.465000 ;
      RECT 2.465000 1.665000 2.715000 2.465000 ;
      RECT 3.305000 1.665000 3.555000 2.465000 ;
      RECT 4.145000 1.665000 4.395000 2.465000 ;
      RECT 4.985000 1.665000 5.235000 2.295000 ;
      RECT 4.985000 2.295000 8.595000 2.465000 ;
      RECT 5.825000 1.785000 6.075000 2.295000 ;
      RECT 6.665000 1.785000 6.915000 2.295000 ;
      RECT 7.505000 1.785000 7.755000 2.295000 ;
      RECT 8.345000 1.785000 8.595000 2.295000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_8

* File: sky130_fd_sc_hd__dfbbp_1.spice.pex
* Created: Thu Aug 27 14:14:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFBBP_1%CLK 4 5 7 8 10 13 17 19 20 24 26
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.262 $Y=1.19
+ $X2=0.262 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_27_47# 1 2 9 13 15 17 20 26 28 29 32 36 40
+ 41 42 45 47 51 52 55 56 57 58 59 68 73 80 81 85 86 87
c249 85 0 2.05666e-19 $X=6.15 $Y=1.74
c250 52 0 2.66835e-19 $X=2.415 $Y=0.87
c251 51 0 1.79319e-19 $X=2.415 $Y=0.87
c252 45 0 1.81794e-19 $X=0.725 $Y=1.795
c253 42 0 3.29888e-20 $X=0.61 $Y=1.88
c254 26 0 3.84972e-20 $X=6.21 $Y=2.275
r255 85 88 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.15 $Y=1.74
+ $X2=6.15 $Y2=1.905
r256 85 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.15 $Y=1.74
+ $X2=6.15 $Y2=1.575
r257 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.15
+ $Y=1.74 $X2=6.15 $Y2=1.74
r258 80 83 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.745 $Y=1.74
+ $X2=2.745 $Y2=1.875
r259 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.745
+ $Y=1.74 $X2=2.745 $Y2=1.74
r260 68 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=1.87
+ $X2=6.215 $Y2=1.87
r261 66 81 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=2.535 $Y=1.765
+ $X2=2.745 $Y2=1.765
r262 66 93 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.535 $Y=1.765
+ $X2=2.44 $Y2=1.765
r263 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.535 $Y=1.87
+ $X2=2.535 $Y2=1.87
r264 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.87
+ $X2=0.695 $Y2=1.87
r265 59 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.68 $Y=1.87
+ $X2=2.535 $Y2=1.87
r266 58 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.07 $Y=1.87
+ $X2=6.215 $Y2=1.87
r267 58 59 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=6.07 $Y=1.87
+ $X2=2.68 $Y2=1.87
r268 57 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.87
+ $X2=0.695 $Y2=1.87
r269 56 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.39 $Y=1.87
+ $X2=2.535 $Y2=1.87
r270 56 57 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.39 $Y=1.87
+ $X2=0.84 $Y2=1.87
r271 52 75 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.415 $Y=0.87
+ $X2=2.305 $Y2=0.87
r272 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=0.87 $X2=2.415 $Y2=0.87
r273 49 93 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.44 $Y=1.575
+ $X2=2.44 $Y2=1.765
r274 49 51 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.44 $Y=1.575
+ $X2=2.44 $Y2=0.87
r275 48 73 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r276 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r277 45 62 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r278 45 47 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r279 44 47 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r280 43 55 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r281 42 62 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r282 42 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r283 40 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r284 40 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r285 34 41 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r286 34 36 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r287 30 32 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=6.745 $Y=1.245
+ $X2=6.745 $Y2=0.415
r288 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.67 $Y=1.32
+ $X2=6.745 $Y2=1.245
r289 28 29 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.67 $Y=1.32
+ $X2=6.285 $Y2=1.32
r290 26 88 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.21 $Y=2.275
+ $X2=6.21 $Y2=1.905
r291 22 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.21 $Y=1.395
+ $X2=6.285 $Y2=1.32
r292 22 87 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.21 $Y=1.395
+ $X2=6.21 $Y2=1.575
r293 20 83 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.715 $Y=2.275
+ $X2=2.715 $Y2=1.875
r294 15 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r295 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r296 11 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r297 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r298 7 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r299 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r300 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r301 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%D 3 7 9 10 14 15
c40 7 0 1.79319e-19 $X=1.83 $Y=2.275
r41 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.17
+ $X2=1.835 $Y2=1.335
r42 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.17
+ $X2=1.835 $Y2=1.005
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=1.17 $X2=1.835 $Y2=1.17
r44 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.955 $Y=1.19
+ $X2=1.955 $Y2=1.53
r45 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.955 $Y=1.19
+ $X2=1.955 $Y2=1.17
r46 7 17 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.83 $Y=2.275 $X2=1.83
+ $Y2=1.335
r47 3 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.83 $Y=0.445
+ $X2=1.83 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_193_47# 1 2 9 11 12 15 18 19 21 24 28 29
+ 31 33 34 36 37 39 40 41 48 49 52 56 68
c216 39 0 9.15927e-20 $X=3.022 $Y=1.12
c217 31 0 1.20913e-19 $X=6.642 $Y=1.305
c218 29 0 1.7288e-19 $X=6.325 $Y=0.87
c219 9 0 4.43992e-20 $X=2.295 $Y=2.275
r220 56 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.895 $Y=0.93
+ $X2=2.895 $Y2=1.095
r221 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.895 $Y=0.93
+ $X2=2.895 $Y2=0.765
r222 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.215 $Y=1.19
+ $X2=6.215 $Y2=1.19
r223 49 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.895
+ $Y=0.93 $X2=2.895 $Y2=0.93
r224 48 50 0.0716299 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=2.975 $Y=0.85
+ $X2=2.975 $Y2=0.965
r225 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.975 $Y=0.85
+ $X2=2.975 $Y2=0.85
r226 44 72 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.96
r227 44 68 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.51
r228 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=0.85
+ $X2=1.155 $Y2=0.85
r229 40 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.07 $Y=1.19
+ $X2=6.215 $Y2=1.19
r230 40 41 3.65098 $w=1.4e-07 $l=2.95e-06 $layer=MET1_cond $X=6.07 $Y=1.19
+ $X2=3.12 $Y2=1.19
r231 39 41 0.0723178 $w=1.4e-07 $l=1.28312e-07 $layer=MET1_cond $X=3.022 $Y=1.12
+ $X2=3.12 $Y2=1.19
r232 39 50 0.12202 $w=1.95e-07 $l=1.55e-07 $layer=MET1_cond $X=3.022 $Y=1.12
+ $X2=3.022 $Y2=0.965
r233 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=0.85
+ $X2=1.155 $Y2=0.85
r234 36 48 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.83 $Y=0.85
+ $X2=2.975 $Y2=0.85
r235 36 37 1.89356 $w=1.4e-07 $l=1.53e-06 $layer=MET1_cond $X=2.83 $Y=0.85
+ $X2=1.3 $Y2=0.85
r236 34 66 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.66 $Y=1.74
+ $X2=6.66 $Y2=1.875
r237 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.74 $X2=6.66 $Y2=1.74
r238 31 53 26.3101 $w=1.78e-07 $l=4.27e-07 $layer=LI1_cond $X=6.642 $Y=1.215
+ $X2=6.215 $Y2=1.215
r239 31 33 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=6.642 $Y=1.305
+ $X2=6.642 $Y2=1.74
r240 29 60 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.325 $Y=0.87
+ $X2=6.2 $Y2=0.87
r241 28 53 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=6.267 $Y=0.87
+ $X2=6.267 $Y2=1.125
r242 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.325
+ $Y=0.87 $X2=6.325 $Y2=0.87
r243 24 66 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.63 $Y=2.275
+ $X2=6.63 $Y2=1.875
r244 19 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.2 $Y=0.705
+ $X2=6.2 $Y2=0.87
r245 19 21 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.2 $Y=0.705
+ $X2=6.2 $Y2=0.415
r246 18 59 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.835 $Y=1.245
+ $X2=2.835 $Y2=1.095
r247 15 58 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.835 $Y=0.415
+ $X2=2.835 $Y2=0.765
r248 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.76 $Y=1.32
+ $X2=2.835 $Y2=1.245
r249 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.76 $Y=1.32
+ $X2=2.37 $Y2=1.32
r250 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.295 $Y=1.395
+ $X2=2.37 $Y2=1.32
r251 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.295 $Y=1.395
+ $X2=2.295 $Y2=2.275
r252 2 72 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r253 1 68 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_648_21# 1 2 9 13 17 19 21 22 26 28 30 31
+ 32 35 36 41 45 49
c146 9 0 7.56837e-20 $X=3.315 $Y=0.445
r147 49 56 10.4783 $w=2.76e-07 $l=6e-08 $layer=POLY_cond $X=5.665 $Y=1.15
+ $X2=5.725 $Y2=1.15
r148 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.665
+ $Y=1.15 $X2=5.665 $Y2=1.15
r149 45 48 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.665 $Y=0.98
+ $X2=5.665 $Y2=1.15
r150 43 44 14.1313 $w=2.59e-07 $l=3e-07 $layer=LI1_cond $X=4.575 $Y=0.68
+ $X2=4.575 $Y2=0.98
r151 36 53 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.74
+ $X2=3.4 $Y2=1.905
r152 36 52 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.74
+ $X2=3.4 $Y2=1.575
r153 35 38 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.465 $Y=1.74
+ $X2=3.465 $Y2=1.91
r154 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.74 $X2=3.425 $Y2=1.74
r155 33 44 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=0.98
+ $X2=4.575 $Y2=0.98
r156 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.5 $Y=0.98
+ $X2=5.665 $Y2=0.98
r157 32 33 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.5 $Y=0.98
+ $X2=4.74 $Y2=0.98
r158 30 44 5.44435 $w=2.59e-07 $l=9.88686e-08 $layer=LI1_cond $X=4.605 $Y=1.065
+ $X2=4.575 $Y2=0.98
r159 30 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.605 $Y=1.065
+ $X2=4.605 $Y2=1.785
r160 29 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=1.91
+ $X2=4.175 $Y2=1.91
r161 28 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.52 $Y=1.91
+ $X2=4.605 $Y2=1.785
r162 28 29 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=4.52 $Y=1.91
+ $X2=4.26 $Y2=1.91
r163 24 41 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.175 $Y=2.035
+ $X2=4.175 $Y2=1.91
r164 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.175 $Y=2.035
+ $X2=4.175 $Y2=2.21
r165 23 38 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.59 $Y=1.91
+ $X2=3.465 $Y2=1.91
r166 22 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=1.91
+ $X2=4.175 $Y2=1.91
r167 22 23 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=4.09 $Y=1.91 $X2=3.59
+ $Y2=1.91
r168 19 56 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=0.985
+ $X2=5.725 $Y2=1.15
r169 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.725 $Y=0.985
+ $X2=5.725 $Y2=0.555
r170 15 49 30.5616 $w=2.76e-07 $l=2.43926e-07 $layer=POLY_cond $X=5.49 $Y=1.315
+ $X2=5.665 $Y2=1.15
r171 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.49 $Y=1.315
+ $X2=5.49 $Y2=2.065
r172 13 53 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.315 $Y=2.275
+ $X2=3.315 $Y2=1.905
r173 9 52 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.315 $Y=0.445
+ $X2=3.315 $Y2=1.575
r174 2 41 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=2.065 $X2=4.175 $Y2=1.87
r175 2 26 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=2.065 $X2=4.175 $Y2=2.21
r176 1 43 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=4.44
+ $Y=0.235 $X2=4.575 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%SET_B 1 3 7 11 15 17 19 20 26 27 33
c131 33 0 1.0279e-19 $X=7.64 $Y=0.98
c132 19 0 1.0411e-19 $X=7.45 $Y=0.85
c133 15 0 1.0852e-19 $X=7.76 $Y=2.275
r134 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=0.98
+ $X2=7.67 $Y2=1.145
r135 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=0.98
+ $X2=7.67 $Y2=0.815
r136 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.64
+ $Y=0.98 $X2=7.64 $Y2=0.98
r137 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.595 $Y=0.85
+ $X2=7.595 $Y2=0.85
r138 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=0.85
+ $X2=3.915 $Y2=0.85
r139 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.45 $Y=0.85
+ $X2=7.595 $Y2=0.85
r140 19 20 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=7.45 $Y=0.85
+ $X2=4.06 $Y2=0.85
r141 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.755
+ $Y=0.98 $X2=3.755 $Y2=0.98
r142 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.915 $Y=0.85
+ $X2=3.915 $Y2=0.85
r143 15 36 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.76 $Y=2.275
+ $X2=7.76 $Y2=1.145
r144 11 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.65 $Y=0.445
+ $X2=7.65 $Y2=0.815
r145 5 30 38.532 $w=3.09e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.865 $Y=0.815
+ $X2=3.78 $Y2=0.98
r146 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.865 $Y=0.815
+ $X2=3.865 $Y2=0.445
r147 1 30 38.532 $w=3.09e-07 $l=1.94808e-07 $layer=POLY_cond $X=3.845 $Y=1.145
+ $X2=3.78 $Y2=0.98
r148 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.845 $Y=1.145
+ $X2=3.845 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_474_413# 1 2 9 13 15 19 24 26 27 32 35
c105 35 0 1.0411e-19 $X=4.265 $Y=1.32
c106 32 0 4.43992e-20 $X=3.4 $Y=1.3
r107 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.32
+ $X2=4.295 $Y2=1.485
r108 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.32
+ $X2=4.295 $Y2=1.155
r109 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=1.32 $X2=4.265 $Y2=1.32
r110 31 32 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=1.3
+ $X2=3.4 $Y2=1.3
r111 29 31 12.1472 $w=2.08e-07 $l=2.3e-07 $layer=LI1_cond $X=3.085 $Y=1.3
+ $X2=3.315 $Y2=1.3
r112 27 34 8.9562 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=1.32
+ $X2=4.265 $Y2=1.32
r113 27 32 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.1 $Y=1.32 $X2=3.4
+ $Y2=1.32
r114 26 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.315 $Y=1.195
+ $X2=3.315 $Y2=1.3
r115 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.315 $Y=0.465
+ $X2=3.315 $Y2=1.195
r116 23 29 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.085 $Y=1.405
+ $X2=3.085 $Y2=1.3
r117 23 24 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.085 $Y=1.405
+ $X2=3.085 $Y2=2.25
r118 19 25 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.23 $Y=0.365
+ $X2=3.315 $Y2=0.465
r119 19 21 36.6 $w=1.98e-07 $l=6.6e-07 $layer=LI1_cond $X=3.23 $Y=0.365 $X2=2.57
+ $Y2=0.365
r120 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3 $Y=2.335
+ $X2=3.085 $Y2=2.25
r121 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3 $Y=2.335
+ $X2=2.505 $Y2=2.335
r122 13 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.385 $Y=2.065
+ $X2=4.385 $Y2=1.485
r123 9 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.365 $Y=0.555
+ $X2=4.365 $Y2=1.155
r124 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=2.065 $X2=2.505 $Y2=2.335
r125 1 21 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.57 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_942_21# 1 2 9 13 17 21 23 24 25 27 31 34
+ 35 42 43 46 49 58 61
c160 58 0 1.89563e-19 $X=8.66 $Y=1.32
c161 42 0 2.58372e-20 $X=8.83 $Y=1.53
c162 27 0 1.511e-19 $X=9.38 $Y=1.66
r163 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.32 $X2=8.87 $Y2=1.32
r164 58 60 32.9707 $w=3.07e-07 $l=2.1e-07 $layer=POLY_cond $X=8.66 $Y=1.32
+ $X2=8.87 $Y2=1.32
r165 57 58 9.4202 $w=3.07e-07 $l=6e-08 $layer=POLY_cond $X=8.6 $Y=1.32 $X2=8.66
+ $Y2=1.32
r166 52 54 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.785 $Y=1.32
+ $X2=4.805 $Y2=1.32
r167 50 61 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=8.922 $Y=1.53
+ $X2=8.922 $Y2=1.32
r168 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.975 $Y=1.53
+ $X2=8.975 $Y2=1.53
r169 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.755 $Y=1.53
+ $X2=5.755 $Y2=1.53
r170 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.9 $Y=1.53
+ $X2=5.755 $Y2=1.53
r171 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.83 $Y=1.53
+ $X2=8.975 $Y2=1.53
r172 42 43 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=8.83 $Y=1.53
+ $X2=5.9 $Y2=1.53
r173 41 50 1.88582 $w=2.73e-07 $l=4.5e-08 $layer=LI1_cond $X=8.922 $Y=1.575
+ $X2=8.922 $Y2=1.53
r174 40 61 16.5533 $w=2.73e-07 $l=3.95e-07 $layer=LI1_cond $X=8.922 $Y=0.925
+ $X2=8.922 $Y2=1.32
r175 38 46 27.1304 $w=2.38e-07 $l=5.65e-07 $layer=LI1_cond $X=5.19 $Y=1.535
+ $X2=5.755 $Y2=1.535
r176 37 38 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=1.535
+ $X2=5.19 $Y2=1.535
r177 35 54 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.025 $Y=1.32
+ $X2=4.805 $Y2=1.32
r178 34 37 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.025 $Y=1.32
+ $X2=5.025 $Y2=1.535
r179 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.025
+ $Y=1.32 $X2=5.025 $Y2=1.32
r180 29 31 15.938 $w=2.33e-07 $l=3.25e-07 $layer=LI1_cond $X=9.357 $Y=0.755
+ $X2=9.357 $Y2=0.43
r181 25 41 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=9.06 $Y=1.66
+ $X2=8.922 $Y2=1.575
r182 25 27 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.06 $Y=1.66
+ $X2=9.38 $Y2=1.66
r183 24 40 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=9.06 $Y=0.84
+ $X2=8.922 $Y2=0.925
r184 23 29 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=9.24 $Y=0.84
+ $X2=9.357 $Y2=0.755
r185 23 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=9.24 $Y=0.84
+ $X2=9.06 $Y2=0.84
r186 19 58 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.66 $Y=1.155
+ $X2=8.66 $Y2=1.32
r187 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.66 $Y=1.155 $X2=8.66
+ $Y2=0.555
r188 15 57 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.6 $Y=1.485
+ $X2=8.6 $Y2=1.32
r189 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.6 $Y=1.485
+ $X2=8.6 $Y2=2.065
r190 11 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.485
+ $X2=4.805 $Y2=1.32
r191 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.805 $Y=1.485
+ $X2=4.805 $Y2=2.065
r192 7 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.155
+ $X2=4.785 $Y2=1.32
r193 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.785 $Y=1.155 $X2=4.785
+ $Y2=0.555
r194 2 27 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=9.255
+ $Y=1.505 $X2=9.38 $Y2=1.66
r195 1 31 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=9.265
+ $Y=0.235 $X2=9.39 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_1429_21# 1 2 9 13 15 17 20 22 23 25 27 28
+ 30 31 33 36 38 41 45 46 48 49 52 54 57 58 61 62 66 68 70
c178 70 0 1.15237e-19 $X=10.025 $Y=1.16
c179 66 0 1.22108e-19 $X=8.525 $Y=0.687
c180 20 0 1.511e-19 $X=10.075 $Y=1.985
c181 9 0 8.81272e-20 $X=7.22 $Y=0.445
r182 71 79 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=10.025 $Y=1.16
+ $X2=10.075 $Y2=1.16
r183 70 73 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.985 $Y=1.16
+ $X2=9.985 $Y2=1.325
r184 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.025
+ $Y=1.16 $X2=10.025 $Y2=1.16
r185 64 66 4.49631 $w=1.83e-07 $l=7.5e-08 $layer=LI1_cond $X=8.45 $Y=0.687
+ $X2=8.525 $Y2=0.687
r186 61 73 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.945 $Y=1.915
+ $X2=9.945 $Y2=1.325
r187 59 68 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.615 $Y=2 $X2=8.525
+ $Y2=2
r188 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.86 $Y=2
+ $X2=9.945 $Y2=1.915
r189 58 59 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=9.86 $Y=2
+ $X2=8.615 $Y2=2
r190 57 68 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=1.915
+ $X2=8.525 $Y2=2
r191 56 66 0.88302 $w=1.8e-07 $l=9.3e-08 $layer=LI1_cond $X=8.525 $Y=0.78
+ $X2=8.525 $Y2=0.687
r192 56 57 69.9343 $w=1.78e-07 $l=1.135e-06 $layer=LI1_cond $X=8.525 $Y=0.78
+ $X2=8.525 $Y2=1.915
r193 55 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=2 $X2=8.03
+ $Y2=2
r194 54 68 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.435 $Y=2 $X2=8.525
+ $Y2=2
r195 54 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.435 $Y=2 $X2=8.115
+ $Y2=2
r196 50 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.03 $Y=2.085
+ $X2=8.03 $Y2=2
r197 50 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.03 $Y=2.085
+ $X2=8.03 $Y2=2.21
r198 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.945 $Y=2 $X2=8.03
+ $Y2=2
r199 48 49 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.945 $Y=2
+ $X2=7.505 $Y2=2
r200 46 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=1.74
+ $X2=7.31 $Y2=1.905
r201 46 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=1.74
+ $X2=7.31 $Y2=1.575
r202 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.74 $X2=7.34 $Y2=1.74
r203 43 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.38 $Y=1.915
+ $X2=7.505 $Y2=2
r204 43 45 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=7.38 $Y=1.915
+ $X2=7.38 $Y2=1.74
r205 39 41 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=10.885 $Y=1.61
+ $X2=11.015 $Y2=1.61
r206 34 36 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=10.885 $Y=0.805
+ $X2=11.015 $Y2=0.805
r207 31 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=1.685
+ $X2=11.015 $Y2=1.61
r208 31 33 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=11.015 $Y=1.685
+ $X2=11.015 $Y2=2.085
r209 28 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=0.73
+ $X2=11.015 $Y2=0.805
r210 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.015 $Y=0.73
+ $X2=11.015 $Y2=0.445
r211 27 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.885 $Y=1.535
+ $X2=10.885 $Y2=1.61
r212 26 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.885 $Y=1.295
+ $X2=10.885 $Y2=1.16
r213 26 27 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.885 $Y=1.295
+ $X2=10.885 $Y2=1.535
r214 25 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.885 $Y=1.025
+ $X2=10.885 $Y2=1.16
r215 24 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.885 $Y=0.88
+ $X2=10.885 $Y2=0.805
r216 24 25 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=10.885 $Y=0.88
+ $X2=10.885 $Y2=1.025
r217 23 79 15.1926 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.15 $Y=1.16
+ $X2=10.075 $Y2=1.16
r218 22 38 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=10.81 $Y=1.16
+ $X2=10.885 $Y2=1.16
r219 22 23 146.635 $w=2.7e-07 $l=6.6e-07 $layer=POLY_cond $X=10.81 $Y=1.16
+ $X2=10.15 $Y2=1.16
r220 18 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.075 $Y=1.325
+ $X2=10.075 $Y2=1.16
r221 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.075 $Y=1.325
+ $X2=10.075 $Y2=1.985
r222 15 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.075 $Y=0.995
+ $X2=10.075 $Y2=1.16
r223 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.075 $Y=0.995
+ $X2=10.075 $Y2=0.56
r224 13 76 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.22 $Y=2.275
+ $X2=7.22 $Y2=1.905
r225 9 75 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.22 $Y=0.445
+ $X2=7.22 $Y2=1.575
r226 2 52 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=7.835
+ $Y=2.065 $X2=8.03 $Y2=2.21
r227 1 64 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=8.315
+ $Y=0.235 $X2=8.45 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_1255_47# 1 2 9 13 15 19 24 26 27 29 31 32
c99 32 0 2.58372e-20 $X=8.18 $Y=1.24
c100 31 0 1.75976e-19 $X=8.18 $Y=1.24
c101 26 0 3.84972e-20 $X=7 $Y=2.25
r102 32 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.18 $Y=1.24
+ $X2=8.18 $Y2=1.405
r103 32 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.18 $Y=1.24
+ $X2=8.18 $Y2=1.075
r104 31 34 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=8.155 $Y=1.24
+ $X2=8.155 $Y2=1.32
r105 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.18
+ $Y=1.24 $X2=8.18 $Y2=1.24
r106 28 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.085 $Y=1.32 $X2=7
+ $Y2=1.32
r107 27 34 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=8.045 $Y=1.32
+ $X2=8.155 $Y2=1.32
r108 27 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.045 $Y=1.32
+ $X2=7.085 $Y2=1.32
r109 25 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=1.405 $X2=7
+ $Y2=1.32
r110 25 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=7 $Y=1.405 $X2=7
+ $Y2=2.25
r111 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=1.235 $X2=7
+ $Y2=1.32
r112 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7 $Y=0.465 $X2=7
+ $Y2=1.235
r113 19 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.915 $Y=0.365
+ $X2=7 $Y2=0.465
r114 19 21 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=6.915 $Y=0.365
+ $X2=6.485 $Y2=0.365
r115 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.915 $Y=2.335
+ $X2=7 $Y2=2.25
r116 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.915 $Y=2.335
+ $X2=6.42 $Y2=2.335
r117 13 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.24 $Y=2.065
+ $X2=8.24 $Y2=1.405
r118 9 37 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.24 $Y=0.555
+ $X2=8.24 $Y2=1.075
r119 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=2.065 $X2=6.42 $Y2=2.335
r120 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.275
+ $Y=0.235 $X2=6.485 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%RESET_B 3 7 9 12 17
r38 12 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=9.52 $Y=1.18
+ $X2=9.52 $Y2=1.345
r39 12 14 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=9.52 $Y=1.18
+ $X2=9.52 $Y2=1.015
r40 9 17 4.76009 $w=2.28e-07 $l=9.5e-08 $layer=LI1_cond $X=9.525 $Y=1.21
+ $X2=9.43 $Y2=1.21
r41 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.525
+ $Y=1.18 $X2=9.525 $Y2=1.18
r42 7 14 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=9.6 $Y=0.445 $X2=9.6
+ $Y2=1.015
r43 3 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.59 $Y=1.825
+ $X2=9.59 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_2136_47# 1 2 9 12 16 20 24 25 27 29
c50 27 0 1.4681e-19 $X=10.812 $Y=1.16
r51 25 30 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.417 $Y=1.16
+ $X2=11.417 $Y2=1.325
r52 25 29 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.417 $Y=1.16
+ $X2=11.417 $Y2=0.995
r53 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.405
+ $Y=1.16 $X2=11.405 $Y2=1.16
r54 22 27 1.17559 $w=3.3e-07 $l=1.58e-07 $layer=LI1_cond $X=10.97 $Y=1.16
+ $X2=10.812 $Y2=1.16
r55 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=10.97 $Y=1.16
+ $X2=11.405 $Y2=1.16
r56 18 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=10.812 $Y=1.325
+ $X2=10.812 $Y2=1.16
r57 18 20 21.4025 $w=3.13e-07 $l=5.85e-07 $layer=LI1_cond $X=10.812 $Y=1.325
+ $X2=10.812 $Y2=1.91
r58 14 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=10.812 $Y=0.995
+ $X2=10.812 $Y2=1.16
r59 14 16 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=10.812 $Y=0.995
+ $X2=10.812 $Y2=0.51
r60 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.49 $Y=1.985
+ $X2=11.49 $Y2=1.325
r61 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.49 $Y=0.56
+ $X2=11.49 $Y2=0.995
r62 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.68
+ $Y=1.765 $X2=10.805 $Y2=1.91
r63 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=10.68
+ $Y=0.235 $X2=10.805 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 46 47 48
+ 52 53 55 57 63 68 80 91 95 102 103 106 109 112 115 126 128
c184 103 0 1.81794e-19 $X=11.73 $Y=2.72
c185 1 0 3.29888e-20 $X=0.545 $Y=1.815
r186 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r187 124 126 9.28831 $w=5.48e-07 $l=1.4e-07 $layer=LI1_cond $X=9.89 $Y=2.53
+ $X2=10.03 $Y2=2.53
r188 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r189 122 124 0.543672 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=9.865 $Y=2.53
+ $X2=9.89 $Y2=2.53
r190 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r191 115 118 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=7.515 $Y=2.34
+ $X2=7.515 $Y2=2.72
r192 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r193 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r194 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r195 103 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r196 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r197 100 128 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=11.445 $Y=2.72
+ $X2=11.297 $Y2=2.72
r198 100 102 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.445 $Y=2.72
+ $X2=11.73 $Y2=2.72
r199 99 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r200 99 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=9.89 $Y2=2.72
r201 98 126 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=10.03 $Y2=2.72
r202 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r203 95 128 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=11.15 $Y=2.72
+ $X2=11.297 $Y2=2.72
r204 95 98 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.15 $Y=2.72
+ $X2=10.81 $Y2=2.72
r205 94 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r206 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r207 91 122 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=9.755 $Y=2.53
+ $X2=9.865 $Y2=2.53
r208 91 93 17.0713 $w=5.48e-07 $l=7.85e-07 $layer=LI1_cond $X=9.755 $Y=2.53
+ $X2=8.97 $Y2=2.53
r209 90 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r210 90 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=7.59 $Y2=2.72
r211 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r212 87 118 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=7.515 $Y2=2.72
r213 87 89 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=8.51 $Y2=2.72
r214 86 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r215 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r216 83 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r217 82 85 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r218 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r219 80 118 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.325 $Y=2.72
+ $X2=7.515 $Y2=2.72
r220 80 85 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.325 $Y=2.72
+ $X2=7.13 $Y2=2.72
r221 79 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r222 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r223 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r224 76 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r225 75 78 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r226 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r227 73 112 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.79 $Y=2.72
+ $X2=3.6 $Y2=2.72
r228 73 75 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.79 $Y=2.72
+ $X2=3.91 $Y2=2.72
r229 72 113 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r230 72 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r231 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r232 69 109 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.61 $Y2=2.72
r233 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r234 68 112 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.41 $Y=2.72
+ $X2=3.6 $Y2=2.72
r235 68 71 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=3.41 $Y=2.72
+ $X2=2.07 $Y2=2.72
r236 67 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r237 67 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r238 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r239 64 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r240 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r241 63 109 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.61 $Y2=2.72
r242 63 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r243 57 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r244 55 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r245 53 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r246 53 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r247 52 89 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=8.645 $Y=2.72
+ $X2=8.51 $Y2=2.72
r248 51 52 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.81 $Y=2.53
+ $X2=8.645 $Y2=2.53
r249 48 93 1.08734 $w=5.48e-07 $l=5e-08 $layer=LI1_cond $X=8.92 $Y=2.53 $X2=8.97
+ $Y2=2.53
r250 48 51 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=8.92 $Y=2.53
+ $X2=8.81 $Y2=2.53
r251 46 78 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.88 $Y=2.72 $X2=4.83
+ $Y2=2.72
r252 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=2.72
+ $X2=5.045 $Y2=2.72
r253 45 82 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=5.21 $Y=2.72 $X2=5.29
+ $Y2=2.72
r254 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=2.72
+ $X2=5.045 $Y2=2.72
r255 41 128 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=11.297 $Y=2.635
+ $X2=11.297 $Y2=2.72
r256 41 43 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=11.297 $Y=2.635
+ $X2=11.297 $Y2=1.94
r257 37 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=2.635
+ $X2=5.045 $Y2=2.72
r258 37 39 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.045 $Y=2.635
+ $X2=5.045 $Y2=2
r259 33 112 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2.72
r260 33 35 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2.29
r261 29 109 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=2.635
+ $X2=1.61 $Y2=2.72
r262 29 31 13.6647 $w=3.48e-07 $l=4.15e-07 $layer=LI1_cond $X=1.61 $Y=2.635
+ $X2=1.61 $Y2=2.22
r263 25 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r264 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r265 8 43 300 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=2 $X=11.09
+ $Y=1.765 $X2=11.28 $Y2=1.94
r266 7 122 600 $w=1.7e-07 $l=9.29637e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.505 $X2=9.865 $Y2=2.34
r267 6 51 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=8.675
+ $Y=1.645 $X2=8.81 $Y2=2.34
r268 5 115 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=2.065 $X2=7.49 $Y2=2.34
r269 4 39 300 $w=1.7e-07 $l=4.29651e-07 $layer=licon1_PDIFF $count=2 $X=4.88
+ $Y=1.645 $X2=5.045 $Y2=2
r270 3 35 600 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=2.065 $X2=3.575 $Y2=2.29
r271 2 31 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.065 $X2=1.62 $Y2=2.22
r272 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_381_47# 1 2 8 9 10 11 12 15 19
r58 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=1.965
+ $X2=2.04 $Y2=2.3
r59 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r60 11 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.965
r61 11 12 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.58 $Y2=1.88
r62 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r63 9 10 21.89 $w=1.88e-07 $l=3.75e-07 $layer=LI1_cond $X=1.955 $Y=0.73 $X2=1.58
+ $Y2=0.73
r64 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=1.795
+ $X2=1.58 $Y2=1.88
r65 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.495 $Y=0.825
+ $X2=1.58 $Y2=0.73
r66 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.495 $Y=0.825
+ $X2=1.495 $Y2=1.795
r67 2 19 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.065 $X2=2.04 $Y2=2.3
r68 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%Q_N 1 2 9 10 11 12 13 18 21
r30 18 21 2.69684 $w=2.85e-07 $l=6.3e-08 $layer=LI1_cond $X=10.342 $Y=0.573
+ $X2=10.342 $Y2=0.51
r31 12 13 15.9725 $w=2.83e-07 $l=3.95e-07 $layer=LI1_cond $X=10.342 $Y=1.815
+ $X2=10.342 $Y2=2.21
r32 11 30 6.22369 $w=2.83e-07 $l=1.31e-07 $layer=LI1_cond $X=10.342 $Y=0.584
+ $X2=10.342 $Y2=0.715
r33 11 18 0.444803 $w=2.83e-07 $l=1.1e-08 $layer=LI1_cond $X=10.342 $Y=0.584
+ $X2=10.342 $Y2=0.573
r34 11 21 0.470877 $w=2.85e-07 $l=1.1e-08 $layer=LI1_cond $X=10.342 $Y=0.499
+ $X2=10.342 $Y2=0.51
r35 10 30 49.5033 $w=2.03e-07 $l=9.15e-07 $layer=LI1_cond $X=10.382 $Y=1.63
+ $X2=10.382 $Y2=0.715
r36 9 12 1.73877 $w=2.83e-07 $l=4.3e-08 $layer=LI1_cond $X=10.342 $Y=1.772
+ $X2=10.342 $Y2=1.815
r37 9 10 6.6685 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=10.342 $Y=1.772
+ $X2=10.342 $Y2=1.63
r38 2 12 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=10.15
+ $Y=1.485 $X2=10.285 $Y2=1.815
r39 1 21 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=10.15
+ $Y=0.235 $X2=10.285 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%Q 1 2 10 11 12 13 14 15
r16 14 15 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=11.745 $Y=1.82
+ $X2=11.745 $Y2=2.21
r17 11 14 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=11.745 $Y=1.575
+ $X2=11.745 $Y2=1.82
r18 11 12 6.14153 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=11.745 $Y=1.575
+ $X2=11.745 $Y2=1.445
r19 10 12 33.2332 $w=2.13e-07 $l=6.2e-07 $layer=LI1_cond $X=11.767 $Y=0.825
+ $X2=11.767 $Y2=1.445
r20 9 13 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=11.745 $Y=0.695
+ $X2=11.745 $Y2=0.51
r21 9 10 6.14153 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=11.745 $Y=0.695
+ $X2=11.745 $Y2=0.825
r22 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=11.565
+ $Y=1.485 $X2=11.7 $Y2=1.82
r23 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=11.565
+ $Y=0.235 $X2=11.7 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 48 51
+ 52 54 55 57 58 59 61 63 69 93 100 107 108 111 114 117 120
c185 108 0 2.71124e-20 $X=11.73 $Y=0
c186 51 0 1.75242e-19 $X=3.57 $Y=0
c187 40 0 1.0279e-19 $X=7.44 $Y=0.36
r188 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r189 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r190 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r191 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r192 108 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r193 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r194 105 120 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=11.445 $Y=0
+ $X2=11.297 $Y2=0
r195 105 107 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.445 $Y=0
+ $X2=11.73 $Y2=0
r196 104 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r197 104 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=9.89 $Y2=0
r198 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r199 101 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.03 $Y=0
+ $X2=9.865 $Y2=0
r200 101 103 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=10.03 $Y=0
+ $X2=10.81 $Y2=0
r201 100 120 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=11.297 $Y2=0
r202 100 103 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=10.81 $Y2=0
r203 99 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r204 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r205 96 99 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r206 95 98 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=0 $X2=9.43
+ $Y2=0
r207 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r208 93 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.7 $Y=0 $X2=9.865
+ $Y2=0
r209 93 98 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.7 $Y=0 $X2=9.43
+ $Y2=0
r210 92 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r211 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r212 89 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=7.13 $Y2=0
r213 88 91 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=7.13
+ $Y2=0
r214 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r215 86 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r216 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r217 83 86 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r218 82 85 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r219 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r220 80 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r221 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r222 77 80 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r223 77 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r224 76 79 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r225 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r226 74 114 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.61
+ $Y2=0
r227 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r228 73 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r229 73 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r230 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r231 70 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r232 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r233 69 114 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.61
+ $Y2=0
r234 69 72 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0
+ $X2=1.15 $Y2=0
r235 63 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r236 61 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r237 59 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r238 59 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r239 57 91 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.265 $Y=0
+ $X2=7.13 $Y2=0
r240 57 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.265 $Y=0 $X2=7.395
+ $Y2=0
r241 56 95 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.525 $Y=0 $X2=7.59
+ $Y2=0
r242 56 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.525 $Y=0 $X2=7.395
+ $Y2=0
r243 54 85 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.29
+ $Y2=0
r244 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.515
+ $Y2=0
r245 53 88 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.68 $Y=0 $X2=5.75
+ $Y2=0
r246 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=5.515
+ $Y2=0
r247 51 79 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.45
+ $Y2=0
r248 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.655
+ $Y2=0
r249 50 82 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.91
+ $Y2=0
r250 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.655
+ $Y2=0
r251 46 120 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=11.297 $Y=0.085
+ $X2=11.297 $Y2=0
r252 46 48 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=11.297 $Y=0.085
+ $X2=11.297 $Y2=0.38
r253 42 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.865 $Y=0.085
+ $X2=9.865 $Y2=0
r254 42 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.865 $Y=0.085
+ $X2=9.865 $Y2=0.38
r255 38 58 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=0.085
+ $X2=7.395 $Y2=0
r256 38 40 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=7.395 $Y=0.085
+ $X2=7.395 $Y2=0.36
r257 34 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0
r258 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0.38
r259 30 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0
r260 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0.36
r261 26 114 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0
r262 26 28 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0.38
r263 22 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r264 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r265 7 48 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=11.09
+ $Y=0.235 $X2=11.28 $Y2=0.38
r266 6 44 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=9.675
+ $Y=0.235 $X2=9.865 $Y2=0.38
r267 5 40 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.295
+ $Y=0.235 $X2=7.44 $Y2=0.36
r268 4 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.235 $X2=5.515 $Y2=0.38
r269 3 32 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=3.39
+ $Y=0.235 $X2=3.655 $Y2=0.36
r270 2 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r271 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_788_47# 1 2 7 11 13
c26 13 0 7.56837e-20 $X=4.075 $Y=0.34
r27 13 16 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.075 $Y=0.34
+ $X2=4.075 $Y2=0.46
r28 9 11 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.995 $Y=0.425
+ $X2=4.995 $Y2=0.55
r29 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.24 $Y=0.34
+ $X2=4.075 $Y2=0.34
r30 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.91 $Y=0.34
+ $X2=4.995 $Y2=0.425
r31 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.91 $Y=0.34 $X2=4.24
+ $Y2=0.34
r32 2 11 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.235 $X2=4.995 $Y2=0.55
r33 1 16 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=3.94
+ $Y=0.235 $X2=4.075 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBP_1%A_1545_47# 1 2 7 9 16
r22 9 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.95 $Y=0.34 $X2=7.95
+ $Y2=0.46
r23 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.115 $Y=0.34 $X2=7.95
+ $Y2=0.34
r24 7 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.34
+ $X2=8.87 $Y2=0.34
r25 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.785 $Y=0.34
+ $X2=8.115 $Y2=0.34
r26 2 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.235 $X2=8.87 $Y2=0.42
r27 1 12 182 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=1 $X=7.725
+ $Y=0.235 $X2=7.95 $Y2=0.46
.ends


* File: sky130_fd_sc_hd__xor2_2.spice.pex
* Created: Thu Aug 27 14:49:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XOR2_2%A 1 3 6 8 10 13 15 17 20 22 24 27 30 32 33 35
+ 42 44 45 46 51 56
c131 56 0 1.33666e-19 $X=3.105 $Y=1.16
c132 42 0 1.52981e-19 $X=0.79 $Y=1.175
r133 45 46 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.71 $Y=1.53
+ $X2=1.15 $Y2=1.53
r134 44 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=1.53
+ $X2=1.15 $Y2=1.53
r135 40 51 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.71 $Y=1.16
+ $X2=0.905 $Y2=1.16
r136 40 48 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.71 $Y=1.16
+ $X2=0.485 $Y2=1.16
r137 39 42 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=0.71 $Y=1.175
+ $X2=0.79 $Y2=1.175
r138 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.16 $X2=0.71 $Y2=1.16
r139 36 56 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.065 $Y=1.16
+ $X2=3.105 $Y2=1.16
r140 36 53 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.065 $Y=1.16
+ $X2=2.685 $Y2=1.16
r141 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.065
+ $Y=1.16 $X2=3.065 $Y2=1.16
r142 33 35 65.7136 $w=1.98e-07 $l=1.185e-06 $layer=LI1_cond $X=1.88 $Y=1.175
+ $X2=3.065 $Y2=1.175
r143 32 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=1.445
+ $X2=1.71 $Y2=1.53
r144 31 33 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.795 $Y=1.275
+ $X2=1.88 $Y2=1.175
r145 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.795 $Y=1.275
+ $X2=1.795 $Y2=1.445
r146 30 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.79 $Y=1.445
+ $X2=0.875 $Y2=1.53
r147 29 42 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.79 $Y=1.275 $X2=0.79
+ $Y2=1.175
r148 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.79 $Y=1.275
+ $X2=0.79 $Y2=1.445
r149 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.325
+ $X2=3.105 $Y2=1.16
r150 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.105 $Y=1.325
+ $X2=3.105 $Y2=1.985
r151 22 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=0.995
+ $X2=3.105 $Y2=1.16
r152 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.105 $Y=0.995
+ $X2=3.105 $Y2=0.56
r153 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.685 $Y=1.325
+ $X2=2.685 $Y2=1.16
r154 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.685 $Y=1.325
+ $X2=2.685 $Y2=1.985
r155 15 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.685 $Y=0.995
+ $X2=2.685 $Y2=1.16
r156 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.685 $Y=0.995
+ $X2=2.685 $Y2=0.56
r157 11 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r158 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r159 8 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r160 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r161 4 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.16
r162 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.985
r163 1 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.16
r164 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%B 1 3 6 8 10 13 15 17 20 22 24 27 29 31 32 38
+ 45 46 53
c120 46 0 1.52981e-19 $X=1.745 $Y=1.16
c121 38 0 1.33666e-19 $X=3.91 $Y=1.19
c122 15 0 1.92258e-19 $X=3.525 $Y=0.995
r123 51 53 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=1.16 $X2=4
+ $Y2=1.16
r124 48 51 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=3.525 $Y=1.16
+ $X2=3.925 $Y2=1.16
r125 44 46 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.375 $Y=1.16
+ $X2=1.745 $Y2=1.16
r126 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.375
+ $Y=1.16 $X2=1.375 $Y2=1.16
r127 41 44 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.325 $Y=1.16
+ $X2=1.375 $Y2=1.16
r128 35 45 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=1.375 $Y2=1.175
r129 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.19
+ $X2=1.15 $Y2=1.19
r130 32 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.19
+ $X2=1.15 $Y2=1.19
r131 31 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.765 $Y=1.19
+ $X2=3.91 $Y2=1.19
r132 31 32 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=3.765 $Y=1.19
+ $X2=1.295 $Y2=1.19
r133 29 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.925
+ $Y=1.16 $X2=3.925 $Y2=1.16
r134 29 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=1.19
+ $X2=3.91 $Y2=1.19
r135 25 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=1.325 $X2=4
+ $Y2=1.16
r136 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4 $Y=1.325 $X2=4
+ $Y2=1.985
r137 22 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=0.995 $X2=4
+ $Y2=1.16
r138 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4 $Y=0.995 $X2=4
+ $Y2=0.56
r139 18 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.325
+ $X2=3.525 $Y2=1.16
r140 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.525 $Y=1.325
+ $X2=3.525 $Y2=1.985
r141 15 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=0.995
+ $X2=3.525 $Y2=1.16
r142 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.525 $Y=0.995
+ $X2=3.525 $Y2=0.56
r143 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=1.325
+ $X2=1.745 $Y2=1.16
r144 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.745 $Y=1.325
+ $X2=1.745 $Y2=1.985
r145 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=1.16
r146 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=0.56
r147 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.325
+ $X2=1.325 $Y2=1.16
r148 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.325 $Y=1.325
+ $X2=1.325 $Y2=1.985
r149 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=0.995
+ $X2=1.325 $Y2=1.16
r150 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.325 $Y=0.995
+ $X2=1.325 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%A_112_47# 1 2 3 10 12 15 17 19 22 25 26 27 28
+ 29 32 34 38 40 43 44 45 47 48 50 53 54 62
r169 54 57 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.535 $Y=1.87
+ $X2=1.535 $Y2=1.96
r170 51 62 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.11 $Y=1.16
+ $X2=5.36 $Y2=1.16
r171 51 59 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=5.11 $Y=1.16
+ $X2=4.94 $Y2=1.16
r172 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.11
+ $Y=1.16 $X2=5.11 $Y2=1.16
r173 48 50 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.785 $Y=1.16
+ $X2=5.11 $Y2=1.16
r174 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.7 $Y=1.245
+ $X2=4.785 $Y2=1.16
r175 46 47 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.7 $Y=1.245 $X2=4.7
+ $Y2=1.445
r176 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.615 $Y=1.53
+ $X2=4.7 $Y2=1.445
r177 44 45 156.251 $w=1.68e-07 $l=2.395e-06 $layer=LI1_cond $X=4.615 $Y=1.53
+ $X2=2.22 $Y2=1.53
r178 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=1.615
+ $X2=2.22 $Y2=1.53
r179 42 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.135 $Y=1.615
+ $X2=2.135 $Y2=1.785
r180 41 54 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.66 $Y=1.87
+ $X2=1.535 $Y2=1.87
r181 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=1.87
+ $X2=2.135 $Y2=1.785
r182 40 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.05 $Y=1.87
+ $X2=1.66 $Y2=1.87
r183 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0.725
+ $X2=1.535 $Y2=0.39
r184 35 53 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=0.815
+ $X2=0.695 $Y2=0.815
r185 34 36 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.37 $Y=0.815
+ $X2=1.535 $Y2=0.725
r186 34 35 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.37 $Y=0.815
+ $X2=0.86 $Y2=0.815
r187 30 53 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.695 $Y=0.725
+ $X2=0.695 $Y2=0.815
r188 30 32 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.695 $Y=0.725
+ $X2=0.695 $Y2=0.39
r189 28 54 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.41 $Y=1.87
+ $X2=1.535 $Y2=1.87
r190 28 29 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=1.41 $Y=1.87
+ $X2=0.29 $Y2=1.87
r191 26 53 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=0.815
+ $X2=0.695 $Y2=0.815
r192 26 27 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.53 $Y=0.815
+ $X2=0.29 $Y2=0.815
r193 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.205 $Y=1.785
+ $X2=0.29 $Y2=1.87
r194 24 27 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.205 $Y=0.905
+ $X2=0.29 $Y2=0.815
r195 24 25 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.205 $Y=0.905
+ $X2=0.205 $Y2=1.785
r196 20 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.36 $Y=1.325
+ $X2=5.36 $Y2=1.16
r197 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.36 $Y=1.325
+ $X2=5.36 $Y2=1.985
r198 17 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.36 $Y=0.995
+ $X2=5.36 $Y2=1.16
r199 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.36 $Y=0.995
+ $X2=5.36 $Y2=0.56
r200 13 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.94 $Y=1.325
+ $X2=4.94 $Y2=1.16
r201 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.94 $Y=1.325
+ $X2=4.94 $Y2=1.985
r202 10 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.94 $Y=0.995
+ $X2=4.94 $Y2=1.16
r203 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.94 $Y=0.995
+ $X2=4.94 $Y2=0.56
r204 3 57 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.4
+ $Y=1.485 $X2=1.535 $Y2=1.96
r205 2 38 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.4
+ $Y=0.235 $X2=1.535 $Y2=0.39
r206 1 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.235 $X2=0.695 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%A_27_297# 1 2 3 10 13 17 18 21 24 25
c56 24 0 1.9698e-19 $X=1.15 $Y=2.21
r57 25 31 8.39676 $w=2.47e-07 $l=1.7e-07 $layer=LI1_cond $X=1.115 $Y=2.21
+ $X2=1.115 $Y2=2.38
r58 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.21
+ $X2=1.15 $Y2=2.21
r59 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.21
+ $X2=0.23 $Y2=2.21
r60 18 20 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.375 $Y=2.21
+ $X2=0.23 $Y2=2.21
r61 17 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.005 $Y=2.21
+ $X2=1.15 $Y2=2.21
r62 17 18 0.779701 $w=1.4e-07 $l=6.3e-07 $layer=MET1_cond $X=1.005 $Y=2.21
+ $X2=0.375 $Y2=2.21
r63 13 15 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.955 $Y=2.3 $X2=1.955
+ $Y2=2.38
r64 11 31 2.92482 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.24 $Y=2.38
+ $X2=1.115 $Y2=2.38
r65 10 15 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=2.38
+ $X2=1.955 $Y2=2.38
r66 10 11 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.83 $Y=2.38 $X2=1.24
+ $Y2=2.38
r67 3 13 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=1.485 $X2=1.955 $Y2=2.3
r68 2 25 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.485 $X2=1.115 $Y2=2.3
r69 1 21 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%VPWR 1 2 3 12 16 20 23 24 25 27 39 45 46 49
+ 52
c89 23 0 1.9698e-19 $X=2.77 $Y=2.72
r90 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r91 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r92 46 53 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r93 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r94 43 52 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.915 $Y=2.72
+ $X2=3.762 $Y2=2.72
r95 43 45 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=3.915 $Y=2.72
+ $X2=5.75 $Y2=2.72
r96 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r97 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r98 39 52 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.762 $Y2=2.72
r99 39 41 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r100 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r101 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r102 35 38 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 35 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r104 34 37 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r106 32 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=0.695 $Y2=2.72
r107 32 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=1.15 $Y2=2.72
r108 27 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.57 $Y=2.72
+ $X2=0.695 $Y2=2.72
r109 27 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.57 $Y=2.72
+ $X2=0.23 $Y2=2.72
r110 25 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r112 23 37 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.77 $Y=2.72
+ $X2=2.53 $Y2=2.72
r113 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.77 $Y=2.72
+ $X2=2.895 $Y2=2.72
r114 22 41 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=3.45 $Y2=2.72
r115 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=2.895 $Y2=2.72
r116 18 52 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.762 $Y=2.635
+ $X2=3.762 $Y2=2.72
r117 18 20 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=3.762 $Y=2.635
+ $X2=3.762 $Y2=2.3
r118 14 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=2.635
+ $X2=2.895 $Y2=2.72
r119 14 16 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.895 $Y=2.635
+ $X2=2.895 $Y2=2.3
r120 10 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r121 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.3
r122 3 20 600 $w=1.7e-07 $l=9.05028e-07 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=1.485 $X2=3.79 $Y2=2.3
r123 2 16 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=1.485 $X2=2.895 $Y2=2.3
r124 1 12 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.485 $X2=0.695 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%A_470_297# 1 2 3 4 5 19 20 21 24 28 32 35 38
+ 41 44
r47 43 44 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=4.73 $Y=2.125
+ $X2=4.855 $Y2=2.125
r48 40 43 9.14648 $w=6.78e-07 $l=5.2e-07 $layer=LI1_cond $X=4.21 $Y=2.125
+ $X2=4.73 $Y2=2.125
r49 40 41 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=4.21 $Y=2.125
+ $X2=4.085 $Y2=2.125
r50 35 36 7.68595 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=2.442 $Y=2.3
+ $X2=2.442 $Y2=2.125
r51 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.57 $Y=2.295
+ $X2=5.57 $Y2=1.96
r52 28 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.445 $Y=2.38
+ $X2=5.57 $Y2=2.295
r53 28 44 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.445 $Y=2.38
+ $X2=4.855 $Y2=2.38
r54 27 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.44 $Y=1.87
+ $X2=3.315 $Y2=1.87
r55 27 41 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.44 $Y=1.87
+ $X2=4.085 $Y2=1.87
r56 22 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=1.955
+ $X2=3.315 $Y2=1.87
r57 22 24 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.315 $Y=1.955
+ $X2=3.315 $Y2=1.96
r58 20 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.19 $Y=1.87
+ $X2=3.315 $Y2=1.87
r59 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.19 $Y=1.87 $X2=2.6
+ $Y2=1.87
r60 19 36 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=1.96
+ $X2=2.495 $Y2=2.125
r61 16 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.495 $Y=1.955
+ $X2=2.6 $Y2=1.87
r62 16 19 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=2.495 $Y=1.955
+ $X2=2.495 $Y2=1.96
r63 5 32 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.435
+ $Y=1.485 $X2=5.57 $Y2=1.96
r64 4 43 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.605
+ $Y=1.485 $X2=4.73 $Y2=1.96
r65 3 40 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.075
+ $Y=1.485 $X2=4.21 $Y2=1.96
r66 2 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.18
+ $Y=1.485 $X2=3.315 $Y2=1.96
r67 1 35 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.485 $X2=2.475 $Y2=2.3
r68 1 19 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.485 $X2=2.475 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%X 1 2 3 10 15 19 21 23 26
c51 19 0 1.92258e-19 $X=3.955 $Y=0.775
r52 17 19 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=0.775
+ $X2=3.955 $Y2=0.775
r53 15 23 3.16883 $w=2.08e-07 $l=6e-08 $layer=LI1_cond $X=5.69 $Y=1.52 $X2=5.75
+ $Y2=1.52
r54 15 26 28.5195 $w=2.08e-07 $l=5.4e-07 $layer=LI1_cond $X=5.69 $Y=1.52
+ $X2=5.15 $Y2=1.52
r55 14 21 31.5215 $w=2.09e-07 $l=5.4e-07 $layer=LI1_cond $X=5.69 $Y=0.775
+ $X2=5.15 $Y2=0.775
r56 14 15 14.3353 $w=4.08e-07 $l=5.1e-07 $layer=LI1_cond $X=5.69 $Y=0.905
+ $X2=5.69 $Y2=1.415
r57 10 21 9.90026 $w=2.09e-07 $l=1.83916e-07 $layer=LI1_cond $X=4.985 $Y=0.815
+ $X2=5.15 $Y2=0.775
r58 10 19 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=4.985 $Y=0.815
+ $X2=3.955 $Y2=0.815
r59 3 26 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.015
+ $Y=1.485 $X2=5.15 $Y2=1.62
r60 2 21 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.15 $Y2=0.73
r61 1 17 182 $w=1.7e-07 $l=5.82301e-07 $layer=licon1_NDIFF $count=1 $X=3.6
+ $Y=0.235 $X2=3.79 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 56 57 58 80 81
r99 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r100 78 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r101 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r102 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r103 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r104 72 75 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=4.37 $Y2=0
r105 71 74 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.37
+ $Y2=0
r106 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r107 69 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r108 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r109 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r110 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r111 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r112 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r113 60 84 3.40825 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r114 60 62 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.69
+ $Y2=0
r115 58 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r116 58 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r117 56 77 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.485 $Y=0
+ $X2=5.29 $Y2=0
r118 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.57
+ $Y2=0
r119 55 80 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.75
+ $Y2=0
r120 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.57
+ $Y2=0
r121 53 74 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.645 $Y=0
+ $X2=4.37 $Y2=0
r122 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=0 $X2=4.73
+ $Y2=0
r123 52 77 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.815 $Y=0
+ $X2=5.29 $Y2=0
r124 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=0 $X2=4.73
+ $Y2=0
r125 50 68 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.53
+ $Y2=0
r126 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.895
+ $Y2=0
r127 49 71 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.98 $Y=0 $X2=2.99
+ $Y2=0
r128 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0 $X2=2.895
+ $Y2=0
r129 47 65 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.61
+ $Y2=0
r130 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.955
+ $Y2=0
r131 46 68 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.53
+ $Y2=0
r132 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.955
+ $Y2=0
r133 44 62 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.69
+ $Y2=0
r134 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.115
+ $Y2=0
r135 43 65 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.61
+ $Y2=0
r136 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.115
+ $Y2=0
r137 39 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=0.085
+ $X2=5.57 $Y2=0
r138 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.57 $Y=0.085
+ $X2=5.57 $Y2=0.39
r139 35 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=0.085
+ $X2=4.73 $Y2=0
r140 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.73 $Y=0.085
+ $X2=4.73 $Y2=0.39
r141 31 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0
r142 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0.39
r143 27 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0
r144 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0.39
r145 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r146 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.39
r147 19 84 3.40825 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.18 $Y2=0
r148 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.39
r149 6 41 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.235 $X2=5.57 $Y2=0.39
r150 5 37 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.605
+ $Y=0.235 $X2=4.73 $Y2=0.39
r151 4 33 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.76
+ $Y=0.235 $X2=2.895 $Y2=0.39
r152 3 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.235 $X2=1.955 $Y2=0.39
r153 2 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.115 $Y2=0.39
r154 1 21 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_2%A_470_47# 1 2 3 12 14 15 19 20 22
r48 20 22 42.4309 $w=2.18e-07 $l=8.1e-07 $layer=LI1_cond $X=3.4 $Y=0.365
+ $X2=4.21 $Y2=0.365
r49 17 19 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=3.275 $Y=0.725
+ $X2=3.275 $Y2=0.54
r50 16 20 6.85268 $w=2.2e-07 $l=1.71391e-07 $layer=LI1_cond $X=3.275 $Y=0.475
+ $X2=3.4 $Y2=0.365
r51 16 19 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=3.275 $Y=0.475
+ $X2=3.275 $Y2=0.54
r52 14 17 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=3.15 $Y=0.815
+ $X2=3.275 $Y2=0.725
r53 14 15 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.15 $Y=0.815
+ $X2=2.64 $Y2=0.815
r54 10 15 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.475 $Y=0.725
+ $X2=2.64 $Y2=0.815
r55 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.475 $Y=0.725
+ $X2=2.475 $Y2=0.39
r56 3 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.235 $X2=4.21 $Y2=0.39
r57 2 19 182 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.235 $X2=3.315 $Y2=0.54
r58 1 12 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=2.35
+ $Y=0.235 $X2=2.475 $Y2=0.39
.ends


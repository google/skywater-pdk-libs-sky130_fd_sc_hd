* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s25_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
M1000 X a_331_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=5.287e+11p ps=5.41e+06u
M1001 VPWR a_225_47# a_331_47# VPB phighvt w=820000u l=250000u
+  ad=9.58e+11p pd=7.97e+06u as=2.132e+11p ps=2.16e+06u
M1002 X a_331_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
M1003 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1005 VPWR a_331_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_225_47# a_27_47# VPWR VPB phighvt w=820000u l=250000u
+  ad=2.132e+11p pd=2.16e+06u as=0p ps=0u
M1007 a_225_47# a_27_47# VGND VNB nshort w=650000u l=250000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1008 VGND a_225_47# a_331_47# VNB nshort w=650000u l=250000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1009 VGND a_331_47# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__dfsbp_1.spice.pex
* Created: Thu Aug 27 14:15:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFSBP_1%CLK 4 5 7 8 10 13 17 19 20 24 26
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r47 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.265 $Y=1.19
+ $X2=0.265 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_27_47# 1 2 9 13 15 17 20 24 28 31 35 36 37
+ 40 42 46 47 50 51 52 54 55 59 61 62 63 64 73 78 85 86 92 93 96
c273 92 0 3.28258e-19 $X=5.155 $Y=1.74
c274 86 0 3.30612e-20 $X=2.765 $Y=1.74
c275 85 0 2.53448e-20 $X=2.765 $Y=1.74
c276 73 0 1.81067e-19 $X=5.29 $Y=1.87
c277 63 0 1.39518e-19 $X=5.145 $Y=1.87
c278 61 0 1.01003e-19 $X=2.385 $Y=1.87
c279 52 0 3.16972e-20 $X=5.07 $Y=0.81
c280 51 0 1.753e-19 $X=5.82 $Y=0.81
c281 47 0 9.52104e-20 $X=2.435 $Y=0.87
c282 46 0 1.76471e-19 $X=2.435 $Y=0.87
c283 40 0 1.81794e-19 $X=0.725 $Y=1.795
c284 37 0 3.29888e-20 $X=0.61 $Y=1.88
c285 24 0 7.27138e-20 $X=5.065 $Y=2.275
r286 93 104 6.31985 $w=3.08e-07 $l=1.7e-07 $layer=LI1_cond $X=5.155 $Y=1.81
+ $X2=4.985 $Y2=1.81
r287 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.74 $X2=5.155 $Y2=1.74
r288 89 92 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.065 $Y=1.74
+ $X2=5.155 $Y2=1.74
r289 85 88 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.765 $Y=1.74
+ $X2=2.765 $Y2=1.875
r290 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.74 $X2=2.765 $Y2=1.74
r291 73 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r292 71 86 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.765 $Y2=1.765
r293 71 99 2.12292 $w=3.78e-07 $l=7e-08 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.46 $Y2=1.765
r294 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=1.87
r295 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=1.87
+ $X2=0.73 $Y2=1.87
r296 64 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.87
+ $X2=2.53 $Y2=1.87
r297 63 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r298 63 64 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=2.675 $Y2=1.87
r299 62 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=1.87
+ $X2=0.73 $Y2=1.87
r300 61 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=2.53 $Y2=1.87
r301 61 62 1.86881 $w=1.4e-07 $l=1.51e-06 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=0.875 $Y2=1.87
r302 59 96 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.985 $Y=0.93
+ $X2=5.985 $Y2=0.765
r303 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=0.93 $X2=5.985 $Y2=0.93
r304 55 58 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.985 $Y=0.81
+ $X2=5.985 $Y2=0.93
r305 51 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.985 $Y2=0.81
r306 51 52 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.07 $Y2=0.81
r307 50 104 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.985 $Y=1.655
+ $X2=4.985 $Y2=1.81
r308 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.985 $Y=0.895
+ $X2=5.07 $Y2=0.81
r309 49 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.985 $Y=0.895
+ $X2=4.985 $Y2=1.655
r310 47 80 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.435 $Y=0.87
+ $X2=2.305 $Y2=0.87
r311 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=0.87 $X2=2.435 $Y2=0.87
r312 44 99 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=1.765
r313 44 46 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=0.87
r314 43 78 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r315 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r316 40 67 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r317 40 42 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r318 39 42 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r319 38 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r320 37 67 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r321 37 38 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r322 35 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r323 35 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r324 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r325 29 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r326 28 96 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.045 $Y=0.445
+ $X2=6.045 $Y2=0.765
r327 22 89 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=1.74
r328 22 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=2.275
r329 20 88 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.875
r330 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r331 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r332 11 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r333 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r334 7 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r335 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r336 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r337 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%D 3 7 9 10 14 15
c39 14 0 1.34441e-19 $X=1.855 $Y=1.17
c40 7 0 1.76471e-19 $X=1.83 $Y=2.065
r41 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.335
r42 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.005
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.17 $X2=1.855 $Y2=1.17
r44 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.53
r45 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.17
r46 7 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.83 $Y=2.065
+ $X2=1.83 $Y2=1.335
r47 3 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.83 $Y=0.555
+ $X2=1.83 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_193_47# 1 2 9 11 12 15 18 21 23 25 28 29
+ 30 32 33 34 41 42 45 46 53 58
c196 46 0 4.72633e-20 $X=5.33 $Y=1.19
c197 45 0 2.56901e-19 $X=5.33 $Y=1.19
c198 41 0 3.30612e-20 $X=2.99 $Y=0.85
c199 34 0 2.53448e-20 $X=3.135 $Y=1.19
c200 33 0 1.51904e-19 $X=5.185 $Y=1.19
c201 32 0 9.52104e-20 $X=3.027 $Y=1.12
c202 25 0 1.67681e-19 $X=5.605 $Y=2.275
c203 23 0 1.753e-19 $X=5.605 $Y=1.455
c204 9 0 4.43992e-20 $X=2.315 $Y=2.275
r205 53 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=1.095
r206 53 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=0.765
r207 46 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.335
+ $Y=1.26 $X2=5.335 $Y2=1.26
r208 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.33 $Y=1.19
+ $X2=5.33 $Y2=1.19
r209 42 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=0.93 $X2=2.915 $Y2=0.93
r210 41 43 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.965
r211 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.85
r212 37 62 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.96
r213 37 58 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.51
r214 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0.85
+ $X2=1.15 $Y2=0.85
r215 33 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.19
+ $X2=5.33 $Y2=1.19
r216 33 34 2.53712 $w=1.4e-07 $l=2.05e-06 $layer=MET1_cond $X=5.185 $Y=1.19
+ $X2=3.135 $Y2=1.19
r217 32 34 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.135 $Y2=1.19
r218 32 43 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.027 $Y2=0.965
r219 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=0.85
+ $X2=1.15 $Y2=0.85
r220 29 41 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=2.99 $Y2=0.85
r221 29 30 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=1.295 $Y2=0.85
r222 28 49 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=5.47 $Y=1.26
+ $X2=5.335 $Y2=1.26
r223 23 28 52.102 $w=1.88e-07 $l=2.09464e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.575 $Y2=1.26
r224 23 25 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.605 $Y2=2.275
r225 19 28 36.719 $w=1.88e-07 $l=1.39911e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.575 $Y2=1.26
r226 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.565 $Y2=0.445
r227 18 56 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.855 $Y=1.245
+ $X2=2.855 $Y2=1.095
r228 15 55 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.855 $Y=0.415
+ $X2=2.855 $Y2=0.765
r229 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.855 $Y2=1.245
r230 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.39 $Y2=1.32
r231 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.39 $Y2=1.32
r232 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.315 $Y2=2.275
r233 2 62 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r234 1 58 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_652_21# 1 2 9 13 15 19 21 25 28 30 31 35
+ 38
c115 38 0 1.32054e-19 $X=4.625 $Y=0.895
c116 35 0 2.11834e-19 $X=4.075 $Y=1.96
c117 28 0 3.22473e-19 $X=4.625 $Y=1.835
c118 21 0 1.87283e-19 $X=4.54 $Y=1.96
r119 36 38 6.44012 $w=3.38e-07 $l=1.9e-07 $layer=LI1_cond $X=4.435 $Y=0.895
+ $X2=4.625 $Y2=0.895
r120 31 42 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.905
r121 31 41 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.575
r122 30 33 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=3.485 $Y=1.74
+ $X2=3.485 $Y2=1.96
r123 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.74 $X2=3.445 $Y2=1.74
r124 27 38 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=0.895
r125 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=1.835
r126 23 36 2.53954 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.895
r127 23 25 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.46
r128 22 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.96
+ $X2=4.075 $Y2=1.96
r129 21 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.625 $Y2=1.835
r130 21 22 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.16 $Y2=1.96
r131 17 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=1.96
r132 17 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=2.21
r133 16 33 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.61 $Y=1.96
+ $X2=3.485 $Y2=1.96
r134 15 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=4.075 $Y2=1.96
r135 15 16 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=3.61 $Y2=1.96
r136 13 42 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.335 $Y=2.275
+ $X2=3.335 $Y2=1.905
r137 9 41 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.335 $Y=0.445
+ $X2=3.335 $Y2=1.575
r138 2 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.065 $X2=4.075 $Y2=2.21
r139 1 25 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.235 $X2=4.475 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%SET_B 1 3 7 11 17 19 20 24 26 27 29 30 36 37
c135 37 0 1.72331e-19 $X=7.13 $Y=0.85
c136 29 0 2.95874e-19 $X=6.985 $Y=0.85
c137 26 0 1.49785e-19 $X=6.99 $Y=0.9
c138 19 0 1.94282e-20 $X=6.895 $Y=1.535
c139 1 0 9.39349e-20 $X=3.865 $Y=1.145
r140 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0.85
+ $X2=7.13 $Y2=0.85
r141 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=0.85
+ $X2=3.91 $Y2=0.85
r142 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=7.13 $Y2=0.85
r143 29 30 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=4.055 $Y2=0.85
r144 27 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=0.98 $X2=3.775 $Y2=0.98
r145 27 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0.85
+ $X2=3.91 $Y2=0.85
r146 26 37 5.97563 $w=2.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.99 $Y=0.87
+ $X2=7.13 $Y2=0.87
r147 24 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=0.98
+ $X2=6.825 $Y2=1.145
r148 24 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=0.98
+ $X2=6.825 $Y2=0.815
r149 23 26 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=0.9
+ $X2=6.99 $Y2=0.9
r150 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.825
+ $Y=0.98 $X2=6.825 $Y2=0.98
r151 19 20 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=6.895 $Y=1.535
+ $X2=6.895 $Y2=1.685
r152 19 44 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.885 $Y=1.535
+ $X2=6.885 $Y2=1.145
r153 17 20 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.905 $Y=2.275
+ $X2=6.905 $Y2=1.685
r154 11 43 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.765 $Y=0.445
+ $X2=6.765 $Y2=0.815
r155 5 40 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.81 $Y2=0.98
r156 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.905 $Y2=0.445
r157 1 40 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.81 $Y2=0.98
r158 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.865 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_476_47# 1 2 7 9 11 14 16 20 22 24 25 26 30
+ 35 37 38 43 44 53
c157 53 0 1.95729e-19 $X=4.705 $Y=1.4
c158 43 0 4.43992e-20 $X=3.44 $Y=1.3
c159 26 0 1.01003e-19 $X=3.02 $Y=2.335
c160 22 0 3.81194e-20 $X=5.205 $Y=0.735
c161 16 0 1.15925e-19 $X=5.13 $Y=0.825
c162 7 0 3.16972e-20 $X=4.265 $Y=0.735
r163 48 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.705 $Y2=1.4
r164 48 50 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.265 $Y2=1.4
r165 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.285
+ $Y=1.4 $X2=4.285 $Y2=1.4
r166 44 47 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.245 $Y=1.32
+ $X2=4.245 $Y2=1.4
r167 42 43 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=1.3
+ $X2=3.44 $Y2=1.3
r168 40 42 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=3.105 $Y=1.3
+ $X2=3.355 $Y2=1.3
r169 38 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=4.245 $Y2=1.32
r170 38 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=3.44 $Y2=1.32
r171 37 42 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.355 $Y=1.195
+ $X2=3.355 $Y2=1.3
r172 36 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.355 $Y=0.465
+ $X2=3.355 $Y2=1.195
r173 34 40 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=1.3
r174 34 35 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=2.25
r175 30 36 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=3.355 $Y2=0.465
r176 30 32 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=2.59 $Y2=0.365
r177 26 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=3.105 $Y2=2.25
r178 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=2.525 $Y2=2.335
r179 22 24 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.205 $Y=0.735
+ $X2=5.205 $Y2=0.445
r180 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=1.4
r181 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=2.275
r182 17 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.34 $Y=0.825
+ $X2=4.265 $Y2=0.825
r183 16 22 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=5.205 $Y2=0.735
r184 16 17 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=4.34 $Y2=0.825
r185 12 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=1.4
r186 12 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=2.275
r187 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.235
+ $X2=4.265 $Y2=1.4
r188 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=0.825
r189 10 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=1.235
r190 7 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.825
r191 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.445
r192 2 28 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.065 $X2=2.525 $Y2=2.335
r193 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.59 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_1178_261# 1 2 8 11 15 19 24 28 31 35 38 39
c76 38 0 1.67681e-19 $X=7.51 $Y=1.67
c77 31 0 1.94282e-20 $X=7.735 $Y=1.575
c78 19 0 6.59327e-20 $X=6.405 $Y=1.38
r79 37 39 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.735 $Y2=1.67
r80 37 38 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.51 $Y2=1.67
r81 33 35 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.595 $Y=0.515
+ $X2=7.735 $Y2=0.515
r82 31 39 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=7.735 $Y=1.575
+ $X2=7.735 $Y2=1.67
r83 30 35 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.735 $Y=0.68
+ $X2=7.735 $Y2=0.515
r84 30 31 52.244 $w=1.88e-07 $l=8.95e-07 $layer=LI1_cond $X=7.735 $Y=0.68
+ $X2=7.735 $Y2=1.575
r85 26 37 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.67
r86 26 28 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.87
r87 24 42 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=6.06 $Y=1.66
+ $X2=6.06 $Y2=1.825
r88 23 38 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=6.095 $Y=1.66
+ $X2=7.51 $Y2=1.66
r89 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.095
+ $Y=1.66 $X2=6.095 $Y2=1.66
r90 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=1.38
r91 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=0.445
r92 11 42 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.965 $Y=2.275
+ $X2=5.965 $Y2=1.825
r93 8 24 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=6.06 $Y=1.655 $X2=6.06
+ $Y2=1.66
r94 7 19 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.06 $Y=1.38
+ $X2=6.405 $Y2=1.38
r95 7 8 33.9437 $w=3.4e-07 $l=2e-07 $layer=POLY_cond $X=6.06 $Y=1.455 $X2=6.06
+ $Y2=1.655
r96 2 28 300 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=2 $X=7.46
+ $Y=1.645 $X2=7.595 $Y2=1.87
r97 1 33 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_1028_413# 1 2 3 12 16 18 19 22 26 28 31 33
+ 34 36 37 39 40 43 45 48 50 55 56 60 61 62 65 70 72 75 77 79
c189 75 0 9.39049e-20 $X=6.405 $Y=1.32
c190 55 0 7.27138e-20 $X=5.675 $Y=1.915
c191 50 0 1.39518e-19 $X=5.59 $Y=2.29
c192 26 0 7.85839e-20 $X=8.325 $Y=1.985
c193 22 0 7.85839e-20 $X=8.325 $Y=0.56
r194 78 82 10.5355 $w=3.66e-07 $l=8e-08 $layer=POLY_cond $X=7.305 $Y=1.225
+ $X2=7.385 $Y2=1.225
r195 77 79 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=1.29
+ $X2=7.14 $Y2=1.29
r196 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.305
+ $Y=1.26 $X2=7.305 $Y2=1.26
r197 68 70 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=2.085
+ $X2=6.66 $Y2=2.21
r198 67 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=6.405 $Y2=1.32
r199 67 79 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=7.14 $Y2=1.32
r200 65 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.235
+ $X2=6.405 $Y2=1.32
r201 64 65 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.405 $Y=0.475
+ $X2=6.405 $Y2=1.235
r202 63 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2 $X2=5.675
+ $Y2=2
r203 62 68 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=6.54 $Y=2
+ $X2=6.66 $Y2=2.085
r204 62 63 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.54 $Y=2 $X2=5.76
+ $Y2=2
r205 60 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=6.405 $Y2=1.32
r206 60 61 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=5.76 $Y2=1.32
r207 56 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=6.405 $Y2=0.475
r208 56 58 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=5.805 $Y2=0.39
r209 55 72 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=1.915
+ $X2=5.675 $Y2=2
r210 54 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.675 $Y=1.405
+ $X2=5.76 $Y2=1.32
r211 54 55 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.675 $Y=1.405
+ $X2=5.675 $Y2=1.915
r212 50 72 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.675 $Y=2.29
+ $X2=5.675 $Y2=2
r213 50 52 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=5.59 $Y=2.29
+ $X2=5.275 $Y2=2.29
r214 46 48 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=9.135 $Y=1.695
+ $X2=9.265 $Y2=1.695
r215 41 43 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=9.135 $Y=0.805
+ $X2=9.265 $Y2=0.805
r216 37 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.265 $Y=1.77
+ $X2=9.265 $Y2=1.695
r217 37 39 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.265 $Y=1.77
+ $X2=9.265 $Y2=2.165
r218 34 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.265 $Y=0.73
+ $X2=9.265 $Y2=0.805
r219 34 36 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.265 $Y=0.73
+ $X2=9.265 $Y2=0.445
r220 33 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.135 $Y=1.62
+ $X2=9.135 $Y2=1.695
r221 32 45 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.135 $Y=1.295
+ $X2=9.135 $Y2=1.16
r222 32 33 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=9.135 $Y=1.295
+ $X2=9.135 $Y2=1.62
r223 31 45 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.135 $Y=1.025
+ $X2=9.135 $Y2=1.16
r224 30 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.135 $Y=0.88
+ $X2=9.135 $Y2=0.805
r225 30 31 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=9.135 $Y=0.88
+ $X2=9.135 $Y2=1.025
r226 29 40 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=8.4 $Y=1.16
+ $X2=8.325 $Y2=1.16
r227 28 45 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=9.06 $Y=1.16
+ $X2=9.135 $Y2=1.16
r228 28 29 146.635 $w=2.7e-07 $l=6.6e-07 $layer=POLY_cond $X=9.06 $Y=1.16
+ $X2=8.4 $Y2=1.16
r229 24 40 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.325 $Y=1.295
+ $X2=8.325 $Y2=1.16
r230 24 26 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.325 $Y=1.295
+ $X2=8.325 $Y2=1.985
r231 20 40 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.325 $Y=1.025
+ $X2=8.325 $Y2=1.16
r232 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.325 $Y=1.025
+ $X2=8.325 $Y2=0.56
r233 19 82 13.2898 $w=3.66e-07 $l=1.0247e-07 $layer=POLY_cond $X=7.46 $Y=1.16
+ $X2=7.385 $Y2=1.225
r234 18 40 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=8.25 $Y=1.16
+ $X2=8.325 $Y2=1.16
r235 18 19 175.517 $w=2.7e-07 $l=7.9e-07 $layer=POLY_cond $X=8.25 $Y=1.16
+ $X2=7.46 $Y2=1.16
r236 14 82 23.7042 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.385 $Y=1.425
+ $X2=7.385 $Y2=1.225
r237 14 16 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.385 $Y=1.425
+ $X2=7.385 $Y2=2.065
r238 10 82 23.7042 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.385 $Y=1.025
+ $X2=7.385 $Y2=1.225
r239 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.385 $Y=1.025
+ $X2=7.385 $Y2=0.505
r240 3 70 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=2.065 $X2=6.695 $Y2=2.21
r241 2 52 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=2.065 $X2=5.275 $Y2=2.33
r242 1 58 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=5.64
+ $Y=0.235 $X2=5.805 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_1786_47# 1 2 9 12 16 20 24 25 27 29
c53 27 0 3.0812e-19 $X=9.055 $Y=1.16
r54 25 30 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=9.667 $Y=1.16
+ $X2=9.667 $Y2=1.325
r55 25 29 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=9.667 $Y=1.16
+ $X2=9.667 $Y2=0.995
r56 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.655
+ $Y=1.16 $X2=9.655 $Y2=1.16
r57 22 27 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.22 $Y=1.16
+ $X2=9.055 $Y2=1.16
r58 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=9.22 $Y=1.16
+ $X2=9.655 $Y2=1.16
r59 18 27 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.055 $Y=1.325
+ $X2=9.055 $Y2=1.16
r60 18 20 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.055 $Y=1.325
+ $X2=9.055 $Y2=2
r61 14 27 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.055 $Y=0.995
+ $X2=9.055 $Y2=1.16
r62 14 16 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=9.055 $Y=0.995
+ $X2=9.055 $Y2=0.51
r63 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.74 $Y=1.985
+ $X2=9.74 $Y2=1.325
r64 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.74 $Y=0.56 $X2=9.74
+ $Y2=0.995
r65 2 20 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=8.93
+ $Y=1.845 $X2=9.055 $Y2=2
r66 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=8.93
+ $Y=0.235 $X2=9.055 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 43 47 53
+ 56 57 58 60 62 68 73 78 86 99 100 103 106 109 116 119 126 129
c180 100 0 1.81794e-19 $X=10.35 $Y=2.72
c181 1 0 3.29888e-20 $X=0.545 $Y=1.815
r182 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r183 127 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r184 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r185 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r186 119 122 10.6812 $w=4.08e-07 $l=3.8e-07 $layer=LI1_cond $X=6.135 $Y=2.34
+ $X2=6.135 $Y2=2.72
r187 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r188 113 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r189 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r190 109 112 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.62 $Y=2.34
+ $X2=3.62 $Y2=2.72
r191 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r192 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r193 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r194 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r195 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r196 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r197 94 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r198 93 96 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r199 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r200 91 129 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.2 $Y=2.72 $X2=8.11
+ $Y2=2.72
r201 91 93 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.2 $Y=2.72
+ $X2=8.51 $Y2=2.72
r202 90 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r203 90 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r204 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r205 87 122 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.135 $Y2=2.72
r206 87 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.67 $Y2=2.72
r207 86 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=7.175 $Y2=2.72
r208 86 89 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=6.67 $Y2=2.72
r209 85 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r210 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r211 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r212 82 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r213 81 84 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r214 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r215 79 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.495 $Y2=2.72
r216 79 81 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.83 $Y2=2.72
r217 78 122 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.93 $Y=2.72
+ $X2=6.135 $Y2=2.72
r218 78 84 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.93 $Y=2.72
+ $X2=5.75 $Y2=2.72
r219 77 113 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r220 77 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r221 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r222 74 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r223 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r224 73 112 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=3.62 $Y2=2.72
r225 73 76 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=2.07 $Y2=2.72
r226 72 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r227 72 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r228 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r229 69 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r230 69 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r231 68 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r232 68 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r233 62 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r234 60 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r235 58 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r236 58 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r237 56 96 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=9.445 $Y=2.72
+ $X2=9.43 $Y2=2.72
r238 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.445 $Y=2.72
+ $X2=9.53 $Y2=2.72
r239 55 99 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=9.615 $Y=2.72
+ $X2=10.35 $Y2=2.72
r240 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.615 $Y=2.72
+ $X2=9.53 $Y2=2.72
r241 51 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.53 $Y=2.635
+ $X2=9.53 $Y2=2.72
r242 51 53 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.53 $Y=2.635
+ $X2=9.53 $Y2=2
r243 47 50 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=8.11 $Y=1.66
+ $X2=8.11 $Y2=2.34
r244 45 129 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=2.635
+ $X2=8.11 $Y2=2.72
r245 45 50 18.1768 $w=1.78e-07 $l=2.95e-07 $layer=LI1_cond $X=8.11 $Y=2.635
+ $X2=8.11 $Y2=2.34
r246 44 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.175 $Y2=2.72
r247 43 129 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.02 $Y=2.72 $X2=8.11
+ $Y2=2.72
r248 43 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.02 $Y=2.72
+ $X2=7.34 $Y2=2.72
r249 39 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.72
r250 39 41 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.21
r251 35 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.72
r252 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.34
r253 34 112 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.81 $Y=2.72
+ $X2=3.62 $Y2=2.72
r254 33 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=4.495 $Y2=2.72
r255 33 34 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=3.81 $Y2=2.72
r256 29 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r257 29 31 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.22
r258 25 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r259 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r260 8 53 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=9.34
+ $Y=1.845 $X2=9.53 $Y2=2
r261 7 50 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=1.485 $X2=8.115 $Y2=2.34
r262 7 47 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=1.485 $X2=8.115 $Y2=1.66
r263 6 41 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=2.065 $X2=7.175 $Y2=2.21
r264 5 119 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.04
+ $Y=2.065 $X2=6.175 $Y2=2.34
r265 4 37 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.065 $X2=4.495 $Y2=2.34
r266 3 109 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.065 $X2=3.595 $Y2=2.34
r267 2 31 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.645 $X2=1.62 $Y2=2.22
r268 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%A_381_47# 1 2 8 9 10 11 12 15 20
c59 20 0 1.34441e-19 $X=2.04 $Y=1.96
r60 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r61 11 20 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.88
r62 11 12 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.6 $Y2=1.88
r63 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r64 9 10 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=1.6 $Y2=0.73
r65 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.795
+ $X2=1.6 $Y2=1.88
r66 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.6 $Y2=0.73
r67 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.515 $Y2=1.795
r68 2 20 300 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.645 $X2=2.04 $Y2=1.96
r69 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%Q_N 1 2 7 8 9 10 11 12 20
r22 12 37 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.535 $Y=2.21
+ $X2=8.535 $Y2=2.34
r23 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=1.87
+ $X2=8.535 $Y2=2.21
r24 11 31 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8.535 $Y=1.87
+ $X2=8.535 $Y2=1.66
r25 10 31 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.535 $Y=1.53
+ $X2=8.535 $Y2=1.66
r26 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=1.19
+ $X2=8.535 $Y2=1.53
r27 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=0.85
+ $X2=8.535 $Y2=1.19
r28 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=0.51
+ $X2=8.535 $Y2=0.85
r29 7 20 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=8.535 $Y=0.51
+ $X2=8.535 $Y2=0.4
r30 2 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.4
+ $Y=1.485 $X2=8.535 $Y2=2.34
r31 2 31 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.4
+ $Y=1.485 $X2=8.535 $Y2=1.66
r32 1 20 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.4
+ $Y=0.235 $X2=8.535 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%Q 1 2 10 11 12 13 14 15
r16 14 15 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=9.995 $Y=1.82
+ $X2=9.995 $Y2=2.21
r17 11 14 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=9.995 $Y=1.575
+ $X2=9.995 $Y2=1.82
r18 11 12 6.14153 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=9.995 $Y=1.575
+ $X2=9.995 $Y2=1.445
r19 10 12 33.2332 $w=2.13e-07 $l=6.2e-07 $layer=LI1_cond $X=10.017 $Y=0.825
+ $X2=10.017 $Y2=1.445
r20 9 13 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=9.995 $Y=0.695
+ $X2=9.995 $Y2=0.51
r21 9 10 6.14153 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=9.995 $Y=0.695
+ $X2=9.995 $Y2=0.825
r22 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=9.815
+ $Y=1.485 $X2=9.95 $Y2=1.82
r23 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=9.815
+ $Y=0.235 $X2=9.95 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 38 42 46 49
+ 50 51 53 55 61 66 74 92 93 96 99 102 105 110 116 118
c163 110 0 1.49785e-19 $X=6.67 $Y=0.24
c164 93 0 1.99443e-19 $X=10.35 $Y=0
r165 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r166 115 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r167 114 116 11.126 $w=6.48e-07 $l=2e-07 $layer=LI1_cond $X=7.13 $Y=0.24
+ $X2=7.33 $Y2=0.24
r168 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r169 112 114 1.01207 $w=6.48e-07 $l=5.5e-08 $layer=LI1_cond $X=7.075 $Y=0.24
+ $X2=7.13 $Y2=0.24
r170 109 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r171 108 112 7.45249 $w=6.48e-07 $l=4.05e-07 $layer=LI1_cond $X=6.67 $Y=0.24
+ $X2=7.075 $Y2=0.24
r172 108 110 7.44573 $w=6.48e-07 $l=4.45988e-08 $layer=LI1_cond $X=6.67 $Y=0.24
+ $X2=6.67 $Y2=0.24
r173 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r174 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r175 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r176 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r177 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r178 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r179 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r180 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r181 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r182 87 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r183 86 89 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r184 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r185 84 118 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.2 $Y=0 $X2=8.11
+ $Y2=0
r186 84 86 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.2 $Y=0 $X2=8.51
+ $Y2=0
r187 83 109 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r188 83 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r189 82 110 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r190 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r191 80 105 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.91
+ $Y2=0
r192 80 82 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.29
+ $Y2=0
r193 78 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r194 78 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r195 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r196 75 102 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.02 $Y=0
+ $X2=3.815 $Y2=0
r197 75 77 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.37
+ $Y2=0
r198 74 105 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.91
+ $Y2=0
r199 74 77 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.37
+ $Y2=0
r200 73 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r201 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r202 70 73 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r203 70 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r204 69 72 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r205 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r206 67 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r207 67 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r208 66 102 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.61 $Y=0
+ $X2=3.815 $Y2=0
r209 66 72 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.45
+ $Y2=0
r210 65 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r211 65 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r212 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r213 62 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r214 62 64 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r215 61 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r216 61 64 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r217 55 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r218 53 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r219 51 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r220 51 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r221 49 89 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=9.445 $Y=0 $X2=9.43
+ $Y2=0
r222 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.445 $Y=0 $X2=9.53
+ $Y2=0
r223 48 92 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=9.615 $Y=0
+ $X2=10.35 $Y2=0
r224 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.615 $Y=0 $X2=9.53
+ $Y2=0
r225 44 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.53 $Y=0.085
+ $X2=9.53 $Y2=0
r226 44 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.53 $Y=0.085
+ $X2=9.53 $Y2=0.38
r227 40 118 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=0.085
+ $X2=8.11 $Y2=0
r228 40 42 19.4091 $w=1.78e-07 $l=3.15e-07 $layer=LI1_cond $X=8.11 $Y=0.085
+ $X2=8.11 $Y2=0.4
r229 38 118 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.02 $Y=0 $X2=8.11
+ $Y2=0
r230 38 116 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.02 $Y=0 $X2=7.33
+ $Y2=0
r231 34 105 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=0.085
+ $X2=4.91 $Y2=0
r232 34 36 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=4.91 $Y=0.085
+ $X2=4.91 $Y2=0.38
r233 30 102 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r234 30 32 7.7298 $w=4.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.36
r235 26 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r236 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.38
r237 22 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r238 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r239 7 46 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=9.34
+ $Y=0.235 $X2=9.53 $Y2=0.38
r240 6 42 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=7.99
+ $Y=0.235 $X2=8.115 $Y2=0.4
r241 5 112 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=6.84
+ $Y=0.235 $X2=7.075 $Y2=0.48
r242 4 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=4.995 $Y2=0.38
r243 3 32 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.235 $X2=3.695 $Y2=0.36
r244 2 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r245 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


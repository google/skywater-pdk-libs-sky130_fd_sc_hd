* File: sky130_fd_sc_hd__nor3_4.pex.spice
* Created: Thu Aug 27 14:32:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR3_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r74 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.6 $Y=1.16 $X2=1.75
+ $Y2=1.16
r75 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.6 $Y=1.16
+ $X2=1.6 $Y2=1.16
r76 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.33 $Y=1.16 $X2=1.6
+ $Y2=1.16
r77 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r78 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=0.58 $Y=1.16
+ $X2=0.91 $Y2=1.16
r79 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.16 $X2=0.58 $Y2=1.16
r80 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.49 $Y=1.16 $X2=0.58
+ $Y2=1.16
r81 29 40 47.7965 $w=2.08e-07 $l=9.05e-07 $layer=LI1_cond $X=0.695 $Y=1.18
+ $X2=1.6 $Y2=1.18
r82 29 35 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=0.695 $Y=1.18
+ $X2=0.58 $Y2=1.18
r83 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r85 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r87 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r89 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r91 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r93 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r95 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r97 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_4%B 1 3 6 8 10 13 15 17 20 24 27 30 31 32 34 35
+ 39 40 42 50 53
r134 48 50 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=2.6 $Y=1.16
+ $X2=3.01 $Y2=1.16
r135 46 48 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.59 $Y=1.16 $X2=2.6
+ $Y2=1.16
r136 44 46 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.17 $Y=1.16
+ $X2=2.59 $Y2=1.16
r137 42 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.6
+ $Y=1.16 $X2=2.6 $Y2=1.16
r138 40 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.16 $Y=1.16
+ $X2=5.16 $Y2=1.325
r139 40 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.16 $Y=1.16
+ $X2=5.16 $Y2=0.995
r140 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.16
+ $Y=1.16 $X2=5.16 $Y2=1.16
r141 36 39 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=5.08 $Y=1.18 $X2=5.16
+ $Y2=1.18
r142 35 42 51.7576 $w=2.08e-07 $l=9.8e-07 $layer=LI1_cond $X=3.515 $Y=1.18
+ $X2=2.535 $Y2=1.18
r143 33 36 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.08 $Y=1.285
+ $X2=5.08 $Y2=1.18
r144 33 34 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.08 $Y=1.285
+ $X2=5.08 $Y2=1.445
r145 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.995 $Y=1.53
+ $X2=5.08 $Y2=1.445
r146 31 32 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=4.995 $Y=1.53
+ $X2=3.685 $Y2=1.53
r147 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.6 $Y=1.445
+ $X2=3.685 $Y2=1.53
r148 29 35 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.6 $Y=1.285
+ $X2=3.515 $Y2=1.18
r149 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.6 $Y=1.285
+ $X2=3.6 $Y2=1.445
r150 27 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.11 $Y=1.985
+ $X2=5.11 $Y2=1.325
r151 24 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.11 $Y=0.56
+ $X2=5.11 $Y2=0.995
r152 18 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.16
r153 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.985
r154 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=1.16
r155 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r156 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.16
r157 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.985
r158 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.16
r159 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r160 4 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.16
r161 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.985
r162 1 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r163 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 37 38
r89 36 38 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.54 $Y=1.16
+ $X2=4.69 $Y2=1.16
r90 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.54
+ $Y=1.16 $X2=4.54 $Y2=1.16
r91 34 36 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.27 $Y=1.16
+ $X2=4.54 $Y2=1.16
r92 33 34 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.85 $Y=1.16
+ $X2=4.27 $Y2=1.16
r93 31 33 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.43 $Y=1.16
+ $X2=3.85 $Y2=1.16
r94 29 37 0.402198 $w=9.08e-07 $l=3e-08 $layer=LI1_cond $X=4.31 $Y=1.19 $X2=4.31
+ $Y2=1.16
r95 25 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.69 $Y2=1.16
r96 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.69 $Y2=1.985
r97 22 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=0.995
+ $X2=4.69 $Y2=1.16
r98 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.69 $Y=0.995
+ $X2=4.69 $Y2=0.56
r99 18 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.325
+ $X2=4.27 $Y2=1.16
r100 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.27 $Y=1.325
+ $X2=4.27 $Y2=1.985
r101 15 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=0.995
+ $X2=4.27 $Y2=1.16
r102 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.27 $Y=0.995
+ $X2=4.27 $Y2=0.56
r103 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=1.325
+ $X2=3.85 $Y2=1.16
r104 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.85 $Y=1.325
+ $X2=3.85 $Y2=1.985
r105 8 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=0.995
+ $X2=3.85 $Y2=1.16
r106 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.85 $Y=0.995
+ $X2=3.85 $Y2=0.56
r107 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.16
r108 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.985
r109 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.16
r110 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 32 37 43 52 54 55 56
c93 56 0 1.98853e-19 $X=5.145 $Y=2.2
r94 54 56 0.113326 $w=2.7e-07 $l=1.45e-07 $layer=MET1_cond $X=5.29 $Y=2.2
+ $X2=5.145 $Y2=2.2
r95 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.21
+ $X2=5.29 $Y2=2.21
r96 52 56 3.05074 $w=1.4e-07 $l=2.465e-06 $layer=MET1_cond $X=2.68 $Y=2.21
+ $X2=5.145 $Y2=2.21
r97 49 52 0.116059 $w=2.7e-07 $l=1.5e-07 $layer=MET1_cond $X=2.53 $Y=2.2
+ $X2=2.68 $Y2=2.2
r98 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.21
+ $X2=2.53 $Y2=2.21
r99 43 50 4.39748 $w=3.78e-07 $l=1.45e-07 $layer=LI1_cond $X=2.675 $Y=2.275
+ $X2=2.53 $Y2=2.275
r100 43 45 2.85751 $w=3.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.675 $Y=2.275
+ $X2=2.8 $Y2=2.275
r101 40 50 13.4957 $w=3.78e-07 $l=4.45e-07 $layer=LI1_cond $X=2.085 $Y=2.275
+ $X2=2.53 $Y2=2.275
r102 40 42 2.85751 $w=3.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=2.275
+ $X2=1.96 $Y2=2.275
r103 30 45 4.34342 $w=2.5e-07 $l=1.9e-07 $layer=LI1_cond $X=2.8 $Y=2.085 $X2=2.8
+ $Y2=2.275
r104 30 32 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.8 $Y=2.085
+ $X2=2.8 $Y2=1.96
r105 29 42 4.34342 $w=2.5e-07 $l=1.9e-07 $layer=LI1_cond $X=1.96 $Y=2.085
+ $X2=1.96 $Y2=2.275
r106 28 39 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=1.625
+ $X2=1.96 $Y2=1.54
r107 28 29 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.96 $Y=1.625
+ $X2=1.96 $Y2=2.085
r108 27 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=1.54
+ $X2=1.12 $Y2=1.54
r109 26 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.96 $Y2=1.54
r110 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=1.54
+ $X2=1.245 $Y2=1.54
r111 22 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=1.54
r112 22 24 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.12 $Y=1.625
+ $X2=1.12 $Y2=2.3
r113 21 35 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r114 20 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=1.12 $Y2=1.54
r115 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.54
+ $X2=0.405 $Y2=1.54
r116 16 35 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r117 16 18 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r118 5 55 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.485 $X2=5.32 $Y2=2.3
r119 4 45 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=2.3
r120 4 32 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=1.96
r121 3 42 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.3
r122 3 39 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r123 2 37 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r124 2 24 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r125 1 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r126 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_4%VPWR 1 2 9 13 15 17 22 29 30 33 36
r83 36 37 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r84 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r85 30 37 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=2.72 $X2=1.61
+ $Y2=2.72
r86 29 30 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r87 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.54 $Y2=2.72
r88 27 29 266.508 $w=1.68e-07 $l=4.085e-06 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=5.75 $Y2=2.72
r89 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r90 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r92 23 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r93 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 22 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.54 $Y2=2.72
r95 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.15 $Y2=2.72
r96 17 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r97 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r98 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r99 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r100 11 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2.72
r101 11 13 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=1.96
r102 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r103 7 9 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=1.96
r104 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.96
r105 1 9 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_4%A_449_297# 1 2 3 4 15 17 18 19 21 24 30 35
c65 3 0 1.98853e-19 $X=3.925 $Y=1.485
r66 35 37 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.9 $Y=2.3 $X2=4.9
+ $Y2=2.38
r67 30 32 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.06 $Y=2.3 $X2=4.06
+ $Y2=2.38
r68 22 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=2.38
+ $X2=4.06 $Y2=2.38
r69 21 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.775 $Y=2.38
+ $X2=4.9 $Y2=2.38
r70 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.775 $Y=2.38
+ $X2=4.185 $Y2=2.38
r71 20 28 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=2.38
+ $X2=3.22 $Y2=2.38
r72 19 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.935 $Y=2.38
+ $X2=4.06 $Y2=2.38
r73 19 20 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.935 $Y=2.38
+ $X2=3.345 $Y2=2.38
r74 18 28 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.295
+ $X2=3.22 $Y2=2.38
r75 17 26 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=1.625
+ $X2=3.22 $Y2=1.54
r76 17 18 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.22 $Y=1.625
+ $X2=3.22 $Y2=2.295
r77 16 24 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=1.54
+ $X2=2.38 $Y2=1.54
r78 15 26 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=1.54
+ $X2=3.22 $Y2=1.54
r79 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.095 $Y=1.54
+ $X2=2.505 $Y2=1.54
r80 4 35 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=1.485 $X2=4.9 $Y2=2.3
r81 3 30 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.06 $Y2=2.3
r82 2 28 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=2.3
r83 2 26 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.62
r84 1 24 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_4%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 41 45 47
+ 49 53 55 57 61 63 69 70 71 72 77 78 84 86 88 89
r194 87 89 10.1336 $w=2.88e-07 $l=2.55e-07 $layer=LI1_cond $X=5.75 $Y=1.785
+ $X2=5.75 $Y2=1.53
r195 87 88 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.75 $Y=1.785
+ $X2=5.75 $Y2=1.87
r196 85 89 24.8371 $w=2.88e-07 $l=6.25e-07 $layer=LI1_cond $X=5.75 $Y=0.905
+ $X2=5.75 $Y2=1.53
r197 85 86 3.41797 $w=2.9e-07 $l=9e-08 $layer=LI1_cond $X=5.75 $Y=0.905 $X2=5.75
+ $Y2=0.815
r198 80 82 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=1.875
+ $X2=4.48 $Y2=1.96
r199 78 80 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.48 $Y=1.87
+ $X2=4.48 $Y2=1.875
r200 72 75 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=1.875
+ $X2=3.64 $Y2=1.96
r201 64 84 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=0.815
+ $X2=4.9 $Y2=0.815
r202 63 86 3.10432 $w=1.8e-07 $l=1.45e-07 $layer=LI1_cond $X=5.605 $Y=0.815
+ $X2=5.75 $Y2=0.815
r203 63 64 33.2727 $w=1.78e-07 $l=5.4e-07 $layer=LI1_cond $X=5.605 $Y=0.815
+ $X2=5.065 $Y2=0.815
r204 59 84 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.9 $Y=0.725 $X2=4.9
+ $Y2=0.815
r205 59 61 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.9 $Y=0.725
+ $X2=4.9 $Y2=0.39
r206 58 78 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.605 $Y=1.87
+ $X2=4.48 $Y2=1.87
r207 57 88 3.25423 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.605 $Y=1.87
+ $X2=5.75 $Y2=1.87
r208 57 58 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=5.605 $Y=1.87
+ $X2=4.605 $Y2=1.87
r209 56 77 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.225 $Y=0.815
+ $X2=4.06 $Y2=0.815
r210 55 84 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=0.815
+ $X2=4.9 $Y2=0.815
r211 55 56 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.735 $Y=0.815
+ $X2=4.225 $Y2=0.815
r212 51 77 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.06 $Y=0.725
+ $X2=4.06 $Y2=0.815
r213 51 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.06 $Y=0.725
+ $X2=4.06 $Y2=0.39
r214 50 72 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.765 $Y=1.875
+ $X2=3.64 $Y2=1.875
r215 49 80 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.355 $Y=1.875
+ $X2=4.48 $Y2=1.875
r216 49 50 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=4.355 $Y=1.875
+ $X2=3.765 $Y2=1.875
r217 48 71 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.815
+ $X2=3.22 $Y2=0.815
r218 47 77 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=0.815
+ $X2=4.06 $Y2=0.815
r219 47 48 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.895 $Y=0.815
+ $X2=3.385 $Y2=0.815
r220 43 71 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.815
r221 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.39
r222 42 70 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0.815
+ $X2=2.38 $Y2=0.815
r223 41 71 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=3.22 $Y2=0.815
r224 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=2.545 $Y2=0.815
r225 37 70 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.815
r226 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.39
r227 36 69 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r228 35 70 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=2.38 $Y2=0.815
r229 35 36 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=1.705 $Y2=0.815
r230 31 69 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.815
r231 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r232 29 69 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r233 29 30 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r234 25 30 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r235 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.7 $Y2=0.39
r236 8 82 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.48 $Y2=1.96
r237 7 75 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=1.96
r238 6 61 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.765
+ $Y=0.235 $X2=4.9 $Y2=0.39
r239 5 53 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.925
+ $Y=0.235 $X2=4.06 $Y2=0.39
r240 4 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.39
r241 3 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.39
r242 2 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r243 1 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46 50
+ 53 54 56 57 59 60 62 63 64 65 66 86 87 93
r111 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r112 87 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r113 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r114 84 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=0 $X2=5.32
+ $Y2=0
r115 84 86 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.405 $Y=0 $X2=5.75
+ $Y2=0
r116 83 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r117 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r118 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r119 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r120 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r121 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r122 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r123 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r124 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r125 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r126 68 90 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r127 68 70 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.69 $Y2=0
r128 66 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r129 66 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r130 64 82 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.37
+ $Y2=0
r131 64 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.48
+ $Y2=0
r132 62 79 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.45 $Y2=0
r133 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.64
+ $Y2=0
r134 61 82 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.725 $Y=0
+ $X2=4.37 $Y2=0
r135 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0 $X2=3.64
+ $Y2=0
r136 59 76 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0
+ $X2=2.53 $Y2=0
r137 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.8
+ $Y2=0
r138 58 79 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.45
+ $Y2=0
r139 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.8
+ $Y2=0
r140 56 73 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r141 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r142 55 76 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.53 $Y2=0
r143 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r144 53 70 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r145 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r146 52 73 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.61 $Y2=0
r147 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r148 48 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.32 $Y=0.085
+ $X2=5.32 $Y2=0
r149 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.32 $Y=0.085
+ $X2=5.32 $Y2=0.39
r150 47 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0 $X2=4.48
+ $Y2=0
r151 46 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.32
+ $Y2=0
r152 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.235 $Y=0
+ $X2=4.565 $Y2=0
r153 42 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0
r154 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0.39
r155 38 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0
r156 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0.39
r157 34 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r158 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.39
r159 30 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r160 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r161 26 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r162 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r163 22 90 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r164 22 24 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r165 7 50 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.185
+ $Y=0.235 $X2=5.32 $Y2=0.39
r166 6 44 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.345
+ $Y=0.235 $X2=4.48 $Y2=0.39
r167 5 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.39
r168 4 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.39
r169 3 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r170 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r171 1 24 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__a32o_4.spice.SKY130_FD_SC_HD__A32O_4.pxi
* Created: Thu Aug 27 14:05:31 2020
* 
x_PM_SKY130_FD_SC_HD__A32O_4%A_79_21# N_A_79_21#_M1010_d N_A_79_21#_M1005_d
+ N_A_79_21#_M1007_d N_A_79_21#_M1013_s N_A_79_21#_c_104_n N_A_79_21#_M1009_g
+ N_A_79_21#_M1000_g N_A_79_21#_c_105_n N_A_79_21#_M1015_g N_A_79_21#_M1001_g
+ N_A_79_21#_c_106_n N_A_79_21#_M1016_g N_A_79_21#_M1017_g N_A_79_21#_c_107_n
+ N_A_79_21#_M1026_g N_A_79_21#_M1025_g N_A_79_21#_c_108_n N_A_79_21#_c_118_n
+ N_A_79_21#_c_119_n N_A_79_21#_c_175_p N_A_79_21#_c_109_n N_A_79_21#_c_110_n
+ N_A_79_21#_c_142_p N_A_79_21#_c_143_p N_A_79_21#_c_157_p N_A_79_21#_c_111_n
+ N_A_79_21#_c_153_p N_A_79_21#_c_154_p N_A_79_21#_c_155_p N_A_79_21#_c_112_n
+ PM_SKY130_FD_SC_HD__A32O_4%A_79_21#
x_PM_SKY130_FD_SC_HD__A32O_4%A3 N_A3_c_270_n N_A3_M1019_g N_A3_M1002_g
+ N_A3_c_271_n N_A3_M1024_g N_A3_M1021_g A3 A3 N_A3_c_273_n
+ PM_SKY130_FD_SC_HD__A32O_4%A3
x_PM_SKY130_FD_SC_HD__A32O_4%A2 N_A2_c_314_n N_A2_M1003_g N_A2_M1014_g
+ N_A2_c_315_n N_A2_M1004_g N_A2_M1023_g A2 A2 N_A2_c_317_n
+ PM_SKY130_FD_SC_HD__A32O_4%A2
x_PM_SKY130_FD_SC_HD__A32O_4%A1 N_A1_M1010_g N_A1_M1006_g N_A1_M1020_g
+ N_A1_M1008_g A1 A1 N_A1_c_362_n PM_SKY130_FD_SC_HD__A32O_4%A1
x_PM_SKY130_FD_SC_HD__A32O_4%B1 N_B1_M1005_g N_B1_M1007_g N_B1_M1011_g
+ N_B1_M1027_g B1 B1 B1 N_B1_c_406_n PM_SKY130_FD_SC_HD__A32O_4%B1
x_PM_SKY130_FD_SC_HD__A32O_4%B2 N_B2_M1012_g N_B2_M1013_g N_B2_M1022_g
+ N_B2_M1018_g B2 B2 B2 N_B2_c_457_n N_B2_c_473_n PM_SKY130_FD_SC_HD__A32O_4%B2
x_PM_SKY130_FD_SC_HD__A32O_4%VPWR N_VPWR_M1000_s N_VPWR_M1001_s N_VPWR_M1025_s
+ N_VPWR_M1021_d N_VPWR_M1014_s N_VPWR_M1006_s N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n
+ N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n VPWR N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_493_n N_VPWR_c_512_n PM_SKY130_FD_SC_HD__A32O_4%VPWR
x_PM_SKY130_FD_SC_HD__A32O_4%X N_X_M1009_s N_X_M1016_s N_X_M1000_d N_X_M1017_d
+ N_X_c_619_n N_X_c_620_n N_X_c_655_p N_X_c_638_n N_X_c_621_n N_X_c_625_n
+ N_X_c_653_p N_X_c_642_n N_X_c_629_n N_X_c_631_n X X X N_X_c_615_n N_X_c_617_n
+ X PM_SKY130_FD_SC_HD__A32O_4%X
x_PM_SKY130_FD_SC_HD__A32O_4%A_445_297# N_A_445_297#_M1002_s
+ N_A_445_297#_M1014_d N_A_445_297#_M1023_d N_A_445_297#_M1008_d
+ N_A_445_297#_M1027_s N_A_445_297#_M1018_d N_A_445_297#_c_710_n
+ N_A_445_297#_c_664_n N_A_445_297#_c_678_n N_A_445_297#_c_691_n
+ N_A_445_297#_c_679_n N_A_445_297#_c_725_n N_A_445_297#_c_680_n
+ N_A_445_297#_c_682_n N_A_445_297#_c_734_n N_A_445_297#_c_665_n
+ N_A_445_297#_c_666_n N_A_445_297#_c_688_n N_A_445_297#_c_689_n
+ PM_SKY130_FD_SC_HD__A32O_4%A_445_297#
x_PM_SKY130_FD_SC_HD__A32O_4%VGND N_VGND_M1009_d N_VGND_M1015_d N_VGND_M1026_d
+ N_VGND_M1024_d N_VGND_M1012_d N_VGND_c_738_n N_VGND_c_739_n N_VGND_c_740_n
+ N_VGND_c_741_n N_VGND_c_742_n N_VGND_c_743_n N_VGND_c_744_n N_VGND_c_745_n
+ N_VGND_c_746_n N_VGND_c_747_n VGND N_VGND_c_748_n N_VGND_c_749_n
+ N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n N_VGND_c_753_n
+ PM_SKY130_FD_SC_HD__A32O_4%VGND
x_PM_SKY130_FD_SC_HD__A32O_4%A_445_47# N_A_445_47#_M1019_s N_A_445_47#_M1003_s
+ N_A_445_47#_c_865_n N_A_445_47#_c_853_n N_A_445_47#_c_850_n
+ PM_SKY130_FD_SC_HD__A32O_4%A_445_47#
x_PM_SKY130_FD_SC_HD__A32O_4%A_635_47# N_A_635_47#_M1003_d N_A_635_47#_M1004_d
+ N_A_635_47#_M1020_s N_A_635_47#_c_875_n PM_SKY130_FD_SC_HD__A32O_4%A_635_47#
x_PM_SKY130_FD_SC_HD__A32O_4%A_1142_47# N_A_1142_47#_M1005_s
+ N_A_1142_47#_M1011_s N_A_1142_47#_M1022_s N_A_1142_47#_c_895_n
+ N_A_1142_47#_c_917_n N_A_1142_47#_c_899_n N_A_1142_47#_c_907_n
+ N_A_1142_47#_c_900_n N_A_1142_47#_c_924_n
+ PM_SKY130_FD_SC_HD__A32O_4%A_1142_47#
cc_1 VNB N_A_79_21#_c_104_n 0.0182736f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_105_n 0.0157735f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_106_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_107_n 0.0159773f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_108_n 0.00499804f $X=-0.19 $Y=-0.24 $X2=1.8 $Y2=1.16
cc_6 VNB N_A_79_21#_c_109_n 0.00911532f $X=-0.19 $Y=-0.24 $X2=5.28 $Y2=0.72
cc_7 VNB N_A_79_21#_c_110_n 0.0133347f $X=-0.19 $Y=-0.24 $X2=5.365 $Y2=1.495
cc_8 VNB N_A_79_21#_c_111_n 0.0155981f $X=-0.19 $Y=-0.24 $X2=6.255 $Y2=0.72
cc_9 VNB N_A_79_21#_c_112_n 0.0647252f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_10 VNB N_A3_c_270_n 0.0159773f $X=-0.19 $Y=-0.24 $X2=4.425 $Y2=0.235
cc_11 VNB N_A3_c_271_n 0.0210871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A3 0.00646996f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_13 VNB N_A3_c_273_n 0.047138f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_14 VNB N_A2_c_314_n 0.0219813f $X=-0.19 $Y=-0.24 $X2=4.425 $Y2=0.235
cc_15 VNB N_A2_c_315_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB A2 0.00392777f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_17 VNB N_A2_c_317_n 0.0406958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_M1010_g 0.017802f $X=-0.19 $Y=-0.24 $X2=6.165 $Y2=1.485
cc_19 VNB N_A1_M1020_g 0.0209838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB A1 0.00229759f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_21 VNB N_A1_c_362_n 0.045811f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_22 VNB N_B1_M1005_g 0.0218177f $X=-0.19 $Y=-0.24 $X2=6.165 $Y2=1.485
cc_23 VNB N_B1_M1011_g 0.0182654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB B1 0.00990395f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_25 VNB N_B1_c_406_n 0.0400083f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_26 VNB N_B2_M1012_g 0.0180382f $X=-0.19 $Y=-0.24 $X2=6.165 $Y2=1.485
cc_27 VNB N_B2_M1022_g 0.0233553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB B2 0.00887859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_B2_c_457_n 0.0524594f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_30 VNB N_VPWR_c_493_n 0.326667f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_31 VNB N_X_c_615_n 0.0071443f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.16
cc_32 VNB X 0.0236638f $X=-0.19 $Y=-0.24 $X2=1.885 $Y2=1.495
cc_33 VNB N_VGND_c_738_n 0.010303f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_34 VNB N_VGND_c_739_n 0.0125988f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_35 VNB N_VGND_c_740_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_36 VNB N_VGND_c_741_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_742_n 0.00552505f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_38 VNB N_VGND_c_743_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_39 VNB N_VGND_c_744_n 0.0117278f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_40 VNB N_VGND_c_745_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_41 VNB N_VGND_c_746_n 0.0117571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_747_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=1.8 $Y2=1.16
cc_43 VNB N_VGND_c_748_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_44 VNB N_VGND_c_749_n 0.0958249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_750_n 0.0151555f $X=-0.19 $Y=-0.24 $X2=6.3 $Y2=2
cc_46 VNB N_VGND_c_751_n 0.381807f $X=-0.19 $Y=-0.24 $X2=7.14 $Y2=2
cc_47 VNB N_VGND_c_752_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_753_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=6.2 $Y2=1.995
cc_49 VNB N_A_445_47#_c_850_n 0.00815884f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_50 VNB N_A_635_47#_c_875_n 0.00569209f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_51 VNB N_A_1142_47#_c_895_n 0.00348834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VPB N_A_79_21#_M1000_g 0.0209859f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_53 VPB N_A_79_21#_M1001_g 0.0182726f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_54 VPB N_A_79_21#_M1017_g 0.0182693f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_55 VPB N_A_79_21#_M1025_g 0.0176229f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_56 VPB N_A_79_21#_c_108_n 2.19146e-19 $X=-0.19 $Y=1.305 $X2=1.8 $Y2=1.16
cc_57 VPB N_A_79_21#_c_118_n 0.00147022f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=1.495
cc_58 VPB N_A_79_21#_c_119_n 0.00765505f $X=-0.19 $Y=1.305 $X2=5.28 $Y2=1.58
cc_59 VPB N_A_79_21#_c_110_n 0.00455514f $X=-0.19 $Y=1.305 $X2=5.365 $Y2=1.495
cc_60 VPB N_A_79_21#_c_112_n 0.0102726f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_61 VPB N_A3_M1002_g 0.0185179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A3_M1021_g 0.0250853f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_63 VPB N_A3_c_273_n 0.0102564f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_64 VPB N_A2_M1014_g 0.0241559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A2_M1023_g 0.0175748f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_66 VPB A2 0.00161583f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_67 VPB N_A2_c_317_n 0.00691477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A1_M1006_g 0.0175748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A1_M1008_g 0.0213557f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_70 VPB A1 0.00231767f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_71 VPB N_A1_c_362_n 0.0131097f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_72 VPB N_B1_M1007_g 0.0223275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B1_M1027_g 0.0172006f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_74 VPB B1 0.00377203f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_75 VPB N_B1_c_406_n 0.00460987f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_76 VPB N_B2_M1013_g 0.0187391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_B2_M1018_g 0.0259373f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_78 VPB B2 0.00250551f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_79 VPB N_B2_c_457_n 0.0146286f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_80 VPB N_VPWR_c_494_n 0.0103102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_495_n 0.0257969f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_82 VPB N_VPWR_c_496_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_83 VPB N_VPWR_c_497_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_84 VPB N_VPWR_c_498_n 0.00479212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_499_n 3.18775e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_86 VPB N_VPWR_c_500_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.8 $Y2=1.16
cc_87 VPB N_VPWR_c_501_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_88 VPB N_VPWR_c_502_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_503_n 0.0117278f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_90 VPB N_VPWR_c_504_n 0.00507168f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_91 VPB N_VPWR_c_505_n 0.0147489f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=1.495
cc_92 VPB N_VPWR_c_506_n 0.00436154f $X=-0.19 $Y=1.305 $X2=5.28 $Y2=1.58
cc_93 VPB N_VPWR_c_507_n 0.0109642f $X=-0.19 $Y=1.305 $X2=5.28 $Y2=0.72
cc_94 VPB N_VPWR_c_508_n 0.00436154f $X=-0.19 $Y=1.305 $X2=4.56 $Y2=0.72
cc_95 VPB N_VPWR_c_509_n 0.0124915f $X=-0.19 $Y=1.305 $X2=5.365 $Y2=0.805
cc_96 VPB N_VPWR_c_510_n 0.074246f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_97 VPB N_VPWR_c_493_n 0.047947f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_98 VPB N_VPWR_c_512_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_X_c_617_n 0.00716948f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_100 VPB X 0.00899487f $X=-0.19 $Y=1.305 $X2=1.885 $Y2=1.495
cc_101 VPB N_A_445_297#_c_664_n 0.00782002f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_102 VPB N_A_445_297#_c_665_n 0.00747984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_445_297#_c_666_n 0.0195224f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.16
cc_104 N_A_79_21#_c_107_n N_A3_c_270_n 0.0232192f $X=1.73 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_79_21#_M1025_g N_A3_M1002_g 0.0232192f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_118_n N_A3_M1002_g 0.00374792f $X=1.885 $Y=1.495 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_119_n N_A3_M1002_g 0.0182499f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_119_n N_A3_M1021_g 0.0131218f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_108_n A3 0.0149831f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_119_n A3 0.0517887f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_108_n N_A3_c_273_n 0.00567593f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_119_n N_A3_c_273_n 0.0070684f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_112_n N_A3_c_273_n 0.0232192f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_119_n N_A2_M1014_g 0.0129401f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_109_n N_A2_c_315_n 5.30585e-19 $X=5.28 $Y=0.72 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_119_n N_A2_M1023_g 0.0107929f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_119_n A2 0.0428809f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_119_n N_A2_c_317_n 0.00262383f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_109_n N_A1_M1010_g 0.00388163f $X=5.28 $Y=0.72 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_119_n N_A1_M1006_g 0.0109456f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_109_n N_A1_M1020_g 0.0110355f $X=5.28 $Y=0.72 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_110_n N_A1_M1020_g 0.00542314f $X=5.365 $Y=1.495 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_119_n N_A1_M1008_g 0.0128075f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_142_p N_A1_M1008_g 0.00618626f $X=5.365 $Y=1.905 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_143_p N_A1_M1008_g 0.00110818f $X=5.45 $Y=1.99 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_119_n A1 0.0514443f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_109_n A1 0.0295632f $X=5.28 $Y=0.72 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_110_n A1 0.0172865f $X=5.365 $Y=1.495 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_119_n N_A1_c_362_n 0.00346913f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_109_n N_A1_c_362_n 0.00684703f $X=5.28 $Y=0.72 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_110_n N_A1_c_362_n 0.00851252f $X=5.365 $Y=1.495 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_110_n N_B1_M1005_g 0.00521041f $X=5.365 $Y=1.495 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_111_n N_B1_M1005_g 0.0110355f $X=6.255 $Y=0.72 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_142_p N_B1_M1007_g 0.00542196f $X=5.365 $Y=1.905 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_153_p N_B1_M1007_g 0.00158666f $X=5.365 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_154_p N_B1_M1007_g 0.00971969f $X=6.135 $Y=1.995 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_155_p N_B1_M1007_g 0.00180292f $X=6.2 $Y=1.995 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_111_n N_B1_M1011_g 0.00303024f $X=6.255 $Y=0.72 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_157_p N_B1_M1027_g 0.00899492f $X=7.14 $Y=2 $X2=0 $Y2=0
cc_140 N_A_79_21#_M1007_d B1 0.00220353f $X=6.165 $Y=1.485 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_110_n B1 0.0339162f $X=5.365 $Y=1.495 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_157_p B1 0.0230654f $X=7.14 $Y=2 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_111_n B1 0.0393341f $X=6.255 $Y=0.72 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_153_p B1 0.0111411f $X=5.365 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_154_p B1 0.0255414f $X=6.135 $Y=1.995 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_110_n N_B1_c_406_n 0.00298573f $X=5.365 $Y=1.495 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_157_p N_B1_c_406_n 3.26393e-19 $X=7.14 $Y=2 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_111_n N_B1_c_406_n 0.00214736f $X=6.255 $Y=0.72 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_154_p N_B1_c_406_n 2.56482e-19 $X=6.135 $Y=1.995 $X2=0 $Y2=0
cc_150 N_A_79_21#_c_157_p N_B2_M1013_g 0.0128635f $X=7.14 $Y=2 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_157_p N_B2_M1018_g 0.00305176f $X=7.14 $Y=2 $X2=0 $Y2=0
cc_152 N_A_79_21#_M1013_s B2 0.00328554f $X=7.005 $Y=1.485 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_157_p B2 0.00863901f $X=7.14 $Y=2 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_157_p B2 0.00128826f $X=7.14 $Y=2 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_157_p N_B2_c_457_n 3.23036e-19 $X=7.14 $Y=2 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_119_n N_VPWR_M1025_s 0.00238703f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_175_p N_VPWR_M1025_s 0.00140883f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_119_n N_VPWR_M1021_d 0.00519517f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_119_n N_VPWR_M1014_s 0.00342606f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A_79_21#_c_119_n N_VPWR_M1006_s 0.00342606f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_161 N_A_79_21#_M1000_g N_VPWR_c_495_n 0.0113889f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_79_21#_M1001_g N_VPWR_c_495_n 6.0901e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_79_21#_M1000_g N_VPWR_c_496_n 6.0901e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_79_21#_M1001_g N_VPWR_c_496_n 0.0102874f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_79_21#_M1017_g N_VPWR_c_496_n 0.0102874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_79_21#_M1025_g N_VPWR_c_496_n 6.0901e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_79_21#_M1017_g N_VPWR_c_497_n 6.0901e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_79_21#_M1025_g N_VPWR_c_497_n 0.0104458f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_108_n N_VPWR_c_497_n 6.69973e-19 $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_119_n N_VPWR_c_497_n 0.0044972f $X=5.28 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A_79_21#_c_175_p N_VPWR_c_497_n 0.00754369f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A_79_21#_M1017_g N_VPWR_c_501_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_79_21#_M1025_g N_VPWR_c_501_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_79_21#_M1000_g N_VPWR_c_509_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_79_21#_M1001_g N_VPWR_c_509_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_79_21#_M1007_d N_VPWR_c_493_n 0.00219239f $X=6.165 $Y=1.485 $X2=0
+ $Y2=0
cc_177 N_A_79_21#_M1013_s N_VPWR_c_493_n 0.00219239f $X=7.005 $Y=1.485 $X2=0
+ $Y2=0
cc_178 N_A_79_21#_M1000_g N_VPWR_c_493_n 0.00789179f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_79_21#_M1001_g N_VPWR_c_493_n 0.00789179f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_79_21#_M1017_g N_VPWR_c_493_n 0.00789179f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_79_21#_M1025_g N_VPWR_c_493_n 0.00789179f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_79_21#_c_104_n N_X_c_619_n 0.0174029f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_79_21#_M1000_g N_X_c_620_n 0.0201041f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_79_21#_c_105_n N_X_c_621_n 0.0114852f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_79_21#_c_106_n N_X_c_621_n 0.0110971f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_79_21#_c_108_n N_X_c_621_n 0.049617f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_79_21#_c_112_n N_X_c_621_n 0.00405004f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_79_21#_M1001_g N_X_c_625_n 0.0140645f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_79_21#_M1017_g N_X_c_625_n 0.0136764f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_108_n N_X_c_625_n 0.0543828f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_112_n N_X_c_625_n 0.00411446f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_108_n N_X_c_629_n 0.0121035f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_112_n N_X_c_629_n 0.00205824f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_79_21#_c_108_n N_X_c_631_n 0.0134105f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_112_n N_X_c_631_n 0.00209661f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_104_n X 0.0227969f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_79_21#_c_108_n X 0.0212528f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_79_21#_c_119_n N_A_445_297#_M1002_s 0.00352632f $X=5.28 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_199 N_A_79_21#_c_119_n N_A_445_297#_M1014_d 0.00704963f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_200 N_A_79_21#_c_119_n N_A_445_297#_M1023_d 0.0079229f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_201 N_A_79_21#_c_119_n N_A_445_297#_M1008_d 0.017885f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_202 N_A_79_21#_c_110_n N_A_445_297#_M1008_d 3.03179e-19 $X=5.365 $Y=1.495
+ $X2=0 $Y2=0
cc_203 N_A_79_21#_c_142_p N_A_445_297#_M1008_d 0.00954918f $X=5.365 $Y=1.905
+ $X2=0 $Y2=0
cc_204 N_A_79_21#_c_143_p N_A_445_297#_M1008_d 0.00529247f $X=5.45 $Y=1.99 $X2=0
+ $Y2=0
cc_205 N_A_79_21#_c_153_p N_A_445_297#_M1008_d 0.00371171f $X=5.365 $Y=1.58
+ $X2=0 $Y2=0
cc_206 N_A_79_21#_c_154_p N_A_445_297#_M1008_d 0.0200581f $X=6.135 $Y=1.995
+ $X2=0 $Y2=0
cc_207 N_A_79_21#_c_157_p N_A_445_297#_M1027_s 0.00416331f $X=7.14 $Y=2 $X2=0
+ $Y2=0
cc_208 N_A_79_21#_c_119_n N_A_445_297#_c_664_n 0.036268f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_209 N_A_79_21#_c_119_n N_A_445_297#_c_678_n 0.0093748f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_210 N_A_79_21#_c_119_n N_A_445_297#_c_679_n 0.0234696f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_211 N_A_79_21#_c_119_n N_A_445_297#_c_680_n 0.0332057f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_212 N_A_79_21#_c_143_p N_A_445_297#_c_680_n 0.0121023f $X=5.45 $Y=1.99 $X2=0
+ $Y2=0
cc_213 N_A_79_21#_M1007_d N_A_445_297#_c_682_n 0.00325828f $X=6.165 $Y=1.485
+ $X2=0 $Y2=0
cc_214 N_A_79_21#_M1013_s N_A_445_297#_c_682_n 0.00325828f $X=7.005 $Y=1.485
+ $X2=0 $Y2=0
cc_215 N_A_79_21#_c_119_n N_A_445_297#_c_682_n 0.00613779f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_216 N_A_79_21#_c_143_p N_A_445_297#_c_682_n 0.0123638f $X=5.45 $Y=1.99 $X2=0
+ $Y2=0
cc_217 N_A_79_21#_c_154_p N_A_445_297#_c_682_n 0.0406236f $X=6.135 $Y=1.995
+ $X2=0 $Y2=0
cc_218 N_A_79_21#_c_155_p N_A_445_297#_c_682_n 0.0552336f $X=6.2 $Y=1.995 $X2=0
+ $Y2=0
cc_219 N_A_79_21#_c_119_n N_A_445_297#_c_688_n 0.00979651f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_220 N_A_79_21#_c_119_n N_A_445_297#_c_689_n 0.0093748f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_221 N_A_79_21#_c_104_n N_VGND_c_739_n 0.00774571f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_79_21#_c_105_n N_VGND_c_739_n 5.08801e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_79_21#_c_104_n N_VGND_c_740_n 5.08801e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_79_21#_c_105_n N_VGND_c_740_n 0.00664421f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_c_106_n N_VGND_c_740_n 0.00664421f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_79_21#_c_107_n N_VGND_c_740_n 5.08801e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_79_21#_c_106_n N_VGND_c_741_n 5.08801e-19 $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_79_21#_c_107_n N_VGND_c_741_n 0.00685487f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_229 N_A_79_21#_c_108_n N_VGND_c_741_n 0.00637759f $X=1.8 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_79_21#_c_106_n N_VGND_c_744_n 0.00339367f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_79_21#_c_107_n N_VGND_c_744_n 0.0046653f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_79_21#_c_104_n N_VGND_c_748_n 0.00339367f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_79_21#_c_105_n N_VGND_c_748_n 0.00339367f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_c_109_n N_VGND_c_749_n 0.00958638f $X=5.28 $Y=0.72 $X2=0 $Y2=0
cc_235 N_A_79_21#_M1010_d N_VGND_c_751_n 0.00219239f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_M1005_d N_VGND_c_751_n 0.00219239f $X=6.12 $Y=0.235 $X2=0
+ $Y2=0
cc_237 N_A_79_21#_c_104_n N_VGND_c_751_n 0.00394406f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_79_21#_c_105_n N_VGND_c_751_n 0.00394406f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_79_21#_c_106_n N_VGND_c_751_n 0.00394406f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_79_21#_c_107_n N_VGND_c_751_n 0.00789179f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_79_21#_c_109_n N_VGND_c_751_n 0.0176492f $X=5.28 $Y=0.72 $X2=0 $Y2=0
cc_242 N_A_79_21#_c_119_n N_A_445_47#_c_850_n 0.00615854f $X=5.28 $Y=1.58 $X2=0
+ $Y2=0
cc_243 N_A_79_21#_c_109_n N_A_445_47#_c_850_n 0.00507639f $X=5.28 $Y=0.72 $X2=0
+ $Y2=0
cc_244 N_A_79_21#_c_109_n N_A_635_47#_M1020_s 0.00573919f $X=5.28 $Y=0.72 $X2=0
+ $Y2=0
cc_245 N_A_79_21#_M1010_d N_A_635_47#_c_875_n 0.0031669f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_246 N_A_79_21#_c_109_n N_A_635_47#_c_875_n 0.0390874f $X=5.28 $Y=0.72 $X2=0
+ $Y2=0
cc_247 N_A_79_21#_c_111_n N_A_1142_47#_M1005_s 0.00549112f $X=6.255 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_248 N_A_79_21#_M1005_d N_A_1142_47#_c_895_n 0.0031669f $X=6.12 $Y=0.235 $X2=0
+ $Y2=0
cc_249 N_A_79_21#_c_111_n N_A_1142_47#_c_895_n 0.0394091f $X=6.255 $Y=0.72 $X2=0
+ $Y2=0
cc_250 N_A_79_21#_c_111_n N_A_1142_47#_c_899_n 5.69174e-19 $X=6.255 $Y=0.72
+ $X2=0 $Y2=0
cc_251 N_A_79_21#_c_111_n N_A_1142_47#_c_900_n 0.011791f $X=6.255 $Y=0.72 $X2=0
+ $Y2=0
cc_252 A3 A2 0.0154972f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_253 N_A3_c_273_n A2 9.92259e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_254 A3 N_A2_c_317_n 0.00102695f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_255 N_A3_c_273_n N_A2_c_317_n 0.0076518f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A3_M1002_g N_VPWR_c_497_n 0.0102341f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A3_M1021_g N_VPWR_c_497_n 6.87435e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A3_M1002_g N_VPWR_c_498_n 5.08801e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A3_M1021_g N_VPWR_c_498_n 0.00774571f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A3_M1002_g N_VPWR_c_503_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A3_M1021_g N_VPWR_c_503_n 0.00339367f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A3_M1002_g N_VPWR_c_493_n 0.00789179f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A3_M1021_g N_VPWR_c_493_n 0.00394406f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A3_M1021_g N_A_445_297#_c_664_n 0.0135476f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A3_M1021_g N_A_445_297#_c_691_n 0.00260065f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_A3_c_270_n N_VGND_c_741_n 0.00762683f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A3_c_271_n N_VGND_c_741_n 5.08801e-19 $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A3_c_270_n N_VGND_c_742_n 5.08801e-19 $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A3_c_271_n N_VGND_c_742_n 0.00776975f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A3_c_270_n N_VGND_c_746_n 0.0046653f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A3_c_271_n N_VGND_c_746_n 0.00341689f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A3_c_270_n N_VGND_c_751_n 0.00789179f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A3_c_271_n N_VGND_c_751_n 0.0039829f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_274 A3 N_A_445_47#_c_853_n 0.00954402f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_275 N_A3_c_273_n N_A_445_47#_c_853_n 0.00219251f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A3_c_271_n N_A_445_47#_c_850_n 0.0136404f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_277 A3 N_A_445_47#_c_850_n 0.0330443f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_278 N_A3_c_273_n N_A_445_47#_c_850_n 0.00511673f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A2_c_315_n N_A1_M1010_g 0.0300535f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A2_M1023_g N_A1_M1006_g 0.0300535f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_281 A2 A1 0.0165684f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_282 N_A2_c_317_n A1 2.97858e-19 $X=3.93 $Y=1.17 $X2=0 $Y2=0
cc_283 A2 N_A1_c_362_n 0.00191046f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_284 N_A2_c_317_n N_A1_c_362_n 0.0300535f $X=3.93 $Y=1.17 $X2=0 $Y2=0
cc_285 N_A2_M1014_g N_VPWR_c_498_n 0.00186705f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A2_M1014_g N_VPWR_c_499_n 0.00703031f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A2_M1023_g N_VPWR_c_499_n 0.00664421f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A2_M1023_g N_VPWR_c_500_n 5.08801e-19 $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A2_M1014_g N_VPWR_c_505_n 0.00339367f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_290 N_A2_M1023_g N_VPWR_c_507_n 0.00339367f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A2_M1014_g N_VPWR_c_493_n 0.00527013f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A2_M1023_g N_VPWR_c_493_n 0.00397127f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_293 N_A2_M1014_g N_A_445_297#_c_679_n 0.014024f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A2_M1023_g N_A_445_297#_c_679_n 0.0118769f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_295 N_A2_c_314_n N_VGND_c_742_n 0.00294182f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A2_c_314_n N_VGND_c_749_n 0.00366111f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A2_c_315_n N_VGND_c_749_n 0.00366111f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A2_c_314_n N_VGND_c_751_n 0.00656615f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A2_c_315_n N_VGND_c_751_n 0.00526729f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A2_c_314_n N_A_445_47#_c_850_n 0.0110467f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_301 N_A2_c_315_n N_A_445_47#_c_850_n 0.0038838f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_302 A2 N_A_445_47#_c_850_n 0.0244044f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_303 N_A2_c_317_n N_A_445_47#_c_850_n 0.00412269f $X=3.93 $Y=1.17 $X2=0 $Y2=0
cc_304 N_A2_c_314_n N_A_635_47#_c_875_n 0.00801257f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A2_c_315_n N_A_635_47#_c_875_n 0.00956283f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_306 A2 N_A_635_47#_c_875_n 0.00330756f $X=3.85 $Y=1.105 $X2=0 $Y2=0
cc_307 N_A1_M1006_g N_VPWR_c_499_n 5.08801e-19 $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A1_M1006_g N_VPWR_c_500_n 0.00664421f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A1_M1008_g N_VPWR_c_500_n 0.00965315f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A1_M1006_g N_VPWR_c_507_n 0.00339367f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A1_M1008_g N_VPWR_c_510_n 0.00339367f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A1_M1006_g N_VPWR_c_493_n 0.00397127f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A1_M1008_g N_VPWR_c_493_n 0.00536411f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A1_M1006_g N_A_445_297#_c_680_n 0.0118327f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A1_M1008_g N_A_445_297#_c_680_n 0.0131292f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A1_M1010_g N_VGND_c_749_n 0.00366111f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A1_M1020_g N_VGND_c_749_n 0.00366111f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_318 N_A1_M1010_g N_VGND_c_751_n 0.00526729f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_319 N_A1_M1020_g N_VGND_c_751_n 0.00656615f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_320 N_A1_M1010_g N_A_445_47#_c_850_n 5.30585e-19 $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_321 N_A1_M1010_g N_A_635_47#_c_875_n 0.00942834f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_322 N_A1_M1020_g N_A_635_47#_c_875_n 0.00789149f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_323 A1 N_A_635_47#_c_875_n 0.00278778f $X=4.77 $Y=1.105 $X2=0 $Y2=0
cc_324 N_B1_M1011_g N_B2_M1012_g 0.0219887f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_325 N_B1_M1027_g N_B2_M1013_g 0.0304268f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_326 B1 B2 0.0168586f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_327 B1 N_B2_c_457_n 0.00543153f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_328 N_B1_c_406_n N_B2_c_457_n 0.0304268f $X=6.465 $Y=1.175 $X2=0 $Y2=0
cc_329 B1 N_B2_c_473_n 0.014598f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_330 N_B1_M1007_g N_VPWR_c_510_n 0.00366111f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_331 N_B1_M1027_g N_VPWR_c_510_n 0.00366111f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_332 N_B1_M1007_g N_VPWR_c_493_n 0.00656615f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_333 N_B1_M1027_g N_VPWR_c_493_n 0.00526729f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_334 B1 N_A_445_297#_M1008_d 0.00770625f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_335 B1 N_A_445_297#_M1027_s 0.00344244f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_336 N_B1_M1007_g N_A_445_297#_c_682_n 0.00794015f $X=6.09 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_B1_M1027_g N_A_445_297#_c_682_n 0.00789149f $X=6.51 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_B1_M1011_g N_VGND_c_743_n 0.00104498f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_339 N_B1_M1005_g N_VGND_c_749_n 0.00366111f $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_340 N_B1_M1011_g N_VGND_c_749_n 0.00366111f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_341 N_B1_M1005_g N_VGND_c_751_n 0.00656615f $X=6.045 $Y=0.56 $X2=0 $Y2=0
cc_342 N_B1_M1011_g N_VGND_c_751_n 0.00537416f $X=6.465 $Y=0.56 $X2=0 $Y2=0
cc_343 N_B1_M1005_g N_A_1142_47#_c_895_n 0.00784733f $X=6.045 $Y=0.56 $X2=0
+ $Y2=0
cc_344 N_B1_M1011_g N_A_1142_47#_c_895_n 0.00946925f $X=6.465 $Y=0.56 $X2=0
+ $Y2=0
cc_345 B1 N_A_1142_47#_c_895_n 0.00503476f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_346 N_B1_M1011_g N_A_1142_47#_c_899_n 0.00335185f $X=6.465 $Y=0.56 $X2=0
+ $Y2=0
cc_347 N_B1_M1011_g N_A_1142_47#_c_900_n 0.00170325f $X=6.465 $Y=0.56 $X2=0
+ $Y2=0
cc_348 B1 N_A_1142_47#_c_900_n 0.00948197f $X=6.58 $Y=1.105 $X2=0 $Y2=0
cc_349 N_B2_M1013_g N_VPWR_c_510_n 0.00366111f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_350 N_B2_M1018_g N_VPWR_c_510_n 0.00366111f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_351 N_B2_M1013_g N_VPWR_c_493_n 0.00526729f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_352 N_B2_M1018_g N_VPWR_c_493_n 0.00619429f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_353 N_B2_M1013_g N_A_445_297#_c_682_n 0.00789149f $X=6.93 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_B2_M1018_g N_A_445_297#_c_682_n 0.0115259f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_355 B2 N_A_445_297#_c_666_n 0.00861518f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_356 N_B2_c_457_n N_A_445_297#_c_666_n 0.0044264f $X=7.35 $Y=1.17 $X2=0 $Y2=0
cc_357 N_B2_M1012_g N_VGND_c_743_n 0.00787515f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_358 N_B2_M1022_g N_VGND_c_743_n 0.00835959f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_359 N_B2_M1012_g N_VGND_c_749_n 0.00340533f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_360 N_B2_M1022_g N_VGND_c_750_n 0.00340533f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_361 N_B2_M1012_g N_VGND_c_751_n 0.00409751f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_362 N_B2_M1022_g N_VGND_c_751_n 0.00491764f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_363 N_B2_M1012_g N_A_1142_47#_c_907_n 0.0157323f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_364 N_B2_M1022_g N_A_1142_47#_c_907_n 0.0131871f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_365 B2 N_A_1142_47#_c_907_n 0.0193451f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_366 N_B2_c_457_n N_A_1142_47#_c_907_n 0.00586263f $X=7.35 $Y=1.17 $X2=0 $Y2=0
cc_367 N_B2_c_473_n N_A_1142_47#_c_907_n 0.0098263f $X=7.127 $Y=1.295 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_493_n N_X_M1000_d 0.00562358f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_c_493_n N_X_M1017_d 0.00562358f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_370 N_VPWR_c_495_n N_X_c_620_n 0.00158991f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_371 N_VPWR_c_509_n N_X_c_638_n 0.0113958f $X=0.935 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_c_493_n N_X_c_638_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_373 N_VPWR_M1001_s N_X_c_625_n 0.00342716f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_374 N_VPWR_c_496_n N_X_c_625_n 0.0127176f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_375 N_VPWR_c_501_n N_X_c_642_n 0.0113958f $X=1.775 $Y=2.72 $X2=0 $Y2=0
cc_376 N_VPWR_c_493_n N_X_c_642_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_377 N_VPWR_M1000_s N_X_c_617_n 0.00342683f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_378 N_VPWR_c_495_n N_X_c_617_n 0.0147696f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_379 N_VPWR_c_493_n N_A_445_297#_M1002_s 0.00405853f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_380 N_VPWR_c_493_n N_A_445_297#_M1014_d 0.00240182f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_493_n N_A_445_297#_M1023_d 0.00249348f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_493_n N_A_445_297#_M1008_d 0.00980575f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_493_n N_A_445_297#_M1027_s 0.00217615f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_493_n N_A_445_297#_M1018_d 0.00211581f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_503_n N_A_445_297#_c_710_n 0.0112274f $X=2.615 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_493_n N_A_445_297#_c_710_n 0.00643448f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_VPWR_M1021_d N_A_445_297#_c_664_n 0.00517998f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_498_n N_A_445_297#_c_664_n 0.0206068f $X=2.78 $Y=2.34 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_503_n N_A_445_297#_c_664_n 0.00244309f $X=2.615 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_505_n N_A_445_297#_c_664_n 0.0048861f $X=3.555 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_493_n N_A_445_297#_c_664_n 0.0133342f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_498_n N_A_445_297#_c_691_n 0.0117639f $X=2.78 $Y=2.34 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_505_n N_A_445_297#_c_691_n 0.01143f $X=3.555 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_c_493_n N_A_445_297#_c_691_n 0.00643448f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_M1014_s N_A_445_297#_c_679_n 0.0034528f $X=3.585 $Y=1.485 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_499_n N_A_445_297#_c_679_n 0.0159625f $X=3.72 $Y=2.34 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_505_n N_A_445_297#_c_679_n 0.00244309f $X=3.555 $Y=2.72 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_507_n N_A_445_297#_c_679_n 0.00244309f $X=4.395 $Y=2.72 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_493_n N_A_445_297#_c_679_n 0.00984256f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_507_n N_A_445_297#_c_725_n 0.0112274f $X=4.395 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_493_n N_A_445_297#_c_725_n 0.00643448f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_M1006_s N_A_445_297#_c_680_n 0.0034528f $X=4.425 $Y=1.485 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_500_n N_A_445_297#_c_680_n 0.0159625f $X=4.56 $Y=2.34 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_507_n N_A_445_297#_c_680_n 0.00244309f $X=4.395 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_510_n N_A_445_297#_c_680_n 0.00244309f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_493_n N_A_445_297#_c_680_n 0.00988417f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_510_n N_A_445_297#_c_682_n 0.110877f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_493_n N_A_445_297#_c_682_n 0.0845075f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_510_n N_A_445_297#_c_734_n 0.00912819f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_493_n N_A_445_297#_c_734_n 0.00636368f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_510_n N_A_445_297#_c_665_n 0.0138224f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_493_n N_A_445_297#_c_665_n 0.00943351f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_X_c_615_n N_VGND_M1009_d 0.00291379f $X=0.23 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_414 X N_VGND_M1009_d 3.49814e-19 $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_415 N_X_c_621_n N_VGND_M1015_d 0.00312394f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_416 N_X_c_619_n N_VGND_c_739_n 0.0020301f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_417 N_X_c_615_n N_VGND_c_739_n 0.018421f $X=0.23 $Y=0.805 $X2=0 $Y2=0
cc_418 N_X_c_621_n N_VGND_c_740_n 0.0159625f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_419 N_X_c_621_n N_VGND_c_744_n 0.00244309f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_420 N_X_c_653_p N_VGND_c_744_n 0.0112274f $X=1.52 $Y=0.42 $X2=0 $Y2=0
cc_421 N_X_c_619_n N_VGND_c_748_n 0.00244309f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_422 N_X_c_655_p N_VGND_c_748_n 0.0112274f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_423 N_X_c_621_n N_VGND_c_748_n 0.00244309f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_424 N_X_M1009_s N_VGND_c_751_n 0.00249348f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_425 N_X_M1016_s N_VGND_c_751_n 0.00405853f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_426 N_X_c_619_n N_VGND_c_751_n 0.00456408f $X=0.595 $Y=0.72 $X2=0 $Y2=0
cc_427 N_X_c_655_p N_VGND_c_751_n 0.00643448f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_428 N_X_c_621_n N_VGND_c_751_n 0.00984256f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_429 N_X_c_653_p N_VGND_c_751_n 0.00643448f $X=1.52 $Y=0.42 $X2=0 $Y2=0
cc_430 N_X_c_615_n N_VGND_c_751_n 0.00110403f $X=0.23 $Y=0.805 $X2=0 $Y2=0
cc_431 N_VGND_c_751_n N_A_445_47#_M1019_s 0.00407273f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_432 N_VGND_c_751_n N_A_445_47#_M1003_s 0.00219239f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_c_746_n N_A_445_47#_c_865_n 0.0112554f $X=2.615 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_751_n N_A_445_47#_c_865_n 0.00644035f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_M1024_d N_A_445_47#_c_850_n 0.00498884f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_436 N_VGND_c_742_n N_A_445_47#_c_850_n 0.0187846f $X=2.78 $Y=0.38 $X2=0 $Y2=0
cc_437 N_VGND_c_746_n N_A_445_47#_c_850_n 0.0023303f $X=2.615 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_749_n N_A_445_47#_c_850_n 0.00332039f $X=6.975 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_751_n N_A_445_47#_c_850_n 0.0124182f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_751_n N_A_635_47#_M1003_d 0.00211652f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_441 N_VGND_c_751_n N_A_635_47#_M1004_d 0.00217615f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_442 N_VGND_c_751_n N_A_635_47#_M1020_s 0.00211652f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_742_n N_A_635_47#_c_875_n 0.0137364f $X=2.78 $Y=0.38 $X2=0 $Y2=0
cc_444 N_VGND_c_749_n N_A_635_47#_c_875_n 0.0906008f $X=6.975 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_751_n N_A_635_47#_c_875_n 0.0699807f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_751_n N_A_1142_47#_M1005_s 0.00211652f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_447 N_VGND_c_751_n N_A_1142_47#_M1011_s 0.00270767f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_448 N_VGND_c_751_n N_A_1142_47#_M1022_s 0.00369435f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_749_n N_A_1142_47#_c_895_n 0.043256f $X=6.975 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_751_n N_A_1142_47#_c_895_n 0.0335323f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_749_n N_A_1142_47#_c_917_n 0.0115494f $X=6.975 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_751_n N_A_1142_47#_c_917_n 0.00651407f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_M1012_d N_A_1142_47#_c_907_n 0.00338961f $X=7.005 $Y=0.235 $X2=0
+ $Y2=0
cc_454 N_VGND_c_743_n N_A_1142_47#_c_907_n 0.0152077f $X=7.14 $Y=0.38 $X2=0
+ $Y2=0
cc_455 N_VGND_c_749_n N_A_1142_47#_c_907_n 0.00238578f $X=6.975 $Y=0 $X2=0 $Y2=0
cc_456 N_VGND_c_750_n N_A_1142_47#_c_907_n 0.00238578f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_457 N_VGND_c_751_n N_A_1142_47#_c_907_n 0.0097758f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_750_n N_A_1142_47#_c_924_n 0.0114446f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_751_n N_A_1142_47#_c_924_n 0.00643744f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_460 N_A_445_47#_c_850_n N_A_635_47#_M1003_d 0.00672949f $X=3.72 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_461 N_A_445_47#_M1003_s N_A_635_47#_c_875_n 0.00323216f $X=3.585 $Y=0.235
+ $X2=0 $Y2=0
cc_462 N_A_445_47#_c_850_n N_A_635_47#_c_875_n 0.0355575f $X=3.72 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_635_47#_c_875_n N_A_1142_47#_c_895_n 0.00716889f $X=4.98 $Y=0.38
+ $X2=0 $Y2=0

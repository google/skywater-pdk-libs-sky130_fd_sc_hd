* File: sky130_fd_sc_hd__and2b_4.spice.SKY130_FD_SC_HD__AND2B_4.pxi
* Created: Thu Aug 27 14:07:27 2020
* 
x_PM_SKY130_FD_SC_HD__AND2B_4%A_33_199# N_A_33_199#_M1004_d N_A_33_199#_M1002_d
+ N_A_33_199#_M1012_g N_A_33_199#_M1010_g N_A_33_199#_c_75_n N_A_33_199#_c_76_n
+ N_A_33_199#_c_113_p N_A_33_199#_c_77_n N_A_33_199#_c_69_n N_A_33_199#_c_70_n
+ N_A_33_199#_c_71_n N_A_33_199#_c_72_n N_A_33_199#_c_73_n
+ PM_SKY130_FD_SC_HD__AND2B_4%A_33_199#
x_PM_SKY130_FD_SC_HD__AND2B_4%B N_B_M1011_g N_B_M1006_g B N_B_c_139_n
+ N_B_c_140_n N_B_c_141_n PM_SKY130_FD_SC_HD__AND2B_4%B
x_PM_SKY130_FD_SC_HD__AND2B_4%A_27_47# N_A_27_47#_M1012_s N_A_27_47#_M1010_d
+ N_A_27_47#_c_174_n N_A_27_47#_M1003_g N_A_27_47#_M1000_g N_A_27_47#_c_175_n
+ N_A_27_47#_M1005_g N_A_27_47#_M1001_g N_A_27_47#_c_176_n N_A_27_47#_M1008_g
+ N_A_27_47#_M1007_g N_A_27_47#_c_177_n N_A_27_47#_M1009_g N_A_27_47#_M1013_g
+ N_A_27_47#_c_178_n N_A_27_47#_c_196_n N_A_27_47#_c_179_n N_A_27_47#_c_200_n
+ N_A_27_47#_c_180_n N_A_27_47#_c_181_n N_A_27_47#_c_188_n N_A_27_47#_c_182_n
+ PM_SKY130_FD_SC_HD__AND2B_4%A_27_47#
x_PM_SKY130_FD_SC_HD__AND2B_4%A_N N_A_N_M1004_g N_A_N_M1002_g A_N N_A_N_c_288_n
+ N_A_N_c_289_n N_A_N_c_290_n PM_SKY130_FD_SC_HD__AND2B_4%A_N
x_PM_SKY130_FD_SC_HD__AND2B_4%VPWR N_VPWR_M1010_s N_VPWR_M1006_d N_VPWR_M1001_s
+ N_VPWR_M1013_s N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n
+ N_VPWR_c_328_n VPWR N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n
+ N_VPWR_c_332_n N_VPWR_c_323_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n
+ PM_SKY130_FD_SC_HD__AND2B_4%VPWR
x_PM_SKY130_FD_SC_HD__AND2B_4%X N_X_M1003_d N_X_M1008_d N_X_M1000_d N_X_M1007_d
+ N_X_c_387_n N_X_c_393_n N_X_c_388_n X N_X_c_400_n X
+ PM_SKY130_FD_SC_HD__AND2B_4%X
x_PM_SKY130_FD_SC_HD__AND2B_4%VGND N_VGND_M1011_d N_VGND_M1005_s N_VGND_M1009_s
+ N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n VGND N_VGND_c_431_n
+ N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n N_VGND_c_436_n
+ N_VGND_c_437_n N_VGND_c_438_n PM_SKY130_FD_SC_HD__AND2B_4%VGND
cc_1 VNB N_A_33_199#_c_69_n 0.00601813f $X=-0.19 $Y=-0.24 $X2=3.46 $Y2=0.845
cc_2 VNB N_A_33_199#_c_70_n 0.0111949f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=1.16
cc_3 VNB N_A_33_199#_c_71_n 0.0320811f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=1.16
cc_4 VNB N_A_33_199#_c_72_n 0.0194216f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.53
cc_5 VNB N_A_33_199#_c_73_n 0.0217282f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=0.995
cc_6 VNB N_B_c_139_n 0.0213454f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_7 VNB N_B_c_140_n 0.0032562f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_8 VNB N_B_c_141_n 0.017206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_174_n 0.0169506f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_10 VNB N_A_27_47#_c_175_n 0.0159671f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.325
cc_11 VNB N_A_27_47#_c_176_n 0.016002f $X=-0.19 $Y=-0.24 $X2=3.46 $Y2=1.53
cc_12 VNB N_A_27_47#_c_177_n 0.0179086f $X=-0.19 $Y=-0.24 $X2=3.437 $Y2=0.68
cc_13 VNB N_A_27_47#_c_178_n 0.0143075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_179_n 0.00980077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_180_n 0.00112303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_181_n 0.00185646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_182_n 0.0646727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_N_c_288_n 0.024155f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.915
cc_19 VNB N_A_N_c_289_n 0.0024888f $X=-0.19 $Y=-0.24 $X2=3.335 $Y2=2
cc_20 VNB N_A_N_c_290_n 0.0209342f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=2
cc_21 VNB N_VPWR_c_323_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB X 0.00108133f $X=-0.19 $Y=-0.24 $X2=3.44 $Y2=1.53
cc_23 VNB N_VGND_c_428_n 0.00500766f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_24 VNB N_VGND_c_429_n 3.20903e-19 $X=-0.19 $Y=-0.24 $X2=3.335 $Y2=2
cc_25 VNB N_VGND_c_430_n 0.00770873f $X=-0.19 $Y=-0.24 $X2=3.46 $Y2=0.845
cc_26 VNB N_VGND_c_431_n 0.026813f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=1.16
cc_27 VNB N_VGND_c_432_n 0.0157647f $X=-0.19 $Y=-0.24 $X2=3.415 $Y2=0.68
cc_28 VNB N_VGND_c_433_n 0.0123295f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_29 VNB N_VGND_c_434_n 0.0198578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_435_n 0.208357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_436_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_437_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_438_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_33_199#_M1010_g 0.0213171f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_35 VPB N_A_33_199#_c_75_n 0.00695159f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.915
cc_36 VPB N_A_33_199#_c_76_n 0.0153435f $X=-0.19 $Y=1.305 $X2=3.335 $Y2=2
cc_37 VPB N_A_33_199#_c_77_n 3.96483e-19 $X=-0.19 $Y=1.305 $X2=3.42 $Y2=1.915
cc_38 VPB N_A_33_199#_c_70_n 6.88357e-19 $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_39 VPB N_A_33_199#_c_71_n 0.00841841f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_40 VPB N_A_33_199#_c_72_n 0.00837891f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.53
cc_41 VPB N_B_M1006_g 0.020144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B_c_139_n 0.00418065f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_43 VPB N_B_c_140_n 0.00147473f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_A_27_47#_M1000_g 0.019888f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_45 VPB N_A_27_47#_M1001_g 0.0183712f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=1.915
cc_46 VPB N_A_27_47#_M1007_g 0.0181173f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_47 VPB N_A_27_47#_M1013_g 0.0202446f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.7
cc_48 VPB N_A_27_47#_c_181_n 0.0036561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_188_n 0.0054084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_182_n 0.0122453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_N_M1002_g 0.0198345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB A_N 9.44539e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_53 VPB N_A_N_c_288_n 0.00639398f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.915
cc_54 VPB N_VPWR_c_324_n 0.0102396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_325_n 0.0133481f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.915
cc_56 VPB N_VPWR_c_326_n 0.00433352f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=1.915
cc_57 VPB N_VPWR_c_327_n 3.1483e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_328_n 0.0107613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_329_n 0.0143676f $X=-0.19 $Y=1.305 $X2=3.42 $Y2=1.695
cc_60 VPB N_VPWR_c_330_n 0.0149152f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.325
cc_61 VPB N_VPWR_c_331_n 0.011815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_332_n 0.0194881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_323_n 0.0511583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_334_n 0.00631318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_335_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_336_n 0.00507043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB X 0.00145578f $X=-0.19 $Y=1.305 $X2=3.44 $Y2=1.53
cc_68 N_A_33_199#_M1010_g N_B_M1006_g 0.0437006f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A_33_199#_c_76_n N_B_M1006_g 0.0121939f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_70 N_A_33_199#_c_70_n N_B_c_139_n 2.63582e-19 $X=0.34 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_33_199#_c_71_n N_B_c_139_n 0.0205885f $X=0.34 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_33_199#_c_70_n N_B_c_140_n 0.0243633f $X=0.34 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_33_199#_c_71_n N_B_c_140_n 0.00243572f $X=0.34 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_33_199#_c_73_n N_B_c_141_n 0.0530016f $X=0.355 $Y=0.995 $X2=0 $Y2=0
cc_75 N_A_33_199#_c_76_n N_A_27_47#_M1010_d 0.00435118f $X=3.335 $Y=2 $X2=0
+ $Y2=0
cc_76 N_A_33_199#_c_76_n N_A_27_47#_M1000_g 0.0143148f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_77 N_A_33_199#_c_76_n N_A_27_47#_M1001_g 0.0116569f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_78 N_A_33_199#_c_76_n N_A_27_47#_M1007_g 0.0114745f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_79 N_A_33_199#_c_76_n N_A_27_47#_M1013_g 0.0137414f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_80 N_A_33_199#_c_73_n N_A_27_47#_c_178_n 0.00657339f $X=0.355 $Y=0.995 $X2=0
+ $Y2=0
cc_81 N_A_33_199#_c_73_n N_A_27_47#_c_196_n 0.0118531f $X=0.355 $Y=0.995 $X2=0
+ $Y2=0
cc_82 N_A_33_199#_c_70_n N_A_27_47#_c_179_n 0.0169686f $X=0.34 $Y=1.16 $X2=0
+ $Y2=0
cc_83 N_A_33_199#_c_71_n N_A_27_47#_c_179_n 0.00508593f $X=0.34 $Y=1.16 $X2=0
+ $Y2=0
cc_84 N_A_33_199#_c_73_n N_A_27_47#_c_179_n 9.45079e-19 $X=0.355 $Y=0.995 $X2=0
+ $Y2=0
cc_85 N_A_33_199#_M1010_g N_A_27_47#_c_200_n 0.00448628f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_86 N_A_33_199#_c_75_n N_A_27_47#_c_200_n 0.0182669f $X=0.25 $Y=1.915 $X2=0
+ $Y2=0
cc_87 N_A_33_199#_c_76_n N_A_27_47#_c_200_n 0.030664f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_88 N_A_33_199#_c_76_n N_A_27_47#_c_181_n 0.0143706f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_89 N_A_33_199#_c_76_n N_A_27_47#_c_188_n 0.00349389f $X=3.335 $Y=2 $X2=0
+ $Y2=0
cc_90 N_A_33_199#_c_76_n N_A_27_47#_c_182_n 2.68063e-19 $X=3.335 $Y=2 $X2=0
+ $Y2=0
cc_91 N_A_33_199#_c_76_n N_A_N_M1002_g 0.0128628f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_92 N_A_33_199#_c_77_n N_A_N_M1002_g 6.3613e-19 $X=3.42 $Y=1.915 $X2=0 $Y2=0
cc_93 N_A_33_199#_c_76_n A_N 0.0180009f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_94 N_A_33_199#_c_72_n A_N 0.0123027f $X=3.44 $Y=1.53 $X2=0 $Y2=0
cc_95 N_A_33_199#_c_76_n N_A_N_c_288_n 4.42296e-19 $X=3.335 $Y=2 $X2=0 $Y2=0
cc_96 N_A_33_199#_c_76_n N_A_N_c_289_n 0.00125482f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_97 N_A_33_199#_c_72_n N_A_N_c_289_n 0.0336485f $X=3.44 $Y=1.53 $X2=0 $Y2=0
cc_98 N_A_33_199#_c_72_n N_A_N_c_290_n 0.0144599f $X=3.44 $Y=1.53 $X2=0 $Y2=0
cc_99 N_A_33_199#_c_75_n N_VPWR_M1010_s 0.0230719f $X=0.25 $Y=1.915 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_33_199#_c_113_p N_VPWR_M1010_s 0.0099277f $X=0.335 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_33_199#_c_76_n N_VPWR_M1006_d 0.00552345f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_102 N_A_33_199#_c_76_n N_VPWR_M1001_s 0.00324696f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_103 N_A_33_199#_c_76_n N_VPWR_M1013_s 0.00658751f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_104 N_A_33_199#_M1010_g N_VPWR_c_325_n 0.00954136f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_105 N_A_33_199#_c_76_n N_VPWR_c_325_n 0.00216057f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_106 N_A_33_199#_c_113_p N_VPWR_c_325_n 0.0142454f $X=0.335 $Y=2 $X2=0 $Y2=0
cc_107 N_A_33_199#_c_76_n N_VPWR_c_326_n 0.0176844f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_108 N_A_33_199#_c_76_n N_VPWR_c_327_n 0.0144274f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_109 N_A_33_199#_c_76_n N_VPWR_c_328_n 0.0185984f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_110 N_A_33_199#_M1010_g N_VPWR_c_329_n 0.00339367f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_33_199#_c_76_n N_VPWR_c_329_n 0.00848923f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_112 N_A_33_199#_c_76_n N_VPWR_c_330_n 0.00891648f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_113 N_A_33_199#_c_76_n N_VPWR_c_331_n 0.0077537f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_114 N_A_33_199#_c_76_n N_VPWR_c_332_n 0.0081729f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_115 N_A_33_199#_M1010_g N_VPWR_c_323_n 0.00401529f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_33_199#_c_76_n N_VPWR_c_323_n 0.0606048f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_117 N_A_33_199#_c_113_p N_VPWR_c_323_n 8.51964e-19 $X=0.335 $Y=2 $X2=0 $Y2=0
cc_118 N_A_33_199#_c_76_n N_X_M1000_d 0.00511359f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_119 N_A_33_199#_c_76_n N_X_M1007_d 0.00424264f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_120 N_A_33_199#_c_76_n N_X_c_387_n 0.0478692f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_121 N_A_33_199#_c_76_n N_X_c_388_n 0.0182832f $X=3.335 $Y=2 $X2=0 $Y2=0
cc_122 N_A_33_199#_c_73_n N_VGND_c_431_n 0.00410742f $X=0.355 $Y=0.995 $X2=0
+ $Y2=0
cc_123 N_A_33_199#_c_69_n N_VGND_c_434_n 0.00526302f $X=3.46 $Y=0.845 $X2=0
+ $Y2=0
cc_124 N_A_33_199#_c_69_n N_VGND_c_435_n 0.00693229f $X=3.46 $Y=0.845 $X2=0
+ $Y2=0
cc_125 N_A_33_199#_c_73_n N_VGND_c_435_n 0.00651603f $X=0.355 $Y=0.995 $X2=0
+ $Y2=0
cc_126 N_B_c_141_n N_A_27_47#_c_174_n 0.0228172f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_M1006_g N_A_27_47#_M1000_g 0.0307733f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_128 N_B_c_141_n N_A_27_47#_c_178_n 0.00140175f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B_c_139_n N_A_27_47#_c_196_n 0.00324796f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B_c_140_n N_A_27_47#_c_196_n 0.0212986f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B_c_141_n N_A_27_47#_c_196_n 0.0129179f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B_M1006_g N_A_27_47#_c_200_n 0.0107643f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_133 N_B_c_139_n N_A_27_47#_c_200_n 0.00267363f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B_c_140_n N_A_27_47#_c_200_n 0.0247547f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B_c_141_n N_A_27_47#_c_180_n 0.00401133f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B_M1006_g N_A_27_47#_c_181_n 0.0040715f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B_c_139_n N_A_27_47#_c_181_n 0.00267591f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_138 N_B_c_140_n N_A_27_47#_c_181_n 0.0279866f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B_c_139_n N_A_27_47#_c_182_n 0.0121499f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B_c_140_n N_A_27_47#_c_182_n 2.82297e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B_M1006_g N_VPWR_c_325_n 0.00117943f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B_M1006_g N_VPWR_c_326_n 0.00167244f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B_M1006_g N_VPWR_c_329_n 0.00425094f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B_M1006_g N_VPWR_c_323_n 0.00593012f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B_c_141_n N_VGND_c_428_n 0.00443612f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B_c_141_n N_VGND_c_431_n 0.00422112f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B_c_141_n N_VGND_c_435_n 0.00594019f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_27_47#_M1013_g N_A_N_M1002_g 0.0218739f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_27_47#_M1013_g A_N 0.00260841f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_182_n N_A_N_c_288_n 0.0225707f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_177_n N_A_N_c_289_n 0.00260841f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_182_n N_A_N_c_289_n 0.00260841f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_177_n N_A_N_c_290_n 0.0167986f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_200_n N_VPWR_M1006_d 0.00428751f $X=1.11 $Y=1.622 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_181_n N_VPWR_M1006_d 0.00353162f $X=1.355 $Y=1.175 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_M1000_g N_VPWR_c_326_n 0.00174557f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_M1000_g N_VPWR_c_327_n 0.00108373f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_M1001_g N_VPWR_c_327_n 0.00822055f $X=1.86 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_M1007_g N_VPWR_c_327_n 0.00778395f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_M1013_g N_VPWR_c_327_n 0.0010441f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_27_47#_M1007_g N_VPWR_c_328_n 0.0010441f $X=2.28 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_27_47#_M1013_g N_VPWR_c_328_n 0.00888545f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1000_g N_VPWR_c_330_n 0.00425094f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1001_g N_VPWR_c_330_n 0.00339367f $X=1.86 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_M1007_g N_VPWR_c_331_n 0.00339367f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_M1013_g N_VPWR_c_331_n 0.00339367f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_27_47#_M1010_d N_VPWR_c_323_n 0.00315309f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_M1000_g N_VPWR_c_323_n 0.0059574f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_27_47#_M1001_g N_VPWR_c_323_n 0.00406766f $X=1.86 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_M1007_g N_VPWR_c_323_n 0.00398704f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_M1013_g N_VPWR_c_323_n 0.00398704f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1001_g N_X_c_387_n 0.00950374f $X=1.86 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_27_47#_M1007_g N_X_c_387_n 0.0124269f $X=2.28 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_188_n N_X_c_387_n 0.0496512f $X=2.175 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_182_n N_X_c_387_n 0.00136917f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_188_n N_X_c_393_n 0.0138754f $X=2.175 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_182_n N_X_c_393_n 0.00227989f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_27_47#_M1013_g N_X_c_388_n 0.00476177f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_175_n X 0.0105076f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_176_n X 0.0131838f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_188_n X 0.0344384f $X=2.175 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_182_n X 0.00252546f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_177_n N_X_c_400_n 0.00567041f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_176_n X 0.00401795f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1007_g X 0.00457037f $X=2.28 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_177_n X 0.00350566f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_27_47#_M1013_g X 0.00447851f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_188_n X 0.027114f $X=2.175 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_182_n X 0.0194051f $X=2.7 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_196_n A_109_47# 0.00322045f $X=1.145 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_191 N_A_27_47#_c_196_n N_VGND_M1011_d 0.00832189f $X=1.145 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_192 N_A_27_47#_c_180_n N_VGND_M1011_d 9.82356e-19 $X=1.25 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_193 N_A_27_47#_c_174_n N_VGND_c_428_n 0.00293602f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_196_n N_VGND_c_428_n 0.0243121f $X=1.145 $Y=0.71 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_174_n N_VGND_c_429_n 0.00109956f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_175_n N_VGND_c_429_n 0.0082981f $X=1.84 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_176_n N_VGND_c_429_n 0.0073705f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_177_n N_VGND_c_429_n 0.00103247f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_176_n N_VGND_c_430_n 0.00105539f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_177_n N_VGND_c_430_n 0.009994f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_178_n N_VGND_c_431_n 0.0210984f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_196_n N_VGND_c_431_n 0.00818831f $X=1.145 $Y=0.71 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_174_n N_VGND_c_432_n 0.00563595f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_175_n N_VGND_c_432_n 0.00337001f $X=1.84 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_196_n N_VGND_c_432_n 8.83096e-19 $X=1.145 $Y=0.71 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_176_n N_VGND_c_433_n 0.00365142f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_177_n N_VGND_c_433_n 0.00352135f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1012_s N_VGND_c_435_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_174_n N_VGND_c_435_n 0.0104168f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_175_n N_VGND_c_435_n 0.00397572f $X=1.84 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_176_n N_VGND_c_435_n 0.00425782f $X=2.27 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_177_n N_VGND_c_435_n 0.00450554f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_178_n N_VGND_c_435_n 0.0125495f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_196_n N_VGND_c_435_n 0.0175956f $X=1.145 $Y=0.71 $X2=0 $Y2=0
cc_215 A_N N_VPWR_M1013_s 0.00453898f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A_N_M1002_g N_VPWR_c_332_n 5.36286e-19 $X=3.205 $Y=1.695 $X2=0 $Y2=0
cc_217 A_N N_X_c_388_n 0.0169853f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_218 N_A_N_c_289_n N_X_c_400_n 0.0161764f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_N_c_290_n N_X_c_400_n 2.06071e-19 $X=3.132 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_N_c_288_n X 3.40899e-19 $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_N_c_289_n X 0.0545107f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_N_c_289_n N_VGND_M1009_s 0.00445213f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_N_c_288_n N_VGND_c_430_n 3.1887e-19 $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_N_c_289_n N_VGND_c_430_n 0.0137913f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_N_c_290_n N_VGND_c_430_n 0.00308742f $X=3.132 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_N_c_289_n N_VGND_c_434_n 9.85095e-19 $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_N_c_290_n N_VGND_c_434_n 0.0049127f $X=3.132 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_N_c_289_n N_VGND_c_435_n 0.00332621f $X=3.12 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_N_c_290_n N_VGND_c_435_n 0.00512902f $X=3.132 $Y=0.995 $X2=0 $Y2=0
cc_230 N_VPWR_c_323_n N_X_M1000_d 0.00350343f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_231 N_VPWR_c_323_n N_X_M1007_d 0.00315309f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_M1001_s N_X_c_387_n 0.00318416f $X=1.935 $Y=1.485 $X2=0 $Y2=0
cc_233 X N_VGND_M1005_s 0.0032524f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_234 X N_VGND_c_429_n 0.0161306f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_235 N_X_c_393_n N_VGND_c_432_n 0.00459233f $X=1.62 $Y=0.66 $X2=0 $Y2=0
cc_236 X N_VGND_c_432_n 0.00258359f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_237 X N_VGND_c_433_n 0.00352663f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_238 N_X_c_400_n N_VGND_c_433_n 0.0051409f $X=2.585 $Y=0.825 $X2=0 $Y2=0
cc_239 N_X_M1003_d N_VGND_c_435_n 0.00416103f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_240 N_X_M1008_d N_VGND_c_435_n 0.00318706f $X=2.345 $Y=0.235 $X2=0 $Y2=0
cc_241 N_X_c_393_n N_VGND_c_435_n 0.00607819f $X=1.62 $Y=0.66 $X2=0 $Y2=0
cc_242 X N_VGND_c_435_n 0.0117695f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_243 N_X_c_400_n N_VGND_c_435_n 0.00830293f $X=2.585 $Y=0.825 $X2=0 $Y2=0
cc_244 A_109_47# N_VGND_c_435_n 0.00250619f $X=0.545 $Y=0.235 $X2=0.68 $Y2=1.622

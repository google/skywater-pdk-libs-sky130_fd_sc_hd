* File: sky130_fd_sc_hd__dfxbp_2.pex.spice
* Created: Tue Sep  1 19:04:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFXBP_2%CLK 1 2 3 5 6 8 11 13
c40 1 0 2.71124e-20 $X=0.305 $Y=1.325
r41 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r42 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r43 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r44 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r45 3 16 88.7086 $w=2.58e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r46 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r47 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r48 1 16 39.2009 $w=2.58e-07 $l=1.75656e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.327 $Y2=1.16
r49 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_27_47# 1 2 9 13 17 21 25 27 31 35 39 40 41
+ 44 46 48 51 54 56 57 58 59 60 67 69 74 82 85 89
c239 89 0 1.92554e-19 $X=4.375 $Y=1.41
c240 60 0 3.69553e-20 $X=2.96 $Y=1.87
c241 59 0 8.81722e-20 $X=4.24 $Y=1.87
c242 51 0 1.91737e-19 $X=2.38 $Y=0.87
c243 44 0 1.81794e-19 $X=0.725 $Y=1.795
c244 41 0 3.29888e-20 $X=0.61 $Y=1.88
r245 88 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.41
+ $X2=4.375 $Y2=1.575
r246 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.375
+ $Y=1.41 $X2=4.375 $Y2=1.41
r247 85 88 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=4.375 $Y=1.32
+ $X2=4.375 $Y2=1.41
r248 79 82 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.73 $Y=1.74
+ $X2=2.825 $Y2=1.74
r249 70 89 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=4.385 $Y=1.87
+ $X2=4.385 $Y2=1.41
r250 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.385 $Y=1.87
+ $X2=4.385 $Y2=1.87
r251 67 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.74 $X2=2.825 $Y2=1.74
r252 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.815 $Y=1.87
+ $X2=2.815 $Y2=1.87
r253 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.715 $Y=1.87
+ $X2=0.715 $Y2=1.87
r254 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.96 $Y=1.87
+ $X2=2.815 $Y2=1.87
r255 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.24 $Y=1.87
+ $X2=4.385 $Y2=1.87
r256 59 60 1.58416 $w=1.4e-07 $l=1.28e-06 $layer=MET1_cond $X=4.24 $Y=1.87
+ $X2=2.96 $Y2=1.87
r257 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.86 $Y=1.87
+ $X2=0.715 $Y2=1.87
r258 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.67 $Y=1.87
+ $X2=2.815 $Y2=1.87
r259 57 58 2.24009 $w=1.4e-07 $l=1.81e-06 $layer=MET1_cond $X=2.67 $Y=1.87
+ $X2=0.86 $Y2=1.87
r260 54 67 5.05181 $w=3.63e-07 $l=1.6e-07 $layer=LI1_cond $X=2.655 $Y=1.837
+ $X2=2.815 $Y2=1.837
r261 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.655 $Y=0.955
+ $X2=2.655 $Y2=1.655
r262 51 77 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.38 $Y=0.87
+ $X2=2.38 $Y2=0.735
r263 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=0.87 $X2=2.38 $Y2=0.87
r264 48 53 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.57 $Y=0.845
+ $X2=2.655 $Y2=0.955
r265 48 50 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=2.57 $Y=0.845
+ $X2=2.38 $Y2=0.845
r266 47 74 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r267 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r268 44 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r269 44 46 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r270 43 46 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r271 42 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r272 41 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r273 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r274 39 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r275 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r276 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r277 33 35 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r278 29 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=5.01 $Y=1.245
+ $X2=5.01 $Y2=0.415
r279 28 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.51 $Y=1.32
+ $X2=4.375 $Y2=1.32
r280 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.935 $Y=1.32
+ $X2=5.01 $Y2=1.245
r281 27 28 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.935 $Y=1.32
+ $X2=4.51 $Y2=1.32
r282 25 90 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.38 $Y=2.275
+ $X2=4.38 $Y2=1.575
r283 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.905
+ $X2=2.73 $Y2=1.74
r284 19 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.73 $Y=1.905
+ $X2=2.73 $Y2=2.275
r285 17 77 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.39 $Y=0.415
+ $X2=2.39 $Y2=0.735
r286 11 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r287 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r288 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r289 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r290 2 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r291 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%D 3 7 9 15
r45 12 15 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.565 $Y=1.5
+ $X2=1.83 $Y2=1.5
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.5 $X2=1.565 $Y2=1.5
r47 9 13 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.51 $Y=1.19 $X2=1.51
+ $Y2=1.5
r48 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.665
+ $X2=1.83 $Y2=1.5
r49 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.83 $Y=1.665 $X2=1.83
+ $Y2=2.275
r50 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.335
+ $X2=1.83 $Y2=1.5
r51 1 3 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.83 $Y=1.335 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_193_47# 1 2 9 11 15 17 19 22 26 27 30 31
+ 32 33 42 43 45 49 58 62
c179 45 0 1.74123e-19 $X=2.28 $Y=1.29
c180 43 0 2.06462e-20 $X=4.82 $Y=1.53
c181 22 0 1.92554e-19 $X=4.8 $Y=2.275
r182 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.74 $X2=4.885 $Y2=1.74
r183 55 58 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=4.8 $Y=1.74
+ $X2=4.885 $Y2=1.74
r184 48 50 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.28 $Y=1.35
+ $X2=2.28 $Y2=1.485
r185 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.35 $X2=2.28 $Y2=1.35
r186 45 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.28 $Y=1.29 $X2=2.28
+ $Y2=1.35
r187 43 59 7.56291 $w=3.18e-07 $l=2.1e-07 $layer=LI1_cond $X=4.81 $Y=1.53
+ $X2=4.81 $Y2=1.74
r188 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.82 $Y=1.53
+ $X2=4.82 $Y2=1.53
r189 40 49 8.64332 $w=2.38e-07 $l=1.8e-07 $layer=LI1_cond $X=2.28 $Y=1.53
+ $X2=2.28 $Y2=1.35
r190 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.3 $Y=1.53 $X2=2.3
+ $Y2=1.53
r191 36 66 25.7789 $w=1.83e-07 $l=4.3e-07 $layer=LI1_cond $X=1.107 $Y=1.53
+ $X2=1.107 $Y2=1.96
r192 36 62 61.1499 $w=1.83e-07 $l=1.02e-06 $layer=LI1_cond $X=1.107 $Y=1.53
+ $X2=1.107 $Y2=0.51
r193 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.11 $Y=1.53
+ $X2=1.11 $Y2=1.53
r194 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.445 $Y=1.53
+ $X2=2.3 $Y2=1.53
r195 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.675 $Y=1.53
+ $X2=4.82 $Y2=1.53
r196 32 33 2.7599 $w=1.4e-07 $l=2.23e-06 $layer=MET1_cond $X=4.675 $Y=1.53
+ $X2=2.445 $Y2=1.53
r197 31 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.255 $Y=1.53
+ $X2=1.11 $Y2=1.53
r198 30 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.155 $Y=1.53
+ $X2=2.3 $Y2=1.53
r199 30 31 1.11386 $w=1.4e-07 $l=9e-07 $layer=MET1_cond $X=2.155 $Y=1.53
+ $X2=1.255 $Y2=1.53
r200 29 43 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=4.81 $Y=1.035
+ $X2=4.81 $Y2=1.53
r201 27 51 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.59 $Y=0.87
+ $X2=4.48 $Y2=0.87
r202 26 29 5.41706 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=4.737 $Y=0.87
+ $X2=4.737 $Y2=1.035
r203 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.59
+ $Y=0.87 $X2=4.59 $Y2=0.87
r204 20 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.8 $Y=1.875
+ $X2=4.8 $Y2=1.74
r205 20 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.8 $Y=1.875 $X2=4.8
+ $Y2=2.275
r206 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=0.705
+ $X2=4.48 $Y2=0.87
r207 17 19 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.48 $Y=0.705
+ $X2=4.48 $Y2=0.415
r208 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.885 $Y=1.215
+ $X2=2.885 $Y2=0.415
r209 12 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=1.29
+ $X2=2.28 $Y2=1.29
r210 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=1.29
+ $X2=2.885 $Y2=1.215
r211 11 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.81 $Y=1.29
+ $X2=2.445 $Y2=1.29
r212 9 50 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.255 $Y=2.275
+ $X2=2.255 $Y2=1.485
r213 2 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r214 1 62 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_634_159# 1 2 9 13 15 18 25 29 31 33 34 39
r90 33 34 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.3
+ $X2=4.075 $Y2=2.135
r91 26 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.035 $Y=0.45
+ $X2=4.19 $Y2=0.45
r92 23 39 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=3.375 $Y=0.93 $X2=3.38
+ $Y2=0.93
r93 23 36 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=3.375 $Y=0.93
+ $X2=3.245 $Y2=0.93
r94 22 25 4.13427 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.375 $Y=0.93
+ $X2=3.49 $Y2=0.93
r95 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.375
+ $Y=0.93 $X2=3.375 $Y2=0.93
r96 19 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.035 $Y=1.065
+ $X2=4.035 $Y2=0.915
r97 19 34 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.035 $Y=1.065
+ $X2=4.035 $Y2=2.135
r98 18 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.035 $Y=0.765
+ $X2=4.035 $Y2=0.915
r99 17 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.535
+ $X2=4.035 $Y2=0.45
r100 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.035 $Y=0.535
+ $X2=4.035 $Y2=0.765
r101 15 31 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=0.915
+ $X2=4.035 $Y2=0.915
r102 15 25 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.95 $Y=0.915
+ $X2=3.49 $Y2=0.915
r103 11 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.38 $Y=0.795
+ $X2=3.38 $Y2=0.93
r104 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.38 $Y=0.795
+ $X2=3.38 $Y2=0.445
r105 7 36 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.245 $Y=1.065
+ $X2=3.245 $Y2=0.93
r106 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=3.245 $Y=1.065
+ $X2=3.245 $Y2=2.275
r107 2 33 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.735 $X2=4.115 $Y2=2.3
r108 1 29 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.05
+ $Y=0.235 $X2=4.19 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_466_413# 1 2 8 11 15 16 17 18 19 20 24 29
+ 30 31 33 34
c120 31 0 1.25128e-19 $X=3.08 $Y=1.4
c121 29 0 2.60836e-19 $X=2.995 $Y=1.315
r122 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.41 $X2=3.695 $Y2=1.41
r123 34 36 14.6572 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=3.355 $Y=1.41
+ $X2=3.695 $Y2=1.41
r124 32 34 3.71884 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=1.575
+ $X2=3.355 $Y2=1.41
r125 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.355 $Y=1.575
+ $X2=3.355 $Y2=2.19
r126 30 34 5.59441 $w=2.83e-07 $l=8.9861e-08 $layer=LI1_cond $X=3.27 $Y=1.4
+ $X2=3.355 $Y2=1.41
r127 30 31 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.27 $Y=1.4
+ $X2=3.08 $Y2=1.4
r128 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=1.315
+ $X2=3.08 $Y2=1.4
r129 28 29 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.995 $Y=0.535
+ $X2=2.995 $Y2=1.315
r130 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.91 $Y=0.45
+ $X2=2.995 $Y2=0.535
r131 24 26 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.91 $Y=0.45
+ $X2=2.6 $Y2=0.45
r132 20 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=2.275
+ $X2=3.355 $Y2=2.19
r133 20 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.27 $Y=2.275
+ $X2=2.5 $Y2=2.275
r134 18 37 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.41
+ $X2=3.695 $Y2=1.41
r135 18 19 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.83 $Y=1.41
+ $X2=3.905 $Y2=1.41
r136 16 17 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.94 $Y=0.95
+ $X2=3.94 $Y2=1.1
r137 15 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.975 $Y=0.555
+ $X2=3.975 $Y2=0.95
r138 9 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.905 $Y=1.545
+ $X2=3.905 $Y2=1.41
r139 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.905 $Y=1.545
+ $X2=3.905 $Y2=2.11
r140 8 19 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.905 $Y=1.275
+ $X2=3.905 $Y2=1.41
r141 8 17 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.905 $Y=1.275
+ $X2=3.905 $Y2=1.1
r142 2 22 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=2.065 $X2=2.5 $Y2=2.275
r143 1 26 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.6 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_1059_315# 1 2 9 13 17 19 21 24 26 28 29 30
+ 32 37 40 42 43 44 45 46 47 50 54 58 61 63 66 70 71 72
c147 45 0 1.49613e-19 $X=8.257 $Y=1.515
c148 44 0 1.20328e-19 $X=8.235 $Y=1.16
c149 30 0 2.70314e-19 $X=7.35 $Y=1.16
c150 13 0 2.06462e-20 $X=5.485 $Y=0.445
r151 81 82 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=7.265 $Y=1.16
+ $X2=7.275 $Y2=1.16
r152 73 75 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.37 $Y=1.74
+ $X2=5.485 $Y2=1.74
r153 67 81 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=6.855 $Y=1.16
+ $X2=7.265 $Y2=1.16
r154 67 78 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.855 $Y=1.16
+ $X2=6.845 $Y2=1.16
r155 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.855
+ $Y=1.16 $X2=6.855 $Y2=1.16
r156 64 72 0.463323 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=6.39 $Y=1.16 $X2=6.29
+ $Y2=1.16
r157 64 66 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.39 $Y=1.16
+ $X2=6.855 $Y2=1.16
r158 63 70 6.82437 $w=2.65e-07 $l=2.21346e-07 $layer=LI1_cond $X=6.285 $Y=1.53
+ $X2=6.21 $Y2=1.717
r159 62 72 7.80489 $w=1.95e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.285 $Y=1.325
+ $X2=6.29 $Y2=1.16
r160 62 63 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=6.285 $Y=1.325
+ $X2=6.285 $Y2=1.53
r161 61 72 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=6.29 $Y=0.995
+ $X2=6.29 $Y2=1.16
r162 61 71 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=6.29 $Y=0.995
+ $X2=6.29 $Y2=0.825
r163 56 71 7.53752 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=0.66
+ $X2=6.225 $Y2=0.825
r164 56 58 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.225 $Y=0.66
+ $X2=6.225 $Y2=0.385
r165 52 70 6.82437 $w=2.65e-07 $l=1.88e-07 $layer=LI1_cond $X=6.21 $Y=1.905
+ $X2=6.21 $Y2=1.717
r166 52 54 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=6.21 $Y=1.905
+ $X2=6.21 $Y2=2.34
r167 50 75 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.565 $Y=1.74
+ $X2=5.485 $Y2=1.74
r168 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.565
+ $Y=1.74 $X2=5.565 $Y2=1.74
r169 47 70 0.127723 $w=3.75e-07 $l=1.7e-07 $layer=LI1_cond $X=6.04 $Y=1.717
+ $X2=6.21 $Y2=1.717
r170 47 49 14.5976 $w=3.73e-07 $l=4.75e-07 $layer=LI1_cond $X=6.04 $Y=1.717
+ $X2=5.565 $Y2=1.717
r171 45 46 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=8.257 $Y=1.515
+ $X2=8.257 $Y2=1.665
r172 42 43 40.8095 $w=1.95e-07 $l=1.2e-07 $layer=POLY_cond $X=8.257 $Y=0.73
+ $X2=8.257 $Y2=0.85
r173 40 46 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=8.28 $Y=2.165
+ $X2=8.28 $Y2=1.665
r174 37 42 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.28 $Y=0.445
+ $X2=8.28 $Y2=0.73
r175 33 44 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=1.325
+ $X2=8.235 $Y2=1.16
r176 33 45 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.235 $Y=1.325
+ $X2=8.235 $Y2=1.515
r177 32 44 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=0.995
+ $X2=8.235 $Y2=1.16
r178 32 43 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.235 $Y=0.995
+ $X2=8.235 $Y2=0.85
r179 30 82 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.35 $Y=1.16
+ $X2=7.275 $Y2=1.16
r180 29 44 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.16 $Y=1.16
+ $X2=8.235 $Y2=1.16
r181 29 30 141.638 $w=3.3e-07 $l=8.1e-07 $layer=POLY_cond $X=8.16 $Y=1.16
+ $X2=7.35 $Y2=1.16
r182 26 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.275 $Y=0.995
+ $X2=7.275 $Y2=1.16
r183 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.275 $Y=0.995
+ $X2=7.275 $Y2=0.56
r184 22 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.265 $Y=1.325
+ $X2=7.265 $Y2=1.16
r185 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.265 $Y=1.325
+ $X2=7.265 $Y2=1.985
r186 19 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.855 $Y=0.995
+ $X2=6.855 $Y2=1.16
r187 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.855 $Y=0.995
+ $X2=6.855 $Y2=0.56
r188 15 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=1.325
+ $X2=6.845 $Y2=1.16
r189 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.845 $Y=1.325
+ $X2=6.845 $Y2=1.985
r190 11 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=1.575
+ $X2=5.485 $Y2=1.74
r191 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=5.485 $Y=1.575
+ $X2=5.485 $Y2=0.445
r192 7 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.37 $Y=1.905
+ $X2=5.37 $Y2=1.74
r193 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.37 $Y=1.905
+ $X2=5.37 $Y2=2.275
r194 2 70 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.08
+ $Y=1.485 $X2=6.205 $Y2=1.63
r195 2 54 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=6.08
+ $Y=1.485 $X2=6.205 $Y2=2.34
r196 1 58 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=6.1
+ $Y=0.235 $X2=6.225 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_891_413# 1 2 9 11 13 14 15 16 20 25 27 30
+ 33
c82 33 0 1.78258e-19 $X=5.225 $Y=1.16
c83 30 0 9.97377e-20 $X=5.935 $Y=1.16
c84 15 0 1.26047e-19 $X=6.43 $Y=1.16
c85 11 0 1.81857e-19 $X=6.435 $Y=0.995
r86 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.935
+ $Y=1.16 $X2=5.935 $Y2=1.16
r87 28 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=1.16
+ $X2=5.225 $Y2=1.16
r88 28 30 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=5.31 $Y=1.16
+ $X2=5.935 $Y2=1.16
r89 26 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=1.325
+ $X2=5.225 $Y2=1.16
r90 26 27 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.225 $Y=1.325
+ $X2=5.225 $Y2=2.165
r91 25 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0.995
+ $X2=5.225 $Y2=1.16
r92 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.225 $Y=0.535
+ $X2=5.225 $Y2=0.995
r93 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=0.45
+ $X2=5.225 $Y2=0.535
r94 20 22 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.14 $Y=0.45
+ $X2=4.705 $Y2=0.45
r95 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.14 $Y=2.25
+ $X2=5.225 $Y2=2.165
r96 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.14 $Y=2.25
+ $X2=4.59 $Y2=2.25
r97 14 31 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=6.35 $Y=1.16
+ $X2=5.935 $Y2=1.16
r98 14 15 5.03009 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=6.35 $Y=1.16 $X2=6.43
+ $Y2=1.16
r99 11 15 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=6.435 $Y=0.995
+ $X2=6.43 $Y2=1.16
r100 11 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.435 $Y=0.995
+ $X2=6.435 $Y2=0.56
r101 7 15 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=6.425 $Y=1.325
+ $X2=6.43 $Y2=1.16
r102 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.425 $Y=1.325
+ $X2=6.425 $Y2=1.985
r103 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=2.065 $X2=4.59 $Y2=2.25
r104 1 22 182 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_NDIFF $count=1 $X=4.555
+ $Y=0.235 $X2=4.705 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_1589_47# 1 2 7 9 12 14 16 19 21 23 26 31
+ 35 38 39 43
r77 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.765 $Y=1.16
+ $X2=9.185 $Y2=1.16
r78 35 37 5.29728 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=8.035 $Y=0.51
+ $X2=8.035 $Y2=0.615
r79 32 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.675 $Y=1.16
+ $X2=8.765 $Y2=1.16
r80 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.675
+ $Y=1.16 $X2=8.675 $Y2=1.16
r81 29 39 0.153733 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=8.235 $Y=1.16
+ $X2=8.1 $Y2=1.16
r82 29 31 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=8.235 $Y=1.16
+ $X2=8.675 $Y2=1.16
r83 27 39 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=8.1 $Y=1.325 $X2=8.1
+ $Y2=1.16
r84 27 38 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.1 $Y=1.325 $X2=8.1
+ $Y2=1.715
r85 26 39 6.7841 $w=2.35e-07 $l=1.81659e-07 $layer=LI1_cond $X=8.065 $Y=0.995
+ $X2=8.1 $Y2=1.16
r86 26 37 21.0727 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=8.065 $Y=0.995
+ $X2=8.065 $Y2=0.615
r87 21 38 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=1.88
+ $X2=8.07 $Y2=1.715
r88 21 23 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=8.07 $Y=1.88 $X2=8.07
+ $Y2=2
r89 17 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.185 $Y=1.325
+ $X2=9.185 $Y2=1.16
r90 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.185 $Y=1.325
+ $X2=9.185 $Y2=1.985
r91 14 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.185 $Y=0.995
+ $X2=9.185 $Y2=1.16
r92 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.185 $Y=0.995
+ $X2=9.185 $Y2=0.56
r93 10 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=1.325
+ $X2=8.765 $Y2=1.16
r94 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.765 $Y=1.325
+ $X2=8.765 $Y2=1.985
r95 7 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=0.995
+ $X2=8.765 $Y2=1.16
r96 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.765 $Y=0.995
+ $X2=8.765 $Y2=0.56
r97 2 23 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=7.945
+ $Y=1.845 $X2=8.07 $Y2=2
r98 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=7.945
+ $Y=0.235 $X2=8.07 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 55
+ 57 62 63 65 66 68 69 71 72 73 75 80 104 108 114 117 120 124
c147 124 0 1.81794e-19 $X=9.43 $Y=2.72
c148 51 0 1.49613e-19 $X=8.555 $Y=1.66
c149 1 0 3.29888e-20 $X=0.545 $Y=1.815
r150 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r151 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r152 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r153 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 112 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r155 112 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r156 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r157 109 120 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=8.64 $Y=2.72
+ $X2=8.532 $Y2=2.72
r158 109 111 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.64 $Y=2.72
+ $X2=8.97 $Y2=2.72
r159 108 123 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=9.315 $Y=2.72
+ $X2=9.487 $Y2=2.72
r160 108 111 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.315 $Y=2.72
+ $X2=8.97 $Y2=2.72
r161 107 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r162 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r163 104 120 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=8.425 $Y=2.72
+ $X2=8.532 $Y2=2.72
r164 104 106 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.425 $Y=2.72
+ $X2=8.05 $Y2=2.72
r165 103 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r166 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r167 100 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r168 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r169 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r170 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r171 94 97 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r172 93 96 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r173 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r174 91 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r175 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r176 88 91 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r177 88 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r178 87 90 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r179 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r180 85 117 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.572 $Y2=2.72
r181 85 87 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=2.07 $Y2=2.72
r182 84 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r183 84 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r185 81 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r186 81 83 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r187 80 117 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.572 $Y2=2.72
r188 80 83 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.15 $Y2=2.72
r189 75 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r190 75 77 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r191 73 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r192 73 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r193 71 102 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.39 $Y=2.72
+ $X2=7.13 $Y2=2.72
r194 71 72 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=7.39 $Y=2.72
+ $X2=7.477 $Y2=2.72
r195 70 106 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=7.565 $Y=2.72
+ $X2=8.05 $Y2=2.72
r196 70 72 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=7.565 $Y=2.72
+ $X2=7.477 $Y2=2.72
r197 68 99 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.55 $Y=2.72
+ $X2=6.21 $Y2=2.72
r198 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=2.72
+ $X2=6.635 $Y2=2.72
r199 67 102 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.72 $Y=2.72
+ $X2=7.13 $Y2=2.72
r200 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.72 $Y=2.72
+ $X2=6.635 $Y2=2.72
r201 65 96 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.49 $Y=2.72 $X2=5.29
+ $Y2=2.72
r202 65 66 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=5.49 $Y=2.72
+ $X2=5.647 $Y2=2.72
r203 64 99 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.805 $Y=2.72
+ $X2=6.21 $Y2=2.72
r204 64 66 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=5.805 $Y=2.72
+ $X2=5.647 $Y2=2.72
r205 62 90 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r206 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=2.72
+ $X2=3.695 $Y2=2.72
r207 61 93 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.91 $Y2=2.72
r208 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=2.72
+ $X2=3.695 $Y2=2.72
r209 57 60 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=9.44 $Y=1.66
+ $X2=9.44 $Y2=2.34
r210 55 123 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=9.44 $Y=2.635
+ $X2=9.487 $Y2=2.72
r211 55 60 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.44 $Y=2.635
+ $X2=9.44 $Y2=2.34
r212 51 54 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=8.532 $Y=1.66
+ $X2=8.532 $Y2=2
r213 49 120 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.532 $Y=2.635
+ $X2=8.532 $Y2=2.72
r214 49 54 34.0373 $w=2.13e-07 $l=6.35e-07 $layer=LI1_cond $X=8.532 $Y=2.635
+ $X2=8.532 $Y2=2
r215 45 72 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.477 $Y=2.635
+ $X2=7.477 $Y2=2.72
r216 45 47 47.5325 $w=1.73e-07 $l=7.5e-07 $layer=LI1_cond $X=7.477 $Y=2.635
+ $X2=7.477 $Y2=1.885
r217 41 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.635 $Y=2.635
+ $X2=6.635 $Y2=2.72
r218 41 43 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=6.635 $Y=2.635
+ $X2=6.635 $Y2=1.79
r219 37 66 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.647 $Y=2.635
+ $X2=5.647 $Y2=2.72
r220 37 39 12.2561 $w=3.13e-07 $l=3.35e-07 $layer=LI1_cond $X=5.647 $Y=2.635
+ $X2=5.647 $Y2=2.3
r221 33 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2.72
r222 33 35 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.695 $Y=2.635
+ $X2=3.695 $Y2=2
r223 29 117 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.572 $Y=2.635
+ $X2=1.572 $Y2=2.72
r224 29 31 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.572 $Y=2.635
+ $X2=1.572 $Y2=2.34
r225 25 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r226 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r227 8 60 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.26
+ $Y=1.485 $X2=9.4 $Y2=2.34
r228 8 57 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=9.26
+ $Y=1.485 $X2=9.4 $Y2=1.66
r229 7 54 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=8.355
+ $Y=1.845 $X2=8.555 $Y2=2
r230 7 51 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=8.355
+ $Y=1.845 $X2=8.555 $Y2=1.66
r231 6 47 300 $w=1.7e-07 $l=4.62601e-07 $layer=licon1_PDIFF $count=2 $X=7.34
+ $Y=1.485 $X2=7.475 $Y2=1.885
r232 5 43 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=6.5
+ $Y=1.485 $X2=6.635 $Y2=1.79
r233 4 39 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=2.065 $X2=5.585 $Y2=2.3
r234 3 35 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=3.32
+ $Y=2.065 $X2=3.695 $Y2=2
r235 2 31 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.065 $X2=1.62 $Y2=2.34
r236 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%A_381_47# 1 2 13 15 16 17 18 21
c49 18 0 1.74123e-19 $X=1.972 $Y=2.04
c50 15 0 1.97281e-19 $X=1.932 $Y=0.675
r51 17 18 7.17986 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.972 $Y=1.91
+ $X2=1.972 $Y2=2.04
r52 16 17 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=1.905 $Y=0.805
+ $X2=1.905 $Y2=1.91
r53 15 16 6.65856 $w=2.23e-07 $l=1.3e-07 $layer=LI1_cond $X=1.932 $Y=0.675
+ $X2=1.932 $Y2=0.805
r54 13 18 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2 $Y=2.3 $X2=2
+ $Y2=2.04
r55 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.535
+ $X2=1.96 $Y2=0.45
r56 9 15 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.96 $Y=0.535
+ $X2=1.96 $Y2=0.675
r57 2 13 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.065 $X2=2.04 $Y2=2.3
r58 1 21 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.045 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%Q 1 2 9 14 15 16 19
c38 19 0 1.81857e-19 $X=7.065 $Y=0.395
c39 14 0 1.26047e-19 $X=7.205 $Y=1.445
r40 16 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.065 $Y=0.51
+ $X2=7.065 $Y2=0.395
r41 15 16 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=7.065 $Y=0.74
+ $X2=7.065 $Y2=0.51
r42 13 15 4.35714 $w=3.5e-07 $l=1.92614e-07 $layer=LI1_cond $X=7.205 $Y=0.865
+ $X2=7.065 $Y2=0.74
r43 13 14 33.8565 $w=1.88e-07 $l=5.8e-07 $layer=LI1_cond $X=7.205 $Y=0.865
+ $X2=7.205 $Y2=1.445
r44 9 11 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.055 $Y=1.63
+ $X2=7.055 $Y2=2.31
r45 7 14 4.63743 $w=3.42e-07 $l=2.04939e-07 $layer=LI1_cond $X=7.055 $Y=1.575
+ $X2=7.205 $Y2=1.445
r46 7 9 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=7.055 $Y=1.575
+ $X2=7.055 $Y2=1.63
r47 2 11 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.485 $X2=7.055 $Y2=2.31
r48 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.485 $X2=7.055 $Y2=1.63
r49 1 19 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=6.93
+ $Y=0.235 $X2=7.065 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%Q_N 1 2 9 13 14 23 25
c20 23 0 1.20328e-19 $X=8.977 $Y=1.495
r21 17 25 1.78887 $w=3.33e-07 $l=5.2e-08 $layer=LI1_cond $X=8.977 $Y=1.662
+ $X2=8.977 $Y2=1.61
r22 14 25 0.653624 $w=3.33e-07 $l=1.9e-08 $layer=LI1_cond $X=8.977 $Y=1.591
+ $X2=8.977 $Y2=1.61
r23 14 23 4.77693 $w=3.33e-07 $l=9.6e-08 $layer=LI1_cond $X=8.977 $Y=1.591
+ $X2=8.977 $Y2=1.495
r24 14 20 22.8425 $w=3.33e-07 $l=6.64e-07 $layer=LI1_cond $X=8.977 $Y=1.676
+ $X2=8.977 $Y2=2.34
r25 14 17 0.481618 $w=3.33e-07 $l=1.4e-08 $layer=LI1_cond $X=8.977 $Y=1.676
+ $X2=8.977 $Y2=1.662
r26 13 23 32.6972 $w=2.13e-07 $l=6.1e-07 $layer=LI1_cond $X=9.037 $Y=0.885
+ $X2=9.037 $Y2=1.495
r27 7 13 6.05672 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=9.017 $Y=0.758
+ $X2=9.017 $Y2=0.885
r28 7 9 8.49644 $w=2.53e-07 $l=1.88e-07 $layer=LI1_cond $X=9.017 $Y=0.758
+ $X2=9.017 $Y2=0.57
r29 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.84
+ $Y=1.485 $X2=8.975 $Y2=1.63
r30 2 20 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.84
+ $Y=1.485 $X2=8.975 $Y2=2.34
r31 1 9 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=8.84
+ $Y=0.235 $X2=8.975 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HD__DFXBP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 53
+ 55 58 59 61 62 64 65 66 68 73 78 96 100 106 109 112 115 119
c148 119 0 2.71124e-20 $X=9.43 $Y=0
c149 43 0 1.70577e-19 $X=6.645 $Y=0.53
r150 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r151 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r152 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r153 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r154 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r155 104 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r156 104 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=8.51 $Y2=0
r157 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r158 101 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.72 $Y=0
+ $X2=8.555 $Y2=0
r159 101 103 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.72 $Y=0
+ $X2=8.97 $Y2=0
r160 100 118 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=9.315 $Y=0
+ $X2=9.487 $Y2=0
r161 100 103 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.315 $Y=0
+ $X2=8.97 $Y2=0
r162 99 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r163 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r164 96 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.39 $Y=0
+ $X2=8.555 $Y2=0
r165 96 98 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.39 $Y=0 $X2=8.05
+ $Y2=0
r166 95 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r167 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r168 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r169 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r170 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r171 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r172 86 89 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r173 86 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=3.45 $Y2=0
r174 85 88 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r175 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r176 83 112 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.77 $Y=0
+ $X2=3.585 $Y2=0
r177 83 85 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.77 $Y=0 $X2=3.91
+ $Y2=0
r178 82 113 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r179 82 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r180 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r181 79 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=1.58 $Y2=0
r182 79 81 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r183 78 112 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.585
+ $Y2=0
r184 78 81 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.4 $Y=0 $X2=2.07
+ $Y2=0
r185 77 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r186 77 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r187 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r188 74 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r189 74 76 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r190 73 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.58 $Y2=0
r191 73 76 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r192 68 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r193 68 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r194 66 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r195 66 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r196 64 94 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.4 $Y=0 $X2=7.13
+ $Y2=0
r197 64 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0 $X2=7.485
+ $Y2=0
r198 63 98 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=7.57 $Y=0 $X2=8.05
+ $Y2=0
r199 63 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.57 $Y=0 $X2=7.485
+ $Y2=0
r200 61 91 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.21
+ $Y2=0
r201 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.645
+ $Y2=0
r202 60 94 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.73 $Y=0 $X2=7.13
+ $Y2=0
r203 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.73 $Y=0 $X2=6.645
+ $Y2=0
r204 58 88 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.585 $Y=0 $X2=5.29
+ $Y2=0
r205 58 59 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.585 $Y=0 $X2=5.69
+ $Y2=0
r206 57 91 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.795 $Y=0
+ $X2=6.21 $Y2=0
r207 57 59 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.69
+ $Y2=0
r208 53 118 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=9.44 $Y=0.085
+ $X2=9.487 $Y2=0
r209 53 55 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.44 $Y=0.085
+ $X2=9.44 $Y2=0.38
r210 49 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=0.085
+ $X2=8.555 $Y2=0
r211 49 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.555 $Y=0.085
+ $X2=8.555 $Y2=0.38
r212 45 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0
r213 45 47 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0.435
r214 41 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=0.085
+ $X2=6.645 $Y2=0
r215 41 43 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.645 $Y=0.085
+ $X2=6.645 $Y2=0.53
r216 37 59 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.69 $Y=0.085
+ $X2=5.69 $Y2=0
r217 37 39 19.2771 $w=2.08e-07 $l=3.65e-07 $layer=LI1_cond $X=5.69 $Y=0.085
+ $X2=5.69 $Y2=0.45
r218 33 112 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0
r219 33 35 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0.42
r220 29 109 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r221 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.38
r222 25 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r223 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r224 8 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.26
+ $Y=0.235 $X2=9.4 $Y2=0.38
r225 7 51 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=8.355
+ $Y=0.235 $X2=8.555 $Y2=0.38
r226 6 47 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=7.35
+ $Y=0.235 $X2=7.485 $Y2=0.435
r227 5 43 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=6.51
+ $Y=0.235 $X2=6.645 $Y2=0.53
r228 4 39 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.235 $X2=5.695 $Y2=0.45
r229 3 35 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.235 $X2=3.595 $Y2=0.42
r230 2 31 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r231 1 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__fa_1.pex.spice
* Created: Thu Aug 27 14:21:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__FA_1%A_76_199# 1 2 9 12 16 20 25 26 27 30 33 34 35
+ 38 39 42 45 49 52 53
c168 52 0 5.62553e-20 $X=4.96 $Y=1.04
c169 45 0 3.78383e-20 $X=5.315 $Y=0.85
c170 42 0 2.631e-19 $X=1.615 $Y=0.85
c171 39 0 3.35934e-19 $X=1.76 $Y=0.85
c172 33 0 1.32337e-19 $X=0.515 $Y=1.16
c173 25 0 1.92424e-19 $X=0.6 $Y=1.625
r174 52 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.96 $Y=1.04
+ $X2=4.96 $Y2=1.205
r175 52 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.96 $Y=1.04
+ $X2=4.96 $Y2=0.875
r176 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.96
+ $Y=1.04 $X2=4.96 $Y2=1.04
r177 46 53 13.926 $w=3.11e-07 $l=3.99687e-07 $layer=LI1_cond $X=5.315 $Y=0.945
+ $X2=4.96 $Y2=1.04
r178 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.315 $Y=0.85
+ $X2=5.315 $Y2=0.85
r179 42 58 0.202658 $w=6.02e-07 $l=1e-08 $layer=LI1_cond $X=1.615 $Y=0.595
+ $X2=1.625 $Y2=0.595
r180 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.615 $Y=0.85
+ $X2=1.615 $Y2=0.85
r181 39 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.76 $Y=0.85
+ $X2=1.615 $Y2=0.85
r182 38 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.17 $Y=0.85
+ $X2=5.315 $Y2=0.85
r183 38 39 4.22029 $w=1.4e-07 $l=3.41e-06 $layer=MET1_cond $X=5.17 $Y=0.85
+ $X2=1.76 $Y2=0.85
r184 34 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r185 34 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r186 33 36 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.557 $Y=1.16
+ $X2=0.557 $Y2=1.325
r187 33 35 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.557 $Y=1.16
+ $X2=0.557 $Y2=0.995
r188 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r189 28 30 14.9818 $w=3.98e-07 $l=5.2e-07 $layer=LI1_cond $X=1.105 $Y=2.265
+ $X2=1.625 $Y2=2.265
r190 26 42 17.2629 $w=6.02e-07 $l=5.64048e-07 $layer=LI1_cond $X=1.11 $Y=0.72
+ $X2=1.615 $Y2=0.595
r191 26 27 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.11 $Y=0.72
+ $X2=0.685 $Y2=0.72
r192 25 28 26.5188 $w=3.3e-07 $l=8.56037e-07 $layer=LI1_cond $X=0.6 $Y=1.625
+ $X2=1.105 $Y2=2.265
r193 25 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.6 $Y=1.625 $X2=0.6
+ $Y2=1.325
r194 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=0.805
+ $X2=0.685 $Y2=0.72
r195 22 35 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.6 $Y=0.805
+ $X2=0.6 $Y2=0.995
r196 20 55 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=4.9 $Y=2.275
+ $X2=4.9 $Y2=1.205
r197 16 54 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.9 $Y=0.445
+ $X2=4.9 $Y2=0.875
r198 12 50 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r199 9 49 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
r200 2 30 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=2.065 $X2=1.625 $Y2=2.275
r201 1 58 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.235 $X2=1.625 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%A 3 7 11 15 19 23 27 31 33 35 36 37 38 39 40 47
+ 52 56 61 66 67 71 72
c242 67 0 3.78383e-20 $X=4.46 $Y=1.04
c243 56 0 1.52202e-19 $X=0.995 $Y=1.16
c244 38 0 3.10095e-19 $X=2.68 $Y=1.19
c245 37 0 1.34551e-19 $X=4.25 $Y=1.19
c246 11 0 1.9888e-19 $X=2.255 $Y=0.445
c247 7 0 1.39992e-19 $X=0.965 $Y=2.275
c248 3 0 1.37054e-19 $X=0.965 $Y=0.445
r249 71 74 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.12
+ $X2=6.16 $Y2=1.285
r250 71 73 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.12
+ $X2=6.16 $Y2=0.955
r251 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.16
+ $Y=1.12 $X2=6.16 $Y2=1.12
r252 66 69 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.46 $Y=1.04
+ $X2=4.46 $Y2=1.205
r253 66 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.46 $Y=1.04
+ $X2=4.46 $Y2=0.875
r254 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.46
+ $Y=1.04 $X2=4.46 $Y2=1.04
r255 61 64 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.195
+ $X2=2.315 $Y2=1.36
r256 61 63 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.195
+ $X2=2.315 $Y2=1.03
r257 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.315
+ $Y=1.195 $X2=2.315 $Y2=1.195
r258 56 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=1.325
r259 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=0.995
r260 52 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.235 $Y=1.19
+ $X2=6.235 $Y2=1.19
r261 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.395 $Y=1.19
+ $X2=4.395 $Y2=1.19
r262 47 62 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.535 $Y=1.195
+ $X2=2.315 $Y2=1.195
r263 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.535 $Y=1.19
+ $X2=2.535 $Y2=1.19
r264 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.54 $Y=1.19
+ $X2=4.395 $Y2=1.19
r265 39 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.09 $Y=1.19
+ $X2=6.235 $Y2=1.19
r266 39 40 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=6.09 $Y=1.19
+ $X2=4.54 $Y2=1.19
r267 38 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.68 $Y=1.19
+ $X2=2.535 $Y2=1.19
r268 37 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.25 $Y=1.19
+ $X2=4.395 $Y2=1.19
r269 37 38 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=4.25 $Y=1.19
+ $X2=2.68 $Y2=1.19
r270 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.19
+ $X2=1.155 $Y2=1.19
r271 35 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.39 $Y=1.19
+ $X2=2.535 $Y2=1.19
r272 35 36 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=2.39 $Y=1.19
+ $X2=1.3 $Y2=1.19
r273 33 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.16 $X2=0.995 $Y2=1.16
r274 33 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.19
+ $X2=1.155 $Y2=1.19
r275 31 74 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=6.22 $Y=2.275
+ $X2=6.22 $Y2=1.285
r276 27 73 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.22 $Y=0.445
+ $X2=6.22 $Y2=0.955
r277 23 69 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=4.455 $Y=2.275
+ $X2=4.455 $Y2=1.205
r278 19 68 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.455 $Y=0.445
+ $X2=4.455 $Y2=0.875
r279 15 64 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.255 $Y=2.275
+ $X2=2.255 $Y2=1.36
r280 11 63 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=2.255 $Y=0.445
+ $X2=2.255 $Y2=1.03
r281 7 59 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.965 $Y=2.275
+ $X2=0.965 $Y2=1.325
r282 3 58 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.965 $Y=0.445
+ $X2=0.965 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%B 3 7 9 11 12 14 15 16 17 18 23 24 26 29 33 35
+ 36 38 40 42 44 45 46 47 54 56 57 60 63 68
c223 63 0 2.96357e-19 $X=1.385 $Y=1.715
c224 45 0 2.54181e-19 $X=1.76 $Y=1.53
r225 68 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=1.68
+ $X2=5.8 $Y2=1.845
r226 68 70 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=1.68
+ $X2=5.8 $Y2=1.515
r227 63 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.715
+ $X2=1.385 $Y2=1.88
r228 63 65 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.715
+ $X2=1.385 $Y2=1.55
r229 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=1.715 $X2=1.385 $Y2=1.715
r230 57 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.8
+ $Y=1.68 $X2=5.8 $Y2=1.68
r231 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.775 $Y=1.53
+ $X2=5.775 $Y2=1.53
r232 54 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=1.6 $X2=3.45 $Y2=1.6
r233 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.475 $Y=1.53
+ $X2=3.475 $Y2=1.53
r234 47 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.62 $Y=1.53
+ $X2=3.475 $Y2=1.53
r235 46 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.63 $Y=1.53
+ $X2=5.775 $Y2=1.53
r236 46 47 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=5.63 $Y=1.53
+ $X2=3.62 $Y2=1.53
r237 45 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.76 $Y=1.53
+ $X2=1.615 $Y2=1.53
r238 44 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.33 $Y=1.53
+ $X2=3.475 $Y2=1.53
r239 44 45 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=3.33 $Y=1.53
+ $X2=1.76 $Y2=1.53
r240 42 64 6.09338 $w=4.33e-07 $l=2.3e-07 $layer=LI1_cond $X=1.615 $Y=1.662
+ $X2=1.385 $Y2=1.662
r241 42 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.615 $Y=1.53
+ $X2=1.615 $Y2=1.53
r242 37 60 43.2782 $w=3.2e-07 $l=2.4e-07 $layer=POLY_cond $X=3.475 $Y=1.84
+ $X2=3.475 $Y2=1.6
r243 37 38 13.8458 $w=2.35e-07 $l=8.74643e-08 $layer=POLY_cond $X=3.475 $Y=1.84
+ $X2=3.502 $Y2=1.915
r244 36 41 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.56 $Y=1.435
+ $X2=3.56 $Y2=0.955
r245 35 60 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=3.475 $Y=1.595
+ $X2=3.475 $Y2=1.6
r246 35 36 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=3.475 $Y=1.595
+ $X2=3.475 $Y2=1.435
r247 33 71 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.74 $Y=2.275
+ $X2=5.74 $Y2=1.845
r248 29 70 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=5.74 $Y=0.445
+ $X2=5.74 $Y2=1.515
r249 24 38 13.8458 $w=2.35e-07 $l=1.45753e-07 $layer=POLY_cond $X=3.615 $Y=1.99
+ $X2=3.502 $Y2=1.915
r250 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.615 $Y=1.99
+ $X2=3.615 $Y2=2.275
r251 23 40 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.615 $Y=0.445
+ $X2=3.615 $Y2=0.73
r252 17 38 11.8488 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.315 $Y=1.915
+ $X2=3.502 $Y2=1.915
r253 17 18 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.315 $Y=1.915
+ $X2=2.75 $Y2=1.915
r254 15 41 53.4216 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=3.587 $Y=0.805
+ $X2=3.587 $Y2=0.955
r255 15 40 29.1598 $w=2.05e-07 $l=7.5e-08 $layer=POLY_cond $X=3.587 $Y=0.805
+ $X2=3.587 $Y2=0.73
r256 15 16 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=3.485 $Y=0.805
+ $X2=2.75 $Y2=0.805
r257 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.675 $Y=1.99
+ $X2=2.75 $Y2=1.915
r258 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.675 $Y=1.99
+ $X2=2.675 $Y2=2.275
r259 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.675 $Y=0.73
+ $X2=2.75 $Y2=0.805
r260 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.675 $Y=0.73
+ $X2=2.675 $Y2=0.445
r261 7 66 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.415 $Y=2.275
+ $X2=1.415 $Y2=1.88
r262 3 65 566.606 $w=1.5e-07 $l=1.105e-06 $layer=POLY_cond $X=1.415 $Y=0.445
+ $X2=1.415 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%CIN 3 7 11 14 20 24 26 27 29 30 31 33 34 35 37
+ 38 39 42 45 47 49 53 55 59
c225 47 0 1.55247e-19 $X=1.955 $Y=1.19
c226 45 0 3.34578e-20 $X=1.835 $Y=1.19
c227 42 0 2.4081e-20 $X=4.035 $Y=1.6
c228 31 0 1.34126e-19 $X=2.04 $Y=1.68
c229 29 0 2.06181e-19 $X=1.955 $Y=1.595
c230 27 0 1.32582e-20 $X=4.037 $Y=0.88
r231 56 59 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.28 $Y=1.68 $X2=5.28
+ $Y2=1.6
r232 55 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.68
+ $X2=5.32 $Y2=1.845
r233 55 57 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.68
+ $X2=5.32 $Y2=1.515
r234 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.32
+ $Y=1.68 $X2=5.32 $Y2=1.68
r235 49 56 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=5.28 $Y=1.87
+ $X2=5.28 $Y2=1.68
r236 44 47 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.835 $Y=1.19
+ $X2=1.955 $Y2=1.19
r237 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=1.19 $X2=1.835 $Y2=1.19
r238 42 53 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.035 $Y=1.6
+ $X2=4.035 $Y2=1.435
r239 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=1.6 $X2=4.035 $Y2=1.6
r240 39 41 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.955 $Y=1.6
+ $X2=4.035 $Y2=1.6
r241 38 59 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=1.6
+ $X2=5.28 $Y2=1.6
r242 38 41 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=5.155 $Y=1.6
+ $X2=4.035 $Y2=1.6
r243 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.87 $Y=1.515
+ $X2=3.955 $Y2=1.6
r244 36 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.87 $Y=1.25
+ $X2=3.87 $Y2=1.515
r245 34 36 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.785 $Y=1.107
+ $X2=3.87 $Y2=1.25
r246 34 35 33.3602 $w=2.83e-07 $l=8.25e-07 $layer=LI1_cond $X=3.785 $Y=1.107
+ $X2=2.96 $Y2=1.107
r247 32 35 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=2.875 $Y=1.25
+ $X2=2.96 $Y2=1.107
r248 32 33 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=1.25
+ $X2=2.875 $Y2=1.595
r249 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.79 $Y=1.68
+ $X2=2.875 $Y2=1.595
r250 30 31 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.79 $Y=1.68
+ $X2=2.04 $Y2=1.68
r251 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=1.595
+ $X2=2.04 $Y2=1.68
r252 28 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.275
+ $X2=1.955 $Y2=1.19
r253 28 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.955 $Y=1.275
+ $X2=1.955 $Y2=1.595
r254 27 53 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.04 $Y=0.88
+ $X2=4.04 $Y2=1.435
r255 26 27 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=4.037 $Y=0.73
+ $X2=4.037 $Y2=0.88
r256 24 58 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.38 $Y=2.275
+ $X2=5.38 $Y2=1.845
r257 20 57 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=5.38 $Y=0.445
+ $X2=5.38 $Y2=1.515
r258 12 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.035 $Y=1.765
+ $X2=4.035 $Y2=1.6
r259 12 14 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.035 $Y=1.765
+ $X2=4.035 $Y2=2.275
r260 11 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.035 $Y=0.445
+ $X2=4.035 $Y2=0.73
r261 5 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.355
+ $X2=1.835 $Y2=1.19
r262 5 7 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.835 $Y=1.355
+ $X2=1.835 $Y2=2.275
r263 1 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.025
+ $X2=1.835 $Y2=1.19
r264 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.835 $Y=1.025
+ $X2=1.835 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%A_995_47# 1 2 9 12 14 18 20 22 27 31 36 41 42
+ 43 46
c95 31 0 5.62553e-20 $X=5.255 $Y=0.425
r96 42 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.655 $Y=1.16
+ $X2=6.655 $Y2=1.325
r97 42 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.655 $Y=1.16
+ $X2=6.655 $Y2=0.995
r98 41 44 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=6.617 $Y=1.16
+ $X2=6.617 $Y2=1.325
r99 41 43 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=6.617 $Y=1.16
+ $X2=6.617 $Y2=0.995
r100 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.655
+ $Y=1.16 $X2=6.655 $Y2=1.16
r101 29 31 3.71115 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=0.425
+ $X2=5.255 $Y2=0.425
r102 27 44 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.58 $Y=1.935
+ $X2=6.58 $Y2=1.325
r103 24 43 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.58 $Y=0.785
+ $X2=6.58 $Y2=0.995
r104 23 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=2.02
+ $X2=6.085 $Y2=2.02
r105 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.495 $Y=2.02
+ $X2=6.58 $Y2=1.935
r106 22 23 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.495 $Y=2.02
+ $X2=6.17 $Y2=2.02
r107 21 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.095 $Y=0.7
+ $X2=6.01 $Y2=0.7
r108 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.495 $Y=0.7
+ $X2=6.58 $Y2=0.785
r109 20 21 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.495 $Y=0.7
+ $X2=6.095 $Y2=0.7
r110 18 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.01 $Y=0.38
+ $X2=6.01 $Y2=0.7
r111 18 31 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.925 $Y=0.38
+ $X2=5.255 $Y2=0.38
r112 14 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.085 $Y=2.295
+ $X2=6.085 $Y2=2.02
r113 14 16 28.1332 $w=3.38e-07 $l=8.3e-07 $layer=LI1_cond $X=6 $Y=2.295 $X2=5.17
+ $Y2=2.295
r114 12 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.715 $Y=1.985
+ $X2=6.715 $Y2=1.325
r115 9 46 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.715 $Y=0.56
+ $X2=6.715 $Y2=0.995
r116 2 16 600 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=2.065 $X2=5.17 $Y2=2.3
r117 1 29 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.235 $X2=5.17 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%COUT 1 2 10 11 12 13 14 15 24
r18 14 15 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=2.21
r19 14 24 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.215 $Y2=1.775
r20 11 24 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=0.215 $Y=1.615
+ $X2=0.215 $Y2=1.775
r21 11 12 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=1.615
+ $X2=0.215 $Y2=1.485
r22 10 12 41.5117 $w=1.73e-07 $l=6.55e-07 $layer=LI1_cond $X=0.172 $Y=0.83
+ $X2=0.172 $Y2=1.485
r23 9 13 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=0.215 $Y=0.7 $X2=0.215
+ $Y2=0.51
r24 9 10 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=0.7
+ $X2=0.215 $Y2=0.83
r25 2 24 300 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.775
r26 1 13 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 39 41 43 48
+ 50 55 60 70 71 74 77 80 83
r114 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r116 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r117 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r119 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r120 68 84 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=4.37 $Y2=2.72
r121 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r122 65 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=2.72
+ $X2=4.245 $Y2=2.72
r123 65 67 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=4.41 $Y=2.72
+ $X2=6.21 $Y2=2.72
r124 64 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r125 64 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r126 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r127 61 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=2.72
+ $X2=3.405 $Y2=2.72
r128 61 63 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.57 $Y=2.72
+ $X2=3.91 $Y2=2.72
r129 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=2.72
+ $X2=4.245 $Y2=2.72
r130 60 63 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.08 $Y=2.72
+ $X2=3.91 $Y2=2.72
r131 59 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r132 59 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r133 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r134 56 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=2.72
+ $X2=2.465 $Y2=2.72
r135 56 58 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.63 $Y=2.72
+ $X2=2.99 $Y2=2.72
r136 55 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=2.72
+ $X2=3.405 $Y2=2.72
r137 55 58 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.24 $Y=2.72
+ $X2=2.99 $Y2=2.72
r138 54 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r139 54 75 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=0.69 $Y2=2.72
r140 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 51 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.64 $Y2=2.72
r142 51 53 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=2.07 $Y2=2.72
r143 50 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=2.72
+ $X2=2.465 $Y2=2.72
r144 50 53 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.3 $Y=2.72
+ $X2=2.07 $Y2=2.72
r145 43 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.64 $Y2=2.72
r146 41 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r147 41 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r148 39 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.515 $Y2=2.72
r149 39 48 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r150 37 67 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.21 $Y2=2.72
r151 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.505 $Y2=2.72
r152 36 70 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r153 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=6.505 $Y2=2.72
r154 32 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=2.635
+ $X2=6.505 $Y2=2.72
r155 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.505 $Y=2.635
+ $X2=6.505 $Y2=2.36
r156 28 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=2.635
+ $X2=4.245 $Y2=2.72
r157 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.245 $Y=2.635
+ $X2=4.245 $Y2=2.36
r158 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.405 $Y2=2.72
r159 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.405 $Y2=2.34
r160 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=2.635
+ $X2=2.465 $Y2=2.72
r161 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.465 $Y=2.635
+ $X2=2.465 $Y2=2.36
r162 16 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=2.635
+ $X2=0.64 $Y2=2.72
r163 16 18 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.64 $Y=2.635
+ $X2=0.64 $Y2=2.32
r164 5 34 600 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=2.065 $X2=6.505 $Y2=2.36
r165 4 30 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=4.11
+ $Y=2.065 $X2=4.245 $Y2=2.36
r166 3 26 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=2.065 $X2=3.405 $Y2=2.34
r167 2 22 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=2.065 $X2=2.465 $Y2=2.36
r168 1 18 600 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%A_382_413# 1 2 9 11 12 15
c27 12 0 3.34578e-20 $X=2.13 $Y=2.02
r28 13 15 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=2.917 $Y=2.105
+ $X2=2.917 $Y2=2.275
r29 11 13 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.8 $Y=2.02
+ $X2=2.917 $Y2=2.105
r30 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.8 $Y=2.02 $X2=2.13
+ $Y2=2.02
r31 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=2.105
+ $X2=2.13 $Y2=2.02
r32 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.045 $Y=2.105
+ $X2=2.045 $Y2=2.275
r33 2 15 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=2.75
+ $Y=2.065 $X2=2.885 $Y2=2.275
r34 1 9 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=2.065 $X2=2.045 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%A_738_413# 1 2 9 11 12 15
r26 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.665 $Y=2.105
+ $X2=4.665 $Y2=2.275
r27 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.58 $Y=2.02
+ $X2=4.665 $Y2=2.105
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.58 $Y=2.02
+ $X2=3.91 $Y2=2.02
r29 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.825 $Y=2.105
+ $X2=3.91 $Y2=2.02
r30 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.825 $Y=2.105
+ $X2=3.825 $Y2=2.275
r31 2 15 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=4.53
+ $Y=2.065 $X2=4.665 $Y2=2.275
r32 1 9 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=3.69
+ $Y=2.065 $X2=3.825 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%SUM 1 2 7 8 9 10 11 12 24 31 45
r15 45 46 1.68354 $w=3.98e-07 $l=4.5e-08 $layer=LI1_cond $X=7.04 $Y=1.53
+ $X2=7.04 $Y2=1.485
r16 29 31 2.16083 $w=3.98e-07 $l=7.5e-08 $layer=LI1_cond $X=7.04 $Y=1.685
+ $X2=7.04 $Y2=1.76
r17 24 43 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=7.075 $Y=0.85 $X2=7.075
+ $Y2=0.81
r18 11 12 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=7.04 $Y=1.87
+ $X2=7.04 $Y2=2.21
r19 11 31 3.16922 $w=3.98e-07 $l=1.1e-07 $layer=LI1_cond $X=7.04 $Y=1.87
+ $X2=7.04 $Y2=1.76
r20 10 29 3.8895 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=7.04 $Y=1.55
+ $X2=7.04 $Y2=1.685
r21 10 45 0.576222 $w=3.98e-07 $l=2e-08 $layer=LI1_cond $X=7.04 $Y=1.55 $X2=7.04
+ $Y2=1.53
r22 10 46 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=7.075 $Y=1.465
+ $X2=7.075 $Y2=1.485
r23 9 10 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.075 $Y=1.19
+ $X2=7.075 $Y2=1.465
r24 8 43 1.04969 $w=3.98e-07 $l=2.3e-08 $layer=LI1_cond $X=7.04 $Y=0.787
+ $X2=7.04 $Y2=0.81
r25 8 41 6.54011 $w=3.98e-07 $l=2.27e-07 $layer=LI1_cond $X=7.04 $Y=0.787
+ $X2=7.04 $Y2=0.56
r26 8 9 11.1054 $w=3.28e-07 $l=3.18e-07 $layer=LI1_cond $X=7.075 $Y=0.872
+ $X2=7.075 $Y2=1.19
r27 8 24 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=7.075 $Y=0.872
+ $X2=7.075 $Y2=0.85
r28 7 41 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=7.04 $Y=0.51 $X2=7.04
+ $Y2=0.56
r29 2 31 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=6.79
+ $Y=1.485 $X2=6.925 $Y2=1.76
r30 1 41 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=6.79
+ $Y=0.235 $X2=6.925 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 39 41 43 48
+ 50 58 63 73 74 77 80 83 86
r127 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r128 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r129 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r130 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r131 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r132 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r133 71 87 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=4.37 $Y2=0
r134 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r135 68 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.245
+ $Y2=0
r136 68 70 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=4.41 $Y=0 $X2=6.21
+ $Y2=0
r137 67 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r138 67 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r139 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r140 64 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.405
+ $Y2=0
r141 64 66 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.91
+ $Y2=0
r142 63 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=4.245
+ $Y2=0
r143 63 66 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.91
+ $Y2=0
r144 62 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r145 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r146 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r147 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.465
+ $Y2=0
r148 59 61 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.99
+ $Y2=0
r149 58 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.405
+ $Y2=0
r150 58 61 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=2.99
+ $Y2=0
r151 57 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r152 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r153 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r154 54 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r155 53 56 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r156 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r157 51 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r158 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r159 50 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=0 $X2=2.465
+ $Y2=0
r160 50 56 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.3 $Y=0 $X2=2.07
+ $Y2=0
r161 43 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r162 41 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r163 41 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r164 39 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.235 $Y=0
+ $X2=0.515 $Y2=0
r165 39 48 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r166 37 70 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.265 $Y=0 $X2=6.21
+ $Y2=0
r167 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=0 $X2=6.43
+ $Y2=0
r168 36 73 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.595 $Y=0
+ $X2=7.13 $Y2=0
r169 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.43
+ $Y2=0
r170 32 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=0.085
+ $X2=6.43 $Y2=0
r171 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.43 $Y=0.085
+ $X2=6.43 $Y2=0.36
r172 28 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.085
+ $X2=4.245 $Y2=0
r173 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.245 $Y=0.085
+ $X2=4.245 $Y2=0.36
r174 24 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=0.085
+ $X2=3.405 $Y2=0
r175 24 26 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.405 $Y=0.085
+ $X2=3.405 $Y2=0.405
r176 20 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.085
+ $X2=2.465 $Y2=0
r177 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.465 $Y=0.085
+ $X2=2.465 $Y2=0.36
r178 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r179 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r180 5 34 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.295
+ $Y=0.235 $X2=6.43 $Y2=0.36
r181 4 30 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.11
+ $Y=0.235 $X2=4.245 $Y2=0.36
r182 3 26 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.235 $X2=3.405 $Y2=0.405
r183 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.235 $X2=2.465 $Y2=0.36
r184 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%A_382_47# 1 2 9 11 12 15
r35 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.885 $Y=0.615
+ $X2=2.885 $Y2=0.445
r36 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.8 $Y=0.7
+ $X2=2.885 $Y2=0.615
r37 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.8 $Y=0.7 $X2=2.13
+ $Y2=0.7
r38 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=0.615
+ $X2=2.13 $Y2=0.7
r39 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.045 $Y=0.615
+ $X2=2.045 $Y2=0.445
r40 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.75
+ $Y=0.235 $X2=2.885 $Y2=0.445
r41 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.235 $X2=2.045 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_1%A_738_47# 1 2 9 11 12 15
c31 12 0 1.45374e-19 $X=3.91 $Y=0.7
r32 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.665 $Y=0.615
+ $X2=4.665 $Y2=0.445
r33 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.58 $Y=0.7
+ $X2=4.665 $Y2=0.615
r34 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.58 $Y=0.7 $X2=3.91
+ $Y2=0.7
r35 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.825 $Y=0.615
+ $X2=3.91 $Y2=0.7
r36 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.825 $Y=0.615
+ $X2=3.825 $Y2=0.445
r37 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.235 $X2=4.665 $Y2=0.445
r38 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.69
+ $Y=0.235 $X2=3.825 $Y2=0.445
.ends


* File: sky130_fd_sc_hd__lpflow_clkinvkapwr_8.pxi.spice
* Created: Thu Aug 27 14:24:15 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%A N_A_c_86_n N_A_M1000_g N_A_c_87_n
+ N_A_M1003_g N_A_c_88_n N_A_M1004_g N_A_M1001_g N_A_c_89_n N_A_M1006_g
+ N_A_M1002_g N_A_c_90_n N_A_M1007_g N_A_M1005_g N_A_c_91_n N_A_M1010_g
+ N_A_M1008_g N_A_c_92_n N_A_M1012_g N_A_M1009_g N_A_c_93_n N_A_M1013_g
+ N_A_M1011_g N_A_c_94_n N_A_M1014_g N_A_M1016_g N_A_c_95_n N_A_M1015_g
+ N_A_M1017_g N_A_c_96_n N_A_M1018_g N_A_c_97_n N_A_M1019_g A A A A A A A A A
+ N_A_c_128_p N_A_c_85_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%KAPWR N_KAPWR_M1000_s N_KAPWR_M1003_s
+ N_KAPWR_M1006_s N_KAPWR_M1010_s N_KAPWR_M1013_s N_KAPWR_M1015_s
+ N_KAPWR_M1019_s N_KAPWR_c_280_n N_KAPWR_c_282_n N_KAPWR_c_283_n
+ N_KAPWR_c_285_n N_KAPWR_c_286_n N_KAPWR_c_288_n N_KAPWR_c_289_n
+ N_KAPWR_c_291_n N_KAPWR_c_292_n N_KAPWR_c_294_n N_KAPWR_c_276_n
+ N_KAPWR_c_295_n KAPWR N_KAPWR_c_278_n N_KAPWR_c_298_n N_KAPWR_c_300_n
+ N_KAPWR_c_302_n N_KAPWR_c_304_n N_KAPWR_c_306_n N_KAPWR_c_279_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%Y N_Y_M1001_d N_Y_M1005_d N_Y_M1009_d
+ N_Y_M1016_d N_Y_M1000_d N_Y_M1004_d N_Y_M1007_d N_Y_M1012_d N_Y_M1014_d
+ N_Y_M1018_d N_Y_c_417_n N_Y_c_418_n N_Y_c_419_n N_Y_c_431_n N_Y_c_432_n
+ N_Y_c_454_n N_Y_c_433_n N_Y_c_460_n N_Y_c_420_n N_Y_c_434_n N_Y_c_421_n
+ N_Y_c_472_n N_Y_c_422_n N_Y_c_435_n N_Y_c_423_n N_Y_c_484_n N_Y_c_424_n
+ N_Y_c_436_n N_Y_c_425_n N_Y_c_496_n N_Y_c_426_n N_Y_c_437_n N_Y_c_427_n
+ N_Y_c_507_n N_Y_c_438_n N_Y_c_439_n N_Y_c_440_n N_Y_c_514_n N_Y_c_441_n
+ N_Y_c_518_n N_Y_c_442_n N_Y_c_522_n N_Y_c_443_n N_Y_c_526_n N_Y_c_444_n Y Y Y
+ N_Y_c_429_n N_Y_c_446_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%Y
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%VGND N_VGND_M1001_s N_VGND_M1002_s
+ N_VGND_M1008_s N_VGND_M1011_s N_VGND_M1017_s N_VGND_c_661_n N_VGND_c_662_n
+ N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ N_VGND_c_668_n N_VGND_c_669_n VGND N_VGND_c_670_n N_VGND_c_671_n
+ N_VGND_c_672_n N_VGND_c_673_n N_VGND_c_674_n N_VGND_c_675_n N_VGND_c_676_n
+ N_VGND_c_677_n VGND PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%VPWR VPWR N_VPWR_c_752_n
+ N_VPWR_c_751_n PM_SKY130_FD_SC_HD__LPFLOW_CLKINVKAPWR_8%VPWR
cc_1 VNB N_A_M1001_g 0.0222492f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=0.445
cc_2 VNB N_A_M1002_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=1.845 $Y2=0.445
cc_3 VNB N_A_M1005_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=2.275 $Y2=0.445
cc_4 VNB N_A_M1008_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.445
cc_5 VNB N_A_M1009_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=3.135 $Y2=0.445
cc_6 VNB N_A_M1011_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.445
cc_7 VNB N_A_M1016_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.445
cc_8 VNB N_A_M1017_g 0.0222492f $X=-0.19 $Y=-0.24 $X2=4.425 $Y2=0.445
cc_9 VNB N_A_c_85_n 0.342075f $X=-0.19 $Y=-0.24 $X2=5.095 $Y2=1.097
cc_10 VNB N_Y_c_417_n 0.0204208f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.445
cc_11 VNB N_Y_c_418_n 0.0150647f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.445
cc_12 VNB N_Y_c_419_n 0.00997812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_Y_c_420_n 6.75361e-19 $X=-0.19 $Y=-0.24 $X2=3.835 $Y2=1.385
cc_14 VNB N_Y_c_421_n 0.0035731f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.445
cc_15 VNB N_Y_c_422_n 6.52615e-19 $X=-0.19 $Y=-0.24 $X2=4.425 $Y2=0.445
cc_16 VNB N_Y_c_423_n 0.0035731f $X=-0.19 $Y=-0.24 $X2=4.675 $Y2=1.985
cc_17 VNB N_Y_c_424_n 6.52615e-19 $X=-0.19 $Y=-0.24 $X2=2.45 $Y2=1.105
cc_18 VNB N_Y_c_425_n 0.0035731f $X=-0.19 $Y=-0.24 $X2=4.29 $Y2=1.105
cc_19 VNB N_Y_c_426_n 6.75361e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_427_n 0.00820216f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.097
cc_21 VNB Y 0.0225443f $X=-0.19 $Y=-0.24 $X2=4.255 $Y2=1.097
cc_22 VNB N_Y_c_429_n 0.0113484f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.162
cc_23 VNB N_VGND_c_661_n 0.0141137f $X=-0.19 $Y=-0.24 $X2=1.845 $Y2=0.445
cc_24 VNB N_VGND_c_662_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=2.155 $Y2=1.985
cc_25 VNB N_VGND_c_663_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=2.275 $Y2=0.445
cc_26 VNB N_VGND_c_664_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=1.985
cc_27 VNB N_VGND_c_665_n 0.0141137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_666_n 0.011666f $X=-0.19 $Y=-0.24 $X2=2.995 $Y2=1.985
cc_29 VNB N_VGND_c_667_n 0.00436502f $X=-0.19 $Y=-0.24 $X2=3.135 $Y2=0.81
cc_30 VNB N_VGND_c_668_n 0.011666f $X=-0.19 $Y=-0.24 $X2=3.135 $Y2=0.445
cc_31 VNB N_VGND_c_669_n 0.00510476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_670_n 0.0314546f $X=-0.19 $Y=-0.24 $X2=3.415 $Y2=1.985
cc_33 VNB N_VGND_c_671_n 0.011666f $X=-0.19 $Y=-0.24 $X2=3.835 $Y2=1.385
cc_34 VNB N_VGND_c_672_n 0.011666f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.445
cc_35 VNB N_VGND_c_673_n 0.0370325f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_36 VNB N_VGND_c_674_n 0.332673f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_37 VNB N_VGND_c_675_n 0.00510476f $X=-0.19 $Y=-0.24 $X2=2.91 $Y2=1.105
cc_38 VNB N_VGND_c_676_n 0.00436502f $X=-0.19 $Y=-0.24 $X2=4.29 $Y2=1.105
cc_39 VNB N_VGND_c_677_n 0.00436502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_751_n 0.250759f $X=-0.19 $Y=-0.24 $X2=1.315 $Y2=1.985
cc_41 VPB N_A_c_86_n 0.0186504f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.385
cc_42 VPB N_A_c_87_n 0.0152912f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.385
cc_43 VPB N_A_c_88_n 0.0153104f $X=-0.19 $Y=1.305 $X2=1.315 $Y2=1.385
cc_44 VPB N_A_c_89_n 0.0152623f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=1.385
cc_45 VPB N_A_c_90_n 0.0152623f $X=-0.19 $Y=1.305 $X2=2.155 $Y2=1.385
cc_46 VPB N_A_c_91_n 0.0152623f $X=-0.19 $Y=1.305 $X2=2.575 $Y2=1.385
cc_47 VPB N_A_c_92_n 0.0152623f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.385
cc_48 VPB N_A_c_93_n 0.0152623f $X=-0.19 $Y=1.305 $X2=3.415 $Y2=1.385
cc_49 VPB N_A_c_94_n 0.0152623f $X=-0.19 $Y=1.305 $X2=3.835 $Y2=1.385
cc_50 VPB N_A_c_95_n 0.0152623f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.385
cc_51 VPB N_A_c_96_n 0.0152408f $X=-0.19 $Y=1.305 $X2=4.675 $Y2=1.385
cc_52 VPB N_A_c_97_n 0.0186132f $X=-0.19 $Y=1.305 $X2=5.095 $Y2=1.385
cc_53 VPB N_A_c_85_n 0.0693676f $X=-0.19 $Y=1.305 $X2=5.095 $Y2=1.097
cc_54 VPB N_KAPWR_c_276_n 0.0300426f $X=-0.19 $Y=1.305 $X2=4.425 $Y2=0.445
cc_55 VPB KAPWR 0.0114777f $X=-0.19 $Y=1.305 $X2=4.675 $Y2=1.985
cc_56 VPB N_KAPWR_c_278_n 0.0206334f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_57 VPB N_KAPWR_c_279_n 0.0209459f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.097
cc_58 VPB N_Y_c_417_n 0.00728169f $X=-0.19 $Y=1.305 $X2=2.705 $Y2=0.445
cc_59 VPB N_Y_c_431_n 0.00198626f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.385
cc_60 VPB N_Y_c_432_n 0.0072865f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.985
cc_61 VPB N_Y_c_433_n 0.00310598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_Y_c_434_n 0.00307692f $X=-0.19 $Y=1.305 $X2=3.835 $Y2=1.985
cc_63 VPB N_Y_c_435_n 0.00307692f $X=-0.19 $Y=1.305 $X2=4.675 $Y2=1.385
cc_64 VPB N_Y_c_436_n 0.00307692f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.105
cc_65 VPB N_Y_c_437_n 0.00307692f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.097
cc_66 VPB N_Y_c_438_n 6.90551e-19 $X=-0.19 $Y=1.305 $X2=1.735 $Y2=1.097
cc_67 VPB N_Y_c_439_n 0.00128591f $X=-0.19 $Y=1.305 $X2=2.155 $Y2=1.097
cc_68 VPB N_Y_c_440_n 0.00128591f $X=-0.19 $Y=1.305 $X2=2.275 $Y2=1.097
cc_69 VPB N_Y_c_441_n 0.00128591f $X=-0.19 $Y=1.305 $X2=2.705 $Y2=1.097
cc_70 VPB N_Y_c_442_n 0.00128591f $X=-0.19 $Y=1.305 $X2=3.135 $Y2=1.097
cc_71 VPB N_Y_c_443_n 0.00128591f $X=-0.19 $Y=1.305 $X2=3.565 $Y2=1.097
cc_72 VPB N_Y_c_444_n 0.00161539f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=1.097
cc_73 VPB Y 0.00758238f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.097
cc_74 VPB N_Y_c_446_n 0.0071387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_752_n 0.162696f $X=-0.19 $Y=1.305 $X2=1.315 $Y2=1.985
cc_76 VPB N_VPWR_c_751_n 0.0463907f $X=-0.19 $Y=1.305 $X2=1.315 $Y2=1.985
cc_77 N_A_c_86_n N_KAPWR_c_280_n 0.00237585f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_78 N_A_c_87_n N_KAPWR_c_280_n 0.00223726f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_79 N_A_c_87_n N_KAPWR_c_282_n 7.03399e-19 $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_80 N_A_c_88_n N_KAPWR_c_283_n 0.00237585f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_81 N_A_c_89_n N_KAPWR_c_283_n 0.00237585f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_82 N_A_c_90_n N_KAPWR_c_285_n 7.00608e-19 $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_83 N_A_c_90_n N_KAPWR_c_286_n 0.00213827f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_84 N_A_c_91_n N_KAPWR_c_286_n 0.00237585f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_85 N_A_c_92_n N_KAPWR_c_288_n 0.0012643f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_86 N_A_c_92_n N_KAPWR_c_289_n 0.00134632f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_87 N_A_c_93_n N_KAPWR_c_289_n 0.00184129f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_88 N_A_c_93_n N_KAPWR_c_291_n 7.95764e-19 $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_89 N_A_c_94_n N_KAPWR_c_292_n 0.00237585f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_90 N_A_c_95_n N_KAPWR_c_292_n 0.00223726f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_91 N_A_c_95_n N_KAPWR_c_294_n 6.07272e-19 $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_92 N_A_c_96_n N_KAPWR_c_295_n 0.00237585f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_93 N_A_c_97_n N_KAPWR_c_295_n 0.00237585f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_94 N_A_c_86_n N_KAPWR_c_278_n 0.00714216f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_95 N_A_c_87_n N_KAPWR_c_298_n 0.00667948f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_96 N_A_c_88_n N_KAPWR_c_298_n 0.00714046f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_97 N_A_c_89_n N_KAPWR_c_300_n 0.00714046f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A_c_90_n N_KAPWR_c_300_n 0.0069478f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A_c_91_n N_KAPWR_c_302_n 0.00713954f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_100 N_A_c_92_n N_KAPWR_c_302_n 0.0069478f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_101 N_A_c_93_n N_KAPWR_c_304_n 0.0069478f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_102 N_A_c_94_n N_KAPWR_c_304_n 0.00713964f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_103 N_A_c_95_n N_KAPWR_c_306_n 0.0069478f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_104 N_A_c_96_n N_KAPWR_c_306_n 0.00714053f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_105 N_A_c_97_n N_KAPWR_c_279_n 0.0071404f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_106 N_A_c_128_p N_Y_c_417_n 0.0202172f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_c_85_n N_Y_c_417_n 0.0216629f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_108 N_A_M1001_g N_Y_c_418_n 0.0090634f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_c_128_p N_Y_c_418_n 0.0755218f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_c_85_n N_Y_c_418_n 0.0388808f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_111 N_A_c_86_n N_Y_c_431_n 0.0135657f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_112 N_A_c_128_p N_Y_c_431_n 0.00994463f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_c_86_n N_Y_c_454_n 6.71917e-19 $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_114 N_A_c_87_n N_Y_c_454_n 6.78346e-19 $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_115 N_A_c_87_n N_Y_c_433_n 0.0114248f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_116 N_A_c_88_n N_Y_c_433_n 0.01144f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_117 N_A_c_128_p N_Y_c_433_n 0.0485548f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_c_85_n N_Y_c_433_n 0.0026718f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_119 N_A_c_88_n N_Y_c_460_n 4.66008e-19 $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_120 N_A_c_89_n N_Y_c_460_n 4.66008e-19 $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_121 N_A_M1001_g N_Y_c_420_n 0.00101119f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_M1002_g N_Y_c_420_n 5.8681e-19 $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A_c_89_n N_Y_c_434_n 0.0114086f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_124 N_A_c_90_n N_Y_c_434_n 0.0113936f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A_c_128_p N_Y_c_434_n 0.0481863f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_c_85_n N_Y_c_434_n 0.00265179f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_127 N_A_M1002_g N_Y_c_421_n 0.0076909f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A_M1005_g N_Y_c_421_n 0.0076909f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_129 N_A_c_128_p N_Y_c_421_n 0.0468048f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_c_85_n N_Y_c_421_n 0.014197f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_131 N_A_c_90_n N_Y_c_472_n 4.66008e-19 $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_132 N_A_c_91_n N_Y_c_472_n 4.66008e-19 $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_133 N_A_M1005_g N_Y_c_422_n 5.8681e-19 $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A_M1008_g N_Y_c_422_n 5.8681e-19 $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_c_91_n N_Y_c_435_n 0.0114086f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_136 N_A_c_92_n N_Y_c_435_n 0.0113431f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_137 N_A_c_128_p N_Y_c_435_n 0.0481863f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_85_n N_Y_c_435_n 0.00265179f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_139 N_A_M1008_g N_Y_c_423_n 0.0076909f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A_M1009_g N_Y_c_423_n 0.0076909f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_c_128_p N_Y_c_423_n 0.0468048f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_c_85_n N_Y_c_423_n 0.0141423f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_143 N_A_c_92_n N_Y_c_484_n 4.66008e-19 $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_144 N_A_c_93_n N_Y_c_484_n 4.66008e-19 $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_145 N_A_M1009_g N_Y_c_424_n 5.8681e-19 $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_M1011_g N_Y_c_424_n 5.8681e-19 $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_c_93_n N_Y_c_436_n 0.0113747f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_148 N_A_c_94_n N_Y_c_436_n 0.0114086f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A_c_128_p N_Y_c_436_n 0.0481863f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_c_85_n N_Y_c_436_n 0.00265179f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_151 N_A_M1011_g N_Y_c_425_n 0.0076909f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_152 N_A_M1016_g N_Y_c_425_n 0.0076909f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A_c_128_p N_Y_c_425_n 0.0468048f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_c_85_n N_Y_c_425_n 0.014197f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_155 N_A_c_94_n N_Y_c_496_n 4.66008e-19 $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A_c_95_n N_Y_c_496_n 4.66008e-19 $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_157 N_A_M1016_g N_Y_c_426_n 5.8681e-19 $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_M1017_g N_Y_c_426_n 0.00101119f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_c_95_n N_Y_c_437_n 0.0113999f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_160 N_A_c_96_n N_Y_c_437_n 0.0113644f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_161 N_A_c_128_p N_Y_c_437_n 0.0481863f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_c_85_n N_Y_c_437_n 0.00263839f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_163 N_A_M1017_g N_Y_c_427_n 0.0090634f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_c_128_p N_Y_c_427_n 0.0391432f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_c_85_n N_Y_c_427_n 0.0310785f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_166 N_A_c_96_n N_Y_c_507_n 4.66008e-19 $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_167 N_A_c_97_n N_Y_c_507_n 4.66008e-19 $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_168 N_A_c_97_n N_Y_c_438_n 0.0113418f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_169 N_A_c_128_p N_Y_c_439_n 0.014089f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_85_n N_Y_c_439_n 0.00262698f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_171 N_A_c_128_p N_Y_c_440_n 0.014089f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_c_85_n N_Y_c_440_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_173 N_A_c_128_p N_Y_c_514_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_c_85_n N_Y_c_514_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_175 N_A_c_128_p N_Y_c_441_n 0.014089f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_c_85_n N_Y_c_441_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_177 N_A_c_128_p N_Y_c_518_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_85_n N_Y_c_518_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_179 N_A_c_128_p N_Y_c_442_n 0.014089f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_c_85_n N_Y_c_442_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_181 N_A_c_128_p N_Y_c_522_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_c_85_n N_Y_c_522_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_183 N_A_c_128_p N_Y_c_443_n 0.014089f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_c_85_n N_Y_c_443_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_185 N_A_c_128_p N_Y_c_526_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_85_n N_Y_c_526_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_187 N_A_c_128_p N_Y_c_444_n 0.00538726f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_c_85_n N_Y_c_444_n 0.00309075f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_189 N_A_c_128_p Y 0.0134731f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_c_85_n Y 0.0260193f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_191 N_A_c_85_n N_Y_c_429_n 0.00106081f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_192 N_A_c_97_n N_Y_c_446_n 0.0033003f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_193 N_A_M1001_g N_VGND_c_661_n 0.00831231f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A_M1002_g N_VGND_c_661_n 5.62611e-19 $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A_c_85_n N_VGND_c_661_n 0.00163226f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_196 N_A_M1001_g N_VGND_c_662_n 5.62611e-19 $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_197 N_A_M1002_g N_VGND_c_662_n 0.00724882f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_198 N_A_M1005_g N_VGND_c_662_n 0.00724882f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A_M1008_g N_VGND_c_662_n 5.62611e-19 $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_200 N_A_c_85_n N_VGND_c_662_n 5.80335e-19 $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_201 N_A_M1005_g N_VGND_c_663_n 5.62611e-19 $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A_M1008_g N_VGND_c_663_n 0.00724882f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_203 N_A_M1009_g N_VGND_c_663_n 0.00724882f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_204 N_A_M1011_g N_VGND_c_663_n 5.62611e-19 $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A_c_85_n N_VGND_c_663_n 5.80335e-19 $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_206 N_A_M1009_g N_VGND_c_664_n 5.62611e-19 $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A_M1011_g N_VGND_c_664_n 0.00724882f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A_M1016_g N_VGND_c_664_n 0.00724882f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A_M1017_g N_VGND_c_664_n 5.62611e-19 $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_210 N_A_c_85_n N_VGND_c_664_n 5.80335e-19 $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_211 N_A_M1016_g N_VGND_c_665_n 5.62611e-19 $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_212 N_A_M1017_g N_VGND_c_665_n 0.00831231f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A_c_85_n N_VGND_c_665_n 0.0016306f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_214 N_A_M1009_g N_VGND_c_666_n 0.00360664f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A_M1011_g N_VGND_c_666_n 0.00360664f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A_M1016_g N_VGND_c_668_n 0.00360664f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A_M1017_g N_VGND_c_668_n 0.00360664f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A_M1001_g N_VGND_c_671_n 0.00360664f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A_M1002_g N_VGND_c_671_n 0.00360664f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_M1005_g N_VGND_c_672_n 0.00360664f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_221 N_A_M1008_g N_VGND_c_672_n 0.00360664f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_M1001_g N_VGND_c_674_n 0.00428048f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A_M1002_g N_VGND_c_674_n 0.00428048f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_224 N_A_M1005_g N_VGND_c_674_n 0.00428048f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_M1008_g N_VGND_c_674_n 0.00428048f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_226 N_A_M1009_g N_VGND_c_674_n 0.00428048f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_227 N_A_M1011_g N_VGND_c_674_n 0.00428048f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_228 N_A_M1016_g N_VGND_c_674_n 0.00428048f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_M1017_g N_VGND_c_674_n 0.00428048f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A_c_86_n N_VPWR_c_752_n 0.00541359f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_231 N_A_c_87_n N_VPWR_c_752_n 0.0054895f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_232 N_A_c_88_n N_VPWR_c_752_n 0.00541359f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_233 N_A_c_89_n N_VPWR_c_752_n 0.00541359f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_234 N_A_c_90_n N_VPWR_c_752_n 0.00541359f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_235 N_A_c_91_n N_VPWR_c_752_n 0.00541359f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_236 N_A_c_92_n N_VPWR_c_752_n 0.00541359f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_237 N_A_c_93_n N_VPWR_c_752_n 0.00541359f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_238 N_A_c_94_n N_VPWR_c_752_n 0.00541359f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_239 N_A_c_95_n N_VPWR_c_752_n 0.00541359f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_240 N_A_c_96_n N_VPWR_c_752_n 0.00541359f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_241 N_A_c_97_n N_VPWR_c_752_n 0.00541359f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_242 N_A_c_86_n N_VPWR_c_751_n 0.00604573f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_243 N_A_c_87_n N_VPWR_c_751_n 0.00512384f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_244 N_A_c_88_n N_VPWR_c_751_n 0.00510477f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_245 N_A_c_89_n N_VPWR_c_751_n 0.00509152f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_246 N_A_c_90_n N_VPWR_c_751_n 0.00509152f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_247 N_A_c_91_n N_VPWR_c_751_n 0.00509152f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_248 N_A_c_92_n N_VPWR_c_751_n 0.00509152f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_249 N_A_c_93_n N_VPWR_c_751_n 0.00509152f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_250 N_A_c_94_n N_VPWR_c_751_n 0.00509152f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_251 N_A_c_95_n N_VPWR_c_751_n 0.00509152f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_252 N_A_c_96_n N_VPWR_c_751_n 0.00509152f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_253 N_A_c_97_n N_VPWR_c_751_n 0.00641759f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_254 N_KAPWR_c_280_n N_Y_M1000_d 0.0016492f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_255 N_KAPWR_c_283_n N_Y_M1004_d 0.0016492f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_256 N_KAPWR_c_286_n N_Y_M1007_d 0.0016492f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_257 N_KAPWR_c_289_n N_Y_M1012_d 0.0016492f $X=3.435 $Y=2.21 $X2=0 $Y2=0
cc_258 N_KAPWR_c_292_n N_Y_M1014_d 0.0016492f $X=4.295 $Y=2.21 $X2=0 $Y2=0
cc_259 N_KAPWR_c_295_n N_Y_M1018_d 0.0016492f $X=5.195 $Y=2.21 $X2=0 $Y2=0
cc_260 N_KAPWR_M1000_s N_Y_c_431_n 5.36738e-19 $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_261 N_KAPWR_c_280_n N_Y_c_431_n 0.00513051f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_262 KAPWR N_Y_c_431_n 3.08139e-19 $X=0.17 $Y=2.16 $X2=0 $Y2=0
cc_263 N_KAPWR_c_278_n N_Y_c_431_n 0.00620619f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_264 N_KAPWR_M1000_s N_Y_c_432_n 0.00225375f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_265 KAPWR N_Y_c_432_n 7.93205e-19 $X=0.17 $Y=2.16 $X2=0 $Y2=0
cc_266 N_KAPWR_c_278_n N_Y_c_432_n 0.0146951f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_267 N_KAPWR_c_280_n N_Y_c_454_n 0.0182386f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_268 N_KAPWR_c_282_n N_Y_c_454_n 0.00149834f $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_269 KAPWR N_Y_c_454_n 3.81051e-19 $X=0.17 $Y=2.16 $X2=0 $Y2=0
cc_270 N_KAPWR_c_278_n N_Y_c_454_n 0.0262181f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_271 N_KAPWR_c_298_n N_Y_c_454_n 0.0253869f $X=1.105 $Y=1.965 $X2=0 $Y2=0
cc_272 N_KAPWR_M1003_s N_Y_c_433_n 0.00166182f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_273 N_KAPWR_c_280_n N_Y_c_433_n 0.00472442f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_274 N_KAPWR_c_282_n N_Y_c_433_n 0.00147061f $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_275 N_KAPWR_c_283_n N_Y_c_433_n 0.00507375f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_276 N_KAPWR_c_298_n N_Y_c_433_n 0.0163967f $X=1.105 $Y=1.965 $X2=0 $Y2=0
cc_277 N_KAPWR_c_282_n N_Y_c_460_n 3.95806e-19 $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_278 N_KAPWR_c_283_n N_Y_c_460_n 0.0181896f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_279 N_KAPWR_c_285_n N_Y_c_460_n 3.95806e-19 $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_280 N_KAPWR_c_298_n N_Y_c_460_n 0.0262468f $X=1.105 $Y=1.965 $X2=0 $Y2=0
cc_281 N_KAPWR_c_300_n N_Y_c_460_n 0.0262468f $X=1.945 $Y=1.965 $X2=0 $Y2=0
cc_282 N_KAPWR_M1006_s N_Y_c_434_n 0.00161021f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_283 N_KAPWR_c_283_n N_Y_c_434_n 0.00507375f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_284 N_KAPWR_c_285_n N_Y_c_434_n 0.00146885f $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_285 N_KAPWR_c_286_n N_Y_c_434_n 0.00458945f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_286 N_KAPWR_c_300_n N_Y_c_434_n 0.0163718f $X=1.945 $Y=1.965 $X2=0 $Y2=0
cc_287 N_KAPWR_c_285_n N_Y_c_472_n 0.00150299f $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_288 N_KAPWR_c_286_n N_Y_c_472_n 0.0181896f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_289 N_KAPWR_c_288_n N_Y_c_472_n 3.58876e-19 $X=3 $Y=2.21 $X2=0 $Y2=0
cc_290 N_KAPWR_c_300_n N_Y_c_472_n 0.0260808f $X=1.945 $Y=1.965 $X2=0 $Y2=0
cc_291 N_KAPWR_c_302_n N_Y_c_472_n 0.0262152f $X=2.785 $Y=1.965 $X2=0 $Y2=0
cc_292 N_KAPWR_M1010_s N_Y_c_435_n 0.00157925f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_293 N_KAPWR_c_286_n N_Y_c_435_n 0.00522512f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_294 N_KAPWR_c_288_n N_Y_c_435_n 0.00248978f $X=3 $Y=2.21 $X2=0 $Y2=0
cc_295 N_KAPWR_c_289_n N_Y_c_435_n 0.00350968f $X=3.435 $Y=2.21 $X2=0 $Y2=0
cc_296 N_KAPWR_c_302_n N_Y_c_435_n 0.0163736f $X=2.785 $Y=1.965 $X2=0 $Y2=0
cc_297 N_KAPWR_c_288_n N_Y_c_484_n 6.12705e-19 $X=3 $Y=2.21 $X2=0 $Y2=0
cc_298 N_KAPWR_c_289_n N_Y_c_484_n 0.0181896f $X=3.435 $Y=2.21 $X2=0 $Y2=0
cc_299 N_KAPWR_c_291_n N_Y_c_484_n 5.82753e-19 $X=3.725 $Y=2.21 $X2=0 $Y2=0
cc_300 N_KAPWR_c_302_n N_Y_c_484_n 0.0260808f $X=2.785 $Y=1.965 $X2=0 $Y2=0
cc_301 N_KAPWR_c_304_n N_Y_c_484_n 0.0260808f $X=3.625 $Y=1.965 $X2=0 $Y2=0
cc_302 N_KAPWR_M1013_s N_Y_c_436_n 0.00161021f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_303 N_KAPWR_c_289_n N_Y_c_436_n 0.00418454f $X=3.435 $Y=2.21 $X2=0 $Y2=0
cc_304 N_KAPWR_c_291_n N_Y_c_436_n 0.0018517f $X=3.725 $Y=2.21 $X2=0 $Y2=0
cc_305 N_KAPWR_c_292_n N_Y_c_436_n 0.00513051f $X=4.295 $Y=2.21 $X2=0 $Y2=0
cc_306 N_KAPWR_c_304_n N_Y_c_436_n 0.0163718f $X=3.625 $Y=1.965 $X2=0 $Y2=0
cc_307 N_KAPWR_c_291_n N_Y_c_496_n 3.81051e-19 $X=3.725 $Y=2.21 $X2=0 $Y2=0
cc_308 N_KAPWR_c_292_n N_Y_c_496_n 0.0181896f $X=4.295 $Y=2.21 $X2=0 $Y2=0
cc_309 N_KAPWR_c_294_n N_Y_c_496_n 0.00149354f $X=4.585 $Y=2.21 $X2=0 $Y2=0
cc_310 N_KAPWR_c_304_n N_Y_c_496_n 0.0262181f $X=3.625 $Y=1.965 $X2=0 $Y2=0
cc_311 N_KAPWR_c_306_n N_Y_c_496_n 0.0260808f $X=4.465 $Y=1.965 $X2=0 $Y2=0
cc_312 N_KAPWR_M1015_s N_Y_c_437_n 0.00161021f $X=4.33 $Y=1.485 $X2=0 $Y2=0
cc_313 N_KAPWR_c_292_n N_Y_c_437_n 0.00472442f $X=4.295 $Y=2.21 $X2=0 $Y2=0
cc_314 N_KAPWR_c_294_n N_Y_c_437_n 0.00134123f $X=4.585 $Y=2.21 $X2=0 $Y2=0
cc_315 N_KAPWR_c_295_n N_Y_c_437_n 0.00505483f $X=5.195 $Y=2.21 $X2=0 $Y2=0
cc_316 N_KAPWR_c_306_n N_Y_c_437_n 0.0163718f $X=4.465 $Y=1.965 $X2=0 $Y2=0
cc_317 N_KAPWR_c_294_n N_Y_c_507_n 4.01003e-19 $X=4.585 $Y=2.21 $X2=0 $Y2=0
cc_318 N_KAPWR_c_276_n N_Y_c_507_n 3.90753e-19 $X=5.34 $Y=2.21 $X2=0 $Y2=0
cc_319 N_KAPWR_c_295_n N_Y_c_507_n 0.0181896f $X=5.195 $Y=2.21 $X2=0 $Y2=0
cc_320 N_KAPWR_c_306_n N_Y_c_507_n 0.0262492f $X=4.465 $Y=1.965 $X2=0 $Y2=0
cc_321 N_KAPWR_c_279_n N_Y_c_507_n 0.0262444f $X=5.305 $Y=1.965 $X2=0 $Y2=0
cc_322 N_KAPWR_c_295_n N_Y_c_438_n 0.00499898f $X=5.195 $Y=2.21 $X2=0 $Y2=0
cc_323 N_KAPWR_c_279_n N_Y_c_438_n 0.00206485f $X=5.305 $Y=1.965 $X2=0 $Y2=0
cc_324 N_KAPWR_M1019_s N_Y_c_446_n 0.00283124f $X=5.17 $Y=1.485 $X2=0 $Y2=0
cc_325 N_KAPWR_c_276_n N_Y_c_446_n 0.00114417f $X=5.34 $Y=2.21 $X2=0 $Y2=0
cc_326 N_KAPWR_c_279_n N_Y_c_446_n 0.0183721f $X=5.305 $Y=1.965 $X2=0 $Y2=0
cc_327 N_KAPWR_c_280_n N_VPWR_c_752_n 0.00187854f $X=0.93 $Y=2.21 $X2=0 $Y2=0
cc_328 N_KAPWR_c_282_n N_VPWR_c_752_n 2.2288e-19 $X=1.22 $Y=2.21 $X2=0 $Y2=0
cc_329 N_KAPWR_c_283_n N_VPWR_c_752_n 0.00207717f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_330 N_KAPWR_c_285_n N_VPWR_c_752_n 8.63828e-19 $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_331 N_KAPWR_c_286_n N_VPWR_c_752_n 0.00121299f $X=2.71 $Y=2.21 $X2=0 $Y2=0
cc_332 N_KAPWR_c_288_n N_VPWR_c_752_n 8.67652e-19 $X=3 $Y=2.21 $X2=0 $Y2=0
cc_333 N_KAPWR_c_289_n N_VPWR_c_752_n 9.90738e-19 $X=3.435 $Y=2.21 $X2=0 $Y2=0
cc_334 N_KAPWR_c_291_n N_VPWR_c_752_n 2.22965e-19 $X=3.725 $Y=2.21 $X2=0 $Y2=0
cc_335 N_KAPWR_c_292_n N_VPWR_c_752_n 0.00185323f $X=4.295 $Y=2.21 $X2=0 $Y2=0
cc_336 N_KAPWR_c_294_n N_VPWR_c_752_n 2.22852e-19 $X=4.585 $Y=2.21 $X2=0 $Y2=0
cc_337 N_KAPWR_c_276_n N_VPWR_c_752_n 0.00234274f $X=5.34 $Y=2.21 $X2=0 $Y2=0
cc_338 N_KAPWR_c_295_n N_VPWR_c_752_n 0.00207719f $X=5.195 $Y=2.21 $X2=0 $Y2=0
cc_339 KAPWR N_VPWR_c_752_n 3.63792e-19 $X=0.17 $Y=2.16 $X2=0 $Y2=0
cc_340 N_KAPWR_c_278_n N_VPWR_c_752_n 0.021007f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_341 N_KAPWR_c_298_n N_VPWR_c_752_n 0.0188904f $X=1.105 $Y=1.965 $X2=0 $Y2=0
cc_342 N_KAPWR_c_300_n N_VPWR_c_752_n 0.0188798f $X=1.945 $Y=1.965 $X2=0 $Y2=0
cc_343 N_KAPWR_c_302_n N_VPWR_c_752_n 0.0188798f $X=2.785 $Y=1.965 $X2=0 $Y2=0
cc_344 N_KAPWR_c_304_n N_VPWR_c_752_n 0.0188798f $X=3.625 $Y=1.965 $X2=0 $Y2=0
cc_345 N_KAPWR_c_306_n N_VPWR_c_752_n 0.0188798f $X=4.465 $Y=1.965 $X2=0 $Y2=0
cc_346 N_KAPWR_c_279_n N_VPWR_c_752_n 0.021007f $X=5.305 $Y=1.965 $X2=0 $Y2=0
cc_347 N_KAPWR_M1000_s N_VPWR_c_751_n 0.0010704f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_348 N_KAPWR_M1003_s N_VPWR_c_751_n 0.00111408f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_349 N_KAPWR_M1006_s N_VPWR_c_751_n 0.00109368f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_350 N_KAPWR_M1010_s N_VPWR_c_751_n 0.00109368f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_351 N_KAPWR_M1013_s N_VPWR_c_751_n 0.00109368f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_352 N_KAPWR_M1015_s N_VPWR_c_751_n 0.00109368f $X=4.33 $Y=1.485 $X2=0 $Y2=0
cc_353 N_KAPWR_M1019_s N_VPWR_c_751_n 0.0010704f $X=5.17 $Y=1.485 $X2=0 $Y2=0
cc_354 KAPWR N_VPWR_c_751_n 0.60265f $X=0.17 $Y=2.16 $X2=0 $Y2=0
cc_355 N_KAPWR_c_278_n N_VPWR_c_751_n 0.00298827f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_356 N_KAPWR_c_298_n N_VPWR_c_751_n 0.00294505f $X=1.105 $Y=1.965 $X2=0 $Y2=0
cc_357 N_KAPWR_c_300_n N_VPWR_c_751_n 0.00293968f $X=1.945 $Y=1.965 $X2=0 $Y2=0
cc_358 N_KAPWR_c_302_n N_VPWR_c_751_n 0.00293968f $X=2.785 $Y=1.965 $X2=0 $Y2=0
cc_359 N_KAPWR_c_304_n N_VPWR_c_751_n 0.00293968f $X=3.625 $Y=1.965 $X2=0 $Y2=0
cc_360 N_KAPWR_c_306_n N_VPWR_c_751_n 0.00293968f $X=4.465 $Y=1.965 $X2=0 $Y2=0
cc_361 N_KAPWR_c_279_n N_VPWR_c_751_n 0.00298827f $X=5.305 $Y=1.965 $X2=0 $Y2=0
cc_362 N_Y_c_418_n N_VGND_c_661_n 0.0232314f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_363 N_Y_c_421_n N_VGND_c_662_n 0.020457f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_364 N_Y_c_423_n N_VGND_c_663_n 0.020457f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_365 N_Y_c_425_n N_VGND_c_664_n 0.020457f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_366 N_Y_c_427_n N_VGND_c_665_n 0.0232314f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_367 N_Y_c_423_n N_VGND_c_666_n 0.00249722f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_368 N_Y_c_424_n N_VGND_c_666_n 0.0106278f $X=3.35 $Y=0.445 $X2=0 $Y2=0
cc_369 N_Y_c_425_n N_VGND_c_666_n 0.00249722f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_370 N_Y_c_425_n N_VGND_c_668_n 0.00249722f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_371 N_Y_c_426_n N_VGND_c_668_n 0.0106278f $X=4.21 $Y=0.445 $X2=0 $Y2=0
cc_372 N_Y_c_427_n N_VGND_c_668_n 0.00249722f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_373 N_Y_c_418_n N_VGND_c_670_n 0.0121037f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_374 N_Y_c_419_n N_VGND_c_670_n 0.0030627f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_375 N_Y_c_418_n N_VGND_c_671_n 0.00249722f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_376 N_Y_c_420_n N_VGND_c_671_n 0.0106278f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_377 N_Y_c_421_n N_VGND_c_671_n 0.00249722f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_378 N_Y_c_421_n N_VGND_c_672_n 0.00249722f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_379 N_Y_c_422_n N_VGND_c_672_n 0.0106278f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_380 N_Y_c_423_n N_VGND_c_672_n 0.00249722f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_381 N_Y_c_427_n N_VGND_c_673_n 0.00588215f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_382 N_Y_c_429_n N_VGND_c_673_n 0.0048643f $X=5.305 $Y=0.865 $X2=0 $Y2=0
cc_383 N_Y_M1001_d N_VGND_c_674_n 0.00264766f $X=1.49 $Y=0.235 $X2=0 $Y2=0
cc_384 N_Y_M1005_d N_VGND_c_674_n 0.00264766f $X=2.35 $Y=0.235 $X2=0 $Y2=0
cc_385 N_Y_M1009_d N_VGND_c_674_n 0.00264766f $X=3.21 $Y=0.235 $X2=0 $Y2=0
cc_386 N_Y_M1016_d N_VGND_c_674_n 0.00264766f $X=4.07 $Y=0.235 $X2=0 $Y2=0
cc_387 N_Y_c_418_n N_VGND_c_674_n 0.0256198f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_388 N_Y_c_419_n N_VGND_c_674_n 0.00489372f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_389 N_Y_c_420_n N_VGND_c_674_n 0.00712214f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_390 N_Y_c_421_n N_VGND_c_674_n 0.00929518f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_391 N_Y_c_422_n N_VGND_c_674_n 0.00712214f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_392 N_Y_c_423_n N_VGND_c_674_n 0.00929518f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_393 N_Y_c_424_n N_VGND_c_674_n 0.00712214f $X=3.35 $Y=0.445 $X2=0 $Y2=0
cc_394 N_Y_c_425_n N_VGND_c_674_n 0.00929518f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_395 N_Y_c_426_n N_VGND_c_674_n 0.00712214f $X=4.21 $Y=0.445 $X2=0 $Y2=0
cc_396 N_Y_c_427_n N_VGND_c_674_n 0.0152079f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_397 N_Y_c_429_n N_VGND_c_674_n 0.00777238f $X=5.305 $Y=0.865 $X2=0 $Y2=0
cc_398 N_Y_c_454_n N_VPWR_c_752_n 0.00955594f $X=0.68 $Y=1.93 $X2=0 $Y2=0
cc_399 N_Y_c_460_n N_VPWR_c_752_n 0.00955594f $X=1.525 $Y=1.83 $X2=0 $Y2=0
cc_400 N_Y_c_472_n N_VPWR_c_752_n 0.00955594f $X=2.365 $Y=1.83 $X2=0 $Y2=0
cc_401 N_Y_c_484_n N_VPWR_c_752_n 0.00955594f $X=3.205 $Y=1.83 $X2=0 $Y2=0
cc_402 N_Y_c_496_n N_VPWR_c_752_n 0.00955594f $X=4.045 $Y=1.83 $X2=0 $Y2=0
cc_403 N_Y_c_507_n N_VPWR_c_752_n 0.00955594f $X=4.885 $Y=1.83 $X2=0 $Y2=0
cc_404 N_Y_M1000_d N_VPWR_c_751_n 0.00151665f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_405 N_Y_M1004_d N_VPWR_c_751_n 0.00151665f $X=1.39 $Y=1.485 $X2=0 $Y2=0
cc_406 N_Y_M1007_d N_VPWR_c_751_n 0.00151665f $X=2.23 $Y=1.485 $X2=0 $Y2=0
cc_407 N_Y_M1012_d N_VPWR_c_751_n 0.00151665f $X=3.07 $Y=1.485 $X2=0 $Y2=0
cc_408 N_Y_M1014_d N_VPWR_c_751_n 0.00151665f $X=3.91 $Y=1.485 $X2=0 $Y2=0
cc_409 N_Y_M1018_d N_VPWR_c_751_n 0.00151665f $X=4.75 $Y=1.485 $X2=0 $Y2=0
cc_410 N_Y_c_454_n N_VPWR_c_751_n 0.00159601f $X=0.68 $Y=1.93 $X2=0 $Y2=0
cc_411 N_Y_c_460_n N_VPWR_c_751_n 0.00159601f $X=1.525 $Y=1.83 $X2=0 $Y2=0
cc_412 N_Y_c_472_n N_VPWR_c_751_n 0.00159601f $X=2.365 $Y=1.83 $X2=0 $Y2=0
cc_413 N_Y_c_484_n N_VPWR_c_751_n 0.00159601f $X=3.205 $Y=1.83 $X2=0 $Y2=0
cc_414 N_Y_c_496_n N_VPWR_c_751_n 0.00159601f $X=4.045 $Y=1.83 $X2=0 $Y2=0
cc_415 N_Y_c_507_n N_VPWR_c_751_n 0.00159601f $X=4.885 $Y=1.83 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__clkdlybuf4s15_2.pxi.spice
* Created: Thu Aug 27 14:11:24 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A N_A_M1000_g N_A_M1005_g A A N_A_c_74_n
+ N_A_c_75_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_27_47# N_A_27_47#_M1000_s
+ N_A_27_47#_M1005_s N_A_27_47#_M1003_g N_A_27_47#_M1001_g N_A_27_47#_c_108_n
+ N_A_27_47#_c_109_n N_A_27_47#_c_110_n N_A_27_47#_c_127_n N_A_27_47#_c_111_n
+ N_A_27_47#_c_112_n N_A_27_47#_c_117_n N_A_27_47#_c_113_n N_A_27_47#_c_114_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_228_47# N_A_228_47#_M1003_d
+ N_A_228_47#_M1001_d N_A_228_47#_M1009_g N_A_228_47#_M1004_g
+ N_A_228_47#_c_185_n N_A_228_47#_c_186_n N_A_228_47#_c_187_n
+ N_A_228_47#_c_188_n N_A_228_47#_c_194_n N_A_228_47#_c_195_n
+ N_A_228_47#_c_189_n N_A_228_47#_c_190_n N_A_228_47#_c_191_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_228_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_362_333# N_A_362_333#_M1009_s
+ N_A_362_333#_M1004_s N_A_362_333#_M1006_g N_A_362_333#_M1002_g
+ N_A_362_333#_c_259_n N_A_362_333#_M1008_g N_A_362_333#_M1007_g
+ N_A_362_333#_c_262_n N_A_362_333#_c_274_n N_A_362_333#_c_263_n
+ N_A_362_333#_c_264_n N_A_362_333#_c_283_n N_A_362_333#_c_265_n
+ N_A_362_333#_c_266_n N_A_362_333#_c_322_p N_A_362_333#_c_267_n
+ N_A_362_333#_c_292_n N_A_362_333#_c_268_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%A_362_333#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%VPWR N_VPWR_M1005_d N_VPWR_M1004_d
+ N_VPWR_M1007_d N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n
+ N_VPWR_c_353_n N_VPWR_c_354_n VPWR N_VPWR_c_355_n N_VPWR_c_356_n
+ N_VPWR_c_357_n N_VPWR_c_348_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%X N_X_M1006_d N_X_M1002_s X X X X X X
+ N_X_c_412_n N_X_c_414_n X PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%VGND N_VGND_M1000_d N_VGND_M1009_d
+ N_VGND_M1008_s N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n N_VGND_c_431_n
+ N_VGND_c_432_n N_VGND_c_433_n VGND N_VGND_c_434_n N_VGND_c_435_n
+ N_VGND_c_436_n N_VGND_c_437_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S15_2%VGND
cc_1 VNB N_A_M1000_g 0.0408968f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.445
cc_2 VNB N_A_M1005_g 6.18739e-19 $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.985
cc_3 VNB N_A_c_74_n 0.0343364f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_4 VNB N_A_c_75_n 0.0107864f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_5 VNB N_A_27_47#_M1003_g 0.0221813f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_A_27_47#_M1001_g 5.37909e-19 $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.16
cc_7 VNB N_A_27_47#_c_108_n 0.018703f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.295
cc_8 VNB N_A_27_47#_c_109_n 0.0125816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_110_n 0.0101228f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.53
cc_10 VNB N_A_27_47#_c_111_n 0.00226782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_112_n 7.80269e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_113_n 0.00315383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_114_n 0.0350879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_228_47#_M1009_g 0.0249154f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_228_47#_M1004_g 6.16407e-19 $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.16
cc_16 VNB N_A_228_47#_c_185_n 0.00595696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_228_47#_c_186_n 0.00377212f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.53
cc_18 VNB N_A_228_47#_c_187_n 0.00523688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_228_47#_c_188_n 0.0249206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_228_47#_c_189_n 0.00946197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_228_47#_c_190_n 0.00210576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_228_47#_c_191_n 0.0339223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_362_333#_M1006_g 0.0355433f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB N_A_362_333#_M1002_g 5.64312e-19 $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.16
cc_25 VNB N_A_362_333#_c_259_n 0.0131164f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_26 VNB N_A_362_333#_M1008_g 0.0345971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_362_333#_M1007_g 5.20615e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_362_333#_c_262_n 0.0120052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_362_333#_c_263_n 0.0192805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_362_333#_c_264_n 0.00165257f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_362_333#_c_265_n 0.00303501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_362_333#_c_266_n 5.6245e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_362_333#_c_267_n 0.0176905f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_362_333#_c_268_n 0.00136656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_348_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB X 0.0262155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_428_n 0.00558593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_429_n 0.00558109f $X=-0.19 $Y=-0.24 $X2=0.387 $Y2=1.025
cc_39 VNB N_VGND_c_430_n 0.011356f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_40 VNB N_VGND_c_431_n 0.0235962f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.19
cc_41 VNB N_VGND_c_432_n 0.0435724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_433_n 0.00631673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_434_n 0.0169077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_435_n 0.0216586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_436_n 0.00631594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_437_n 0.22575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VPB N_A_M1005_g 0.0263627f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_48 VPB N_A_c_75_n 0.0132162f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_49 VPB N_A_27_47#_M1001_g 0.0355504f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.16
cc_50 VPB N_A_27_47#_c_112_n 0.00309433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_117_n 0.0276567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_228_47#_M1004_g 0.0404384f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.16
cc_53 VPB N_A_228_47#_c_187_n 0.013277f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_228_47#_c_194_n 0.00926368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_228_47#_c_195_n 0.00691222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_228_47#_c_190_n 0.00219817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_362_333#_M1002_g 0.0234618f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.16
cc_58 VPB N_A_362_333#_M1007_g 0.0236642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_362_333#_c_266_n 0.00311316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_349_n 0.00558649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_350_n 0.00563065f $X=-0.19 $Y=1.305 $X2=0.387 $Y2=1.025
cc_62 VPB N_VPWR_c_351_n 0.0113301f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_63 VPB N_VPWR_c_352_n 0.0582611f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.19
cc_64 VPB N_VPWR_c_353_n 0.042778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_354_n 0.00632108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_355_n 0.0172818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_356_n 0.0218265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_357_n 0.00631775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_348_n 0.0508767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB X 0.00786947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB X 0.00280295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 N_A_c_75_n N_A_27_47#_M1005_s 0.00304124f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_A_27_47#_M1003_g 0.0180629f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_M1005_g N_A_27_47#_M1001_g 0.0180629f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_A_27_47#_c_108_n 0.0082379f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_A_27_47#_c_109_n 0.010303f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_c_75_n N_A_27_47#_c_109_n 0.0103915f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_M1000_g N_A_27_47#_c_110_n 0.00376263f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A_c_74_n N_A_27_47#_c_110_n 0.00430128f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_75_n N_A_27_47#_c_110_n 0.0293359f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_M1005_g N_A_27_47#_c_127_n 0.00956502f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_c_75_n N_A_27_47#_c_127_n 0.00926648f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_A_27_47#_c_111_n 0.00320455f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_c_75_n N_A_27_47#_c_111_n 6.97913e-19 $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_c_74_n N_A_27_47#_c_112_n 0.00560811f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_c_75_n N_A_27_47#_c_112_n 0.0176575f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_M1005_g N_A_27_47#_c_117_n 0.00781784f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_c_74_n N_A_27_47#_c_117_n 6.31831e-19 $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_c_75_n N_A_27_47#_c_117_n 0.0254885f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_c_74_n N_A_27_47#_c_113_n 0.00134854f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_c_75_n N_A_27_47#_c_113_n 0.00843528f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_c_74_n N_A_27_47#_c_114_n 0.0180629f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_c_75_n N_A_27_47#_c_114_n 6.17754e-19 $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_M1005_g N_VPWR_c_349_n 0.00532457f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_M1005_g N_VPWR_c_355_n 0.00429359f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_M1005_g N_VPWR_c_348_n 0.00719626f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_M1000_g N_VGND_c_428_n 0.00323507f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_M1000_g N_VGND_c_434_n 0.00433389f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_M1000_g N_VGND_c_437_n 0.00710934f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_27_47#_M1003_g N_A_228_47#_c_185_n 0.0172775f $X=1.065 $Y=0.56 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_M1003_g N_A_228_47#_c_186_n 0.00208798f $X=1.065 $Y=0.56 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_111_n N_A_228_47#_c_186_n 0.00602797f $X=0.975 $Y=1.075
+ $X2=0 $Y2=0
cc_103 N_A_27_47#_c_114_n N_A_228_47#_c_186_n 5.32093e-19 $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_M1001_g N_A_228_47#_c_194_n 0.0188188f $X=1.065 $Y=2.075 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_127_n N_A_228_47#_c_194_n 0.0142842f $X=0.89 $Y=1.88 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_112_n N_A_228_47#_c_194_n 7.2218e-19 $X=0.975 $Y=1.795 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_113_n N_A_228_47#_c_194_n 0.00285767f $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_c_114_n N_A_228_47#_c_194_n 0.00165105f $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_M1001_g N_A_228_47#_c_195_n 0.00525662f $X=1.065 $Y=2.075
+ $X2=0 $Y2=0
cc_110 N_A_27_47#_c_112_n N_A_228_47#_c_195_n 0.0105254f $X=0.975 $Y=1.795 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_109_n N_A_228_47#_c_189_n 0.0116021f $X=0.89 $Y=0.805 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_c_111_n N_A_228_47#_c_189_n 9.18277e-19 $X=0.975 $Y=1.075
+ $X2=0 $Y2=0
cc_113 N_A_27_47#_c_113_n N_A_228_47#_c_189_n 0.00313414f $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_114_n N_A_228_47#_c_189_n 9.24857e-19 $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1001_g N_A_228_47#_c_190_n 0.00359111f $X=1.065 $Y=2.075
+ $X2=0 $Y2=0
cc_116 N_A_27_47#_c_112_n N_A_228_47#_c_190_n 0.00970162f $X=0.975 $Y=1.795
+ $X2=0 $Y2=0
cc_117 N_A_27_47#_c_113_n N_A_228_47#_c_190_n 0.0144989f $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_c_114_n N_A_228_47#_c_190_n 0.00140835f $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_114_n N_A_228_47#_c_191_n 0.00667289f $X=1.155 $Y=1.16 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_c_127_n N_VPWR_M1005_d 0.0145623f $X=0.89 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_121 N_A_27_47#_c_112_n N_VPWR_M1005_d 0.00171173f $X=0.975 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_27_47#_M1001_g N_VPWR_c_349_n 0.00731985f $X=1.065 $Y=2.075 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_127_n N_VPWR_c_349_n 0.0252566f $X=0.89 $Y=1.88 $X2=0 $Y2=0
cc_124 N_A_27_47#_M1001_g N_VPWR_c_353_n 0.00518352f $X=1.065 $Y=2.075 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_127_n N_VPWR_c_353_n 0.00141724f $X=0.89 $Y=1.88 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_127_n N_VPWR_c_355_n 0.00187601f $X=0.89 $Y=1.88 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_117_n N_VPWR_c_355_n 0.0220955f $X=0.265 $Y=1.96 $X2=0 $Y2=0
cc_128 N_A_27_47#_M1005_s N_VPWR_c_348_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_M1001_g N_VPWR_c_348_n 0.0103194f $X=1.065 $Y=2.075 $X2=0
+ $Y2=0
cc_130 N_A_27_47#_c_127_n N_VPWR_c_348_n 0.00822732f $X=0.89 $Y=1.88 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_117_n N_VPWR_c_348_n 0.0130222f $X=0.265 $Y=1.96 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_109_n N_VGND_M1000_d 0.00359868f $X=0.89 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_27_47#_M1003_g N_VGND_c_428_n 0.00700089f $X=1.065 $Y=0.56 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_109_n N_VGND_c_428_n 0.0246574f $X=0.89 $Y=0.805 $X2=0 $Y2=0
cc_135 N_A_27_47#_M1003_g N_VGND_c_432_n 0.00516154f $X=1.065 $Y=0.56 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_c_109_n N_VGND_c_432_n 0.00171717f $X=0.89 $Y=0.805 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_c_108_n N_VGND_c_434_n 0.0209989f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_109_n N_VGND_c_434_n 0.0023428f $X=0.89 $Y=0.805 $X2=0 $Y2=0
cc_139 N_A_27_47#_M1000_s N_VGND_c_437_n 0.00217517f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_M1003_g N_VGND_c_437_n 0.0103164f $X=1.065 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_108_n N_VGND_c_437_n 0.0124957f $X=0.265 $Y=0.42 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_109_n N_VGND_c_437_n 0.00868894f $X=0.89 $Y=0.805 $X2=0
+ $Y2=0
cc_143 N_A_228_47#_M1009_g N_A_362_333#_M1006_g 0.0109736f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_144 N_A_228_47#_M1004_g N_A_362_333#_M1002_g 0.0145457f $X=2.15 $Y=2.075
+ $X2=0 $Y2=0
cc_145 N_A_228_47#_M1009_g N_A_362_333#_c_274_n 0.0151395f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_146 N_A_228_47#_c_185_n N_A_362_333#_c_274_n 0.0390156f $X=1.42 $Y=0.42 $X2=0
+ $Y2=0
cc_147 N_A_228_47#_M1009_g N_A_362_333#_c_263_n 0.010295f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_148 N_A_228_47#_c_187_n N_A_362_333#_c_263_n 0.0235706f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_228_47#_c_188_n N_A_362_333#_c_263_n 0.00433688f $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_150 N_A_228_47#_M1009_g N_A_362_333#_c_264_n 0.00401422f $X=2.15 $Y=0.56
+ $X2=0 $Y2=0
cc_151 N_A_228_47#_c_187_n N_A_362_333#_c_264_n 0.0228767f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_228_47#_c_189_n N_A_362_333#_c_264_n 0.0149258f $X=1.47 $Y=0.905
+ $X2=0 $Y2=0
cc_153 N_A_228_47#_c_191_n N_A_362_333#_c_264_n 0.00578966f $X=2.075 $Y=1.16
+ $X2=0 $Y2=0
cc_154 N_A_228_47#_M1004_g N_A_362_333#_c_283_n 0.0111533f $X=2.15 $Y=2.075
+ $X2=0 $Y2=0
cc_155 N_A_228_47#_c_187_n N_A_362_333#_c_283_n 0.014291f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_156 N_A_228_47#_c_188_n N_A_362_333#_c_283_n 7.15433e-19 $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_157 N_A_228_47#_M1009_g N_A_362_333#_c_265_n 0.00193853f $X=2.15 $Y=0.56
+ $X2=0 $Y2=0
cc_158 N_A_228_47#_c_188_n N_A_362_333#_c_265_n 9.94107e-19 $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_159 N_A_228_47#_M1004_g N_A_362_333#_c_266_n 0.00551523f $X=2.15 $Y=2.075
+ $X2=0 $Y2=0
cc_160 N_A_228_47#_c_187_n N_A_362_333#_c_266_n 0.0128792f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_161 N_A_228_47#_c_187_n N_A_362_333#_c_267_n 2.32345e-19 $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_162 N_A_228_47#_c_188_n N_A_362_333#_c_267_n 0.00658481f $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_163 N_A_228_47#_M1004_g N_A_362_333#_c_292_n 0.0140516f $X=2.15 $Y=2.075
+ $X2=0 $Y2=0
cc_164 N_A_228_47#_c_187_n N_A_362_333#_c_292_n 0.0137598f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A_228_47#_c_194_n N_A_362_333#_c_292_n 0.056514f $X=1.395 $Y=1.96 $X2=0
+ $Y2=0
cc_166 N_A_228_47#_c_191_n N_A_362_333#_c_292_n 0.00109717f $X=2.075 $Y=1.16
+ $X2=0 $Y2=0
cc_167 N_A_228_47#_c_187_n N_A_362_333#_c_268_n 0.00918792f $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_168 N_A_228_47#_c_188_n N_A_362_333#_c_268_n 7.58904e-19 $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_169 N_A_228_47#_c_194_n N_VPWR_c_349_n 0.0177726f $X=1.395 $Y=1.96 $X2=0
+ $Y2=0
cc_170 N_A_228_47#_M1004_g N_VPWR_c_350_n 0.00570976f $X=2.15 $Y=2.075 $X2=0
+ $Y2=0
cc_171 N_A_228_47#_M1004_g N_VPWR_c_353_n 0.00429359f $X=2.15 $Y=2.075 $X2=0
+ $Y2=0
cc_172 N_A_228_47#_c_194_n N_VPWR_c_353_n 0.0302883f $X=1.395 $Y=1.96 $X2=0
+ $Y2=0
cc_173 N_A_228_47#_M1001_d N_VPWR_c_348_n 0.00624411f $X=1.14 $Y=1.665 $X2=0
+ $Y2=0
cc_174 N_A_228_47#_M1004_g N_VPWR_c_348_n 0.00810568f $X=2.15 $Y=2.075 $X2=0
+ $Y2=0
cc_175 N_A_228_47#_c_194_n N_VPWR_c_348_n 0.016483f $X=1.395 $Y=1.96 $X2=0 $Y2=0
cc_176 N_A_228_47#_c_185_n N_VGND_c_428_n 0.0136181f $X=1.42 $Y=0.42 $X2=0 $Y2=0
cc_177 N_A_228_47#_M1009_g N_VGND_c_429_n 0.00550872f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_178 N_A_228_47#_M1009_g N_VGND_c_432_n 0.00427134f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_179 N_A_228_47#_c_185_n N_VGND_c_432_n 0.0266893f $X=1.42 $Y=0.42 $X2=0 $Y2=0
cc_180 N_A_228_47#_M1003_d N_VGND_c_437_n 0.00818484f $X=1.14 $Y=0.235 $X2=0
+ $Y2=0
cc_181 N_A_228_47#_M1009_g N_VGND_c_437_n 0.00806408f $X=2.15 $Y=0.56 $X2=0
+ $Y2=0
cc_182 N_A_228_47#_c_185_n N_VGND_c_437_n 0.0145479f $X=1.42 $Y=0.42 $X2=0 $Y2=0
cc_183 N_A_362_333#_c_283_n N_VPWR_M1004_d 0.0269203f $X=2.73 $Y=1.877 $X2=0
+ $Y2=0
cc_184 N_A_362_333#_c_266_n N_VPWR_M1004_d 0.00717703f $X=2.815 $Y=1.79 $X2=0
+ $Y2=0
cc_185 N_A_362_333#_M1002_g N_VPWR_c_350_n 0.00651909f $X=3.01 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_362_333#_c_283_n N_VPWR_c_350_n 0.0269595f $X=2.73 $Y=1.877 $X2=0
+ $Y2=0
cc_187 N_A_362_333#_c_292_n N_VPWR_c_350_n 0.0119041f $X=1.935 $Y=1.96 $X2=0
+ $Y2=0
cc_188 N_A_362_333#_M1007_g N_VPWR_c_352_n 0.0108355f $X=3.44 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_362_333#_c_283_n N_VPWR_c_353_n 0.005634f $X=2.73 $Y=1.877 $X2=0
+ $Y2=0
cc_190 N_A_362_333#_c_292_n N_VPWR_c_353_n 0.016768f $X=1.935 $Y=1.96 $X2=0
+ $Y2=0
cc_191 N_A_362_333#_M1002_g N_VPWR_c_356_n 0.00564131f $X=3.01 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_362_333#_M1007_g N_VPWR_c_356_n 0.00357668f $X=3.44 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_362_333#_M1004_s N_VPWR_c_348_n 0.00286321f $X=1.81 $Y=1.665 $X2=0
+ $Y2=0
cc_194 N_A_362_333#_M1002_g N_VPWR_c_348_n 0.0109768f $X=3.01 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_362_333#_M1007_g N_VPWR_c_348_n 0.00640776f $X=3.44 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_362_333#_c_283_n N_VPWR_c_348_n 0.0128489f $X=2.73 $Y=1.877 $X2=0
+ $Y2=0
cc_197 N_A_362_333#_c_292_n N_VPWR_c_348_n 0.010137f $X=1.935 $Y=1.96 $X2=0
+ $Y2=0
cc_198 N_A_362_333#_M1006_g X 0.00363039f $X=3.01 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A_362_333#_M1002_g X 0.00137005f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_362_333#_c_259_n X 0.00487609f $X=3.365 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_362_333#_M1008_g X 0.0131663f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A_362_333#_M1007_g X 0.00599422f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_362_333#_c_262_n X 0.00776074f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_362_333#_c_263_n X 0.00727645f $X=2.73 $Y=0.82 $X2=0 $Y2=0
cc_205 N_A_362_333#_c_265_n X 0.00610516f $X=2.815 $Y=1.075 $X2=0 $Y2=0
cc_206 N_A_362_333#_c_266_n X 0.00876758f $X=2.815 $Y=1.79 $X2=0 $Y2=0
cc_207 N_A_362_333#_c_322_p X 0.0124998f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_362_333#_M1002_g N_X_c_412_n 0.0141381f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_362_333#_M1007_g N_X_c_412_n 0.0231104f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_362_333#_M1006_g N_X_c_414_n 0.00835009f $X=3.01 $Y=0.445 $X2=0 $Y2=0
cc_211 N_A_362_333#_c_259_n N_X_c_414_n 0.00307898f $X=3.365 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_362_333#_M1008_g N_X_c_414_n 0.0130276f $X=3.44 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A_362_333#_c_322_p N_X_c_414_n 0.00363559f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_362_333#_M1002_g X 0.00469352f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_362_333#_c_259_n X 0.00406403f $X=3.365 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_362_333#_M1007_g X 0.00898252f $X=3.44 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_362_333#_c_322_p X 0.00485852f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_362_333#_c_263_n N_VGND_M1009_d 0.00473336f $X=2.73 $Y=0.82 $X2=0
+ $Y2=0
cc_219 N_A_362_333#_M1006_g N_VGND_c_429_n 0.00634021f $X=3.01 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_362_333#_c_274_n N_VGND_c_429_n 0.0111827f $X=1.94 $Y=0.42 $X2=0
+ $Y2=0
cc_221 N_A_362_333#_c_263_n N_VGND_c_429_n 0.0273508f $X=2.73 $Y=0.82 $X2=0
+ $Y2=0
cc_222 N_A_362_333#_M1008_g N_VGND_c_431_n 0.00681007f $X=3.44 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_362_333#_c_274_n N_VGND_c_432_n 0.0167274f $X=1.94 $Y=0.42 $X2=0
+ $Y2=0
cc_224 N_A_362_333#_c_263_n N_VGND_c_432_n 0.0059052f $X=2.73 $Y=0.82 $X2=0
+ $Y2=0
cc_225 N_A_362_333#_M1006_g N_VGND_c_435_n 0.005323f $X=3.01 $Y=0.445 $X2=0
+ $Y2=0
cc_226 N_A_362_333#_M1008_g N_VGND_c_435_n 0.00357877f $X=3.44 $Y=0.445 $X2=0
+ $Y2=0
cc_227 N_A_362_333#_c_263_n N_VGND_c_435_n 3.26665e-19 $X=2.73 $Y=0.82 $X2=0
+ $Y2=0
cc_228 N_A_362_333#_M1009_s N_VGND_c_437_n 0.00264864f $X=1.815 $Y=0.235 $X2=0
+ $Y2=0
cc_229 N_A_362_333#_M1006_g N_VGND_c_437_n 0.0102001f $X=3.01 $Y=0.445 $X2=0
+ $Y2=0
cc_230 N_A_362_333#_M1008_g N_VGND_c_437_n 0.00640792f $X=3.44 $Y=0.445 $X2=0
+ $Y2=0
cc_231 N_A_362_333#_c_274_n N_VGND_c_437_n 0.0101268f $X=1.94 $Y=0.42 $X2=0
+ $Y2=0
cc_232 N_A_362_333#_c_263_n N_VGND_c_437_n 0.0130726f $X=2.73 $Y=0.82 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_348_n N_X_M1002_s 0.00223231f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_234 N_VPWR_c_356_n N_X_c_412_n 0.0280406f $X=3.72 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VPWR_c_348_n N_X_c_412_n 0.0175137f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_236 N_X_c_414_n N_VGND_c_435_n 0.0283548f $X=3.452 $Y=0.447 $X2=0 $Y2=0
cc_237 N_X_M1006_d N_VGND_c_437_n 0.00223258f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_238 N_X_c_414_n N_VGND_c_437_n 0.0179822f $X=3.452 $Y=0.447 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nor3b_4.spice.SKY130_FD_SC_HD__NOR3B_4.pxi
* Created: Thu Aug 27 14:32:34 2020
* 
x_PM_SKY130_FD_SC_HD__NOR3B_4%C_N N_C_N_c_106_n N_C_N_M1017_g N_C_N_M1004_g C_N
+ N_C_N_c_108_n C_N PM_SKY130_FD_SC_HD__NOR3B_4%C_N
x_PM_SKY130_FD_SC_HD__NOR3B_4%A N_A_c_132_n N_A_M1007_g N_A_M1014_g N_A_c_133_n
+ N_A_M1010_g N_A_M1018_g N_A_c_134_n N_A_M1016_g N_A_M1019_g N_A_c_135_n
+ N_A_M1021_g N_A_M1022_g A A A N_A_c_137_n PM_SKY130_FD_SC_HD__NOR3B_4%A
x_PM_SKY130_FD_SC_HD__NOR3B_4%B N_B_c_205_n N_B_M1002_g N_B_M1000_g N_B_c_206_n
+ N_B_M1011_g N_B_M1003_g N_B_c_207_n N_B_M1012_g N_B_M1006_g N_B_c_208_n
+ N_B_M1025_g N_B_M1013_g B N_B_c_209_n N_B_c_210_n
+ PM_SKY130_FD_SC_HD__NOR3B_4%B
x_PM_SKY130_FD_SC_HD__NOR3B_4%A_27_47# N_A_27_47#_M1017_s N_A_27_47#_M1004_s
+ N_A_27_47#_c_280_n N_A_27_47#_M1001_g N_A_27_47#_M1015_g N_A_27_47#_c_281_n
+ N_A_27_47#_M1005_g N_A_27_47#_M1020_g N_A_27_47#_c_282_n N_A_27_47#_M1008_g
+ N_A_27_47#_M1023_g N_A_27_47#_c_283_n N_A_27_47#_M1009_g N_A_27_47#_M1024_g
+ N_A_27_47#_c_284_n N_A_27_47#_c_295_n N_A_27_47#_c_296_n N_A_27_47#_c_297_n
+ N_A_27_47#_c_285_n N_A_27_47#_c_299_n N_A_27_47#_c_286_n N_A_27_47#_c_287_n
+ N_A_27_47#_c_288_n N_A_27_47#_c_289_n N_A_27_47#_c_335_p N_A_27_47#_c_290_n
+ PM_SKY130_FD_SC_HD__NOR3B_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NOR3B_4%VPWR N_VPWR_M1004_d N_VPWR_M1018_d N_VPWR_M1022_d
+ N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n
+ N_VPWR_c_443_n N_VPWR_c_444_n VPWR N_VPWR_c_445_n N_VPWR_c_446_n
+ N_VPWR_c_437_n N_VPWR_c_448_n PM_SKY130_FD_SC_HD__NOR3B_4%VPWR
x_PM_SKY130_FD_SC_HD__NOR3B_4%A_197_297# N_A_197_297#_M1014_s
+ N_A_197_297#_M1019_s N_A_197_297#_M1000_d N_A_197_297#_M1006_d
+ N_A_197_297#_c_534_n N_A_197_297#_c_533_n N_A_197_297#_c_538_n
+ N_A_197_297#_c_547_n N_A_197_297#_c_548_n N_A_197_297#_c_549_n
+ N_A_197_297#_c_550_n PM_SKY130_FD_SC_HD__NOR3B_4%A_197_297#
x_PM_SKY130_FD_SC_HD__NOR3B_4%A_555_297# N_A_555_297#_M1000_s
+ N_A_555_297#_M1003_s N_A_555_297#_M1013_s N_A_555_297#_M1020_s
+ N_A_555_297#_M1024_s N_A_555_297#_c_582_n N_A_555_297#_c_584_n
+ N_A_555_297#_c_590_n N_A_555_297#_c_591_n N_A_555_297#_c_632_p
+ N_A_555_297#_c_581_n N_A_555_297#_c_636_p N_A_555_297#_c_608_n
+ N_A_555_297#_c_611_n N_A_555_297#_c_613_n N_A_555_297#_c_615_n
+ PM_SKY130_FD_SC_HD__NOR3B_4%A_555_297#
x_PM_SKY130_FD_SC_HD__NOR3B_4%Y N_Y_M1007_s N_Y_M1016_s N_Y_M1002_d N_Y_M1012_d
+ N_Y_M1001_s N_Y_M1008_s N_Y_M1015_d N_Y_M1023_d N_Y_c_662_n N_Y_c_641_n
+ N_Y_c_642_n N_Y_c_674_n N_Y_c_643_n N_Y_c_685_n N_Y_c_644_n N_Y_c_692_n
+ N_Y_c_645_n N_Y_c_696_n N_Y_c_655_n N_Y_c_646_n N_Y_c_726_n N_Y_c_656_n
+ N_Y_c_647_n N_Y_c_648_n N_Y_c_649_n N_Y_c_650_n N_Y_c_651_n N_Y_c_652_n
+ N_Y_c_658_n N_Y_c_653_n N_Y_c_659_n N_Y_c_654_n N_Y_c_660_n Y
+ PM_SKY130_FD_SC_HD__NOR3B_4%Y
x_PM_SKY130_FD_SC_HD__NOR3B_4%VGND N_VGND_M1017_d N_VGND_M1010_d N_VGND_M1021_d
+ N_VGND_M1011_s N_VGND_M1025_s N_VGND_M1005_d N_VGND_M1009_d N_VGND_c_821_n
+ N_VGND_c_822_n N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n
+ N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n
+ N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n VGND
+ N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n
+ N_VGND_c_841_n VGND PM_SKY130_FD_SC_HD__NOR3B_4%VGND
cc_1 VNB N_C_N_c_106_n 0.0216587f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB C_N 0.00777182f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_108_n 0.0392772f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_4 VNB N_A_c_132_n 0.0160955f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_5 VNB N_A_c_133_n 0.0157835f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_A_c_134_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_c_135_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB A 0.0120429f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_c_137_n 0.0702338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_c_205_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_11 VNB N_B_c_206_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB N_B_c_207_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B_c_208_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B_c_209_n 0.00258951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B_c_210_n 0.0702655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_280_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_281_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_18 VNB N_A_27_47#_c_282_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_283_n 0.0194103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_284_n 0.0185703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_285_n 0.00785066f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_286_n 3.4592e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_287_n 0.0029651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_288_n 0.00281766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_289_n 0.0101457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_290_n 0.0661726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_437_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_641_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_642_n 0.00253838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_643_n 0.00964455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_644_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_645_n 0.00302181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_646_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_647_n 0.0047059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_648_n 0.0237454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_649_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_650_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_651_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_652_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_653_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_654_n 0.0344618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_821_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_822_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_823_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_824_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_825_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_826_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_827_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_828_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_829_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_830_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_831_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_832_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_833_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_834_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_835_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_836_n 0.0171305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_837_n 0.339005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_838_n 0.02106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_839_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_840_n 0.0197313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_841_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VPB N_C_N_M1004_g 0.0254923f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_64 VPB N_C_N_c_108_n 0.00961737f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_65 VPB N_A_M1014_g 0.0184438f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_66 VPB N_A_M1018_g 0.0181992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_M1019_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_M1022_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_c_137_n 0.010875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B_M1000_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_71 VPB N_B_M1003_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_B_M1006_g 0.0182005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B_M1013_g 0.0184463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B_c_210_n 0.0108754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_M1015_g 0.0187749f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_76 VPB N_A_27_47#_M1020_g 0.0181974f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.18
cc_77 VPB N_A_27_47#_M1023_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_M1024_g 0.0222777f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_295_n 0.00893204f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_296_n 0.0317613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_297_n 7.09682e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_285_n 0.00270308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_299_n 0.030335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_286_n 0.00271274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_290_n 0.0103367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_438_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_87 VPB N_VPWR_c_439_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.18
cc_88 VPB N_VPWR_c_440_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_441_n 0.0157745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_442_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_443_n 0.0151708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_444_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_445_n 0.0176845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_446_n 0.104372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_437_n 0.0591391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_448_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_197_297#_c_533_n 0.0081428f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.18
cc_98 VPB N_A_555_297#_c_581_n 0.00316323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_Y_c_655_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_Y_c_656_n 0.00548674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_Y_c_648_n 0.00915831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_Y_c_658_n 0.00225182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_Y_c_659_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_Y_c_660_n 0.014519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB Y 0.0412233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 N_C_N_c_106_n N_A_c_132_n 0.0215572f $X=0.49 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_107 N_C_N_M1004_g N_A_M1014_g 0.0215572f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_108 N_C_N_c_108_n N_A_c_137_n 0.0215572f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_109 N_C_N_c_106_n N_A_27_47#_c_284_n 0.00658926f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_110 C_N N_A_27_47#_c_295_n 0.0241321f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_111 N_C_N_c_108_n N_A_27_47#_c_295_n 0.00721245f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_112 N_C_N_M1004_g N_A_27_47#_c_297_n 0.0148713f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_113 C_N N_A_27_47#_c_297_n 0.00275577f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_114 N_C_N_c_108_n N_A_27_47#_c_297_n 2.32632e-19 $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C_N_c_106_n N_A_27_47#_c_285_n 0.00996914f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_116 C_N N_A_27_47#_c_285_n 0.0157255f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_117 N_C_N_c_106_n N_A_27_47#_c_289_n 0.0109062f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_118 C_N N_A_27_47#_c_289_n 0.0242211f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_119 N_C_N_c_108_n N_A_27_47#_c_289_n 0.0075174f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C_N_M1004_g N_VPWR_c_438_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_121 N_C_N_M1004_g N_VPWR_c_445_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_122 N_C_N_M1004_g N_VPWR_c_437_n 0.0114368f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_123 N_C_N_c_106_n N_Y_c_662_n 5.22228e-19 $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_124 N_C_N_c_106_n N_VGND_c_821_n 0.00268723f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_125 N_C_N_c_106_n N_VGND_c_837_n 0.00675096f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_126 N_C_N_c_106_n N_VGND_c_838_n 0.00423442f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_127 A N_B_c_209_n 0.0109093f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_128 A N_B_c_210_n 0.0014919f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_129 N_A_c_132_n N_A_27_47#_c_284_n 5.52269e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_132_n N_A_27_47#_c_285_n 0.0104052f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_131 A N_A_27_47#_c_285_n 0.012421f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A_M1014_g N_A_27_47#_c_299_n 0.0189403f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_M1018_g N_A_27_47#_c_299_n 0.0103677f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_M1019_g N_A_27_47#_c_299_n 0.0103677f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1022_g N_A_27_47#_c_299_n 0.0124706f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_136 A N_A_27_47#_c_299_n 0.120277f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A_c_137_n N_A_27_47#_c_299_n 0.00634526f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_132_n N_A_27_47#_c_289_n 7.62115e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_M1014_g N_VPWR_c_438_n 0.00157837f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1018_g N_VPWR_c_439_n 0.00157837f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1019_g N_VPWR_c_439_n 0.00157837f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1022_g N_VPWR_c_440_n 0.00338128f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1014_g N_VPWR_c_441_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1018_g N_VPWR_c_441_n 0.00441875f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1019_g N_VPWR_c_443_n 0.00441875f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1022_g N_VPWR_c_443_n 0.00441875f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1014_g N_VPWR_c_437_n 0.010464f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1018_g N_VPWR_c_437_n 0.00586018f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1019_g N_VPWR_c_437_n 0.00586018f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1022_g N_VPWR_c_437_n 0.00718625f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_M1018_g N_A_197_297#_c_534_n 0.0102286f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1019_g N_A_197_297#_c_534_n 0.0101845f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_M1022_g N_A_197_297#_c_533_n 0.0123316f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_c_132_n N_Y_c_662_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_133_n N_Y_c_662_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_c_134_n N_Y_c_662_n 5.22228e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_133_n N_Y_c_641_n 0.00870364f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_134_n N_Y_c_641_n 0.00870364f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_159 A N_Y_c_641_n 0.0362443f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_160 N_A_c_137_n N_Y_c_641_n 0.00222133f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_c_132_n N_Y_c_642_n 0.00296109f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_133_n N_Y_c_642_n 0.00112129f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_163 A N_Y_c_642_n 0.0202409f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A_c_137_n N_Y_c_642_n 0.00230339f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_c_133_n N_Y_c_674_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_c_134_n N_Y_c_674_n 0.00630972f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_135_n N_Y_c_674_n 0.0109565f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_135_n N_Y_c_643_n 0.0109318f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_169 A N_Y_c_643_n 0.0424717f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_170 N_A_c_134_n N_Y_c_649_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_c_135_n N_Y_c_649_n 0.00113286f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_172 A N_Y_c_649_n 0.0266272f $X=2.45 $Y=1.105 $X2=0 $Y2=0
cc_173 N_A_c_137_n N_Y_c_649_n 0.00230339f $X=2.17 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_c_132_n N_VGND_c_821_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_c_133_n N_VGND_c_822_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_134_n N_VGND_c_822_n 0.00146339f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_132_n N_VGND_c_828_n 0.00541359f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_133_n N_VGND_c_828_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_132_n N_VGND_c_837_n 0.00952874f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_133_n N_VGND_c_837_n 0.0057163f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_134_n N_VGND_c_837_n 0.0057163f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_c_135_n N_VGND_c_837_n 0.0070399f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_134_n N_VGND_c_839_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_c_135_n N_VGND_c_839_n 0.00423334f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_135_n N_VGND_c_840_n 0.00335921f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B_c_208_n N_A_27_47#_c_280_n 0.0228037f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_187 N_B_M1013_g N_A_27_47#_M1015_g 0.0228037f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B_M1000_g N_A_27_47#_c_299_n 0.0124706f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B_M1003_g N_A_27_47#_c_299_n 0.0103677f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_190 N_B_M1006_g N_A_27_47#_c_299_n 0.0103235f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_191 N_B_M1013_g N_A_27_47#_c_299_n 0.0140908f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B_c_209_n N_A_27_47#_c_299_n 0.0901988f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B_c_210_n N_A_27_47#_c_299_n 0.00634526f $X=4.37 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B_c_210_n N_A_27_47#_c_286_n 0.00388409f $X=4.37 $Y=1.16 $X2=0 $Y2=0
cc_195 N_B_c_209_n N_A_27_47#_c_287_n 0.0145223f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B_c_210_n N_A_27_47#_c_287_n 0.0021925f $X=4.37 $Y=1.16 $X2=0 $Y2=0
cc_197 N_B_c_210_n N_A_27_47#_c_290_n 0.0228037f $X=4.37 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B_M1000_g N_VPWR_c_440_n 0.00214938f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B_M1000_g N_VPWR_c_446_n 0.00357877f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B_M1003_g N_VPWR_c_446_n 0.00357877f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_201 N_B_M1006_g N_VPWR_c_446_n 0.00357877f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B_M1013_g N_VPWR_c_446_n 0.00357877f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B_M1000_g N_VPWR_c_437_n 0.00655123f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_204 N_B_M1003_g N_VPWR_c_437_n 0.00522516f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B_M1006_g N_VPWR_c_437_n 0.00522516f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B_M1013_g N_VPWR_c_437_n 0.00525237f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B_M1000_g N_A_197_297#_c_533_n 0.0113377f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B_M1003_g N_A_197_297#_c_538_n 0.00919056f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B_M1006_g N_A_197_297#_c_538_n 0.00919056f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B_M1000_g N_A_555_297#_c_582_n 0.00846708f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B_M1003_g N_A_555_297#_c_582_n 0.00846708f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B_M1006_g N_A_555_297#_c_584_n 0.00851124f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B_M1013_g N_A_555_297#_c_584_n 0.00984328f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B_c_205_n N_Y_c_643_n 0.0109318f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B_c_209_n N_Y_c_643_n 0.00826974f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B_c_205_n N_Y_c_685_n 0.0109565f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B_c_206_n N_Y_c_685_n 0.00630972f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B_c_207_n N_Y_c_685_n 5.22228e-19 $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B_c_206_n N_Y_c_644_n 0.00870364f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B_c_207_n N_Y_c_644_n 0.00870364f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B_c_209_n N_Y_c_644_n 0.0362443f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B_c_210_n N_Y_c_644_n 0.00222133f $X=4.37 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B_c_206_n N_Y_c_692_n 5.22228e-19 $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B_c_207_n N_Y_c_692_n 0.00630972f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B_c_208_n N_Y_c_692_n 0.00630972f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B_c_208_n N_Y_c_645_n 0.0101343f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_227 N_B_c_208_n N_Y_c_696_n 5.22228e-19 $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B_c_205_n N_Y_c_650_n 0.00113286f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B_c_206_n N_Y_c_650_n 0.00113286f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B_c_209_n N_Y_c_650_n 0.0266272f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B_c_210_n N_Y_c_650_n 0.00230339f $X=4.37 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B_c_207_n N_Y_c_651_n 0.00113286f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B_c_208_n N_Y_c_651_n 0.00145053f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B_c_209_n N_Y_c_651_n 0.0247016f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B_c_210_n N_Y_c_651_n 0.00230339f $X=4.37 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B_c_206_n N_VGND_c_823_n 0.00146339f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B_c_207_n N_VGND_c_823_n 0.00146448f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B_c_208_n N_VGND_c_824_n 0.00146448f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B_c_205_n N_VGND_c_830_n 0.00423334f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B_c_206_n N_VGND_c_830_n 0.00423334f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B_c_207_n N_VGND_c_832_n 0.00423334f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B_c_208_n N_VGND_c_832_n 0.00423334f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_243 N_B_c_205_n N_VGND_c_837_n 0.0070399f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_244 N_B_c_206_n N_VGND_c_837_n 0.0057163f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_245 N_B_c_207_n N_VGND_c_837_n 0.0057163f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B_c_208_n N_VGND_c_837_n 0.0057435f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B_c_205_n N_VGND_c_840_n 0.00335921f $X=3.11 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_335_p N_VPWR_M1004_d 0.00172935f $X=0.7 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_249 N_A_27_47#_c_299_n N_VPWR_M1018_d 0.00166235f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_299_n N_VPWR_M1022_d 0.00276803f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_335_p N_VPWR_c_438_n 0.0141251f $X=0.7 $Y=1.54 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_296_n N_VPWR_c_445_n 0.0190343f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1015_g N_VPWR_c_446_n 0.00357877f $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1020_g N_VPWR_c_446_n 0.00357877f $X=5.21 $Y=1.985 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1023_g N_VPWR_c_446_n 0.00357877f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1024_g N_VPWR_c_446_n 0.00357877f $X=6.05 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1004_s N_VPWR_c_437_n 0.00260431f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1015_g N_VPWR_c_437_n 0.00525237f $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1020_g N_VPWR_c_437_n 0.00522516f $X=5.21 $Y=1.985 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1023_g N_VPWR_c_437_n 0.00522516f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_M1024_g N_VPWR_c_437_n 0.00655123f $X=6.05 $Y=1.985 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_296_n N_VPWR_c_437_n 0.0112839f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_299_n N_A_197_297#_M1014_s 0.00165831f $X=4.535 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_264 N_A_27_47#_c_299_n N_A_197_297#_M1019_s 0.00165831f $X=4.535 $Y=1.54
+ $X2=0 $Y2=0
cc_265 N_A_27_47#_c_299_n N_A_197_297#_M1000_d 0.00165831f $X=4.535 $Y=1.54
+ $X2=0 $Y2=0
cc_266 N_A_27_47#_c_299_n N_A_197_297#_M1006_d 0.00165831f $X=4.535 $Y=1.54
+ $X2=0 $Y2=0
cc_267 N_A_27_47#_c_299_n N_A_197_297#_c_534_n 0.0315971f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_299_n N_A_197_297#_c_533_n 0.0700867f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_299_n N_A_197_297#_c_538_n 0.0315971f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_299_n N_A_197_297#_c_547_n 0.0126766f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_299_n N_A_197_297#_c_548_n 0.0126766f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_299_n N_A_197_297#_c_549_n 0.01198f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_299_n N_A_197_297#_c_550_n 0.01198f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_299_n N_A_555_297#_M1000_s 0.00276803f $X=4.535 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_275 N_A_27_47#_c_299_n N_A_555_297#_M1003_s 0.00166235f $X=4.535 $Y=1.54
+ $X2=0 $Y2=0
cc_276 N_A_27_47#_c_299_n N_A_555_297#_M1013_s 0.00194825f $X=4.535 $Y=1.54
+ $X2=0 $Y2=0
cc_277 N_A_27_47#_c_299_n N_A_555_297#_c_584_n 0.00321995f $X=4.535 $Y=1.54
+ $X2=0 $Y2=0
cc_278 N_A_27_47#_c_299_n N_A_555_297#_c_590_n 0.0135511f $X=4.535 $Y=1.54 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1015_g N_A_555_297#_c_591_n 0.0121747f $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1020_g N_A_555_297#_c_591_n 0.00988743f $X=5.21 $Y=1.985
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_M1023_g N_A_555_297#_c_581_n 0.00984328f $X=5.63 $Y=1.985
+ $X2=0 $Y2=0
cc_282 N_A_27_47#_M1024_g N_A_555_297#_c_581_n 0.00988743f $X=6.05 $Y=1.985
+ $X2=0 $Y2=0
cc_283 N_A_27_47#_c_284_n N_Y_c_662_n 0.00519135f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_284_n N_Y_c_642_n 3.24781e-19 $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_299_n N_Y_c_642_n 0.00272444f $X=4.535 $Y=1.54 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_289_n N_Y_c_642_n 0.00795243f $X=0.7 $Y=0.82 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_299_n N_Y_c_643_n 0.0115608f $X=4.535 $Y=1.54 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_280_n N_Y_c_692_n 5.22228e-19 $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_280_n N_Y_c_645_n 0.00865686f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_299_n N_Y_c_645_n 0.00610178f $X=4.535 $Y=1.54 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_287_n N_Y_c_645_n 0.0141654f $X=4.705 $Y=1.18 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_288_n N_Y_c_645_n 0.00899944f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_280_n N_Y_c_696_n 0.00630972f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_281_n N_Y_c_696_n 0.00630972f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_282_n N_Y_c_696_n 5.22228e-19 $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A_27_47#_M1020_g N_Y_c_655_n 0.0109258f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A_27_47#_M1023_g N_Y_c_655_n 0.01094f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_288_n N_Y_c_655_n 0.0416643f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A_27_47#_c_290_n N_Y_c_655_n 0.00211509f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_281_n N_Y_c_646_n 0.00870364f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_282_n N_Y_c_646_n 0.00870364f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_288_n N_Y_c_646_n 0.0362443f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_290_n N_Y_c_646_n 0.00222133f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_281_n N_Y_c_726_n 5.22228e-19 $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_282_n N_Y_c_726_n 0.00630972f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_283_n N_Y_c_726_n 0.00681571f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_27_47#_M1024_g N_Y_c_656_n 0.012984f $X=6.05 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_288_n N_Y_c_656_n 0.0110239f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_309 N_A_27_47#_c_283_n N_Y_c_647_n 0.0108225f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_288_n N_Y_c_647_n 0.00826974f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_283_n N_Y_c_648_n 0.00605338f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_288_n N_Y_c_648_n 0.0115725f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_290_n N_Y_c_648_n 0.0071926f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_27_47#_c_299_n N_Y_c_651_n 7.21395e-19 $X=4.535 $Y=1.54 $X2=0 $Y2=0
cc_315 N_A_27_47#_c_280_n N_Y_c_652_n 0.00113286f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_281_n N_Y_c_652_n 0.00113286f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_288_n N_Y_c_652_n 0.0266272f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_27_47#_c_290_n N_Y_c_652_n 0.00230339f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_27_47#_M1015_g N_Y_c_658_n 2.57315e-19 $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A_27_47#_c_299_n N_Y_c_658_n 0.00271526f $X=4.535 $Y=1.54 $X2=0 $Y2=0
cc_321 N_A_27_47#_c_288_n N_Y_c_658_n 0.0204292f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A_27_47#_c_290_n N_Y_c_658_n 0.00219557f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_27_47#_c_282_n N_Y_c_653_n 0.00113286f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_27_47#_c_283_n N_Y_c_653_n 0.00113286f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_27_47#_c_288_n N_Y_c_653_n 0.0266272f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A_27_47#_c_290_n N_Y_c_653_n 0.00230339f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_27_47#_c_288_n N_Y_c_659_n 0.0204292f $X=5.9 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_27_47#_c_290_n N_Y_c_659_n 0.00219557f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_27_47#_c_283_n N_Y_c_654_n 0.00296375f $X=6.05 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_27_47#_M1024_g Y 0.00322377f $X=6.05 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A_27_47#_c_289_n N_VGND_M1017_d 0.0019056f $X=0.7 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_332 N_A_27_47#_c_289_n N_VGND_c_821_n 0.0116529f $X=0.7 $Y=0.82 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_280_n N_VGND_c_824_n 0.00146448f $X=4.79 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_281_n N_VGND_c_825_n 0.00146448f $X=5.21 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_282_n N_VGND_c_825_n 0.00146448f $X=5.63 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_282_n N_VGND_c_826_n 0.00423334f $X=5.63 $Y=0.995 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_283_n N_VGND_c_826_n 0.00423334f $X=6.05 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_283_n N_VGND_c_827_n 0.00316354f $X=6.05 $Y=0.995 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_280_n N_VGND_c_834_n 0.00423334f $X=4.79 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_281_n N_VGND_c_834_n 0.00423334f $X=5.21 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_M1017_s N_VGND_c_837_n 0.00225715f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_280_n N_VGND_c_837_n 0.0057435f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_343 N_A_27_47#_c_281_n N_VGND_c_837_n 0.0057163f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A_27_47#_c_282_n N_VGND_c_837_n 0.0057163f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A_27_47#_c_283_n N_VGND_c_837_n 0.00704237f $X=6.05 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_284_n N_VGND_c_837_n 0.0125062f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_347 N_A_27_47#_c_289_n N_VGND_c_837_n 0.00451353f $X=0.7 $Y=0.82 $X2=0 $Y2=0
cc_348 N_A_27_47#_c_284_n N_VGND_c_838_n 0.0208864f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_349 N_A_27_47#_c_289_n N_VGND_c_838_n 0.00197124f $X=0.7 $Y=0.82 $X2=0 $Y2=0
cc_350 N_VPWR_c_437_n N_A_197_297#_M1014_s 0.00253991f $X=6.67 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_351 N_VPWR_c_437_n N_A_197_297#_M1019_s 0.0022335f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_437_n N_A_197_297#_M1000_d 0.00215227f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_437_n N_A_197_297#_M1006_d 0.0021603f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_354 N_VPWR_M1018_d N_A_197_297#_c_534_n 0.0031712f $X=1.405 $Y=1.485 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_439_n N_A_197_297#_c_534_n 0.0123012f $X=1.54 $Y=2.3 $X2=0 $Y2=0
cc_356 N_VPWR_c_441_n N_A_197_297#_c_534_n 0.00201582f $X=1.415 $Y=2.72 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_443_n N_A_197_297#_c_534_n 0.00201582f $X=2.255 $Y=2.72 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_437_n N_A_197_297#_c_534_n 0.00800071f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_359 N_VPWR_M1022_d N_A_197_297#_c_533_n 0.00500976f $X=2.245 $Y=1.485 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_440_n N_A_197_297#_c_533_n 0.0159284f $X=2.38 $Y=2.3 $X2=0 $Y2=0
cc_361 N_VPWR_c_443_n N_A_197_297#_c_533_n 0.00201582f $X=2.255 $Y=2.72 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_446_n N_A_197_297#_c_533_n 0.0039015f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_363 N_VPWR_c_437_n N_A_197_297#_c_533_n 0.012288f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_437_n N_A_197_297#_c_538_n 0.00125448f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_441_n N_A_197_297#_c_547_n 0.0142224f $X=1.415 $Y=2.72 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_437_n N_A_197_297#_c_547_n 0.00954719f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_443_n N_A_197_297#_c_548_n 0.0142224f $X=2.255 $Y=2.72 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_437_n N_A_197_297#_c_548_n 0.00954719f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_437_n N_A_555_297#_M1000_s 0.00207714f $X=6.67 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_370 N_VPWR_c_437_n N_A_555_297#_M1003_s 0.00213597f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_437_n N_A_555_297#_M1013_s 0.00215203f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_437_n N_A_555_297#_M1020_s 0.00215203f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_437_n N_A_555_297#_M1024_s 0.0020932f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_446_n N_A_555_297#_c_582_n 0.0330174f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_437_n N_A_555_297#_c_582_n 0.0204707f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_446_n N_A_555_297#_c_584_n 0.0330174f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_437_n N_A_555_297#_c_584_n 0.0204667f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_446_n N_A_555_297#_c_591_n 0.0330174f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_437_n N_A_555_297#_c_591_n 0.0204627f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_446_n N_A_555_297#_c_581_n 0.0489446f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_437_n N_A_555_297#_c_581_n 0.0300869f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_440_n N_A_555_297#_c_608_n 0.0180653f $X=2.38 $Y=2.3 $X2=0 $Y2=0
cc_383 N_VPWR_c_446_n N_A_555_297#_c_608_n 0.0151213f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_437_n N_A_555_297#_c_608_n 0.00938089f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_446_n N_A_555_297#_c_611_n 0.0136817f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_437_n N_A_555_297#_c_611_n 0.00938089f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_446_n N_A_555_297#_c_613_n 0.0142933f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_437_n N_A_555_297#_c_613_n 0.00962421f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_446_n N_A_555_297#_c_615_n 0.0142933f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_437_n N_A_555_297#_c_615_n 0.00962421f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_437_n N_Y_M1015_d 0.00216833f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_c_437_n N_Y_M1023_d 0.00216833f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_446_n Y 0.011051f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_c_437_n Y 0.0076223f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_395 N_A_197_297#_c_533_n N_A_555_297#_M1000_s 0.00500976f $X=3.195 $Y=1.88
+ $X2=-0.19 $Y2=1.305
cc_396 N_A_197_297#_c_538_n N_A_555_297#_M1003_s 0.0031712f $X=4.035 $Y=1.88
+ $X2=0 $Y2=0
cc_397 N_A_197_297#_M1000_d N_A_555_297#_c_582_n 0.00312348f $X=3.185 $Y=1.485
+ $X2=0 $Y2=0
cc_398 N_A_197_297#_c_533_n N_A_555_297#_c_582_n 0.00520504f $X=3.195 $Y=1.88
+ $X2=0 $Y2=0
cc_399 N_A_197_297#_c_538_n N_A_555_297#_c_582_n 0.00520504f $X=4.035 $Y=1.88
+ $X2=0 $Y2=0
cc_400 N_A_197_297#_c_549_n N_A_555_297#_c_582_n 0.0112564f $X=3.32 $Y=1.88
+ $X2=0 $Y2=0
cc_401 N_A_197_297#_M1006_d N_A_555_297#_c_584_n 0.00312348f $X=4.025 $Y=1.485
+ $X2=0 $Y2=0
cc_402 N_A_197_297#_c_538_n N_A_555_297#_c_584_n 0.00520504f $X=4.035 $Y=1.88
+ $X2=0 $Y2=0
cc_403 N_A_197_297#_c_550_n N_A_555_297#_c_584_n 0.0112564f $X=4.16 $Y=1.88
+ $X2=0 $Y2=0
cc_404 N_A_197_297#_c_533_n N_A_555_297#_c_608_n 0.0150265f $X=3.195 $Y=1.88
+ $X2=0 $Y2=0
cc_405 N_A_197_297#_c_538_n N_A_555_297#_c_611_n 0.0116046f $X=4.035 $Y=1.88
+ $X2=0 $Y2=0
cc_406 N_A_555_297#_c_591_n N_Y_M1015_d 0.00312348f $X=5.295 $Y=2.38 $X2=0 $Y2=0
cc_407 N_A_555_297#_c_581_n N_Y_M1023_d 0.00312348f $X=6.135 $Y=2.38 $X2=0 $Y2=0
cc_408 N_A_555_297#_M1020_s N_Y_c_655_n 0.00165831f $X=5.285 $Y=1.485 $X2=0
+ $Y2=0
cc_409 N_A_555_297#_c_591_n N_Y_c_655_n 0.00320918f $X=5.295 $Y=2.38 $X2=0 $Y2=0
cc_410 N_A_555_297#_c_632_p N_Y_c_655_n 0.0126766f $X=5.42 $Y=1.96 $X2=0 $Y2=0
cc_411 N_A_555_297#_c_581_n N_Y_c_655_n 0.00320918f $X=6.135 $Y=2.38 $X2=0 $Y2=0
cc_412 N_A_555_297#_M1024_s N_Y_c_656_n 0.00276279f $X=6.125 $Y=1.485 $X2=0
+ $Y2=0
cc_413 N_A_555_297#_c_581_n N_Y_c_656_n 0.00320918f $X=6.135 $Y=2.38 $X2=0 $Y2=0
cc_414 N_A_555_297#_c_636_p N_Y_c_656_n 0.0164145f $X=6.26 $Y=1.96 $X2=0 $Y2=0
cc_415 N_A_555_297#_c_591_n N_Y_c_658_n 0.0118729f $X=5.295 $Y=2.38 $X2=0 $Y2=0
cc_416 N_A_555_297#_c_581_n N_Y_c_659_n 0.0118729f $X=6.135 $Y=2.38 $X2=0 $Y2=0
cc_417 N_A_555_297#_c_581_n Y 0.0100535f $X=6.135 $Y=2.38 $X2=0 $Y2=0
cc_418 N_A_555_297#_c_636_p Y 0.0385675f $X=6.26 $Y=1.96 $X2=0 $Y2=0
cc_419 N_Y_c_641_n N_VGND_M1010_d 0.00162089f $X=1.795 $Y=0.815 $X2=0 $Y2=0
cc_420 N_Y_c_643_n N_VGND_M1021_d 0.0108248f $X=3.155 $Y=0.815 $X2=0 $Y2=0
cc_421 N_Y_c_644_n N_VGND_M1011_s 0.00162089f $X=3.995 $Y=0.815 $X2=0 $Y2=0
cc_422 N_Y_c_645_n N_VGND_M1025_s 0.00162089f $X=4.835 $Y=0.815 $X2=0 $Y2=0
cc_423 N_Y_c_646_n N_VGND_M1005_d 0.00162089f $X=5.675 $Y=0.815 $X2=0 $Y2=0
cc_424 N_Y_c_647_n N_VGND_M1009_d 0.00315681f $X=6.42 $Y=0.815 $X2=0 $Y2=0
cc_425 N_Y_c_641_n N_VGND_c_822_n 0.0122559f $X=1.795 $Y=0.815 $X2=0 $Y2=0
cc_426 N_Y_c_644_n N_VGND_c_823_n 0.0122559f $X=3.995 $Y=0.815 $X2=0 $Y2=0
cc_427 N_Y_c_645_n N_VGND_c_824_n 0.0122559f $X=4.835 $Y=0.815 $X2=0 $Y2=0
cc_428 N_Y_c_646_n N_VGND_c_825_n 0.0122559f $X=5.675 $Y=0.815 $X2=0 $Y2=0
cc_429 N_Y_c_646_n N_VGND_c_826_n 0.00198695f $X=5.675 $Y=0.815 $X2=0 $Y2=0
cc_430 N_Y_c_726_n N_VGND_c_826_n 0.0188551f $X=5.84 $Y=0.39 $X2=0 $Y2=0
cc_431 N_Y_c_647_n N_VGND_c_826_n 0.00198695f $X=6.42 $Y=0.815 $X2=0 $Y2=0
cc_432 N_Y_c_647_n N_VGND_c_827_n 0.0127273f $X=6.42 $Y=0.815 $X2=0 $Y2=0
cc_433 N_Y_c_654_n N_VGND_c_827_n 0.0182672f $X=6.59 $Y=0.815 $X2=0 $Y2=0
cc_434 N_Y_c_662_n N_VGND_c_828_n 0.0188551f $X=1.12 $Y=0.39 $X2=0 $Y2=0
cc_435 N_Y_c_641_n N_VGND_c_828_n 0.00198695f $X=1.795 $Y=0.815 $X2=0 $Y2=0
cc_436 N_Y_c_643_n N_VGND_c_830_n 0.00198695f $X=3.155 $Y=0.815 $X2=0 $Y2=0
cc_437 N_Y_c_685_n N_VGND_c_830_n 0.0188551f $X=3.32 $Y=0.39 $X2=0 $Y2=0
cc_438 N_Y_c_644_n N_VGND_c_830_n 0.00198695f $X=3.995 $Y=0.815 $X2=0 $Y2=0
cc_439 N_Y_c_644_n N_VGND_c_832_n 0.00198695f $X=3.995 $Y=0.815 $X2=0 $Y2=0
cc_440 N_Y_c_692_n N_VGND_c_832_n 0.0188551f $X=4.16 $Y=0.39 $X2=0 $Y2=0
cc_441 N_Y_c_645_n N_VGND_c_832_n 0.00198695f $X=4.835 $Y=0.815 $X2=0 $Y2=0
cc_442 N_Y_c_645_n N_VGND_c_834_n 0.00198695f $X=4.835 $Y=0.815 $X2=0 $Y2=0
cc_443 N_Y_c_696_n N_VGND_c_834_n 0.0188551f $X=5 $Y=0.39 $X2=0 $Y2=0
cc_444 N_Y_c_646_n N_VGND_c_834_n 0.00198695f $X=5.675 $Y=0.815 $X2=0 $Y2=0
cc_445 N_Y_c_647_n N_VGND_c_836_n 0.00110192f $X=6.42 $Y=0.815 $X2=0 $Y2=0
cc_446 N_Y_c_654_n N_VGND_c_836_n 0.0142348f $X=6.59 $Y=0.815 $X2=0 $Y2=0
cc_447 N_Y_M1007_s N_VGND_c_837_n 0.00215201f $X=0.985 $Y=0.235 $X2=0 $Y2=0
cc_448 N_Y_M1016_s N_VGND_c_837_n 0.00215201f $X=1.825 $Y=0.235 $X2=0 $Y2=0
cc_449 N_Y_M1002_d N_VGND_c_837_n 0.00215201f $X=3.185 $Y=0.235 $X2=0 $Y2=0
cc_450 N_Y_M1012_d N_VGND_c_837_n 0.00215201f $X=4.025 $Y=0.235 $X2=0 $Y2=0
cc_451 N_Y_M1001_s N_VGND_c_837_n 0.00215201f $X=4.865 $Y=0.235 $X2=0 $Y2=0
cc_452 N_Y_M1008_s N_VGND_c_837_n 0.00215201f $X=5.705 $Y=0.235 $X2=0 $Y2=0
cc_453 N_Y_c_662_n N_VGND_c_837_n 0.0122069f $X=1.12 $Y=0.39 $X2=0 $Y2=0
cc_454 N_Y_c_641_n N_VGND_c_837_n 0.00835832f $X=1.795 $Y=0.815 $X2=0 $Y2=0
cc_455 N_Y_c_674_n N_VGND_c_837_n 0.0122069f $X=1.96 $Y=0.39 $X2=0 $Y2=0
cc_456 N_Y_c_643_n N_VGND_c_837_n 0.0103256f $X=3.155 $Y=0.815 $X2=0 $Y2=0
cc_457 N_Y_c_685_n N_VGND_c_837_n 0.0122069f $X=3.32 $Y=0.39 $X2=0 $Y2=0
cc_458 N_Y_c_644_n N_VGND_c_837_n 0.00835832f $X=3.995 $Y=0.815 $X2=0 $Y2=0
cc_459 N_Y_c_692_n N_VGND_c_837_n 0.0122069f $X=4.16 $Y=0.39 $X2=0 $Y2=0
cc_460 N_Y_c_645_n N_VGND_c_837_n 0.00835832f $X=4.835 $Y=0.815 $X2=0 $Y2=0
cc_461 N_Y_c_696_n N_VGND_c_837_n 0.0122069f $X=5 $Y=0.39 $X2=0 $Y2=0
cc_462 N_Y_c_646_n N_VGND_c_837_n 0.00835832f $X=5.675 $Y=0.815 $X2=0 $Y2=0
cc_463 N_Y_c_726_n N_VGND_c_837_n 0.0122069f $X=5.84 $Y=0.39 $X2=0 $Y2=0
cc_464 N_Y_c_647_n N_VGND_c_837_n 0.0065194f $X=6.42 $Y=0.815 $X2=0 $Y2=0
cc_465 N_Y_c_654_n N_VGND_c_837_n 0.0117488f $X=6.59 $Y=0.815 $X2=0 $Y2=0
cc_466 N_Y_c_641_n N_VGND_c_839_n 0.00198695f $X=1.795 $Y=0.815 $X2=0 $Y2=0
cc_467 N_Y_c_674_n N_VGND_c_839_n 0.0188551f $X=1.96 $Y=0.39 $X2=0 $Y2=0
cc_468 N_Y_c_643_n N_VGND_c_839_n 0.00198695f $X=3.155 $Y=0.815 $X2=0 $Y2=0
cc_469 N_Y_c_643_n N_VGND_c_840_n 0.0528344f $X=3.155 $Y=0.815 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a22o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.675000 1.695000 1.075000 ;
        RECT 1.485000 1.075000 1.815000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.040000 2.395000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.075000 1.240000 1.285000 ;
        RECT 1.020000 0.675000 1.240000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 0.255000 3.135000 0.585000 ;
        RECT 2.875000 1.785000 3.135000 2.465000 ;
        RECT 2.965000 0.585000 3.135000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.090000  0.085000 0.545000 0.850000 ;
        RECT 2.375000  0.085000 2.705000 0.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 1.430000 2.255000 1.785000 2.635000 ;
        RECT 2.455000 1.855000 2.705000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 1.455000 1.265000 1.515000 ;
      RECT 0.090000 1.515000 2.795000 1.625000 ;
      RECT 0.090000 1.625000 0.345000 2.245000 ;
      RECT 0.090000 2.245000 0.425000 2.465000 ;
      RECT 0.595000 1.795000 0.780000 1.885000 ;
      RECT 0.595000 1.885000 2.205000 2.085000 ;
      RECT 0.595000 2.085000 0.825000 2.125000 ;
      RECT 0.820000 0.255000 2.120000 0.465000 ;
      RECT 0.935000 1.625000 2.735000 1.685000 ;
      RECT 0.935000 1.685000 1.265000 1.715000 ;
      RECT 1.370000 1.875000 2.205000 1.885000 ;
      RECT 1.950000 0.465000 2.120000 0.615000 ;
      RECT 1.950000 0.615000 2.705000 0.740000 ;
      RECT 1.950000 0.740000 2.795000 0.785000 ;
      RECT 1.955000 2.085000 2.205000 2.465000 ;
      RECT 2.525000 0.785000 2.795000 0.905000 ;
      RECT 2.595000 1.480000 2.795000 1.515000 ;
      RECT 2.625000 0.905000 2.795000 1.480000 ;
  END
END sky130_fd_sc_hd__a22o_1
END LIBRARY

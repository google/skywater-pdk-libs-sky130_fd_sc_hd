* File: sky130_fd_sc_hd__dlygate4sd2_1.pxi.spice
* Created: Thu Aug 27 14:18:45 2020
* 
x_PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A N_A_M1004_g N_A_M1002_g A A N_A_c_65_n
+ N_A_c_66_n PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A
x_PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_49_47# N_A_49_47#_M1004_s
+ N_A_49_47#_M1002_s N_A_49_47#_M1003_g N_A_49_47#_M1006_g N_A_49_47#_c_97_n
+ N_A_49_47#_c_103_n N_A_49_47#_c_98_n N_A_49_47#_c_99_n N_A_49_47#_c_104_n
+ N_A_49_47#_c_105_n N_A_49_47#_c_100_n N_A_49_47#_c_106_n N_A_49_47#_c_101_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_49_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_221_47# N_A_221_47#_M1003_d
+ N_A_221_47#_M1006_d N_A_221_47#_M1001_g N_A_221_47#_M1007_g
+ N_A_221_47#_c_163_n N_A_221_47#_c_169_n N_A_221_47#_c_164_n
+ N_A_221_47#_c_165_n N_A_221_47#_c_171_n N_A_221_47#_c_166_n
+ N_A_221_47#_c_167_n PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_221_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_327_47# N_A_327_47#_M1001_s
+ N_A_327_47#_M1007_s N_A_327_47#_M1005_g N_A_327_47#_M1000_g
+ N_A_327_47#_c_223_n N_A_327_47#_c_230_n N_A_327_47#_c_224_n
+ N_A_327_47#_c_225_n N_A_327_47#_c_231_n N_A_327_47#_c_232_n
+ N_A_327_47#_c_226_n N_A_327_47#_c_233_n N_A_327_47#_c_227_n
+ N_A_327_47#_c_228_n PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%A_327_47#
x_PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%VPWR N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n VPWR
+ N_VPWR_c_295_n N_VPWR_c_290_n N_VPWR_c_297_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%VPWR
x_PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%X N_X_M1005_d N_X_M1000_d X X X X X X X X
+ PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%X
x_PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%VGND N_VGND_M1004_d N_VGND_M1001_d
+ N_VGND_c_347_n N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n VGND
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n
+ PM_SKY130_FD_SC_HD__DLYGATE4SD2_1%VGND
cc_1 VNB N_A_M1004_g 0.0352911f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.445
cc_2 VNB N_A_c_65_n 0.0108204f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_3 VNB N_A_c_66_n 0.0384693f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_4 VNB N_A_49_47#_M1003_g 0.0335659f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_5 VNB N_A_49_47#_c_97_n 0.0221254f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_6 VNB N_A_49_47#_c_98_n 0.00632336f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.53
cc_7 VNB N_A_49_47#_c_99_n 0.0110586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_49_47#_c_100_n 0.00429187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_49_47#_c_101_n 0.0232189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_221_47#_M1001_g 0.0367339f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_11 VNB N_A_221_47#_c_163_n 0.00956033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_221_47#_c_164_n 0.00778299f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.19
cc_13 VNB N_A_221_47#_c_165_n 0.00374017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_221_47#_c_166_n 0.00298146f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_221_47#_c_167_n 0.0328554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_327_47#_c_223_n 0.00461562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_327_47#_c_224_n 0.00358319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_327_47#_c_225_n 0.00346742f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.53
cc_19 VNB N_A_327_47#_c_226_n 0.00313926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_327_47#_c_227_n 0.0227093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_327_47#_c_228_n 0.0193118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_290_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB X 0.031877f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=2.275
cc_24 VNB X 0.0289946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_347_n 0.00527691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_348_n 0.00558565f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.16
cc_27 VNB N_VGND_c_349_n 0.0304046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_350_n 0.00622287f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_29 VNB N_VGND_c_351_n 0.0229408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_352_n 0.19244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_353_n 0.0237548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_M1002_g 0.0613666f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=2.275
cc_33 VPB N_A_c_65_n 0.0171572f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_34 VPB N_A_c_66_n 0.0110519f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_35 VPB N_A_49_47#_M1006_g 0.055353f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_36 VPB N_A_49_47#_c_103_n 0.022127f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.19
cc_37 VPB N_A_49_47#_c_104_n 0.00762252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_49_47#_c_105_n 0.0139826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_49_47#_c_106_n 0.00338034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_49_47#_c_101_n 0.00453682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_221_47#_M1007_g 0.0637134f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_42 VPB N_A_221_47#_c_169_n 0.0108298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_221_47#_c_164_n 0.0114409f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.19
cc_44 VPB N_A_221_47#_c_171_n 0.00374017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_221_47#_c_166_n 0.00392619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_221_47#_c_167_n 0.00940691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_327_47#_M1000_g 0.0237951f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_327_47#_c_230_n 0.0046158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_327_47#_c_231_n 0.00369316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_327_47#_c_232_n 0.0043621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_327_47#_c_233_n 0.00210224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_327_47#_c_227_n 0.00475269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_291_n 0.00527691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_292_n 0.00558565f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.16
cc_55 VPB N_VPWR_c_293_n 0.0304012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_294_n 0.00622287f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_57 VPB N_VPWR_c_295_n 0.0229408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_290_n 0.0555435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_297_n 0.0237548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB X 0.0379359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 0.0114907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB X 0.0146036f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 N_A_M1004_g N_A_49_47#_M1003_g 0.0257692f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_64 N_A_M1002_g N_A_49_47#_M1006_g 0.042978f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_65 N_A_c_65_n N_A_49_47#_M1006_g 2.80519e-19 $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_A_49_47#_c_97_n 0.00383176f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_A_49_47#_c_103_n 0.00383176f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_68 N_A_M1004_g N_A_49_47#_c_98_n 0.0146809f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_69 N_A_c_65_n N_A_49_47#_c_98_n 0.0104548f $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_c_66_n N_A_49_47#_c_98_n 4.78579e-19 $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_65_n N_A_49_47#_c_99_n 0.0353044f $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_66_n N_A_49_47#_c_99_n 0.00747954f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1002_g N_A_49_47#_c_104_n 0.0170987f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_74 N_A_c_65_n N_A_49_47#_c_104_n 0.010736f $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_c_65_n N_A_49_47#_c_105_n 0.0368472f $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_c_66_n N_A_49_47#_c_105_n 0.00125831f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_M1004_g N_A_49_47#_c_100_n 0.0056046f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_78 N_A_c_65_n N_A_49_47#_c_100_n 0.022051f $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_A_49_47#_c_106_n 0.0055615f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_80 N_A_c_65_n N_A_49_47#_c_106_n 0.0231157f $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_c_65_n N_A_49_47#_c_101_n 2.77488e-19 $X=0.32 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_c_66_n N_A_49_47#_c_101_n 0.0210576f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_VPWR_c_291_n 0.00306527f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_84 N_A_M1002_g N_VPWR_c_290_n 0.00688647f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_85 N_A_M1002_g N_VPWR_c_297_n 0.00435702f $X=0.58 $Y=2.275 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_VGND_c_347_n 0.00306527f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_VGND_c_352_n 0.00688647f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_VGND_c_353_n 0.00435702f $X=0.58 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_49_47#_M1003_g N_A_221_47#_c_163_n 0.00994812f $X=1.015 $Y=0.445 $X2=0
+ $Y2=0
cc_90 N_A_49_47#_c_100_n N_A_221_47#_c_163_n 0.0219695f $X=0.912 $Y=1.325 $X2=0
+ $Y2=0
cc_91 N_A_49_47#_c_101_n N_A_221_47#_c_163_n 5.50148e-19 $X=1 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_A_49_47#_M1006_g N_A_221_47#_c_169_n 0.0122684f $X=1.015 $Y=2.275 $X2=0
+ $Y2=0
cc_93 N_A_49_47#_c_104_n N_A_221_47#_c_169_n 0.0142222f $X=0.795 $Y=1.895 $X2=0
+ $Y2=0
cc_94 N_A_49_47#_c_106_n N_A_221_47#_c_169_n 0.0100371f $X=0.912 $Y=1.785 $X2=0
+ $Y2=0
cc_95 N_A_49_47#_M1006_g N_A_221_47#_c_166_n 0.00639748f $X=1.015 $Y=2.275 $X2=0
+ $Y2=0
cc_96 N_A_49_47#_c_100_n N_A_221_47#_c_166_n 0.0226801f $X=0.912 $Y=1.325 $X2=0
+ $Y2=0
cc_97 N_A_49_47#_c_106_n N_A_221_47#_c_166_n 0.0193564f $X=0.912 $Y=1.785 $X2=0
+ $Y2=0
cc_98 N_A_49_47#_c_101_n N_A_221_47#_c_166_n 0.00274356f $X=1 $Y=1.16 $X2=0
+ $Y2=0
cc_99 N_A_49_47#_c_100_n N_A_221_47#_c_167_n 2.10068e-19 $X=0.912 $Y=1.325 $X2=0
+ $Y2=0
cc_100 N_A_49_47#_c_101_n N_A_221_47#_c_167_n 0.0060101f $X=1 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_49_47#_M1006_g N_VPWR_c_291_n 0.00307729f $X=1.015 $Y=2.275 $X2=0
+ $Y2=0
cc_102 N_A_49_47#_c_104_n N_VPWR_c_291_n 0.0175369f $X=0.795 $Y=1.895 $X2=0
+ $Y2=0
cc_103 N_A_49_47#_M1006_g N_VPWR_c_293_n 0.00597353f $X=1.015 $Y=2.275 $X2=0
+ $Y2=0
cc_104 N_A_49_47#_c_104_n N_VPWR_c_293_n 0.00157429f $X=0.795 $Y=1.895 $X2=0
+ $Y2=0
cc_105 N_A_49_47#_M1002_s N_VPWR_c_290_n 0.00218964f $X=0.245 $Y=2.065 $X2=0
+ $Y2=0
cc_106 N_A_49_47#_M1006_g N_VPWR_c_290_n 0.0103249f $X=1.015 $Y=2.275 $X2=0
+ $Y2=0
cc_107 N_A_49_47#_c_103_n N_VPWR_c_290_n 0.0153277f $X=0.37 $Y=2.21 $X2=0 $Y2=0
cc_108 N_A_49_47#_c_104_n N_VPWR_c_290_n 0.00737666f $X=0.795 $Y=1.895 $X2=0
+ $Y2=0
cc_109 N_A_49_47#_c_103_n N_VPWR_c_297_n 0.026952f $X=0.37 $Y=2.21 $X2=0 $Y2=0
cc_110 N_A_49_47#_c_104_n N_VPWR_c_297_n 0.00238773f $X=0.795 $Y=1.895 $X2=0
+ $Y2=0
cc_111 N_A_49_47#_M1003_g N_VGND_c_347_n 0.00307729f $X=1.015 $Y=0.445 $X2=0
+ $Y2=0
cc_112 N_A_49_47#_c_98_n N_VGND_c_347_n 0.00850275f $X=0.795 $Y=0.8 $X2=0 $Y2=0
cc_113 N_A_49_47#_c_100_n N_VGND_c_347_n 0.00884165f $X=0.912 $Y=1.325 $X2=0
+ $Y2=0
cc_114 N_A_49_47#_M1003_g N_VGND_c_349_n 0.00597353f $X=1.015 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A_49_47#_c_100_n N_VGND_c_349_n 0.00157429f $X=0.912 $Y=1.325 $X2=0
+ $Y2=0
cc_116 N_A_49_47#_M1004_s N_VGND_c_352_n 0.00218964f $X=0.245 $Y=0.235 $X2=0
+ $Y2=0
cc_117 N_A_49_47#_M1003_g N_VGND_c_352_n 0.0103249f $X=1.015 $Y=0.445 $X2=0
+ $Y2=0
cc_118 N_A_49_47#_c_97_n N_VGND_c_352_n 0.015297f $X=0.37 $Y=0.51 $X2=0 $Y2=0
cc_119 N_A_49_47#_c_98_n N_VGND_c_352_n 0.0043098f $X=0.795 $Y=0.8 $X2=0 $Y2=0
cc_120 N_A_49_47#_c_100_n N_VGND_c_352_n 0.00301014f $X=0.912 $Y=1.325 $X2=0
+ $Y2=0
cc_121 N_A_49_47#_c_97_n N_VGND_c_353_n 0.0268066f $X=0.37 $Y=0.51 $X2=0 $Y2=0
cc_122 N_A_49_47#_c_98_n N_VGND_c_353_n 0.00234724f $X=0.795 $Y=0.8 $X2=0 $Y2=0
cc_123 N_A_221_47#_M1007_g N_A_327_47#_M1000_g 0.0318699f $X=1.985 $Y=2.275
+ $X2=0 $Y2=0
cc_124 N_A_221_47#_M1001_g N_A_327_47#_c_223_n 0.00379739f $X=1.985 $Y=0.445
+ $X2=0 $Y2=0
cc_125 N_A_221_47#_c_163_n N_A_327_47#_c_223_n 0.00931673f $X=1.34 $Y=1.055
+ $X2=0 $Y2=0
cc_126 N_A_221_47#_c_165_n N_A_327_47#_c_223_n 0.0245355f $X=1.34 $Y=0.42 $X2=0
+ $Y2=0
cc_127 N_A_221_47#_M1007_g N_A_327_47#_c_230_n 0.00379739f $X=1.985 $Y=2.275
+ $X2=0 $Y2=0
cc_128 N_A_221_47#_c_169_n N_A_327_47#_c_230_n 0.00931673f $X=1.34 $Y=2.135
+ $X2=0 $Y2=0
cc_129 N_A_221_47#_c_171_n N_A_327_47#_c_230_n 0.0245355f $X=1.34 $Y=2.3 $X2=0
+ $Y2=0
cc_130 N_A_221_47#_M1001_g N_A_327_47#_c_224_n 0.0167479f $X=1.985 $Y=0.445
+ $X2=0 $Y2=0
cc_131 N_A_221_47#_c_164_n N_A_327_47#_c_224_n 0.0115959f $X=1.76 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_221_47#_c_167_n N_A_327_47#_c_224_n 4.78834e-19 $X=1.985 $Y=1.16
+ $X2=0 $Y2=0
cc_133 N_A_221_47#_c_163_n N_A_327_47#_c_225_n 0.0132713f $X=1.34 $Y=1.055 $X2=0
+ $Y2=0
cc_134 N_A_221_47#_c_164_n N_A_327_47#_c_225_n 0.0226573f $X=1.76 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_221_47#_c_167_n N_A_327_47#_c_225_n 0.00623751f $X=1.985 $Y=1.16
+ $X2=0 $Y2=0
cc_136 N_A_221_47#_M1007_g N_A_327_47#_c_231_n 0.0193272f $X=1.985 $Y=2.275
+ $X2=0 $Y2=0
cc_137 N_A_221_47#_c_164_n N_A_327_47#_c_231_n 0.0118982f $X=1.76 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_221_47#_c_169_n N_A_327_47#_c_232_n 0.0171746f $X=1.34 $Y=2.135 $X2=0
+ $Y2=0
cc_139 N_A_221_47#_c_164_n N_A_327_47#_c_232_n 0.0239038f $X=1.76 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_221_47#_c_167_n N_A_327_47#_c_232_n 0.00105103f $X=1.985 $Y=1.16
+ $X2=0 $Y2=0
cc_141 N_A_221_47#_M1001_g N_A_327_47#_c_226_n 0.00576381f $X=1.985 $Y=0.445
+ $X2=0 $Y2=0
cc_142 N_A_221_47#_c_164_n N_A_327_47#_c_226_n 0.0225506f $X=1.76 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_221_47#_M1007_g N_A_327_47#_c_233_n 0.00591943f $X=1.985 $Y=2.275
+ $X2=0 $Y2=0
cc_144 N_A_221_47#_c_164_n N_A_327_47#_c_233_n 0.0231115f $X=1.76 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_221_47#_c_164_n N_A_327_47#_c_227_n 2.61797e-19 $X=1.76 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_221_47#_c_167_n N_A_327_47#_c_227_n 0.020949f $X=1.985 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A_221_47#_M1001_g N_A_327_47#_c_228_n 0.0204568f $X=1.985 $Y=0.445
+ $X2=0 $Y2=0
cc_148 N_A_221_47#_M1007_g N_VPWR_c_292_n 0.0032307f $X=1.985 $Y=2.275 $X2=0
+ $Y2=0
cc_149 N_A_221_47#_M1007_g N_VPWR_c_293_n 0.00522999f $X=1.985 $Y=2.275 $X2=0
+ $Y2=0
cc_150 N_A_221_47#_c_171_n N_VPWR_c_293_n 0.0177618f $X=1.34 $Y=2.3 $X2=0 $Y2=0
cc_151 N_A_221_47#_M1006_d N_VPWR_c_290_n 0.00379446f $X=1.105 $Y=2.065 $X2=0
+ $Y2=0
cc_152 N_A_221_47#_M1007_g N_VPWR_c_290_n 0.00821351f $X=1.985 $Y=2.275 $X2=0
+ $Y2=0
cc_153 N_A_221_47#_c_171_n N_VPWR_c_290_n 0.0102062f $X=1.34 $Y=2.3 $X2=0 $Y2=0
cc_154 N_A_221_47#_M1001_g N_VGND_c_348_n 0.0032307f $X=1.985 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_A_221_47#_M1001_g N_VGND_c_349_n 0.00522999f $X=1.985 $Y=0.445 $X2=0
+ $Y2=0
cc_156 N_A_221_47#_c_165_n N_VGND_c_349_n 0.0177618f $X=1.34 $Y=0.42 $X2=0 $Y2=0
cc_157 N_A_221_47#_M1003_d N_VGND_c_352_n 0.00379446f $X=1.105 $Y=0.235 $X2=0
+ $Y2=0
cc_158 N_A_221_47#_M1001_g N_VGND_c_352_n 0.00821351f $X=1.985 $Y=0.445 $X2=0
+ $Y2=0
cc_159 N_A_221_47#_c_165_n N_VGND_c_352_n 0.0102062f $X=1.34 $Y=0.42 $X2=0 $Y2=0
cc_160 N_A_327_47#_c_231_n N_VPWR_M1007_d 0.00504323f $X=2.2 $Y=1.895 $X2=0
+ $Y2=0
cc_161 N_A_327_47#_c_233_n N_VPWR_M1007_d 0.00463606f $X=2.3 $Y=1.785 $X2=0
+ $Y2=0
cc_162 N_A_327_47#_M1000_g N_VPWR_c_292_n 0.00321658f $X=2.475 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_327_47#_c_231_n N_VPWR_c_292_n 0.019714f $X=2.2 $Y=1.895 $X2=0 $Y2=0
cc_164 N_A_327_47#_c_230_n N_VPWR_c_293_n 0.0169146f $X=1.76 $Y=2.21 $X2=0 $Y2=0
cc_165 N_A_327_47#_c_231_n N_VPWR_c_293_n 0.00280508f $X=2.2 $Y=1.895 $X2=0
+ $Y2=0
cc_166 N_A_327_47#_M1000_g N_VPWR_c_295_n 0.00583607f $X=2.475 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_327_47#_M1007_s N_VPWR_c_290_n 0.00218964f $X=1.635 $Y=2.065 $X2=0
+ $Y2=0
cc_168 N_A_327_47#_M1000_g N_VPWR_c_290_n 0.0118143f $X=2.475 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_327_47#_c_230_n N_VPWR_c_290_n 0.00993603f $X=1.76 $Y=2.21 $X2=0
+ $Y2=0
cc_170 N_A_327_47#_c_231_n N_VPWR_c_290_n 0.00583597f $X=2.2 $Y=1.895 $X2=0
+ $Y2=0
cc_171 N_A_327_47#_M1000_g X 0.00267098f $X=2.475 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_327_47#_c_226_n X 0.0334268f $X=2.3 $Y=1.325 $X2=0 $Y2=0
cc_173 N_A_327_47#_c_233_n X 0.00703463f $X=2.3 $Y=1.785 $X2=0 $Y2=0
cc_174 N_A_327_47#_c_227_n X 0.00773291f $X=2.42 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_327_47#_c_228_n X 0.00266918f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_327_47#_c_224_n N_VGND_M1001_d 0.00237719f $X=2.2 $Y=0.8 $X2=0 $Y2=0
cc_177 N_A_327_47#_c_226_n N_VGND_M1001_d 0.00202902f $X=2.3 $Y=1.325 $X2=0
+ $Y2=0
cc_178 N_A_327_47#_c_224_n N_VGND_c_348_n 0.00725299f $X=2.2 $Y=0.8 $X2=0 $Y2=0
cc_179 N_A_327_47#_c_226_n N_VGND_c_348_n 0.0123344f $X=2.3 $Y=1.325 $X2=0 $Y2=0
cc_180 N_A_327_47#_c_227_n N_VGND_c_348_n 3.85782e-19 $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_327_47#_c_228_n N_VGND_c_348_n 0.00321658f $X=2.42 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_327_47#_c_223_n N_VGND_c_349_n 0.0168271f $X=1.76 $Y=0.51 $X2=0 $Y2=0
cc_183 N_A_327_47#_c_224_n N_VGND_c_349_n 0.00275765f $X=2.2 $Y=0.8 $X2=0 $Y2=0
cc_184 N_A_327_47#_c_228_n N_VGND_c_351_n 0.00583607f $X=2.42 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_327_47#_M1001_s N_VGND_c_352_n 0.00218964f $X=1.635 $Y=0.235 $X2=0
+ $Y2=0
cc_186 N_A_327_47#_c_223_n N_VGND_c_352_n 0.00991615f $X=1.76 $Y=0.51 $X2=0
+ $Y2=0
cc_187 N_A_327_47#_c_224_n N_VGND_c_352_n 0.00490119f $X=2.2 $Y=0.8 $X2=0 $Y2=0
cc_188 N_A_327_47#_c_226_n N_VGND_c_352_n 8.73954e-19 $X=2.3 $Y=1.325 $X2=0
+ $Y2=0
cc_189 N_A_327_47#_c_228_n N_VGND_c_352_n 0.0118143f $X=2.42 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_290_n N_X_M1000_d 0.00283025f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_295_n X 0.0387817f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_290_n X 0.0216821f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_193 X N_VGND_c_351_n 0.0387205f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_194 N_X_M1005_d N_VGND_c_352_n 0.00283025f $X=2.55 $Y=0.235 $X2=0 $Y2=0
cc_195 X N_VGND_c_352_n 0.0216638f $X=2.905 $Y=0.425 $X2=0 $Y2=0

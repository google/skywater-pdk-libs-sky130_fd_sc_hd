* File: sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.pxi.spice
* Created: Thu Aug 27 14:26:06 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A N_A_c_201_n N_A_M1032_g
+ N_A_M1000_g A N_A_c_202_n N_A_c_203_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_147_47# N_A_147_47#_M1032_d
+ N_A_147_47#_M1000_d N_A_147_47#_c_229_n N_A_147_47#_M1002_g
+ N_A_147_47#_M1005_g N_A_147_47#_c_230_n N_A_147_47#_M1009_g
+ N_A_147_47#_M1017_g N_A_147_47#_c_231_n N_A_147_47#_M1010_g
+ N_A_147_47#_M1029_g N_A_147_47#_c_232_n N_A_147_47#_M1012_g
+ N_A_147_47#_M1052_g N_A_147_47#_c_233_n N_A_147_47#_c_243_n
+ N_A_147_47#_c_234_n N_A_147_47#_c_266_p N_A_147_47#_c_235_n
+ N_A_147_47#_c_244_n N_A_147_47#_c_245_n N_A_147_47#_c_236_n
+ N_A_147_47#_c_237_n N_A_147_47#_c_238_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_147_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%SLEEP N_SLEEP_c_354_n
+ N_SLEEP_M1019_g N_SLEEP_M1006_g N_SLEEP_c_355_n N_SLEEP_M1025_g
+ N_SLEEP_M1034_g N_SLEEP_c_356_n N_SLEEP_M1026_g N_SLEEP_M1039_g
+ N_SLEEP_c_357_n N_SLEEP_M1030_g N_SLEEP_M1053_g SLEEP N_SLEEP_c_358_n
+ N_SLEEP_c_359_n PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%SLEEP
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_341_47# N_A_341_47#_M1002_s
+ N_A_341_47#_M1010_s N_A_341_47#_M1019_s N_A_341_47#_M1026_s
+ N_A_341_47#_M1005_s N_A_341_47#_M1029_s N_A_341_47#_M1003_g
+ N_A_341_47#_c_465_n N_A_341_47#_M1015_g N_A_341_47#_M1007_g
+ N_A_341_47#_c_466_n N_A_341_47#_M1037_g N_A_341_47#_M1028_g
+ N_A_341_47#_c_467_n N_A_341_47#_M1042_g N_A_341_47#_M1038_g
+ N_A_341_47#_c_468_n N_A_341_47#_M1054_g N_A_341_47#_c_475_n
+ N_A_341_47#_c_469_n N_A_341_47#_c_578_p N_A_341_47#_c_470_n
+ N_A_341_47#_c_452_n N_A_341_47#_c_453_n N_A_341_47#_c_496_n
+ N_A_341_47#_c_582_p N_A_341_47#_c_454_n N_A_341_47#_c_499_n
+ N_A_341_47#_c_455_n N_A_341_47#_c_524_n N_A_341_47#_c_472_n
+ N_A_341_47#_c_456_n N_A_341_47#_c_457_n N_A_341_47#_c_458_n
+ N_A_341_47#_c_459_n N_A_341_47#_c_460_n N_A_341_47#_c_461_n
+ N_A_341_47#_c_462_n N_A_341_47#_c_463_n N_A_341_47#_c_464_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_341_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_1122_47# N_A_1122_47#_M1003_d
+ N_A_1122_47#_M1028_d N_A_1122_47#_M1015_d N_A_1122_47#_M1042_d
+ N_A_1122_47#_M1013_g N_A_1122_47#_M1001_g N_A_1122_47#_M1014_g
+ N_A_1122_47#_M1004_g N_A_1122_47#_M1016_g N_A_1122_47#_M1008_g
+ N_A_1122_47#_M1020_g N_A_1122_47#_M1011_g N_A_1122_47#_M1023_g
+ N_A_1122_47#_M1018_g N_A_1122_47#_M1024_g N_A_1122_47#_M1021_g
+ N_A_1122_47#_M1027_g N_A_1122_47#_M1022_g N_A_1122_47#_M1041_g
+ N_A_1122_47#_M1031_g N_A_1122_47#_M1046_g N_A_1122_47#_M1033_g
+ N_A_1122_47#_M1047_g N_A_1122_47#_M1035_g N_A_1122_47#_M1049_g
+ N_A_1122_47#_M1036_g N_A_1122_47#_M1050_g N_A_1122_47#_M1040_g
+ N_A_1122_47#_M1051_g N_A_1122_47#_M1043_g N_A_1122_47#_M1055_g
+ N_A_1122_47#_M1044_g N_A_1122_47#_M1056_g N_A_1122_47#_M1045_g
+ N_A_1122_47#_c_683_n N_A_1122_47#_M1057_g N_A_1122_47#_M1048_g
+ N_A_1122_47#_c_685_n N_A_1122_47#_c_705_n N_A_1122_47#_c_719_n
+ N_A_1122_47#_c_686_n N_A_1122_47#_c_706_n N_A_1122_47#_c_687_n
+ N_A_1122_47#_c_727_n N_A_1122_47#_c_729_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_1122_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%VPWR N_VPWR_M1000_s
+ N_VPWR_M1006_s N_VPWR_M1039_s N_VPWR_c_1005_n N_VPWR_c_1006_n N_VPWR_c_1007_n
+ N_VPWR_c_1008_n VPWR N_VPWR_c_1009_n N_VPWR_c_1010_n N_VPWR_c_1011_n
+ N_VPWR_c_1004_n N_VPWR_c_1013_n N_VPWR_c_1014_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_255_297# N_A_255_297#_M1005_d
+ N_A_255_297#_M1017_d N_A_255_297#_M1052_d N_A_255_297#_M1034_d
+ N_A_255_297#_M1053_d N_A_255_297#_c_1202_n N_A_255_297#_c_1203_n
+ N_A_255_297#_c_1217_n N_A_255_297#_c_1219_n N_A_255_297#_c_1223_n
+ N_A_255_297#_c_1204_n N_A_255_297#_c_1226_n N_A_255_297#_c_1205_n
+ N_A_255_297#_c_1276_n N_A_255_297#_c_1206_n N_A_255_297#_c_1207_n
+ N_A_255_297#_c_1208_n N_A_255_297#_c_1228_n N_A_255_297#_c_1209_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%A_255_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%KAPWR N_KAPWR_M1015_s
+ N_KAPWR_M1037_s N_KAPWR_M1054_s N_KAPWR_M1004_d N_KAPWR_M1011_d
+ N_KAPWR_M1021_d N_KAPWR_M1031_d N_KAPWR_M1035_d N_KAPWR_M1040_d
+ N_KAPWR_M1044_d N_KAPWR_M1048_d N_KAPWR_c_1304_n N_KAPWR_c_1305_n
+ N_KAPWR_c_1338_n N_KAPWR_c_1324_n N_KAPWR_c_1341_n N_KAPWR_c_1326_n
+ N_KAPWR_c_1345_n N_KAPWR_c_1346_n N_KAPWR_c_1348_n N_KAPWR_c_1350_n
+ N_KAPWR_c_1351_n N_KAPWR_c_1353_n N_KAPWR_c_1355_n N_KAPWR_c_1356_n
+ N_KAPWR_c_1358_n N_KAPWR_c_1360_n N_KAPWR_c_1361_n N_KAPWR_c_1363_n
+ N_KAPWR_c_1365_n N_KAPWR_c_1367_n N_KAPWR_c_1369_n N_KAPWR_c_1371_n
+ N_KAPWR_c_1372_n N_KAPWR_c_1374_n N_KAPWR_c_1376_n N_KAPWR_c_1378_n
+ N_KAPWR_c_1381_n N_KAPWR_c_1383_n N_KAPWR_c_1306_n KAPWR N_KAPWR_c_1307_n
+ N_KAPWR_c_1332_n N_KAPWR_c_1335_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%X N_X_M1013_d N_X_M1016_d
+ N_X_M1023_d N_X_M1027_d N_X_M1046_d N_X_M1049_d N_X_M1051_d N_X_M1056_d
+ N_X_M1001_s N_X_M1008_s N_X_M1018_s N_X_M1022_s N_X_M1033_s N_X_M1036_s
+ N_X_M1043_s N_X_M1045_s N_X_c_1543_n N_X_c_1544_n N_X_c_1545_n N_X_c_1579_n
+ N_X_c_1546_n N_X_c_1547_n N_X_c_1589_n N_X_c_1548_n N_X_c_1549_n N_X_c_1599_n
+ N_X_c_1550_n N_X_c_1551_n N_X_c_1610_n N_X_c_1552_n N_X_c_1553_n N_X_c_1620_n
+ N_X_c_1554_n N_X_c_1555_n N_X_c_1630_n N_X_c_1556_n N_X_c_1557_n N_X_c_1558_n
+ N_X_c_1640_n N_X_c_1559_n N_X_c_1646_n N_X_c_1560_n N_X_c_1652_n N_X_c_1561_n
+ N_X_c_1659_n N_X_c_1562_n N_X_c_1666_n N_X_c_1563_n N_X_c_1672_n N_X_c_1564_n
+ X X X X N_X_c_1567_n PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%X
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%VGND N_VGND_M1032_s
+ N_VGND_M1002_d N_VGND_M1009_d N_VGND_M1012_d N_VGND_M1025_d N_VGND_M1030_d
+ N_VGND_M1003_s N_VGND_M1007_s N_VGND_M1038_s N_VGND_M1014_s N_VGND_M1020_s
+ N_VGND_M1024_s N_VGND_M1041_s N_VGND_M1047_s N_VGND_M1050_s N_VGND_M1055_s
+ N_VGND_M1057_s N_VGND_c_1843_n N_VGND_c_1844_n N_VGND_c_1845_n N_VGND_c_1846_n
+ N_VGND_c_1847_n N_VGND_c_1848_n N_VGND_c_1849_n N_VGND_c_1850_n
+ N_VGND_c_1851_n N_VGND_c_1852_n N_VGND_c_1853_n N_VGND_c_1854_n
+ N_VGND_c_1855_n N_VGND_c_1856_n N_VGND_c_1857_n N_VGND_c_1858_n
+ N_VGND_c_1859_n N_VGND_c_1860_n N_VGND_c_1861_n N_VGND_c_1862_n
+ N_VGND_c_1863_n N_VGND_c_1864_n N_VGND_c_1865_n N_VGND_c_1866_n
+ N_VGND_c_1867_n N_VGND_c_1868_n N_VGND_c_1869_n N_VGND_c_1870_n
+ N_VGND_c_1871_n N_VGND_c_1872_n N_VGND_c_1873_n N_VGND_c_1874_n
+ N_VGND_c_1875_n N_VGND_c_1876_n N_VGND_c_1877_n N_VGND_c_1878_n VGND
+ N_VGND_c_1879_n N_VGND_c_1880_n N_VGND_c_1881_n N_VGND_c_1882_n
+ N_VGND_c_1883_n N_VGND_c_1884_n N_VGND_c_1885_n N_VGND_c_1886_n
+ N_VGND_c_1887_n N_VGND_c_1888_n N_VGND_c_1889_n N_VGND_c_1890_n VGND
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRCKAPWR_16%VGND
cc_1 VNB N_A_c_201_n 0.0246248f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.995
cc_2 VNB N_A_c_202_n 0.0153622f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_3 VNB N_A_c_203_n 0.0391805f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_4 VNB N_A_147_47#_c_229_n 0.0197222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_147_47#_c_230_n 0.0157557f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_6 VNB N_A_147_47#_c_231_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_147_47#_c_232_n 0.0153897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_147_47#_c_233_n 0.00335056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_147_47#_c_234_n 0.00362507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_147_47#_c_235_n 0.00134522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_147_47#_c_236_n 0.00117446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_147_47#_c_237_n 0.0442418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_147_47#_c_238_n 0.0592139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_SLEEP_c_354_n 0.0158209f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.995
cc_15 VNB N_SLEEP_c_355_n 0.0156566f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.105
cc_16 VNB N_SLEEP_c_356_n 0.0156747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_SLEEP_c_357_n 0.019609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_SLEEP_c_358_n 0.00316339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_SLEEP_c_359_n 0.0659805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_341_47#_M1003_g 0.027081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_341_47#_M1007_g 0.0229781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_341_47#_M1028_g 0.0229774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_341_47#_M1038_g 0.0234436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_341_47#_c_452_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_341_47#_c_453_n 2.95213e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_341_47#_c_454_n 0.00115298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_341_47#_c_455_n 0.00184455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_341_47#_c_456_n 9.22322e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_341_47#_c_457_n 0.00225983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_341_47#_c_458_n 0.0170632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_341_47#_c_459_n 0.00194781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_341_47#_c_460_n 0.00148995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_341_47#_c_461_n 0.0077932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_341_47#_c_462_n 0.106338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_341_47#_c_463_n 0.00262172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_341_47#_c_464_n 0.00242518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_1122_47#_M1013_g 0.0260664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_1122_47#_M1014_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_1122_47#_M1016_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_1122_47#_M1020_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_1122_47#_M1023_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_1122_47#_M1024_g 0.0241428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_1122_47#_M1027_g 0.0238169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_1122_47#_M1041_g 0.0240545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_1122_47#_M1046_g 0.0240466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1122_47#_M1047_g 0.0241431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_1122_47#_M1049_g 0.0241355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1122_47#_M1050_g 0.0241431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1122_47#_M1051_g 0.0241328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1122_47#_M1055_g 0.0241116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1122_47#_M1056_g 0.0237673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1122_47#_c_683_n 0.300055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1122_47#_M1057_g 0.0320587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1122_47#_c_685_n 0.00409026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1122_47#_c_686_n 0.00481736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1122_47#_c_687_n 0.00429043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_1004_n 0.592346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_X_c_1543_n 0.00160391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_X_c_1544_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_X_c_1545_n 0.00419804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_X_c_1546_n 0.00126237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_X_c_1547_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_X_c_1548_n 0.00125415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_X_c_1549_n 0.00501892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_X_c_1550_n 6.22964e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_X_c_1551_n 0.00491776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_X_c_1552_n 0.00125437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_X_c_1553_n 0.00522562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_X_c_1554_n 0.00126258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_X_c_1555_n 0.00522562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_X_c_1556_n 0.00126798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_X_c_1557_n 4.84646e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_X_c_1558_n 0.00137779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_X_c_1559_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_X_c_1560_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_X_c_1561_n 0.00217463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_X_c_1562_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_X_c_1563_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_X_c_1564_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB X 0.0318745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1843_n 0.0155909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1844_n 0.0335702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1845_n 0.0136791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1846_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1847_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1848_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1849_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1850_n 0.00400874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1851_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1852_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1853_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1854_n 0.00390627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1855_n 0.0157899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1856_n 0.00395785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1857_n 0.0157442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1858_n 0.00397944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1859_n 0.00397944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1860_n 0.00402207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1861_n 0.0135264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1862_n 0.0178379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1863_n 0.0183638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1864_n 0.00557475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1865_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1866_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1867_n 0.0166866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1868_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1869_n 0.0167416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1870_n 0.00500104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1871_n 0.0160902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1872_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1873_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1874_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1875_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1876_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1877_n 0.0157075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1878_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1879_n 0.0169303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1880_n 0.0157442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1881_n 0.0154599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1882_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1883_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1884_n 0.0062357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1885_n 0.0273319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1886_n 0.00497572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1887_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1888_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1889_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1890_n 0.654125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VPB N_A_M1000_g 0.0293544f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.985
cc_130 VPB N_A_c_202_n 0.00365122f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_131 VPB N_A_c_203_n 0.0106215f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_132 VPB N_A_147_47#_M1005_g 0.023038f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_133 VPB N_A_147_47#_M1017_g 0.0181069f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.197
cc_134 VPB N_A_147_47#_M1029_g 0.0176224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_147_47#_M1052_g 0.0185987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_147_47#_c_243_n 0.00550526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_147_47#_c_244_n 0.0013846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_147_47#_c_245_n 0.00513483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_147_47#_c_237_n 0.021667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_147_47#_c_238_n 0.010199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_SLEEP_M1006_g 0.0184925f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.985
cc_142 VPB N_SLEEP_M1034_g 0.0179946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_SLEEP_M1039_g 0.0179946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_SLEEP_M1053_g 0.0233603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_SLEEP_c_359_n 0.0103371f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_341_47#_c_465_n 0.0186661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_341_47#_c_466_n 0.0143984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_341_47#_c_467_n 0.0143984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_341_47#_c_468_n 0.0145807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_341_47#_c_469_n 0.00172897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_341_47#_c_470_n 0.00309212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_341_47#_c_453_n 0.00117101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_341_47#_c_472_n 2.78665e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_341_47#_c_461_n 7.61211e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_341_47#_c_462_n 0.0394256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_1122_47#_M1001_g 0.0190636f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.197
cc_157 VPB N_A_1122_47#_M1004_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_1122_47#_M1008_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_1122_47#_M1011_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_1122_47#_M1018_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_1122_47#_M1021_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_1122_47#_M1022_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_1122_47#_M1031_g 0.0186881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_1122_47#_M1033_g 0.0186881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_1122_47#_M1035_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_1122_47#_M1036_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_1122_47#_M1040_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1122_47#_M1043_g 0.0187387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_1122_47#_M1044_g 0.0186963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1122_47#_M1045_g 0.0173762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_1122_47#_c_683_n 0.0522358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1122_47#_M1048_g 0.0224494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_1122_47#_c_705_n 0.00131518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_1122_47#_c_706_n 0.00131518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1122_47#_c_687_n 0.00258437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1005_n 0.0141086f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_177 VPB N_VPWR_c_1006_n 0.0465776f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_178 VPB N_VPWR_c_1007_n 0.00221708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1008_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1009_n 0.0689736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1010_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1011_n 0.256574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1004_n 0.0490656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1013_n 0.00353635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1014_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_255_297#_c_1202_n 0.00200524f $X=-0.19 $Y=1.305 $X2=0.335
+ $Y2=1.197
cc_187 VPB N_A_255_297#_c_1203_n 0.00694208f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_255_297#_c_1204_n 0.00367521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_255_297#_c_1205_n 0.00252639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_255_297#_c_1206_n 0.00295806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_255_297#_c_1207_n 0.0062088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_255_297#_c_1208_n 0.00682151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_255_297#_c_1209_n 0.00123615f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_KAPWR_c_1304_n 0.0124499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_KAPWR_c_1305_n 0.0249622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_KAPWR_c_1306_n 0.0178729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_KAPWR_c_1307_n 0.00833561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB X 0.0102708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_X_c_1567_n 0.00990633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 N_A_c_201_n N_A_147_47#_c_233_n 0.00457189f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_M1000_g N_A_147_47#_c_243_n 0.00743921f $X=0.66 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_c_201_n N_A_147_47#_c_234_n 0.00617045f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_201_n N_A_147_47#_c_235_n 0.00323581f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_M1000_g N_A_147_47#_c_244_n 0.0032678f $X=0.66 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_c_202_n N_A_147_47#_c_245_n 0.00350706f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_c_203_n N_A_147_47#_c_245_n 0.00696913f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_c_202_n N_A_147_47#_c_236_n 0.0174258f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_c_203_n N_A_147_47#_c_236_n 0.00164603f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_c_203_n N_A_147_47#_c_237_n 0.0209283f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_M1000_g N_VPWR_c_1006_n 0.00490564f $X=0.66 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_c_202_n N_VPWR_c_1006_n 0.0325355f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_c_203_n N_VPWR_c_1006_n 0.00580252f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_M1000_g N_VPWR_c_1009_n 0.00541359f $X=0.66 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_M1000_g N_VPWR_c_1004_n 0.00734932f $X=0.66 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_M1000_g N_KAPWR_c_1305_n 0.00580645f $X=0.66 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_c_201_n N_VGND_c_1844_n 0.00500932f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_c_202_n N_VGND_c_1844_n 0.0239559f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_c_203_n N_VGND_c_1844_n 0.0063933f $X=0.66 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_c_201_n N_VGND_c_1845_n 0.0023653f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_201_n N_VGND_c_1863_n 0.00541359f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_c_201_n N_VGND_c_1890_n 0.0119208f $X=0.66 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_147_47#_c_232_n N_SLEEP_c_354_n 0.0194114f $X=2.89 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_223 N_A_147_47#_M1052_g N_SLEEP_M1006_g 0.0194114f $X=2.89 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_147_47#_c_238_n N_SLEEP_c_358_n 9.19453e-19 $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_225 N_A_147_47#_c_238_n N_SLEEP_c_359_n 0.0194114f $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_226 N_A_147_47#_c_229_n N_A_341_47#_c_475_n 0.00539651f $X=1.63 $Y=0.995
+ $X2=0 $Y2=0
cc_227 N_A_147_47#_c_230_n N_A_341_47#_c_475_n 0.00630972f $X=2.05 $Y=0.995
+ $X2=0 $Y2=0
cc_228 N_A_147_47#_c_231_n N_A_341_47#_c_475_n 5.22228e-19 $X=2.47 $Y=0.995
+ $X2=0 $Y2=0
cc_229 N_A_147_47#_M1005_g N_A_341_47#_c_469_n 0.0012406f $X=1.63 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A_147_47#_c_266_p N_A_341_47#_c_469_n 0.0138639f $X=2.1 $Y=1.16 $X2=0
+ $Y2=0
cc_231 N_A_147_47#_c_238_n N_A_341_47#_c_469_n 0.00222344f $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_232 N_A_147_47#_M1017_g N_A_341_47#_c_470_n 0.0134629f $X=2.05 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_147_47#_M1029_g N_A_341_47#_c_470_n 0.0060983f $X=2.47 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_147_47#_c_266_p N_A_341_47#_c_470_n 0.0251164f $X=2.1 $Y=1.16 $X2=0
+ $Y2=0
cc_235 N_A_147_47#_c_238_n N_A_341_47#_c_470_n 0.00236161f $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_236 N_A_147_47#_c_229_n N_A_341_47#_c_452_n 0.00262807f $X=1.63 $Y=0.995
+ $X2=0 $Y2=0
cc_237 N_A_147_47#_c_230_n N_A_341_47#_c_452_n 0.00113286f $X=2.05 $Y=0.995
+ $X2=0 $Y2=0
cc_238 N_A_147_47#_c_266_p N_A_341_47#_c_452_n 0.0265405f $X=2.1 $Y=1.16 $X2=0
+ $Y2=0
cc_239 N_A_147_47#_c_238_n N_A_341_47#_c_452_n 0.00230339f $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_240 N_A_147_47#_M1017_g N_A_341_47#_c_453_n 6.86349e-19 $X=2.05 $Y=1.985
+ $X2=0 $Y2=0
cc_241 N_A_147_47#_c_231_n N_A_341_47#_c_453_n 0.0010587f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_147_47#_M1029_g N_A_341_47#_c_453_n 0.0039358f $X=2.47 $Y=1.985 $X2=0
+ $Y2=0
cc_243 N_A_147_47#_c_232_n N_A_341_47#_c_453_n 8.10153e-19 $X=2.89 $Y=0.995
+ $X2=0 $Y2=0
cc_244 N_A_147_47#_M1052_g N_A_341_47#_c_453_n 0.00322994f $X=2.89 $Y=1.985
+ $X2=0 $Y2=0
cc_245 N_A_147_47#_c_266_p N_A_341_47#_c_453_n 0.0158053f $X=2.1 $Y=1.16 $X2=0
+ $Y2=0
cc_246 N_A_147_47#_c_238_n N_A_341_47#_c_453_n 0.0283654f $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_247 N_A_147_47#_c_230_n N_A_341_47#_c_496_n 5.23018e-19 $X=2.05 $Y=0.995
+ $X2=0 $Y2=0
cc_248 N_A_147_47#_c_231_n N_A_341_47#_c_496_n 0.00641298f $X=2.47 $Y=0.995
+ $X2=0 $Y2=0
cc_249 N_A_147_47#_c_232_n N_A_341_47#_c_496_n 0.00641298f $X=2.89 $Y=0.995
+ $X2=0 $Y2=0
cc_250 N_A_147_47#_c_232_n N_A_341_47#_c_499_n 5.22228e-19 $X=2.89 $Y=0.995
+ $X2=0 $Y2=0
cc_251 N_A_147_47#_M1029_g N_A_341_47#_c_472_n 0.00629197f $X=2.47 $Y=1.985
+ $X2=0 $Y2=0
cc_252 N_A_147_47#_M1052_g N_A_341_47#_c_472_n 5.53367e-19 $X=2.89 $Y=1.985
+ $X2=0 $Y2=0
cc_253 N_A_147_47#_c_232_n N_A_341_47#_c_457_n 0.00557491f $X=2.89 $Y=0.995
+ $X2=0 $Y2=0
cc_254 N_A_147_47#_c_230_n N_A_341_47#_c_463_n 0.00870364f $X=2.05 $Y=0.995
+ $X2=0 $Y2=0
cc_255 N_A_147_47#_c_231_n N_A_341_47#_c_463_n 0.00468086f $X=2.47 $Y=0.995
+ $X2=0 $Y2=0
cc_256 N_A_147_47#_c_266_p N_A_341_47#_c_463_n 0.018419f $X=2.1 $Y=1.16 $X2=0
+ $Y2=0
cc_257 N_A_147_47#_c_238_n N_A_341_47#_c_463_n 0.00240055f $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_258 N_A_147_47#_c_230_n N_A_341_47#_c_464_n 3.39248e-19 $X=2.05 $Y=0.995
+ $X2=0 $Y2=0
cc_259 N_A_147_47#_c_231_n N_A_341_47#_c_464_n 0.00656662f $X=2.47 $Y=0.995
+ $X2=0 $Y2=0
cc_260 N_A_147_47#_c_232_n N_A_341_47#_c_464_n 0.0133025f $X=2.89 $Y=0.995 $X2=0
+ $Y2=0
cc_261 N_A_147_47#_c_238_n N_A_341_47#_c_464_n 0.00104495f $X=2.89 $Y=1.16 $X2=0
+ $Y2=0
cc_262 N_A_147_47#_c_244_n N_VPWR_c_1006_n 0.0360029f $X=0.87 $Y=1.66 $X2=0
+ $Y2=0
cc_263 N_A_147_47#_M1005_g N_VPWR_c_1009_n 0.00357835f $X=1.63 $Y=1.985 $X2=0
+ $Y2=0
cc_264 N_A_147_47#_M1017_g N_VPWR_c_1009_n 0.00357835f $X=2.05 $Y=1.985 $X2=0
+ $Y2=0
cc_265 N_A_147_47#_M1029_g N_VPWR_c_1009_n 0.00357835f $X=2.47 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_A_147_47#_M1052_g N_VPWR_c_1009_n 0.00357835f $X=2.89 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_A_147_47#_c_243_n N_VPWR_c_1009_n 0.0210244f $X=0.87 $Y=2.34 $X2=0
+ $Y2=0
cc_268 N_A_147_47#_M1000_d N_VPWR_c_1004_n 0.00111289f $X=0.735 $Y=1.485 $X2=0
+ $Y2=0
cc_269 N_A_147_47#_M1005_g N_VPWR_c_1004_n 0.00595613f $X=1.63 $Y=1.985 $X2=0
+ $Y2=0
cc_270 N_A_147_47#_M1017_g N_VPWR_c_1004_n 0.00463006f $X=2.05 $Y=1.985 $X2=0
+ $Y2=0
cc_271 N_A_147_47#_M1029_g N_VPWR_c_1004_n 0.00463006f $X=2.47 $Y=1.985 $X2=0
+ $Y2=0
cc_272 N_A_147_47#_M1052_g N_VPWR_c_1004_n 0.00465727f $X=2.89 $Y=1.985 $X2=0
+ $Y2=0
cc_273 N_A_147_47#_c_243_n N_VPWR_c_1004_n 0.00298519f $X=0.87 $Y=2.34 $X2=0
+ $Y2=0
cc_274 N_A_147_47#_M1005_g N_A_255_297#_c_1202_n 7.12665e-19 $X=1.63 $Y=1.985
+ $X2=0 $Y2=0
cc_275 N_A_147_47#_c_243_n N_A_255_297#_c_1202_n 0.0143557f $X=0.87 $Y=2.34
+ $X2=0 $Y2=0
cc_276 N_A_147_47#_M1005_g N_A_255_297#_c_1203_n 0.00854464f $X=1.63 $Y=1.985
+ $X2=0 $Y2=0
cc_277 N_A_147_47#_M1017_g N_A_255_297#_c_1203_n 6.11469e-19 $X=2.05 $Y=1.985
+ $X2=0 $Y2=0
cc_278 N_A_147_47#_c_266_p N_A_255_297#_c_1203_n 0.0178299f $X=2.1 $Y=1.16 $X2=0
+ $Y2=0
cc_279 N_A_147_47#_c_244_n N_A_255_297#_c_1203_n 0.0586658f $X=0.87 $Y=1.66
+ $X2=0 $Y2=0
cc_280 N_A_147_47#_c_237_n N_A_255_297#_c_1203_n 0.00774573f $X=1.555 $Y=1.16
+ $X2=0 $Y2=0
cc_281 N_A_147_47#_M1005_g N_A_255_297#_c_1217_n 0.00771334f $X=1.63 $Y=1.985
+ $X2=0 $Y2=0
cc_282 N_A_147_47#_M1017_g N_A_255_297#_c_1217_n 0.00705703f $X=2.05 $Y=1.985
+ $X2=0 $Y2=0
cc_283 N_A_147_47#_M1005_g N_A_255_297#_c_1219_n 5.5199e-19 $X=1.63 $Y=1.985
+ $X2=0 $Y2=0
cc_284 N_A_147_47#_M1017_g N_A_255_297#_c_1219_n 0.00467397f $X=2.05 $Y=1.985
+ $X2=0 $Y2=0
cc_285 N_A_147_47#_M1029_g N_A_255_297#_c_1219_n 0.00467397f $X=2.47 $Y=1.985
+ $X2=0 $Y2=0
cc_286 N_A_147_47#_M1052_g N_A_255_297#_c_1219_n 5.5199e-19 $X=2.89 $Y=1.985
+ $X2=0 $Y2=0
cc_287 N_A_147_47#_M1029_g N_A_255_297#_c_1223_n 0.00703675f $X=2.47 $Y=1.985
+ $X2=0 $Y2=0
cc_288 N_A_147_47#_M1052_g N_A_255_297#_c_1223_n 0.00771334f $X=2.89 $Y=1.985
+ $X2=0 $Y2=0
cc_289 N_A_147_47#_M1052_g N_A_255_297#_c_1204_n 0.00328958f $X=2.89 $Y=1.985
+ $X2=0 $Y2=0
cc_290 N_A_147_47#_M1029_g N_A_255_297#_c_1226_n 6.07989e-19 $X=2.47 $Y=1.985
+ $X2=0 $Y2=0
cc_291 N_A_147_47#_M1052_g N_A_255_297#_c_1226_n 0.00775699f $X=2.89 $Y=1.985
+ $X2=0 $Y2=0
cc_292 N_A_147_47#_M1017_g N_A_255_297#_c_1228_n 7.04098e-19 $X=2.05 $Y=1.985
+ $X2=0 $Y2=0
cc_293 N_A_147_47#_M1029_g N_A_255_297#_c_1228_n 7.04098e-19 $X=2.47 $Y=1.985
+ $X2=0 $Y2=0
cc_294 N_A_147_47#_M1005_g N_KAPWR_c_1305_n 0.00597073f $X=1.63 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_A_147_47#_M1017_g N_KAPWR_c_1305_n 0.00233083f $X=2.05 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_147_47#_M1029_g N_KAPWR_c_1305_n 0.00232921f $X=2.47 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_A_147_47#_M1052_g N_KAPWR_c_1305_n 0.00597073f $X=2.89 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_147_47#_c_243_n N_KAPWR_c_1305_n 0.0318893f $X=0.87 $Y=2.34 $X2=0
+ $Y2=0
cc_299 N_A_147_47#_c_234_n N_VGND_c_1844_n 0.00117072f $X=0.91 $Y=1.075 $X2=0
+ $Y2=0
cc_300 N_A_147_47#_c_229_n N_VGND_c_1845_n 0.00367742f $X=1.63 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_A_147_47#_c_233_n N_VGND_c_1845_n 0.0512575f $X=0.87 $Y=0.39 $X2=0
+ $Y2=0
cc_302 N_A_147_47#_c_266_p N_VGND_c_1845_n 0.0234825f $X=2.1 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_147_47#_c_237_n N_VGND_c_1845_n 0.00739466f $X=1.555 $Y=1.16 $X2=0
+ $Y2=0
cc_304 N_A_147_47#_c_230_n N_VGND_c_1846_n 0.00146448f $X=2.05 $Y=0.995 $X2=0
+ $Y2=0
cc_305 N_A_147_47#_c_231_n N_VGND_c_1846_n 0.00146448f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_A_147_47#_c_232_n N_VGND_c_1847_n 0.00146448f $X=2.89 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_147_47#_c_233_n N_VGND_c_1863_n 0.020984f $X=0.87 $Y=0.39 $X2=0 $Y2=0
cc_308 N_A_147_47#_c_229_n N_VGND_c_1865_n 0.00541359f $X=1.63 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_147_47#_c_230_n N_VGND_c_1865_n 0.00423334f $X=2.05 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_A_147_47#_c_231_n N_VGND_c_1867_n 0.0042235f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_A_147_47#_c_232_n N_VGND_c_1867_n 0.0042235f $X=2.89 $Y=0.995 $X2=0
+ $Y2=0
cc_312 N_A_147_47#_M1032_d N_VGND_c_1890_n 0.00225715f $X=0.735 $Y=0.235 $X2=0
+ $Y2=0
cc_313 N_A_147_47#_c_229_n N_VGND_c_1890_n 0.0108276f $X=1.63 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_147_47#_c_230_n N_VGND_c_1890_n 0.0057163f $X=2.05 $Y=0.995 $X2=0
+ $Y2=0
cc_315 N_A_147_47#_c_231_n N_VGND_c_1890_n 0.00555955f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_147_47#_c_232_n N_VGND_c_1890_n 0.00538043f $X=2.89 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_147_47#_c_233_n N_VGND_c_1890_n 0.0124119f $X=0.87 $Y=0.39 $X2=0
+ $Y2=0
cc_318 N_SLEEP_c_358_n N_A_341_47#_c_453_n 0.00659349f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_319 N_SLEEP_c_359_n N_A_341_47#_c_453_n 0.00132221f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_320 N_SLEEP_c_354_n N_A_341_47#_c_496_n 5.23018e-19 $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_SLEEP_c_354_n N_A_341_47#_c_454_n 0.0081969f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_322 N_SLEEP_c_358_n N_A_341_47#_c_454_n 0.00570969f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_SLEEP_c_354_n N_A_341_47#_c_499_n 0.00630972f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_SLEEP_c_355_n N_A_341_47#_c_499_n 0.00630972f $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_SLEEP_c_356_n N_A_341_47#_c_499_n 5.22228e-19 $X=4.15 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_SLEEP_c_355_n N_A_341_47#_c_455_n 0.00796971f $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_SLEEP_c_356_n N_A_341_47#_c_455_n 0.00889955f $X=4.15 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_SLEEP_c_357_n N_A_341_47#_c_455_n 0.00194987f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_329 N_SLEEP_c_358_n N_A_341_47#_c_455_n 0.052811f $X=4.46 $Y=1.16 $X2=0 $Y2=0
cc_330 N_SLEEP_c_359_n N_A_341_47#_c_455_n 0.0043956f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_331 N_SLEEP_c_355_n N_A_341_47#_c_524_n 5.22228e-19 $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_SLEEP_c_356_n N_A_341_47#_c_524_n 0.00630972f $X=4.15 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_SLEEP_c_357_n N_A_341_47#_c_524_n 0.00538019f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_SLEEP_c_354_n N_A_341_47#_c_456_n 9.29836e-19 $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_SLEEP_c_355_n N_A_341_47#_c_456_n 9.29836e-19 $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_SLEEP_c_358_n N_A_341_47#_c_456_n 0.0212739f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_SLEEP_c_359_n N_A_341_47#_c_456_n 0.00221535f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_SLEEP_c_354_n N_A_341_47#_c_458_n 0.0016261f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_339 N_SLEEP_c_355_n N_A_341_47#_c_458_n 0.00150439f $X=3.73 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_SLEEP_c_356_n N_A_341_47#_c_458_n 0.00150439f $X=4.15 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_SLEEP_c_357_n N_A_341_47#_c_458_n 0.0038155f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_342 N_SLEEP_c_358_n N_A_341_47#_c_458_n 0.0374917f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_343 N_SLEEP_c_359_n N_A_341_47#_c_458_n 0.00689377f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_344 N_SLEEP_c_354_n N_A_341_47#_c_459_n 8.79776e-19 $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_SLEEP_c_357_n N_A_341_47#_c_461_n 0.00312483f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_SLEEP_c_358_n N_A_341_47#_c_461_n 0.00894958f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_347 N_SLEEP_c_359_n N_A_341_47#_c_461_n 0.00172293f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_348 N_SLEEP_c_357_n N_A_341_47#_c_462_n 0.0108179f $X=4.57 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_SLEEP_c_358_n N_A_341_47#_c_462_n 9.66026e-19 $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_350 N_SLEEP_c_354_n N_A_341_47#_c_464_n 0.00119908f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_SLEEP_M1006_g N_VPWR_c_1007_n 0.00304729f $X=3.31 $Y=1.985 $X2=0 $Y2=0
cc_352 N_SLEEP_M1034_g N_VPWR_c_1007_n 0.010012f $X=3.73 $Y=1.985 $X2=0 $Y2=0
cc_353 N_SLEEP_M1039_g N_VPWR_c_1007_n 7.00555e-19 $X=4.15 $Y=1.985 $X2=0 $Y2=0
cc_354 N_SLEEP_M1034_g N_VPWR_c_1008_n 7.09046e-19 $X=3.73 $Y=1.985 $X2=0 $Y2=0
cc_355 N_SLEEP_M1039_g N_VPWR_c_1008_n 0.0103803f $X=4.15 $Y=1.985 $X2=0 $Y2=0
cc_356 N_SLEEP_M1053_g N_VPWR_c_1008_n 0.0122081f $X=4.57 $Y=1.985 $X2=0 $Y2=0
cc_357 N_SLEEP_M1006_g N_VPWR_c_1009_n 0.00539841f $X=3.31 $Y=1.985 $X2=0 $Y2=0
cc_358 N_SLEEP_M1034_g N_VPWR_c_1010_n 0.0046653f $X=3.73 $Y=1.985 $X2=0 $Y2=0
cc_359 N_SLEEP_M1039_g N_VPWR_c_1010_n 0.0046653f $X=4.15 $Y=1.985 $X2=0 $Y2=0
cc_360 N_SLEEP_M1053_g N_VPWR_c_1011_n 0.0046653f $X=4.57 $Y=1.985 $X2=0 $Y2=0
cc_361 N_SLEEP_M1006_g N_VPWR_c_1004_n 0.00495344f $X=3.31 $Y=1.985 $X2=0 $Y2=0
cc_362 N_SLEEP_M1034_g N_VPWR_c_1004_n 0.00343211f $X=3.73 $Y=1.985 $X2=0 $Y2=0
cc_363 N_SLEEP_M1039_g N_VPWR_c_1004_n 0.00343211f $X=4.15 $Y=1.985 $X2=0 $Y2=0
cc_364 N_SLEEP_M1053_g N_VPWR_c_1004_n 0.00475818f $X=4.57 $Y=1.985 $X2=0 $Y2=0
cc_365 N_SLEEP_M1006_g N_A_255_297#_c_1204_n 0.00165735f $X=3.31 $Y=1.985 $X2=0
+ $Y2=0
cc_366 N_SLEEP_c_358_n N_A_255_297#_c_1204_n 3.53399e-19 $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_367 N_SLEEP_M1006_g N_A_255_297#_c_1226_n 0.00932833f $X=3.31 $Y=1.985 $X2=0
+ $Y2=0
cc_368 N_SLEEP_M1034_g N_A_255_297#_c_1226_n 4.50937e-19 $X=3.73 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_SLEEP_M1006_g N_A_255_297#_c_1205_n 0.00905509f $X=3.31 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_SLEEP_M1034_g N_A_255_297#_c_1205_n 0.0108273f $X=3.73 $Y=1.985 $X2=0
+ $Y2=0
cc_371 N_SLEEP_c_358_n N_A_255_297#_c_1205_n 0.0389728f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_372 N_SLEEP_c_359_n N_A_255_297#_c_1205_n 0.00213789f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_373 N_SLEEP_M1039_g N_A_255_297#_c_1206_n 0.0108273f $X=4.15 $Y=1.985 $X2=0
+ $Y2=0
cc_374 N_SLEEP_M1053_g N_A_255_297#_c_1206_n 0.0110794f $X=4.57 $Y=1.985 $X2=0
+ $Y2=0
cc_375 N_SLEEP_c_358_n N_A_255_297#_c_1206_n 0.0444806f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_376 N_SLEEP_c_359_n N_A_255_297#_c_1206_n 0.00213789f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_377 N_SLEEP_c_358_n N_A_255_297#_c_1207_n 3.93996e-19 $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_378 N_SLEEP_c_358_n N_A_255_297#_c_1209_n 0.012735f $X=4.46 $Y=1.16 $X2=0
+ $Y2=0
cc_379 N_SLEEP_c_359_n N_A_255_297#_c_1209_n 0.00221654f $X=4.57 $Y=1.16 $X2=0
+ $Y2=0
cc_380 N_SLEEP_M1006_g N_KAPWR_c_1305_n 0.00229224f $X=3.31 $Y=1.985 $X2=0 $Y2=0
cc_381 N_SLEEP_M1034_g N_KAPWR_c_1305_n 0.00230559f $X=3.73 $Y=1.985 $X2=0 $Y2=0
cc_382 N_SLEEP_M1039_g N_KAPWR_c_1305_n 0.00230559f $X=4.15 $Y=1.985 $X2=0 $Y2=0
cc_383 N_SLEEP_M1053_g N_KAPWR_c_1305_n 0.00230559f $X=4.57 $Y=1.985 $X2=0 $Y2=0
cc_384 N_SLEEP_c_354_n N_VGND_c_1847_n 0.00146448f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_385 N_SLEEP_c_354_n N_VGND_c_1848_n 0.00423334f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_386 N_SLEEP_c_355_n N_VGND_c_1848_n 0.00423334f $X=3.73 $Y=0.995 $X2=0 $Y2=0
cc_387 N_SLEEP_c_355_n N_VGND_c_1849_n 0.00146448f $X=3.73 $Y=0.995 $X2=0 $Y2=0
cc_388 N_SLEEP_c_356_n N_VGND_c_1849_n 0.00146339f $X=4.15 $Y=0.995 $X2=0 $Y2=0
cc_389 N_SLEEP_c_356_n N_VGND_c_1883_n 0.00423334f $X=4.15 $Y=0.995 $X2=0 $Y2=0
cc_390 N_SLEEP_c_357_n N_VGND_c_1883_n 0.00541359f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_391 N_SLEEP_c_357_n N_VGND_c_1884_n 4.62653e-19 $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_392 N_SLEEP_c_357_n N_VGND_c_1885_n 0.00336547f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_393 N_SLEEP_c_354_n N_VGND_c_1890_n 0.0054353f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_394 N_SLEEP_c_355_n N_VGND_c_1890_n 0.0054081f $X=3.73 $Y=0.995 $X2=0 $Y2=0
cc_395 N_SLEEP_c_356_n N_VGND_c_1890_n 0.0054081f $X=4.15 $Y=0.995 $X2=0 $Y2=0
cc_396 N_SLEEP_c_357_n N_VGND_c_1890_n 0.00731616f $X=4.57 $Y=0.995 $X2=0 $Y2=0
cc_397 N_A_341_47#_M1038_g N_A_1122_47#_M1013_g 0.0178631f $X=6.825 $Y=0.445
+ $X2=0 $Y2=0
cc_398 N_A_341_47#_c_468_n N_A_1122_47#_M1001_g 0.0178631f $X=6.825 $Y=1.41
+ $X2=0 $Y2=0
cc_399 N_A_341_47#_c_462_n N_A_1122_47#_c_683_n 0.0178631f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_400 N_A_341_47#_M1003_g N_A_1122_47#_c_685_n 0.00335375f $X=5.535 $Y=0.445
+ $X2=0 $Y2=0
cc_401 N_A_341_47#_M1007_g N_A_1122_47#_c_685_n 0.00353563f $X=5.965 $Y=0.445
+ $X2=0 $Y2=0
cc_402 N_A_341_47#_c_460_n N_A_1122_47#_c_685_n 0.00159345f $X=5.295 $Y=0.85
+ $X2=0 $Y2=0
cc_403 N_A_341_47#_c_461_n N_A_1122_47#_c_685_n 0.0217214f $X=5.295 $Y=0.85
+ $X2=0 $Y2=0
cc_404 N_A_341_47#_c_462_n N_A_1122_47#_c_685_n 0.0132485f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_405 N_A_341_47#_c_465_n N_A_1122_47#_c_705_n 0.00207315f $X=5.535 $Y=1.41
+ $X2=0 $Y2=0
cc_406 N_A_341_47#_c_466_n N_A_1122_47#_c_705_n 0.00124674f $X=5.965 $Y=1.41
+ $X2=0 $Y2=0
cc_407 N_A_341_47#_c_462_n N_A_1122_47#_c_705_n 0.00991177f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_408 N_A_341_47#_c_462_n N_A_1122_47#_c_719_n 0.0527608f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_409 N_A_341_47#_M1028_g N_A_1122_47#_c_686_n 0.00352135f $X=6.395 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_341_47#_M1038_g N_A_1122_47#_c_686_n 0.00356184f $X=6.825 $Y=0.445
+ $X2=0 $Y2=0
cc_411 N_A_341_47#_c_462_n N_A_1122_47#_c_686_n 0.0139367f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_412 N_A_341_47#_c_467_n N_A_1122_47#_c_706_n 0.00124674f $X=6.395 $Y=1.41
+ $X2=0 $Y2=0
cc_413 N_A_341_47#_c_468_n N_A_1122_47#_c_706_n 0.00207315f $X=6.825 $Y=1.41
+ $X2=0 $Y2=0
cc_414 N_A_341_47#_c_462_n N_A_1122_47#_c_706_n 0.00774413f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_415 N_A_341_47#_c_462_n N_A_1122_47#_c_687_n 0.0206088f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_416 N_A_341_47#_c_461_n N_A_1122_47#_c_727_n 0.0178087f $X=5.295 $Y=0.85
+ $X2=0 $Y2=0
cc_417 N_A_341_47#_c_462_n N_A_1122_47#_c_727_n 0.010956f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_418 N_A_341_47#_c_462_n N_A_1122_47#_c_729_n 0.00889636f $X=6.825 $Y=1.155
+ $X2=0 $Y2=0
cc_419 N_A_341_47#_c_465_n N_VPWR_c_1011_n 0.0054895f $X=5.535 $Y=1.41 $X2=0
+ $Y2=0
cc_420 N_A_341_47#_c_466_n N_VPWR_c_1011_n 0.0054895f $X=5.965 $Y=1.41 $X2=0
+ $Y2=0
cc_421 N_A_341_47#_c_467_n N_VPWR_c_1011_n 0.0054895f $X=6.395 $Y=1.41 $X2=0
+ $Y2=0
cc_422 N_A_341_47#_c_468_n N_VPWR_c_1011_n 0.0054895f $X=6.825 $Y=1.41 $X2=0
+ $Y2=0
cc_423 N_A_341_47#_M1005_s N_VPWR_c_1004_n 0.00110194f $X=1.705 $Y=1.485 $X2=0
+ $Y2=0
cc_424 N_A_341_47#_M1029_s N_VPWR_c_1004_n 0.00110194f $X=2.545 $Y=1.485 $X2=0
+ $Y2=0
cc_425 N_A_341_47#_c_465_n N_VPWR_c_1004_n 0.00642433f $X=5.535 $Y=1.41 $X2=0
+ $Y2=0
cc_426 N_A_341_47#_c_466_n N_VPWR_c_1004_n 0.00512464f $X=5.965 $Y=1.41 $X2=0
+ $Y2=0
cc_427 N_A_341_47#_c_467_n N_VPWR_c_1004_n 0.00512464f $X=6.395 $Y=1.41 $X2=0
+ $Y2=0
cc_428 N_A_341_47#_c_468_n N_VPWR_c_1004_n 0.00514998f $X=6.825 $Y=1.41 $X2=0
+ $Y2=0
cc_429 N_A_341_47#_c_470_n N_A_255_297#_M1017_d 0.00169861f $X=2.435 $Y=1.595
+ $X2=0 $Y2=0
cc_430 N_A_341_47#_M1005_s N_A_255_297#_c_1217_n 0.00220035f $X=1.705 $Y=1.485
+ $X2=0 $Y2=0
cc_431 N_A_341_47#_c_578_p N_A_255_297#_c_1217_n 0.0110552f $X=1.84 $Y=1.96
+ $X2=0 $Y2=0
cc_432 N_A_341_47#_c_470_n N_A_255_297#_c_1217_n 0.00186348f $X=2.435 $Y=1.595
+ $X2=0 $Y2=0
cc_433 N_A_341_47#_c_470_n N_A_255_297#_c_1219_n 0.0149761f $X=2.435 $Y=1.595
+ $X2=0 $Y2=0
cc_434 N_A_341_47#_M1029_s N_A_255_297#_c_1223_n 0.00220035f $X=2.545 $Y=1.485
+ $X2=0 $Y2=0
cc_435 N_A_341_47#_c_582_p N_A_255_297#_c_1223_n 0.0110552f $X=2.68 $Y=1.96
+ $X2=0 $Y2=0
cc_436 N_A_341_47#_c_472_n N_A_255_297#_c_1223_n 0.00183528f $X=2.68 $Y=1.62
+ $X2=0 $Y2=0
cc_437 N_A_341_47#_c_454_n N_A_255_297#_c_1204_n 0.0034284f $X=3.355 $Y=0.815
+ $X2=0 $Y2=0
cc_438 N_A_341_47#_c_472_n N_A_255_297#_c_1204_n 0.010246f $X=2.68 $Y=1.62 $X2=0
+ $Y2=0
cc_439 N_A_341_47#_c_457_n N_A_255_297#_c_1204_n 0.0041376f $X=3 $Y=0.85 $X2=0
+ $Y2=0
cc_440 N_A_341_47#_c_458_n N_A_255_297#_c_1204_n 0.00302006f $X=5.15 $Y=0.85
+ $X2=0 $Y2=0
cc_441 N_A_341_47#_c_464_n N_A_255_297#_c_1204_n 0.0038236f $X=3.095 $Y=0.845
+ $X2=0 $Y2=0
cc_442 N_A_341_47#_c_465_n N_A_255_297#_c_1207_n 0.00105964f $X=5.535 $Y=1.41
+ $X2=0 $Y2=0
cc_443 N_A_341_47#_c_458_n N_A_255_297#_c_1207_n 0.00597594f $X=5.15 $Y=0.85
+ $X2=0 $Y2=0
cc_444 N_A_341_47#_M1005_s N_KAPWR_c_1305_n 0.00373541f $X=1.705 $Y=1.485 $X2=0
+ $Y2=0
cc_445 N_A_341_47#_M1029_s N_KAPWR_c_1305_n 0.00373477f $X=2.545 $Y=1.485 $X2=0
+ $Y2=0
cc_446 N_A_341_47#_c_578_p N_KAPWR_c_1305_n 0.00559447f $X=1.84 $Y=1.96 $X2=0
+ $Y2=0
cc_447 N_A_341_47#_c_470_n N_KAPWR_c_1305_n 0.00560227f $X=2.435 $Y=1.595 $X2=0
+ $Y2=0
cc_448 N_A_341_47#_c_582_p N_KAPWR_c_1305_n 0.00559447f $X=2.68 $Y=1.96 $X2=0
+ $Y2=0
cc_449 N_A_341_47#_c_472_n N_KAPWR_c_1305_n 0.00365721f $X=2.68 $Y=1.62 $X2=0
+ $Y2=0
cc_450 N_A_341_47#_c_465_n N_KAPWR_c_1324_n 0.00604839f $X=5.535 $Y=1.41 $X2=0
+ $Y2=0
cc_451 N_A_341_47#_c_466_n N_KAPWR_c_1324_n 0.00604839f $X=5.965 $Y=1.41 $X2=0
+ $Y2=0
cc_452 N_A_341_47#_c_467_n N_KAPWR_c_1326_n 0.00604839f $X=6.395 $Y=1.41 $X2=0
+ $Y2=0
cc_453 N_A_341_47#_c_468_n N_KAPWR_c_1326_n 0.00604839f $X=6.825 $Y=1.41 $X2=0
+ $Y2=0
cc_454 N_A_341_47#_c_465_n N_KAPWR_c_1307_n 0.0105462f $X=5.535 $Y=1.41 $X2=0
+ $Y2=0
cc_455 N_A_341_47#_c_460_n N_KAPWR_c_1307_n 0.00117198f $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_456 N_A_341_47#_c_461_n N_KAPWR_c_1307_n 0.0231023f $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_457 N_A_341_47#_c_462_n N_KAPWR_c_1307_n 0.00809407f $X=6.825 $Y=1.155 $X2=0
+ $Y2=0
cc_458 N_A_341_47#_c_466_n N_KAPWR_c_1332_n 0.00968558f $X=5.965 $Y=1.41 $X2=0
+ $Y2=0
cc_459 N_A_341_47#_c_467_n N_KAPWR_c_1332_n 0.00972223f $X=6.395 $Y=1.41 $X2=0
+ $Y2=0
cc_460 N_A_341_47#_c_462_n N_KAPWR_c_1332_n 0.00281536f $X=6.825 $Y=1.155 $X2=0
+ $Y2=0
cc_461 N_A_341_47#_c_468_n N_KAPWR_c_1335_n 0.0097223f $X=6.825 $Y=1.41 $X2=0
+ $Y2=0
cc_462 N_A_341_47#_c_463_n N_VGND_M1009_d 0.00162089f $X=2.435 $Y=0.845 $X2=0
+ $Y2=0
cc_463 N_A_341_47#_c_454_n N_VGND_M1012_d 8.52008e-19 $X=3.355 $Y=0.815 $X2=0
+ $Y2=0
cc_464 N_A_341_47#_c_464_n N_VGND_M1012_d 7.65248e-19 $X=3.095 $Y=0.845 $X2=0
+ $Y2=0
cc_465 N_A_341_47#_c_455_n N_VGND_M1025_d 0.00162089f $X=4.195 $Y=0.815 $X2=0
+ $Y2=0
cc_466 N_A_341_47#_c_458_n N_VGND_M1030_d 6.81311e-19 $X=5.15 $Y=0.85 $X2=0
+ $Y2=0
cc_467 N_A_341_47#_c_452_n N_VGND_c_1845_n 0.00836079f $X=2.005 $Y=0.815 $X2=0
+ $Y2=0
cc_468 N_A_341_47#_c_463_n N_VGND_c_1846_n 0.0122559f $X=2.435 $Y=0.845 $X2=0
+ $Y2=0
cc_469 N_A_341_47#_c_458_n N_VGND_c_1847_n 3.27427e-19 $X=5.15 $Y=0.85 $X2=0
+ $Y2=0
cc_470 N_A_341_47#_c_459_n N_VGND_c_1847_n 5.11134e-19 $X=3.115 $Y=0.85 $X2=0
+ $Y2=0
cc_471 N_A_341_47#_c_464_n N_VGND_c_1847_n 0.0111038f $X=3.095 $Y=0.845 $X2=0
+ $Y2=0
cc_472 N_A_341_47#_c_454_n N_VGND_c_1848_n 0.00198695f $X=3.355 $Y=0.815 $X2=0
+ $Y2=0
cc_473 N_A_341_47#_c_499_n N_VGND_c_1848_n 0.0188551f $X=3.52 $Y=0.39 $X2=0
+ $Y2=0
cc_474 N_A_341_47#_c_455_n N_VGND_c_1848_n 0.00198695f $X=4.195 $Y=0.815 $X2=0
+ $Y2=0
cc_475 N_A_341_47#_c_455_n N_VGND_c_1849_n 0.0111016f $X=4.195 $Y=0.815 $X2=0
+ $Y2=0
cc_476 N_A_341_47#_c_458_n N_VGND_c_1849_n 8.00522e-19 $X=5.15 $Y=0.85 $X2=0
+ $Y2=0
cc_477 N_A_341_47#_M1007_g N_VGND_c_1850_n 0.00167912f $X=5.965 $Y=0.445 $X2=0
+ $Y2=0
cc_478 N_A_341_47#_M1028_g N_VGND_c_1850_n 0.00168046f $X=6.395 $Y=0.445 $X2=0
+ $Y2=0
cc_479 N_A_341_47#_c_462_n N_VGND_c_1850_n 0.00255763f $X=6.825 $Y=1.155 $X2=0
+ $Y2=0
cc_480 N_A_341_47#_M1038_g N_VGND_c_1851_n 0.00170359f $X=6.825 $Y=0.445 $X2=0
+ $Y2=0
cc_481 N_A_341_47#_c_475_n N_VGND_c_1865_n 0.0188551f $X=1.84 $Y=0.39 $X2=0
+ $Y2=0
cc_482 N_A_341_47#_c_463_n N_VGND_c_1865_n 0.00198695f $X=2.435 $Y=0.845 $X2=0
+ $Y2=0
cc_483 N_A_341_47#_c_496_n N_VGND_c_1867_n 0.0185141f $X=2.68 $Y=0.39 $X2=0
+ $Y2=0
cc_484 N_A_341_47#_c_463_n N_VGND_c_1867_n 0.00405835f $X=2.435 $Y=0.845 $X2=0
+ $Y2=0
cc_485 N_A_341_47#_M1028_g N_VGND_c_1869_n 0.00585385f $X=6.395 $Y=0.445 $X2=0
+ $Y2=0
cc_486 N_A_341_47#_M1038_g N_VGND_c_1869_n 0.00585385f $X=6.825 $Y=0.445 $X2=0
+ $Y2=0
cc_487 N_A_341_47#_M1003_g N_VGND_c_1879_n 0.00585385f $X=5.535 $Y=0.445 $X2=0
+ $Y2=0
cc_488 N_A_341_47#_M1007_g N_VGND_c_1879_n 0.00585385f $X=5.965 $Y=0.445 $X2=0
+ $Y2=0
cc_489 N_A_341_47#_c_455_n N_VGND_c_1883_n 0.00198695f $X=4.195 $Y=0.815 $X2=0
+ $Y2=0
cc_490 N_A_341_47#_c_524_n N_VGND_c_1883_n 0.0188551f $X=4.36 $Y=0.39 $X2=0
+ $Y2=0
cc_491 N_A_341_47#_M1003_g N_VGND_c_1884_n 0.00447753f $X=5.535 $Y=0.445 $X2=0
+ $Y2=0
cc_492 N_A_341_47#_c_455_n N_VGND_c_1884_n 0.00904186f $X=4.195 $Y=0.815 $X2=0
+ $Y2=0
cc_493 N_A_341_47#_c_458_n N_VGND_c_1884_n 0.0142417f $X=5.15 $Y=0.85 $X2=0
+ $Y2=0
cc_494 N_A_341_47#_c_460_n N_VGND_c_1884_n 3.50078e-19 $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_495 N_A_341_47#_c_461_n N_VGND_c_1884_n 0.0123196f $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_496 N_A_341_47#_M1003_g N_VGND_c_1885_n 0.00355103f $X=5.535 $Y=0.445 $X2=0
+ $Y2=0
cc_497 N_A_341_47#_c_458_n N_VGND_c_1885_n 0.00656345f $X=5.15 $Y=0.85 $X2=0
+ $Y2=0
cc_498 N_A_341_47#_c_460_n N_VGND_c_1885_n 0.00154076f $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_499 N_A_341_47#_c_461_n N_VGND_c_1885_n 0.020718f $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_500 N_A_341_47#_c_462_n N_VGND_c_1885_n 0.00139917f $X=6.825 $Y=1.155 $X2=0
+ $Y2=0
cc_501 N_A_341_47#_M1002_s N_VGND_c_1890_n 0.00215201f $X=1.705 $Y=0.235 $X2=0
+ $Y2=0
cc_502 N_A_341_47#_M1010_s N_VGND_c_1890_n 0.00170803f $X=2.545 $Y=0.235 $X2=0
+ $Y2=0
cc_503 N_A_341_47#_M1019_s N_VGND_c_1890_n 0.00177024f $X=3.385 $Y=0.235 $X2=0
+ $Y2=0
cc_504 N_A_341_47#_M1026_s N_VGND_c_1890_n 0.00177024f $X=4.225 $Y=0.235 $X2=0
+ $Y2=0
cc_505 N_A_341_47#_M1003_g N_VGND_c_1890_n 0.0118636f $X=5.535 $Y=0.445 $X2=0
+ $Y2=0
cc_506 N_A_341_47#_M1007_g N_VGND_c_1890_n 0.010643f $X=5.965 $Y=0.445 $X2=0
+ $Y2=0
cc_507 N_A_341_47#_M1028_g N_VGND_c_1890_n 0.010643f $X=6.395 $Y=0.445 $X2=0
+ $Y2=0
cc_508 N_A_341_47#_M1038_g N_VGND_c_1890_n 0.0106694f $X=6.825 $Y=0.445 $X2=0
+ $Y2=0
cc_509 N_A_341_47#_c_475_n N_VGND_c_1890_n 0.0122069f $X=1.84 $Y=0.39 $X2=0
+ $Y2=0
cc_510 N_A_341_47#_c_496_n N_VGND_c_1890_n 0.0054329f $X=2.68 $Y=0.39 $X2=0
+ $Y2=0
cc_511 N_A_341_47#_c_454_n N_VGND_c_1890_n 0.00166157f $X=3.355 $Y=0.815 $X2=0
+ $Y2=0
cc_512 N_A_341_47#_c_499_n N_VGND_c_1890_n 0.00580811f $X=3.52 $Y=0.39 $X2=0
+ $Y2=0
cc_513 N_A_341_47#_c_455_n N_VGND_c_1890_n 0.00370618f $X=4.195 $Y=0.815 $X2=0
+ $Y2=0
cc_514 N_A_341_47#_c_524_n N_VGND_c_1890_n 0.00580811f $X=4.36 $Y=0.39 $X2=0
+ $Y2=0
cc_515 N_A_341_47#_c_457_n N_VGND_c_1890_n 0.0317931f $X=3 $Y=0.85 $X2=0 $Y2=0
cc_516 N_A_341_47#_c_458_n N_VGND_c_1890_n 0.0904406f $X=5.15 $Y=0.85 $X2=0
+ $Y2=0
cc_517 N_A_341_47#_c_460_n N_VGND_c_1890_n 0.0131415f $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_518 N_A_341_47#_c_461_n N_VGND_c_1890_n 4.85517e-19 $X=5.295 $Y=0.85 $X2=0
+ $Y2=0
cc_519 N_A_341_47#_c_463_n N_VGND_c_1890_n 0.00942586f $X=2.435 $Y=0.845 $X2=0
+ $Y2=0
cc_520 N_A_341_47#_c_464_n N_VGND_c_1890_n 3.84928e-19 $X=3.095 $Y=0.845 $X2=0
+ $Y2=0
cc_521 N_A_1122_47#_M1001_g N_VPWR_c_1011_n 0.0054895f $X=7.255 $Y=1.985 $X2=0
+ $Y2=0
cc_522 N_A_1122_47#_M1004_g N_VPWR_c_1011_n 0.00585385f $X=7.685 $Y=1.985 $X2=0
+ $Y2=0
cc_523 N_A_1122_47#_M1008_g N_VPWR_c_1011_n 0.00585385f $X=8.115 $Y=1.985 $X2=0
+ $Y2=0
cc_524 N_A_1122_47#_M1011_g N_VPWR_c_1011_n 0.00585385f $X=8.545 $Y=1.985 $X2=0
+ $Y2=0
cc_525 N_A_1122_47#_M1018_g N_VPWR_c_1011_n 0.00585385f $X=8.975 $Y=1.985 $X2=0
+ $Y2=0
cc_526 N_A_1122_47#_M1021_g N_VPWR_c_1011_n 0.00585385f $X=9.405 $Y=1.985 $X2=0
+ $Y2=0
cc_527 N_A_1122_47#_M1022_g N_VPWR_c_1011_n 0.00585385f $X=9.835 $Y=1.985 $X2=0
+ $Y2=0
cc_528 N_A_1122_47#_M1031_g N_VPWR_c_1011_n 0.00585385f $X=10.265 $Y=1.985 $X2=0
+ $Y2=0
cc_529 N_A_1122_47#_M1033_g N_VPWR_c_1011_n 0.00585385f $X=10.69 $Y=1.985 $X2=0
+ $Y2=0
cc_530 N_A_1122_47#_M1035_g N_VPWR_c_1011_n 0.00585385f $X=11.12 $Y=1.985 $X2=0
+ $Y2=0
cc_531 N_A_1122_47#_M1036_g N_VPWR_c_1011_n 0.00585385f $X=11.55 $Y=1.985 $X2=0
+ $Y2=0
cc_532 N_A_1122_47#_M1040_g N_VPWR_c_1011_n 0.00585385f $X=11.98 $Y=1.985 $X2=0
+ $Y2=0
cc_533 N_A_1122_47#_M1043_g N_VPWR_c_1011_n 0.00585385f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_534 N_A_1122_47#_M1044_g N_VPWR_c_1011_n 0.00585385f $X=12.84 $Y=1.985 $X2=0
+ $Y2=0
cc_535 N_A_1122_47#_M1045_g N_VPWR_c_1011_n 0.00585385f $X=13.27 $Y=1.985 $X2=0
+ $Y2=0
cc_536 N_A_1122_47#_M1048_g N_VPWR_c_1011_n 0.00556673f $X=13.7 $Y=1.985 $X2=0
+ $Y2=0
cc_537 N_A_1122_47#_c_705_n N_VPWR_c_1011_n 0.0124538f $X=5.75 $Y=1.62 $X2=0
+ $Y2=0
cc_538 N_A_1122_47#_c_706_n N_VPWR_c_1011_n 0.0120686f $X=6.61 $Y=1.615 $X2=0
+ $Y2=0
cc_539 N_A_1122_47#_M1015_d N_VPWR_c_1004_n 0.00149727f $X=5.61 $Y=1.485 $X2=0
+ $Y2=0
cc_540 N_A_1122_47#_M1042_d N_VPWR_c_1004_n 0.00149767f $X=6.47 $Y=1.485 $X2=0
+ $Y2=0
cc_541 N_A_1122_47#_M1001_g N_VPWR_c_1004_n 0.00514998f $X=7.255 $Y=1.985 $X2=0
+ $Y2=0
cc_542 N_A_1122_47#_M1004_g N_VPWR_c_1004_n 0.00525209f $X=7.685 $Y=1.985 $X2=0
+ $Y2=0
cc_543 N_A_1122_47#_M1008_g N_VPWR_c_1004_n 0.00525209f $X=8.115 $Y=1.985 $X2=0
+ $Y2=0
cc_544 N_A_1122_47#_M1011_g N_VPWR_c_1004_n 0.00525209f $X=8.545 $Y=1.985 $X2=0
+ $Y2=0
cc_545 N_A_1122_47#_M1018_g N_VPWR_c_1004_n 0.00525209f $X=8.975 $Y=1.985 $X2=0
+ $Y2=0
cc_546 N_A_1122_47#_M1021_g N_VPWR_c_1004_n 0.00525209f $X=9.405 $Y=1.985 $X2=0
+ $Y2=0
cc_547 N_A_1122_47#_M1022_g N_VPWR_c_1004_n 0.00525209f $X=9.835 $Y=1.985 $X2=0
+ $Y2=0
cc_548 N_A_1122_47#_M1031_g N_VPWR_c_1004_n 0.00523845f $X=10.265 $Y=1.985 $X2=0
+ $Y2=0
cc_549 N_A_1122_47#_M1033_g N_VPWR_c_1004_n 0.00523845f $X=10.69 $Y=1.985 $X2=0
+ $Y2=0
cc_550 N_A_1122_47#_M1035_g N_VPWR_c_1004_n 0.00525209f $X=11.12 $Y=1.985 $X2=0
+ $Y2=0
cc_551 N_A_1122_47#_M1036_g N_VPWR_c_1004_n 0.00525209f $X=11.55 $Y=1.985 $X2=0
+ $Y2=0
cc_552 N_A_1122_47#_M1040_g N_VPWR_c_1004_n 0.00525209f $X=11.98 $Y=1.985 $X2=0
+ $Y2=0
cc_553 N_A_1122_47#_M1043_g N_VPWR_c_1004_n 0.00525209f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_554 N_A_1122_47#_M1044_g N_VPWR_c_1004_n 0.00525209f $X=12.84 $Y=1.985 $X2=0
+ $Y2=0
cc_555 N_A_1122_47#_M1045_g N_VPWR_c_1004_n 0.00525209f $X=13.27 $Y=1.985 $X2=0
+ $Y2=0
cc_556 N_A_1122_47#_M1048_g N_VPWR_c_1004_n 0.00622573f $X=13.7 $Y=1.985 $X2=0
+ $Y2=0
cc_557 N_A_1122_47#_c_705_n N_VPWR_c_1004_n 0.00174489f $X=5.75 $Y=1.62 $X2=0
+ $Y2=0
cc_558 N_A_1122_47#_c_706_n N_VPWR_c_1004_n 0.00175268f $X=6.61 $Y=1.615 $X2=0
+ $Y2=0
cc_559 N_A_1122_47#_M1045_g N_KAPWR_c_1304_n 0.00272513f $X=13.27 $Y=1.985 $X2=0
+ $Y2=0
cc_560 N_A_1122_47#_M1048_g N_KAPWR_c_1304_n 0.0023812f $X=13.7 $Y=1.985 $X2=0
+ $Y2=0
cc_561 N_A_1122_47#_c_705_n N_KAPWR_c_1338_n 4.33193e-19 $X=5.75 $Y=1.62 $X2=0
+ $Y2=0
cc_562 N_A_1122_47#_M1015_d N_KAPWR_c_1324_n 0.00380222f $X=5.61 $Y=1.485 $X2=0
+ $Y2=0
cc_563 N_A_1122_47#_c_705_n N_KAPWR_c_1324_n 0.0200676f $X=5.75 $Y=1.62 $X2=0
+ $Y2=0
cc_564 N_A_1122_47#_c_705_n N_KAPWR_c_1341_n 4.33193e-19 $X=5.75 $Y=1.62 $X2=0
+ $Y2=0
cc_565 N_A_1122_47#_c_706_n N_KAPWR_c_1341_n 4.33193e-19 $X=6.61 $Y=1.615 $X2=0
+ $Y2=0
cc_566 N_A_1122_47#_M1042_d N_KAPWR_c_1326_n 0.00380222f $X=6.47 $Y=1.485 $X2=0
+ $Y2=0
cc_567 N_A_1122_47#_c_706_n N_KAPWR_c_1326_n 0.0200378f $X=6.61 $Y=1.615 $X2=0
+ $Y2=0
cc_568 N_A_1122_47#_c_706_n N_KAPWR_c_1345_n 4.39484e-19 $X=6.61 $Y=1.615 $X2=0
+ $Y2=0
cc_569 N_A_1122_47#_M1004_g N_KAPWR_c_1346_n 0.00114528f $X=7.685 $Y=1.985 $X2=0
+ $Y2=0
cc_570 N_A_1122_47#_M1008_g N_KAPWR_c_1346_n 0.00114528f $X=8.115 $Y=1.985 $X2=0
+ $Y2=0
cc_571 N_A_1122_47#_M1001_g N_KAPWR_c_1348_n 0.00604839f $X=7.255 $Y=1.985 $X2=0
+ $Y2=0
cc_572 N_A_1122_47#_M1004_g N_KAPWR_c_1348_n 0.00233003f $X=7.685 $Y=1.985 $X2=0
+ $Y2=0
cc_573 N_A_1122_47#_M1004_g N_KAPWR_c_1350_n 6.91139e-19 $X=7.685 $Y=1.985 $X2=0
+ $Y2=0
cc_574 N_A_1122_47#_M1011_g N_KAPWR_c_1351_n 0.00115346f $X=8.545 $Y=1.985 $X2=0
+ $Y2=0
cc_575 N_A_1122_47#_M1018_g N_KAPWR_c_1351_n 0.00115346f $X=8.975 $Y=1.985 $X2=0
+ $Y2=0
cc_576 N_A_1122_47#_M1008_g N_KAPWR_c_1353_n 0.0026941f $X=8.115 $Y=1.985 $X2=0
+ $Y2=0
cc_577 N_A_1122_47#_M1011_g N_KAPWR_c_1353_n 0.0026941f $X=8.545 $Y=1.985 $X2=0
+ $Y2=0
cc_578 N_A_1122_47#_M1018_g N_KAPWR_c_1355_n 6.44793e-19 $X=8.975 $Y=1.985 $X2=0
+ $Y2=0
cc_579 N_A_1122_47#_M1021_g N_KAPWR_c_1356_n 0.00115346f $X=9.405 $Y=1.985 $X2=0
+ $Y2=0
cc_580 N_A_1122_47#_M1022_g N_KAPWR_c_1356_n 0.00115346f $X=9.835 $Y=1.985 $X2=0
+ $Y2=0
cc_581 N_A_1122_47#_M1018_g N_KAPWR_c_1358_n 0.00251207f $X=8.975 $Y=1.985 $X2=0
+ $Y2=0
cc_582 N_A_1122_47#_M1021_g N_KAPWR_c_1358_n 0.0026941f $X=9.405 $Y=1.985 $X2=0
+ $Y2=0
cc_583 N_A_1122_47#_M1022_g N_KAPWR_c_1360_n 6.44793e-19 $X=9.835 $Y=1.985 $X2=0
+ $Y2=0
cc_584 N_A_1122_47#_M1031_g N_KAPWR_c_1361_n 0.00113845f $X=10.265 $Y=1.985
+ $X2=0 $Y2=0
cc_585 N_A_1122_47#_M1033_g N_KAPWR_c_1361_n 0.00111208f $X=10.69 $Y=1.985 $X2=0
+ $Y2=0
cc_586 N_A_1122_47#_M1022_g N_KAPWR_c_1363_n 0.00251207f $X=9.835 $Y=1.985 $X2=0
+ $Y2=0
cc_587 N_A_1122_47#_M1031_g N_KAPWR_c_1363_n 0.00260308f $X=10.265 $Y=1.985
+ $X2=0 $Y2=0
cc_588 N_A_1122_47#_M1031_g N_KAPWR_c_1365_n 4.8879e-19 $X=10.265 $Y=1.985 $X2=0
+ $Y2=0
cc_589 N_A_1122_47#_M1033_g N_KAPWR_c_1365_n 6.40226e-19 $X=10.69 $Y=1.985 $X2=0
+ $Y2=0
cc_590 N_A_1122_47#_M1035_g N_KAPWR_c_1367_n 0.00116608f $X=11.12 $Y=1.985 $X2=0
+ $Y2=0
cc_591 N_A_1122_47#_M1036_g N_KAPWR_c_1367_n 0.00112416f $X=11.55 $Y=1.985 $X2=0
+ $Y2=0
cc_592 N_A_1122_47#_M1033_g N_KAPWR_c_1369_n 0.00251207f $X=10.69 $Y=1.985 $X2=0
+ $Y2=0
cc_593 N_A_1122_47#_M1035_g N_KAPWR_c_1369_n 0.0026941f $X=11.12 $Y=1.985 $X2=0
+ $Y2=0
cc_594 N_A_1122_47#_M1036_g N_KAPWR_c_1371_n 6.40226e-19 $X=11.55 $Y=1.985 $X2=0
+ $Y2=0
cc_595 N_A_1122_47#_M1040_g N_KAPWR_c_1372_n 0.00116608f $X=11.98 $Y=1.985 $X2=0
+ $Y2=0
cc_596 N_A_1122_47#_M1043_g N_KAPWR_c_1372_n 0.00112416f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_597 N_A_1122_47#_M1036_g N_KAPWR_c_1374_n 0.00251207f $X=11.55 $Y=1.985 $X2=0
+ $Y2=0
cc_598 N_A_1122_47#_M1040_g N_KAPWR_c_1374_n 0.00260308f $X=11.98 $Y=1.985 $X2=0
+ $Y2=0
cc_599 N_A_1122_47#_M1040_g N_KAPWR_c_1376_n 4.93728e-19 $X=11.98 $Y=1.985 $X2=0
+ $Y2=0
cc_600 N_A_1122_47#_M1043_g N_KAPWR_c_1376_n 3.61486e-19 $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_601 N_A_1122_47#_M1044_g N_KAPWR_c_1378_n 0.00116801f $X=12.84 $Y=1.985 $X2=0
+ $Y2=0
cc_602 N_A_1122_47#_M1045_g N_KAPWR_c_1378_n 0.00115258f $X=13.27 $Y=1.985 $X2=0
+ $Y2=0
cc_603 N_A_1122_47#_c_683_n N_KAPWR_c_1378_n 3.46041e-19 $X=13.7 $Y=0.95 $X2=0
+ $Y2=0
cc_604 N_A_1122_47#_M1043_g N_KAPWR_c_1381_n 0.00260308f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_605 N_A_1122_47#_M1044_g N_KAPWR_c_1381_n 0.00244893f $X=12.84 $Y=1.985 $X2=0
+ $Y2=0
cc_606 N_A_1122_47#_M1044_g N_KAPWR_c_1383_n 6.11058e-19 $X=12.84 $Y=1.985 $X2=0
+ $Y2=0
cc_607 N_A_1122_47#_M1048_g N_KAPWR_c_1306_n 0.00394183f $X=13.7 $Y=1.985 $X2=0
+ $Y2=0
cc_608 N_A_1122_47#_c_705_n N_KAPWR_c_1307_n 0.0388243f $X=5.75 $Y=1.62 $X2=0
+ $Y2=0
cc_609 N_A_1122_47#_c_705_n N_KAPWR_c_1332_n 0.0388243f $X=5.75 $Y=1.62 $X2=0
+ $Y2=0
cc_610 N_A_1122_47#_c_719_n N_KAPWR_c_1332_n 0.0212385f $X=6.49 $Y=1.2 $X2=0
+ $Y2=0
cc_611 N_A_1122_47#_c_706_n N_KAPWR_c_1332_n 0.0386342f $X=6.61 $Y=1.615 $X2=0
+ $Y2=0
cc_612 N_A_1122_47#_M1001_g N_KAPWR_c_1335_n 0.00962434f $X=7.255 $Y=1.985 $X2=0
+ $Y2=0
cc_613 N_A_1122_47#_c_706_n N_KAPWR_c_1335_n 0.0386367f $X=6.61 $Y=1.615 $X2=0
+ $Y2=0
cc_614 N_A_1122_47#_c_687_n N_KAPWR_c_1335_n 0.0223469f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_615 N_A_1122_47#_M1013_g N_X_c_1543_n 0.00120255f $X=7.255 $Y=0.445 $X2=0
+ $Y2=0
cc_616 N_A_1122_47#_M1014_g N_X_c_1543_n 0.00120255f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_617 N_A_1122_47#_c_686_n N_X_c_1543_n 0.00257148f $X=6.61 $Y=0.445 $X2=0
+ $Y2=0
cc_618 N_A_1122_47#_M1014_g N_X_c_1544_n 0.0119364f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_619 N_A_1122_47#_M1016_g N_X_c_1544_n 0.0122327f $X=8.115 $Y=0.445 $X2=0
+ $Y2=0
cc_620 N_A_1122_47#_c_683_n N_X_c_1544_n 0.00267078f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_621 N_A_1122_47#_c_687_n N_X_c_1544_n 0.0429599f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_622 N_A_1122_47#_M1013_g N_X_c_1545_n 0.00289158f $X=7.255 $Y=0.445 $X2=0
+ $Y2=0
cc_623 N_A_1122_47#_c_683_n N_X_c_1545_n 0.00277135f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_624 N_A_1122_47#_c_686_n N_X_c_1545_n 0.00599637f $X=6.61 $Y=0.445 $X2=0
+ $Y2=0
cc_625 N_A_1122_47#_c_687_n N_X_c_1545_n 0.0213686f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_626 N_A_1122_47#_M1004_g N_X_c_1579_n 0.0113432f $X=7.685 $Y=1.985 $X2=0
+ $Y2=0
cc_627 N_A_1122_47#_M1008_g N_X_c_1579_n 0.0113034f $X=8.115 $Y=1.985 $X2=0
+ $Y2=0
cc_628 N_A_1122_47#_c_683_n N_X_c_1579_n 0.00232005f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_629 N_A_1122_47#_c_687_n N_X_c_1579_n 0.0385727f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_630 N_A_1122_47#_M1016_g N_X_c_1546_n 0.00120255f $X=8.115 $Y=0.445 $X2=0
+ $Y2=0
cc_631 N_A_1122_47#_M1020_g N_X_c_1546_n 0.00120255f $X=8.545 $Y=0.445 $X2=0
+ $Y2=0
cc_632 N_A_1122_47#_M1020_g N_X_c_1547_n 0.0122792f $X=8.545 $Y=0.445 $X2=0
+ $Y2=0
cc_633 N_A_1122_47#_M1023_g N_X_c_1547_n 0.0122792f $X=8.975 $Y=0.445 $X2=0
+ $Y2=0
cc_634 N_A_1122_47#_c_683_n N_X_c_1547_n 0.00267078f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_635 N_A_1122_47#_c_687_n N_X_c_1547_n 0.0429599f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_636 N_A_1122_47#_M1011_g N_X_c_1589_n 0.0113694f $X=8.545 $Y=1.985 $X2=0
+ $Y2=0
cc_637 N_A_1122_47#_M1018_g N_X_c_1589_n 0.0113563f $X=8.975 $Y=1.985 $X2=0
+ $Y2=0
cc_638 N_A_1122_47#_c_683_n N_X_c_1589_n 0.00232005f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_639 N_A_1122_47#_c_687_n N_X_c_1589_n 0.0385727f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_640 N_A_1122_47#_M1023_g N_X_c_1548_n 0.00120255f $X=8.975 $Y=0.445 $X2=0
+ $Y2=0
cc_641 N_A_1122_47#_M1024_g N_X_c_1548_n 0.00118828f $X=9.405 $Y=0.445 $X2=0
+ $Y2=0
cc_642 N_A_1122_47#_M1024_g N_X_c_1549_n 0.0122792f $X=9.405 $Y=0.445 $X2=0
+ $Y2=0
cc_643 N_A_1122_47#_M1027_g N_X_c_1549_n 0.00994201f $X=9.835 $Y=0.445 $X2=0
+ $Y2=0
cc_644 N_A_1122_47#_c_683_n N_X_c_1549_n 0.00267078f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_645 N_A_1122_47#_c_687_n N_X_c_1549_n 0.0418783f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_646 N_A_1122_47#_M1021_g N_X_c_1599_n 0.0113694f $X=9.405 $Y=1.985 $X2=0
+ $Y2=0
cc_647 N_A_1122_47#_M1022_g N_X_c_1599_n 0.0113007f $X=9.835 $Y=1.985 $X2=0
+ $Y2=0
cc_648 N_A_1122_47#_c_683_n N_X_c_1599_n 0.00232005f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_649 N_A_1122_47#_c_687_n N_X_c_1599_n 0.0385727f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_650 N_A_1122_47#_M1024_g N_X_c_1550_n 5.05907e-19 $X=9.405 $Y=0.445 $X2=0
+ $Y2=0
cc_651 N_A_1122_47#_M1027_g N_X_c_1550_n 0.0062908f $X=9.835 $Y=0.445 $X2=0
+ $Y2=0
cc_652 N_A_1122_47#_M1041_g N_X_c_1550_n 0.00119799f $X=10.265 $Y=0.445 $X2=0
+ $Y2=0
cc_653 N_A_1122_47#_M1041_g N_X_c_1551_n 0.0122482f $X=10.265 $Y=0.445 $X2=0
+ $Y2=0
cc_654 N_A_1122_47#_M1046_g N_X_c_1551_n 0.0101865f $X=10.69 $Y=0.445 $X2=0
+ $Y2=0
cc_655 N_A_1122_47#_c_683_n N_X_c_1551_n 0.00253724f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_656 N_A_1122_47#_c_687_n N_X_c_1551_n 0.0418596f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_657 N_A_1122_47#_M1031_g N_X_c_1610_n 0.0113189f $X=10.265 $Y=1.985 $X2=0
+ $Y2=0
cc_658 N_A_1122_47#_M1033_g N_X_c_1610_n 0.0113123f $X=10.69 $Y=1.985 $X2=0
+ $Y2=0
cc_659 N_A_1122_47#_c_683_n N_X_c_1610_n 0.00220405f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_660 N_A_1122_47#_c_687_n N_X_c_1610_n 0.0378421f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_661 N_A_1122_47#_M1046_g N_X_c_1552_n 0.00121272f $X=10.69 $Y=0.445 $X2=0
+ $Y2=0
cc_662 N_A_1122_47#_M1047_g N_X_c_1552_n 0.00117849f $X=11.12 $Y=0.445 $X2=0
+ $Y2=0
cc_663 N_A_1122_47#_M1047_g N_X_c_1553_n 0.0122792f $X=11.12 $Y=0.445 $X2=0
+ $Y2=0
cc_664 N_A_1122_47#_M1049_g N_X_c_1553_n 0.0102175f $X=11.55 $Y=0.445 $X2=0
+ $Y2=0
cc_665 N_A_1122_47#_c_683_n N_X_c_1553_n 0.00267078f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_666 N_A_1122_47#_c_687_n N_X_c_1553_n 0.0429636f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_667 N_A_1122_47#_M1035_g N_X_c_1620_n 0.0113694f $X=11.12 $Y=1.985 $X2=0
+ $Y2=0
cc_668 N_A_1122_47#_M1036_g N_X_c_1620_n 0.0113563f $X=11.55 $Y=1.985 $X2=0
+ $Y2=0
cc_669 N_A_1122_47#_c_683_n N_X_c_1620_n 0.00232005f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_670 N_A_1122_47#_c_687_n N_X_c_1620_n 0.0385727f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_671 N_A_1122_47#_M1049_g N_X_c_1554_n 0.00122723f $X=11.55 $Y=0.445 $X2=0
+ $Y2=0
cc_672 N_A_1122_47#_M1050_g N_X_c_1554_n 0.00117849f $X=11.98 $Y=0.445 $X2=0
+ $Y2=0
cc_673 N_A_1122_47#_M1050_g N_X_c_1555_n 0.0122792f $X=11.98 $Y=0.445 $X2=0
+ $Y2=0
cc_674 N_A_1122_47#_M1051_g N_X_c_1555_n 0.0102175f $X=12.41 $Y=0.445 $X2=0
+ $Y2=0
cc_675 N_A_1122_47#_c_683_n N_X_c_1555_n 0.00267078f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_676 N_A_1122_47#_c_687_n N_X_c_1555_n 0.0429636f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_677 N_A_1122_47#_M1040_g N_X_c_1630_n 0.011359f $X=11.98 $Y=1.985 $X2=0 $Y2=0
cc_678 N_A_1122_47#_M1043_g N_X_c_1630_n 0.0113628f $X=12.41 $Y=1.985 $X2=0
+ $Y2=0
cc_679 N_A_1122_47#_c_683_n N_X_c_1630_n 0.00232005f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_680 N_A_1122_47#_c_687_n N_X_c_1630_n 0.0385727f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_681 N_A_1122_47#_M1051_g N_X_c_1556_n 0.00122723f $X=12.41 $Y=0.445 $X2=0
+ $Y2=0
cc_682 N_A_1122_47#_M1055_g N_X_c_1556_n 0.00118774f $X=12.84 $Y=0.445 $X2=0
+ $Y2=0
cc_683 N_A_1122_47#_M1055_g N_X_c_1557_n 0.0141891f $X=12.84 $Y=0.445 $X2=0
+ $Y2=0
cc_684 N_A_1122_47#_c_687_n N_X_c_1557_n 3.30399e-19 $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_685 N_A_1122_47#_M1056_g N_X_c_1558_n 0.00121196f $X=13.27 $Y=0.445 $X2=0
+ $Y2=0
cc_686 N_A_1122_47#_M1057_g N_X_c_1558_n 0.00221636f $X=13.7 $Y=0.445 $X2=0
+ $Y2=0
cc_687 N_A_1122_47#_M1001_g N_X_c_1640_n 0.00117531f $X=7.255 $Y=1.985 $X2=0
+ $Y2=0
cc_688 N_A_1122_47#_M1004_g N_X_c_1640_n 0.00127033f $X=7.685 $Y=1.985 $X2=0
+ $Y2=0
cc_689 N_A_1122_47#_c_683_n N_X_c_1640_n 0.00238948f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_690 N_A_1122_47#_c_687_n N_X_c_1640_n 0.0155795f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_691 N_A_1122_47#_c_683_n N_X_c_1559_n 0.00277135f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_692 N_A_1122_47#_c_687_n N_X_c_1559_n 0.0213686f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_693 N_A_1122_47#_M1008_g N_X_c_1646_n 0.00127532f $X=8.115 $Y=1.985 $X2=0
+ $Y2=0
cc_694 N_A_1122_47#_M1011_g N_X_c_1646_n 0.00127684f $X=8.545 $Y=1.985 $X2=0
+ $Y2=0
cc_695 N_A_1122_47#_c_683_n N_X_c_1646_n 0.00238948f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_696 N_A_1122_47#_c_687_n N_X_c_1646_n 0.0168441f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_697 N_A_1122_47#_c_683_n N_X_c_1560_n 0.00277135f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_698 N_A_1122_47#_c_687_n N_X_c_1560_n 0.0213686f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_699 N_A_1122_47#_M1018_g N_X_c_1652_n 0.00127684f $X=8.975 $Y=1.985 $X2=0
+ $Y2=0
cc_700 N_A_1122_47#_M1021_g N_X_c_1652_n 0.00127684f $X=9.405 $Y=1.985 $X2=0
+ $Y2=0
cc_701 N_A_1122_47#_c_683_n N_X_c_1652_n 0.00238948f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_702 N_A_1122_47#_c_687_n N_X_c_1652_n 0.0168441f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_703 N_A_1122_47#_M1027_g N_X_c_1561_n 0.00211052f $X=9.835 $Y=0.445 $X2=0
+ $Y2=0
cc_704 N_A_1122_47#_c_683_n N_X_c_1561_n 0.00277135f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_705 N_A_1122_47#_c_687_n N_X_c_1561_n 0.0225791f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_706 N_A_1122_47#_M1022_g N_X_c_1659_n 0.00127684f $X=9.835 $Y=1.985 $X2=0
+ $Y2=0
cc_707 N_A_1122_47#_M1031_g N_X_c_1659_n 0.00127684f $X=10.265 $Y=1.985 $X2=0
+ $Y2=0
cc_708 N_A_1122_47#_c_683_n N_X_c_1659_n 0.00238948f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_709 N_A_1122_47#_c_687_n N_X_c_1659_n 0.0168441f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_710 N_A_1122_47#_M1046_g N_X_c_1562_n 0.00203048f $X=10.69 $Y=0.445 $X2=0
+ $Y2=0
cc_711 N_A_1122_47#_c_683_n N_X_c_1562_n 0.00277135f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_712 N_A_1122_47#_c_687_n N_X_c_1562_n 0.0213686f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_713 N_A_1122_47#_M1035_g N_X_c_1666_n 0.0012701f $X=11.12 $Y=1.985 $X2=0
+ $Y2=0
cc_714 N_A_1122_47#_c_683_n N_X_c_1666_n 0.00238948f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_715 N_A_1122_47#_c_687_n N_X_c_1666_n 0.0168441f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_716 N_A_1122_47#_M1049_g N_X_c_1563_n 0.00203048f $X=11.55 $Y=0.445 $X2=0
+ $Y2=0
cc_717 N_A_1122_47#_c_683_n N_X_c_1563_n 0.00277135f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_718 N_A_1122_47#_c_687_n N_X_c_1563_n 0.0213686f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_719 N_A_1122_47#_M1040_g N_X_c_1672_n 0.0012701f $X=11.98 $Y=1.985 $X2=0
+ $Y2=0
cc_720 N_A_1122_47#_c_683_n N_X_c_1672_n 0.00238948f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_721 N_A_1122_47#_c_687_n N_X_c_1672_n 0.0168441f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_722 N_A_1122_47#_M1051_g N_X_c_1564_n 0.00203048f $X=12.41 $Y=0.445 $X2=0
+ $Y2=0
cc_723 N_A_1122_47#_c_683_n N_X_c_1564_n 0.00277135f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_724 N_A_1122_47#_c_687_n N_X_c_1564_n 0.0213686f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_725 N_A_1122_47#_M1055_g X 0.00147955f $X=12.84 $Y=0.445 $X2=0 $Y2=0
cc_726 N_A_1122_47#_M1044_g X 0.00539328f $X=12.84 $Y=1.985 $X2=0 $Y2=0
cc_727 N_A_1122_47#_M1056_g X 0.011848f $X=13.27 $Y=0.445 $X2=0 $Y2=0
cc_728 N_A_1122_47#_M1045_g X 0.00605481f $X=13.27 $Y=1.985 $X2=0 $Y2=0
cc_729 N_A_1122_47#_c_683_n X 0.0567372f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_730 N_A_1122_47#_M1057_g X 0.0136957f $X=13.7 $Y=0.445 $X2=0 $Y2=0
cc_731 N_A_1122_47#_M1048_g X 0.00773738f $X=13.7 $Y=1.985 $X2=0 $Y2=0
cc_732 N_A_1122_47#_c_687_n X 0.0208936f $X=12.565 $Y=1.16 $X2=0 $Y2=0
cc_733 N_A_1122_47#_M1044_g N_X_c_1567_n 0.0141741f $X=12.84 $Y=1.985 $X2=0
+ $Y2=0
cc_734 N_A_1122_47#_M1045_g N_X_c_1567_n 0.0106923f $X=13.27 $Y=1.985 $X2=0
+ $Y2=0
cc_735 N_A_1122_47#_c_683_n N_X_c_1567_n 0.00238948f $X=13.7 $Y=0.95 $X2=0 $Y2=0
cc_736 N_A_1122_47#_M1048_g N_X_c_1567_n 0.025394f $X=13.7 $Y=1.985 $X2=0 $Y2=0
cc_737 N_A_1122_47#_c_687_n N_X_c_1567_n 0.0170247f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_738 N_A_1122_47#_c_719_n N_VGND_c_1850_n 0.00764914f $X=6.49 $Y=1.2 $X2=0
+ $Y2=0
cc_739 N_A_1122_47#_M1013_g N_VGND_c_1851_n 0.00170359f $X=7.255 $Y=0.445 $X2=0
+ $Y2=0
cc_740 N_A_1122_47#_c_687_n N_VGND_c_1851_n 0.0091835f $X=12.565 $Y=1.16 $X2=0
+ $Y2=0
cc_741 N_A_1122_47#_M1014_g N_VGND_c_1852_n 0.00161372f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_742 N_A_1122_47#_M1016_g N_VGND_c_1852_n 0.00161372f $X=8.115 $Y=0.445 $X2=0
+ $Y2=0
cc_743 N_A_1122_47#_M1020_g N_VGND_c_1853_n 0.00161372f $X=8.545 $Y=0.445 $X2=0
+ $Y2=0
cc_744 N_A_1122_47#_M1023_g N_VGND_c_1853_n 0.00161372f $X=8.975 $Y=0.445 $X2=0
+ $Y2=0
cc_745 N_A_1122_47#_M1024_g N_VGND_c_1854_n 0.00160579f $X=9.405 $Y=0.445 $X2=0
+ $Y2=0
cc_746 N_A_1122_47#_M1027_g N_VGND_c_1854_n 0.0015619f $X=9.835 $Y=0.445 $X2=0
+ $Y2=0
cc_747 N_A_1122_47#_M1027_g N_VGND_c_1855_n 0.00438144f $X=9.835 $Y=0.445 $X2=0
+ $Y2=0
cc_748 N_A_1122_47#_M1041_g N_VGND_c_1855_n 0.00439206f $X=10.265 $Y=0.445 $X2=0
+ $Y2=0
cc_749 N_A_1122_47#_M1041_g N_VGND_c_1856_n 0.00161724f $X=10.265 $Y=0.445 $X2=0
+ $Y2=0
cc_750 N_A_1122_47#_M1046_g N_VGND_c_1856_n 0.00156827f $X=10.69 $Y=0.445 $X2=0
+ $Y2=0
cc_751 N_A_1122_47#_M1046_g N_VGND_c_1857_n 0.00439206f $X=10.69 $Y=0.445 $X2=0
+ $Y2=0
cc_752 N_A_1122_47#_M1047_g N_VGND_c_1857_n 0.00439206f $X=11.12 $Y=0.445 $X2=0
+ $Y2=0
cc_753 N_A_1122_47#_M1047_g N_VGND_c_1858_n 0.00162174f $X=11.12 $Y=0.445 $X2=0
+ $Y2=0
cc_754 N_A_1122_47#_M1049_g N_VGND_c_1858_n 0.00157905f $X=11.55 $Y=0.445 $X2=0
+ $Y2=0
cc_755 N_A_1122_47#_M1050_g N_VGND_c_1859_n 0.00162174f $X=11.98 $Y=0.445 $X2=0
+ $Y2=0
cc_756 N_A_1122_47#_M1051_g N_VGND_c_1859_n 0.00157905f $X=12.41 $Y=0.445 $X2=0
+ $Y2=0
cc_757 N_A_1122_47#_M1055_g N_VGND_c_1860_n 0.00162705f $X=12.84 $Y=0.445 $X2=0
+ $Y2=0
cc_758 N_A_1122_47#_M1056_g N_VGND_c_1860_n 0.00161372f $X=13.27 $Y=0.445 $X2=0
+ $Y2=0
cc_759 N_A_1122_47#_c_683_n N_VGND_c_1860_n 4.7914e-19 $X=13.7 $Y=0.95 $X2=0
+ $Y2=0
cc_760 N_A_1122_47#_M1057_g N_VGND_c_1862_n 0.00341923f $X=13.7 $Y=0.445 $X2=0
+ $Y2=0
cc_761 N_A_1122_47#_c_686_n N_VGND_c_1869_n 0.0137163f $X=6.61 $Y=0.445 $X2=0
+ $Y2=0
cc_762 N_A_1122_47#_M1013_g N_VGND_c_1871_n 0.00585385f $X=7.255 $Y=0.445 $X2=0
+ $Y2=0
cc_763 N_A_1122_47#_M1014_g N_VGND_c_1871_n 0.00439206f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_764 N_A_1122_47#_M1016_g N_VGND_c_1873_n 0.00439206f $X=8.115 $Y=0.445 $X2=0
+ $Y2=0
cc_765 N_A_1122_47#_M1020_g N_VGND_c_1873_n 0.00439206f $X=8.545 $Y=0.445 $X2=0
+ $Y2=0
cc_766 N_A_1122_47#_M1023_g N_VGND_c_1875_n 0.00439206f $X=8.975 $Y=0.445 $X2=0
+ $Y2=0
cc_767 N_A_1122_47#_M1024_g N_VGND_c_1875_n 0.00439206f $X=9.405 $Y=0.445 $X2=0
+ $Y2=0
cc_768 N_A_1122_47#_M1051_g N_VGND_c_1877_n 0.00439206f $X=12.41 $Y=0.445 $X2=0
+ $Y2=0
cc_769 N_A_1122_47#_M1055_g N_VGND_c_1877_n 0.00439206f $X=12.84 $Y=0.445 $X2=0
+ $Y2=0
cc_770 N_A_1122_47#_c_685_n N_VGND_c_1879_n 0.0128787f $X=5.75 $Y=0.445 $X2=0
+ $Y2=0
cc_771 N_A_1122_47#_M1049_g N_VGND_c_1880_n 0.00439206f $X=11.55 $Y=0.445 $X2=0
+ $Y2=0
cc_772 N_A_1122_47#_M1050_g N_VGND_c_1880_n 0.00439206f $X=11.98 $Y=0.445 $X2=0
+ $Y2=0
cc_773 N_A_1122_47#_M1056_g N_VGND_c_1881_n 0.00439071f $X=13.27 $Y=0.445 $X2=0
+ $Y2=0
cc_774 N_A_1122_47#_M1057_g N_VGND_c_1881_n 0.00439071f $X=13.7 $Y=0.445 $X2=0
+ $Y2=0
cc_775 N_A_1122_47#_M1003_d N_VGND_c_1890_n 0.00422994f $X=5.61 $Y=0.235 $X2=0
+ $Y2=0
cc_776 N_A_1122_47#_M1028_d N_VGND_c_1890_n 0.00336236f $X=6.47 $Y=0.235 $X2=0
+ $Y2=0
cc_777 N_A_1122_47#_M1013_g N_VGND_c_1890_n 0.0106694f $X=7.255 $Y=0.445 $X2=0
+ $Y2=0
cc_778 N_A_1122_47#_M1014_g N_VGND_c_1890_n 0.00590932f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_779 N_A_1122_47#_M1016_g N_VGND_c_1890_n 0.00590932f $X=8.115 $Y=0.445 $X2=0
+ $Y2=0
cc_780 N_A_1122_47#_M1020_g N_VGND_c_1890_n 0.00590932f $X=8.545 $Y=0.445 $X2=0
+ $Y2=0
cc_781 N_A_1122_47#_M1023_g N_VGND_c_1890_n 0.00590932f $X=8.975 $Y=0.445 $X2=0
+ $Y2=0
cc_782 N_A_1122_47#_M1024_g N_VGND_c_1890_n 0.00590932f $X=9.405 $Y=0.445 $X2=0
+ $Y2=0
cc_783 N_A_1122_47#_M1027_g N_VGND_c_1890_n 0.00587292f $X=9.835 $Y=0.445 $X2=0
+ $Y2=0
cc_784 N_A_1122_47#_M1041_g N_VGND_c_1890_n 0.00589619f $X=10.265 $Y=0.445 $X2=0
+ $Y2=0
cc_785 N_A_1122_47#_M1046_g N_VGND_c_1890_n 0.00592128f $X=10.69 $Y=0.445 $X2=0
+ $Y2=0
cc_786 N_A_1122_47#_M1047_g N_VGND_c_1890_n 0.00590932f $X=11.12 $Y=0.445 $X2=0
+ $Y2=0
cc_787 N_A_1122_47#_M1049_g N_VGND_c_1890_n 0.00593441f $X=11.55 $Y=0.445 $X2=0
+ $Y2=0
cc_788 N_A_1122_47#_M1050_g N_VGND_c_1890_n 0.00590932f $X=11.98 $Y=0.445 $X2=0
+ $Y2=0
cc_789 N_A_1122_47#_M1051_g N_VGND_c_1890_n 0.00593441f $X=12.41 $Y=0.445 $X2=0
+ $Y2=0
cc_790 N_A_1122_47#_M1055_g N_VGND_c_1890_n 0.00590932f $X=12.84 $Y=0.445 $X2=0
+ $Y2=0
cc_791 N_A_1122_47#_M1056_g N_VGND_c_1890_n 0.00590684f $X=13.27 $Y=0.445 $X2=0
+ $Y2=0
cc_792 N_A_1122_47#_M1057_g N_VGND_c_1890_n 0.00691049f $X=13.7 $Y=0.445 $X2=0
+ $Y2=0
cc_793 N_A_1122_47#_c_685_n N_VGND_c_1890_n 0.00854752f $X=5.75 $Y=0.445 $X2=0
+ $Y2=0
cc_794 N_A_1122_47#_c_686_n N_VGND_c_1890_n 0.00950576f $X=6.61 $Y=0.445 $X2=0
+ $Y2=0
cc_795 N_VPWR_c_1004_n N_A_255_297#_M1005_d 0.00115538f $X=14.03 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_796 N_VPWR_c_1004_n N_A_255_297#_M1017_d 0.00109368f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_797 N_VPWR_c_1004_n N_A_255_297#_M1052_d 0.00109368f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_798 N_VPWR_c_1004_n N_A_255_297#_M1034_d 0.00149677f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_799 N_VPWR_c_1004_n N_A_255_297#_M1053_d 0.00135692f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_800 N_VPWR_c_1009_n N_A_255_297#_c_1202_n 0.0247353f $X=3.435 $Y=2.72 $X2=0
+ $Y2=0
cc_801 N_VPWR_c_1004_n N_A_255_297#_c_1202_n 0.00347719f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_802 N_VPWR_c_1009_n N_A_255_297#_c_1217_n 0.0286211f $X=3.435 $Y=2.72 $X2=0
+ $Y2=0
cc_803 N_VPWR_c_1004_n N_A_255_297#_c_1217_n 0.00384286f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_804 N_VPWR_c_1009_n N_A_255_297#_c_1223_n 0.0286211f $X=3.435 $Y=2.72 $X2=0
+ $Y2=0
cc_805 N_VPWR_c_1004_n N_A_255_297#_c_1223_n 0.00384286f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_806 N_VPWR_c_1007_n N_A_255_297#_c_1226_n 0.0267961f $X=3.52 $Y=2 $X2=0 $Y2=0
cc_807 N_VPWR_c_1009_n N_A_255_297#_c_1226_n 0.0190403f $X=3.435 $Y=2.72 $X2=0
+ $Y2=0
cc_808 N_VPWR_c_1004_n N_A_255_297#_c_1226_n 0.00296342f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_809 N_VPWR_M1006_s N_A_255_297#_c_1205_n 0.00162649f $X=3.385 $Y=1.485 $X2=0
+ $Y2=0
cc_810 N_VPWR_c_1007_n N_A_255_297#_c_1205_n 0.0145488f $X=3.52 $Y=2 $X2=0 $Y2=0
cc_811 N_VPWR_c_1007_n N_A_255_297#_c_1276_n 0.0254999f $X=3.52 $Y=2 $X2=0 $Y2=0
cc_812 N_VPWR_c_1008_n N_A_255_297#_c_1276_n 0.026187f $X=4.36 $Y=2 $X2=0 $Y2=0
cc_813 N_VPWR_c_1010_n N_A_255_297#_c_1276_n 0.0113958f $X=4.195 $Y=2.72 $X2=0
+ $Y2=0
cc_814 N_VPWR_c_1004_n N_A_255_297#_c_1276_n 0.00155926f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_815 N_VPWR_M1039_s N_A_255_297#_c_1206_n 0.00162649f $X=4.225 $Y=1.485 $X2=0
+ $Y2=0
cc_816 N_VPWR_c_1008_n N_A_255_297#_c_1206_n 0.0166706f $X=4.36 $Y=2 $X2=0 $Y2=0
cc_817 N_VPWR_c_1008_n N_A_255_297#_c_1208_n 0.0262428f $X=4.36 $Y=2 $X2=0 $Y2=0
cc_818 N_VPWR_c_1011_n N_A_255_297#_c_1208_n 0.0194075f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_819 N_VPWR_c_1004_n N_A_255_297#_c_1208_n 0.00258021f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_820 N_VPWR_c_1009_n N_A_255_297#_c_1228_n 0.0187749f $X=3.435 $Y=2.72 $X2=0
+ $Y2=0
cc_821 N_VPWR_c_1004_n N_A_255_297#_c_1228_n 0.00288345f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_822 N_VPWR_c_1004_n N_KAPWR_M1015_s 0.00109164f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_823 N_VPWR_c_1004_n N_KAPWR_M1037_s 0.00113449f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_824 N_VPWR_c_1004_n N_KAPWR_M1054_s 0.00113449f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_825 N_VPWR_c_1004_n N_KAPWR_M1004_d 0.00122337f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_826 N_VPWR_c_1004_n N_KAPWR_M1011_d 0.00123133f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_827 N_VPWR_c_1004_n N_KAPWR_M1021_d 0.00123133f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_828 N_VPWR_c_1004_n N_KAPWR_M1031_d 0.00125123f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_829 N_VPWR_c_1004_n N_KAPWR_M1035_d 0.00129179f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_830 N_VPWR_c_1004_n N_KAPWR_M1040_d 0.00129179f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_831 N_VPWR_c_1004_n N_KAPWR_M1044_d 0.00125148f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_832 N_VPWR_c_1004_n N_KAPWR_M1048_d 0.00126099f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_833 N_VPWR_c_1011_n N_KAPWR_c_1304_n 0.00180822f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_834 N_VPWR_M1000_s N_KAPWR_c_1305_n 0.00212217f $X=0.305 $Y=1.485 $X2=0 $Y2=0
cc_835 N_VPWR_M1006_s N_KAPWR_c_1305_n 8.01534e-19 $X=3.385 $Y=1.485 $X2=0 $Y2=0
cc_836 N_VPWR_c_1005_n N_KAPWR_c_1305_n 3.19314e-19 $X=0.332 $Y=2.635 $X2=0
+ $Y2=0
cc_837 N_VPWR_c_1006_n N_KAPWR_c_1305_n 0.0429092f $X=0.45 $Y=1.66 $X2=0 $Y2=0
cc_838 N_VPWR_c_1007_n N_KAPWR_c_1305_n 0.0169826f $X=3.52 $Y=2 $X2=0 $Y2=0
cc_839 N_VPWR_c_1008_n N_KAPWR_c_1305_n 0.0210625f $X=4.36 $Y=2 $X2=0 $Y2=0
cc_840 N_VPWR_c_1009_n N_KAPWR_c_1305_n 0.00425632f $X=3.435 $Y=2.72 $X2=0 $Y2=0
cc_841 N_VPWR_c_1010_n N_KAPWR_c_1305_n 0.00182732f $X=4.195 $Y=2.72 $X2=0 $Y2=0
cc_842 N_VPWR_c_1011_n N_KAPWR_c_1305_n 0.00223609f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_843 N_VPWR_c_1004_n N_KAPWR_c_1305_n 1.43974f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_844 N_VPWR_c_1011_n N_KAPWR_c_1324_n 0.00207669f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_845 N_VPWR_c_1011_n N_KAPWR_c_1326_n 0.00207863f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_846 N_VPWR_c_1011_n N_KAPWR_c_1346_n 0.0147484f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_847 N_VPWR_c_1004_n N_KAPWR_c_1346_n 0.00236391f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_848 N_VPWR_c_1011_n N_KAPWR_c_1348_n 0.00186229f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_849 N_VPWR_c_1011_n N_KAPWR_c_1351_n 0.0147733f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_850 N_VPWR_c_1004_n N_KAPWR_c_1351_n 0.00234462f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_851 N_VPWR_c_1011_n N_KAPWR_c_1353_n 0.00187059f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_852 N_VPWR_c_1011_n N_KAPWR_c_1355_n 0.00102221f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_853 N_VPWR_c_1011_n N_KAPWR_c_1356_n 0.0147733f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_854 N_VPWR_c_1004_n N_KAPWR_c_1356_n 0.00234462f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_855 N_VPWR_c_1011_n N_KAPWR_c_1358_n 0.00102711f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_856 N_VPWR_c_1011_n N_KAPWR_c_1360_n 0.00102221f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_857 N_VPWR_c_1011_n N_KAPWR_c_1361_n 0.0140719f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_858 N_VPWR_c_1004_n N_KAPWR_c_1361_n 0.0022083f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_859 N_VPWR_c_1011_n N_KAPWR_c_1363_n 0.00102587f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_860 N_VPWR_c_1011_n N_KAPWR_c_1365_n 0.001017f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_861 N_VPWR_c_1011_n N_KAPWR_c_1367_n 0.0142411f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_862 N_VPWR_c_1004_n N_KAPWR_c_1367_n 0.0022083f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_863 N_VPWR_c_1011_n N_KAPWR_c_1369_n 0.00110732f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_864 N_VPWR_c_1011_n N_KAPWR_c_1371_n 0.001017f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_865 N_VPWR_c_1011_n N_KAPWR_c_1372_n 0.0142411f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_866 N_VPWR_c_1004_n N_KAPWR_c_1372_n 0.0022083f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_867 N_VPWR_c_1011_n N_KAPWR_c_1374_n 0.00110608f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_868 N_VPWR_c_1011_n N_KAPWR_c_1376_n 0.00101652f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_869 N_VPWR_c_1011_n N_KAPWR_c_1378_n 0.0145959f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_870 N_VPWR_c_1004_n N_KAPWR_c_1378_n 0.00229918f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_871 N_VPWR_c_1011_n N_KAPWR_c_1381_n 0.00110703f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_872 N_VPWR_c_1011_n N_KAPWR_c_1383_n 0.00101719f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_873 N_VPWR_c_1011_n N_KAPWR_c_1306_n 0.0181313f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_874 N_VPWR_c_1004_n N_KAPWR_c_1306_n 0.00244244f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_875 N_VPWR_c_1011_n N_KAPWR_c_1307_n 0.0210489f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_876 N_VPWR_c_1004_n N_KAPWR_c_1307_n 0.00300101f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_877 N_VPWR_c_1011_n N_KAPWR_c_1332_n 0.0189253f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_878 N_VPWR_c_1004_n N_KAPWR_c_1332_n 0.00295774f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_879 N_VPWR_c_1011_n N_KAPWR_c_1335_n 0.0189253f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_880 N_VPWR_c_1004_n N_KAPWR_c_1335_n 0.00295774f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_881 N_VPWR_c_1004_n N_X_M1001_s 0.00135666f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_882 N_VPWR_c_1004_n N_X_M1008_s 0.00121566f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_883 N_VPWR_c_1004_n N_X_M1018_s 0.00121566f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_884 N_VPWR_c_1004_n N_X_M1022_s 0.00121566f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_885 N_VPWR_c_1004_n N_X_M1033_s 0.00121566f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_886 N_VPWR_c_1004_n N_X_M1036_s 0.00121566f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_887 N_VPWR_c_1004_n N_X_M1043_s 0.00121566f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_888 N_VPWR_c_1004_n N_X_M1045_s 0.00117537f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_889 N_VPWR_c_1011_n N_X_c_1640_n 0.0132747f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_890 N_VPWR_c_1004_n N_X_c_1640_n 0.00207897f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_891 N_VPWR_c_1011_n N_X_c_1646_n 0.0144808f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_892 N_VPWR_c_1004_n N_X_c_1646_n 0.00240527f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_893 N_VPWR_c_1011_n N_X_c_1652_n 0.0144808f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_894 N_VPWR_c_1004_n N_X_c_1652_n 0.00240527f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_895 N_VPWR_c_1011_n N_X_c_1659_n 0.0144808f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_896 N_VPWR_c_1004_n N_X_c_1659_n 0.00240527f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_897 N_VPWR_c_1011_n N_X_c_1666_n 0.0144808f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_898 N_VPWR_c_1004_n N_X_c_1666_n 0.00240527f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_899 N_VPWR_c_1011_n N_X_c_1672_n 0.0144808f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_900 N_VPWR_c_1004_n N_X_c_1672_n 0.00240527f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_901 N_VPWR_c_1011_n N_X_c_1567_n 0.0305634f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_902 N_VPWR_c_1004_n N_X_c_1567_n 0.00505204f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_903 N_A_255_297#_M1034_d N_KAPWR_c_1305_n 0.00160307f $X=3.805 $Y=1.485 $X2=0
+ $Y2=0
cc_904 N_A_255_297#_M1053_d N_KAPWR_c_1305_n 8.01534e-19 $X=4.645 $Y=1.485 $X2=0
+ $Y2=0
cc_905 N_A_255_297#_c_1202_n N_KAPWR_c_1305_n 0.00536882f $X=1.395 $Y=2.295
+ $X2=0 $Y2=0
cc_906 N_A_255_297#_c_1203_n N_KAPWR_c_1305_n 0.0321654f $X=1.42 $Y=1.66 $X2=0
+ $Y2=0
cc_907 N_A_255_297#_c_1217_n N_KAPWR_c_1305_n 0.0134771f $X=2.095 $Y=2.38 $X2=0
+ $Y2=0
cc_908 N_A_255_297#_c_1219_n N_KAPWR_c_1305_n 0.0171794f $X=2.26 $Y=2.02 $X2=0
+ $Y2=0
cc_909 N_A_255_297#_c_1223_n N_KAPWR_c_1305_n 0.0134603f $X=2.935 $Y=2.38 $X2=0
+ $Y2=0
cc_910 N_A_255_297#_c_1226_n N_KAPWR_c_1305_n 0.0330753f $X=3.1 $Y=2.295 $X2=0
+ $Y2=0
cc_911 N_A_255_297#_c_1205_n N_KAPWR_c_1305_n 0.0113465f $X=3.855 $Y=1.56 $X2=0
+ $Y2=0
cc_912 N_A_255_297#_c_1276_n N_KAPWR_c_1305_n 0.0183511f $X=3.94 $Y=2.3 $X2=0
+ $Y2=0
cc_913 N_A_255_297#_c_1206_n N_KAPWR_c_1305_n 0.0116372f $X=4.695 $Y=1.56 $X2=0
+ $Y2=0
cc_914 N_A_255_297#_c_1208_n N_KAPWR_c_1305_n 0.0278853f $X=4.78 $Y=2.3 $X2=0
+ $Y2=0
cc_915 N_A_255_297#_c_1228_n N_KAPWR_c_1305_n 0.00427056f $X=2.26 $Y=2.38 $X2=0
+ $Y2=0
cc_916 N_A_255_297#_c_1208_n N_KAPWR_c_1338_n 4.44501e-19 $X=4.78 $Y=2.3 $X2=0
+ $Y2=0
cc_917 N_A_255_297#_c_1207_n N_KAPWR_c_1307_n 0.0144408f $X=4.835 $Y=1.665 $X2=0
+ $Y2=0
cc_918 N_A_255_297#_c_1208_n N_KAPWR_c_1307_n 0.0604757f $X=4.78 $Y=2.3 $X2=0
+ $Y2=0
cc_919 N_A_255_297#_c_1207_n N_VGND_c_1884_n 0.00607409f $X=4.835 $Y=1.665 $X2=0
+ $Y2=0
cc_920 N_KAPWR_c_1348_n N_X_M1001_s 0.00202712f $X=7.74 $Y=2.21 $X2=0 $Y2=0
cc_921 N_KAPWR_c_1353_n N_X_M1008_s 2.52013e-19 $X=8.62 $Y=2.21 $X2=0 $Y2=0
cc_922 N_KAPWR_c_1358_n N_X_M1018_s 2.52013e-19 $X=9.48 $Y=2.21 $X2=0 $Y2=0
cc_923 N_KAPWR_c_1363_n N_X_M1022_s 2.52013e-19 $X=10.335 $Y=2.21 $X2=0 $Y2=0
cc_924 N_KAPWR_c_1369_n N_X_M1033_s 2.83515e-19 $X=11.195 $Y=2.21 $X2=0 $Y2=0
cc_925 N_KAPWR_c_1374_n N_X_M1036_s 2.83515e-19 $X=12.05 $Y=2.21 $X2=0 $Y2=0
cc_926 N_KAPWR_c_1381_n N_X_M1043_s 2.86889e-19 $X=12.9 $Y=2.21 $X2=0 $Y2=0
cc_927 N_KAPWR_M1004_d N_X_c_1579_n 0.00325883f $X=7.76 $Y=1.485 $X2=0 $Y2=0
cc_928 N_KAPWR_c_1346_n N_X_c_1579_n 0.0127908f $X=7.885 $Y=2.21 $X2=0 $Y2=0
cc_929 N_KAPWR_c_1348_n N_X_c_1579_n 0.00434646f $X=7.74 $Y=2.21 $X2=0 $Y2=0
cc_930 N_KAPWR_c_1350_n N_X_c_1579_n 0.0023936f $X=8.03 $Y=2.21 $X2=0 $Y2=0
cc_931 N_KAPWR_c_1353_n N_X_c_1579_n 0.00532372f $X=8.62 $Y=2.21 $X2=0 $Y2=0
cc_932 N_KAPWR_M1011_d N_X_c_1589_n 0.00325489f $X=8.62 $Y=1.485 $X2=0 $Y2=0
cc_933 N_KAPWR_c_1351_n N_X_c_1589_n 0.0128604f $X=8.765 $Y=2.21 $X2=0 $Y2=0
cc_934 N_KAPWR_c_1353_n N_X_c_1589_n 0.00497471f $X=8.62 $Y=2.21 $X2=0 $Y2=0
cc_935 N_KAPWR_c_1355_n N_X_c_1589_n 0.00245411f $X=8.91 $Y=2.21 $X2=0 $Y2=0
cc_936 N_KAPWR_c_1358_n N_X_c_1589_n 0.00466059f $X=9.48 $Y=2.21 $X2=0 $Y2=0
cc_937 N_KAPWR_M1021_d N_X_c_1599_n 0.00325489f $X=9.48 $Y=1.485 $X2=0 $Y2=0
cc_938 N_KAPWR_c_1356_n N_X_c_1599_n 0.0128604f $X=9.625 $Y=2.21 $X2=0 $Y2=0
cc_939 N_KAPWR_c_1358_n N_X_c_1599_n 0.00497471f $X=9.48 $Y=2.21 $X2=0 $Y2=0
cc_940 N_KAPWR_c_1360_n N_X_c_1599_n 0.00245411f $X=9.77 $Y=2.21 $X2=0 $Y2=0
cc_941 N_KAPWR_c_1363_n N_X_c_1599_n 0.00466059f $X=10.335 $Y=2.21 $X2=0 $Y2=0
cc_942 N_KAPWR_M1031_d N_X_c_1610_n 0.00316145f $X=10.34 $Y=1.485 $X2=0 $Y2=0
cc_943 N_KAPWR_c_1361_n N_X_c_1610_n 0.012473f $X=10.48 $Y=2.21 $X2=0 $Y2=0
cc_944 N_KAPWR_c_1363_n N_X_c_1610_n 0.00481765f $X=10.335 $Y=2.21 $X2=0 $Y2=0
cc_945 N_KAPWR_c_1365_n N_X_c_1610_n 0.00295229f $X=10.625 $Y=2.21 $X2=0 $Y2=0
cc_946 N_KAPWR_c_1369_n N_X_c_1610_n 0.00435093f $X=11.195 $Y=2.21 $X2=0 $Y2=0
cc_947 N_KAPWR_M1035_d N_X_c_1620_n 0.00325489f $X=11.195 $Y=1.485 $X2=0 $Y2=0
cc_948 N_KAPWR_c_1367_n N_X_c_1620_n 0.0128604f $X=11.34 $Y=2.21 $X2=0 $Y2=0
cc_949 N_KAPWR_c_1369_n N_X_c_1620_n 0.00536178f $X=11.195 $Y=2.21 $X2=0 $Y2=0
cc_950 N_KAPWR_c_1371_n N_X_c_1620_n 0.00300711f $X=11.485 $Y=2.21 $X2=0 $Y2=0
cc_951 N_KAPWR_c_1374_n N_X_c_1620_n 0.00435093f $X=12.05 $Y=2.21 $X2=0 $Y2=0
cc_952 N_KAPWR_M1040_d N_X_c_1630_n 0.00325489f $X=12.055 $Y=1.485 $X2=0 $Y2=0
cc_953 N_KAPWR_c_1372_n N_X_c_1630_n 0.0128604f $X=12.195 $Y=2.21 $X2=0 $Y2=0
cc_954 N_KAPWR_c_1374_n N_X_c_1630_n 0.00520471f $X=12.05 $Y=2.21 $X2=0 $Y2=0
cc_955 N_KAPWR_c_1376_n N_X_c_1630_n 0.00298967f $X=12.34 $Y=2.21 $X2=0 $Y2=0
cc_956 N_KAPWR_c_1381_n N_X_c_1630_n 0.004508f $X=12.9 $Y=2.21 $X2=0 $Y2=0
cc_957 N_KAPWR_c_1345_n N_X_c_1640_n 2.66244e-19 $X=7.18 $Y=2.21 $X2=0 $Y2=0
cc_958 N_KAPWR_c_1346_n N_X_c_1640_n 0.00825548f $X=7.885 $Y=2.21 $X2=0 $Y2=0
cc_959 N_KAPWR_c_1348_n N_X_c_1640_n 0.0230251f $X=7.74 $Y=2.21 $X2=0 $Y2=0
cc_960 N_KAPWR_c_1350_n N_X_c_1640_n 6.89844e-19 $X=8.03 $Y=2.21 $X2=0 $Y2=0
cc_961 N_KAPWR_c_1335_n N_X_c_1640_n 0.0296427f $X=7.04 $Y=1.66 $X2=0 $Y2=0
cc_962 N_KAPWR_c_1346_n N_X_c_1646_n 0.0082718f $X=7.885 $Y=2.21 $X2=0 $Y2=0
cc_963 N_KAPWR_c_1350_n N_X_c_1646_n 4.70067e-19 $X=8.03 $Y=2.21 $X2=0 $Y2=0
cc_964 N_KAPWR_c_1351_n N_X_c_1646_n 0.00822181f $X=8.765 $Y=2.21 $X2=0 $Y2=0
cc_965 N_KAPWR_c_1353_n N_X_c_1646_n 0.0260214f $X=8.62 $Y=2.21 $X2=0 $Y2=0
cc_966 N_KAPWR_c_1355_n N_X_c_1646_n 0.00175189f $X=8.91 $Y=2.21 $X2=0 $Y2=0
cc_967 N_KAPWR_c_1351_n N_X_c_1652_n 0.00822181f $X=8.765 $Y=2.21 $X2=0 $Y2=0
cc_968 N_KAPWR_c_1355_n N_X_c_1652_n 0.00153797f $X=8.91 $Y=2.21 $X2=0 $Y2=0
cc_969 N_KAPWR_c_1356_n N_X_c_1652_n 0.00822181f $X=9.625 $Y=2.21 $X2=0 $Y2=0
cc_970 N_KAPWR_c_1358_n N_X_c_1652_n 0.0260313f $X=9.48 $Y=2.21 $X2=0 $Y2=0
cc_971 N_KAPWR_c_1360_n N_X_c_1652_n 0.00175189f $X=9.77 $Y=2.21 $X2=0 $Y2=0
cc_972 N_KAPWR_c_1356_n N_X_c_1659_n 0.00822181f $X=9.625 $Y=2.21 $X2=0 $Y2=0
cc_973 N_KAPWR_c_1360_n N_X_c_1659_n 0.00153797f $X=9.77 $Y=2.21 $X2=0 $Y2=0
cc_974 N_KAPWR_c_1361_n N_X_c_1659_n 0.00821313f $X=10.48 $Y=2.21 $X2=0 $Y2=0
cc_975 N_KAPWR_c_1363_n N_X_c_1659_n 0.0260313f $X=10.335 $Y=2.21 $X2=0 $Y2=0
cc_976 N_KAPWR_c_1365_n N_X_c_1659_n 0.00152822f $X=10.625 $Y=2.21 $X2=0 $Y2=0
cc_977 N_KAPWR_c_1361_n N_X_c_1666_n 0.0178876f $X=10.48 $Y=2.21 $X2=0 $Y2=0
cc_978 N_KAPWR_c_1365_n N_X_c_1666_n 0.00155772f $X=10.625 $Y=2.21 $X2=0 $Y2=0
cc_979 N_KAPWR_c_1367_n N_X_c_1666_n 0.00755072f $X=11.34 $Y=2.21 $X2=0 $Y2=0
cc_980 N_KAPWR_c_1369_n N_X_c_1666_n 0.0261776f $X=11.195 $Y=2.21 $X2=0 $Y2=0
cc_981 N_KAPWR_c_1371_n N_X_c_1666_n 0.00174799f $X=11.485 $Y=2.21 $X2=0 $Y2=0
cc_982 N_KAPWR_c_1367_n N_X_c_1672_n 0.0178876f $X=11.34 $Y=2.21 $X2=0 $Y2=0
cc_983 N_KAPWR_c_1371_n N_X_c_1672_n 0.00155772f $X=11.485 $Y=2.21 $X2=0 $Y2=0
cc_984 N_KAPWR_c_1372_n N_X_c_1672_n 0.00755072f $X=12.195 $Y=2.21 $X2=0 $Y2=0
cc_985 N_KAPWR_c_1374_n N_X_c_1672_n 0.0261776f $X=12.05 $Y=2.21 $X2=0 $Y2=0
cc_986 N_KAPWR_c_1376_n N_X_c_1672_n 0.00152454f $X=12.34 $Y=2.21 $X2=0 $Y2=0
cc_987 N_KAPWR_M1044_d N_X_c_1567_n 0.00181589f $X=12.915 $Y=1.485 $X2=0 $Y2=0
cc_988 N_KAPWR_M1048_d N_X_c_1567_n 0.00325733f $X=13.775 $Y=1.485 $X2=0 $Y2=0
cc_989 N_KAPWR_c_1304_n N_X_c_1567_n 0.043721f $X=13.78 $Y=2.24 $X2=0 $Y2=0
cc_990 N_KAPWR_c_1372_n N_X_c_1567_n 0.0178903f $X=12.195 $Y=2.21 $X2=0 $Y2=0
cc_991 N_KAPWR_c_1376_n N_X_c_1567_n 6.89749e-19 $X=12.34 $Y=2.21 $X2=0 $Y2=0
cc_992 N_KAPWR_c_1378_n N_X_c_1567_n 0.0286954f $X=13.045 $Y=2.21 $X2=0 $Y2=0
cc_993 N_KAPWR_c_1381_n N_X_c_1567_n 0.0309849f $X=12.9 $Y=2.21 $X2=0 $Y2=0
cc_994 N_KAPWR_c_1383_n N_X_c_1567_n 0.00521589f $X=13.19 $Y=2.21 $X2=0 $Y2=0
cc_995 N_KAPWR_c_1306_n N_X_c_1567_n 0.0456665f $X=13.925 $Y=2.21 $X2=0 $Y2=0
cc_996 N_X_c_1544_n N_VGND_c_1852_n 0.0164628f $X=8.2 $Y=0.82 $X2=0 $Y2=0
cc_997 N_X_c_1547_n N_VGND_c_1853_n 0.0164628f $X=9.06 $Y=0.82 $X2=0 $Y2=0
cc_998 N_X_c_1549_n N_VGND_c_1854_n 0.015936f $X=9.905 $Y=0.82 $X2=0 $Y2=0
cc_999 N_X_c_1549_n N_VGND_c_1855_n 0.00226107f $X=9.905 $Y=0.82 $X2=0 $Y2=0
cc_1000 N_X_c_1550_n N_VGND_c_1855_n 0.0133875f $X=10.05 $Y=0.445 $X2=0 $Y2=0
cc_1001 N_X_c_1551_n N_VGND_c_1855_n 0.00224999f $X=10.765 $Y=0.82 $X2=0 $Y2=0
cc_1002 N_X_c_1551_n N_VGND_c_1856_n 0.015713f $X=10.765 $Y=0.82 $X2=0 $Y2=0
cc_1003 N_X_c_1551_n N_VGND_c_1857_n 0.00225184f $X=10.765 $Y=0.82 $X2=0 $Y2=0
cc_1004 N_X_c_1552_n N_VGND_c_1857_n 0.0128416f $X=10.905 $Y=0.445 $X2=0 $Y2=0
cc_1005 N_X_c_1553_n N_VGND_c_1857_n 0.00239951f $X=11.625 $Y=0.82 $X2=0 $Y2=0
cc_1006 N_X_c_1553_n N_VGND_c_1858_n 0.0161116f $X=11.625 $Y=0.82 $X2=0 $Y2=0
cc_1007 N_X_c_1555_n N_VGND_c_1859_n 0.0161116f $X=12.485 $Y=0.82 $X2=0 $Y2=0
cc_1008 X N_VGND_c_1860_n 0.0186728f $X=13.025 $Y=0.765 $X2=0 $Y2=0
cc_1009 X N_VGND_c_1862_n 0.0243436f $X=13.025 $Y=0.765 $X2=0 $Y2=0
cc_1010 N_X_c_1543_n N_VGND_c_1871_n 0.0128416f $X=7.47 $Y=0.445 $X2=0 $Y2=0
cc_1011 N_X_c_1544_n N_VGND_c_1871_n 0.00224999f $X=8.2 $Y=0.82 $X2=0 $Y2=0
cc_1012 N_X_c_1544_n N_VGND_c_1873_n 0.00224999f $X=8.2 $Y=0.82 $X2=0 $Y2=0
cc_1013 N_X_c_1546_n N_VGND_c_1873_n 0.0128416f $X=8.33 $Y=0.445 $X2=0 $Y2=0
cc_1014 N_X_c_1547_n N_VGND_c_1873_n 0.00224999f $X=9.06 $Y=0.82 $X2=0 $Y2=0
cc_1015 N_X_c_1547_n N_VGND_c_1875_n 0.00224999f $X=9.06 $Y=0.82 $X2=0 $Y2=0
cc_1016 N_X_c_1548_n N_VGND_c_1875_n 0.0128416f $X=9.19 $Y=0.445 $X2=0 $Y2=0
cc_1017 N_X_c_1549_n N_VGND_c_1875_n 0.00224999f $X=9.905 $Y=0.82 $X2=0 $Y2=0
cc_1018 N_X_c_1555_n N_VGND_c_1877_n 0.00225184f $X=12.485 $Y=0.82 $X2=0 $Y2=0
cc_1019 N_X_c_1556_n N_VGND_c_1877_n 0.0128416f $X=12.625 $Y=0.445 $X2=0 $Y2=0
cc_1020 N_X_c_1557_n N_VGND_c_1877_n 0.00232492f $X=12.92 $Y=0.82 $X2=0 $Y2=0
cc_1021 N_X_c_1553_n N_VGND_c_1880_n 0.00225184f $X=11.625 $Y=0.82 $X2=0 $Y2=0
cc_1022 N_X_c_1554_n N_VGND_c_1880_n 0.0128416f $X=11.765 $Y=0.445 $X2=0 $Y2=0
cc_1023 N_X_c_1555_n N_VGND_c_1880_n 0.00239951f $X=12.485 $Y=0.82 $X2=0 $Y2=0
cc_1024 N_X_c_1558_n N_VGND_c_1881_n 0.0129027f $X=13.485 $Y=0.445 $X2=0 $Y2=0
cc_1025 X N_VGND_c_1881_n 0.00498855f $X=13.025 $Y=0.765 $X2=0 $Y2=0
cc_1026 N_X_M1013_d N_VGND_c_1890_n 0.00268444f $X=7.33 $Y=0.235 $X2=0 $Y2=0
cc_1027 N_X_M1016_d N_VGND_c_1890_n 0.00234574f $X=8.19 $Y=0.235 $X2=0 $Y2=0
cc_1028 N_X_M1023_d N_VGND_c_1890_n 0.00234574f $X=9.05 $Y=0.235 $X2=0 $Y2=0
cc_1029 N_X_M1027_d N_VGND_c_1890_n 0.00230304f $X=9.91 $Y=0.235 $X2=0 $Y2=0
cc_1030 N_X_M1046_d N_VGND_c_1890_n 0.00234574f $X=10.765 $Y=0.235 $X2=0 $Y2=0
cc_1031 N_X_M1049_d N_VGND_c_1890_n 0.00234574f $X=11.625 $Y=0.235 $X2=0 $Y2=0
cc_1032 N_X_M1051_d N_VGND_c_1890_n 0.00234574f $X=12.485 $Y=0.235 $X2=0 $Y2=0
cc_1033 N_X_M1056_d N_VGND_c_1890_n 0.00234544f $X=13.345 $Y=0.235 $X2=0 $Y2=0
cc_1034 N_X_c_1543_n N_VGND_c_1890_n 0.00979224f $X=7.47 $Y=0.445 $X2=0 $Y2=0
cc_1035 N_X_c_1544_n N_VGND_c_1890_n 0.00829353f $X=8.2 $Y=0.82 $X2=0 $Y2=0
cc_1036 N_X_c_1546_n N_VGND_c_1890_n 0.00979224f $X=8.33 $Y=0.445 $X2=0 $Y2=0
cc_1037 N_X_c_1547_n N_VGND_c_1890_n 0.00829353f $X=9.06 $Y=0.82 $X2=0 $Y2=0
cc_1038 N_X_c_1548_n N_VGND_c_1890_n 0.00979224f $X=9.19 $Y=0.445 $X2=0 $Y2=0
cc_1039 N_X_c_1549_n N_VGND_c_1890_n 0.0082634f $X=9.905 $Y=0.82 $X2=0 $Y2=0
cc_1040 N_X_c_1550_n N_VGND_c_1890_n 0.0103326f $X=10.05 $Y=0.445 $X2=0 $Y2=0
cc_1041 N_X_c_1551_n N_VGND_c_1890_n 0.00823851f $X=10.765 $Y=0.82 $X2=0 $Y2=0
cc_1042 N_X_c_1552_n N_VGND_c_1890_n 0.00979224f $X=10.905 $Y=0.445 $X2=0 $Y2=0
cc_1043 N_X_c_1553_n N_VGND_c_1890_n 0.00851943f $X=11.625 $Y=0.82 $X2=0 $Y2=0
cc_1044 N_X_c_1554_n N_VGND_c_1890_n 0.00979224f $X=11.765 $Y=0.445 $X2=0 $Y2=0
cc_1045 N_X_c_1555_n N_VGND_c_1890_n 0.00851943f $X=12.485 $Y=0.82 $X2=0 $Y2=0
cc_1046 N_X_c_1556_n N_VGND_c_1890_n 0.00979224f $X=12.625 $Y=0.445 $X2=0 $Y2=0
cc_1047 N_X_c_1557_n N_VGND_c_1890_n 0.00379347f $X=12.92 $Y=0.82 $X2=0 $Y2=0
cc_1048 N_X_c_1558_n N_VGND_c_1890_n 0.00981584f $X=13.485 $Y=0.445 $X2=0 $Y2=0
cc_1049 X N_VGND_c_1890_n 0.0103915f $X=13.025 $Y=0.765 $X2=0 $Y2=0

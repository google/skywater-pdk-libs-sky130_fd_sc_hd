# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.995000 1.240000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 0.265000 1.770000 0.735000 ;
        RECT 1.440000 0.735000 3.135000 0.905000 ;
        RECT 1.440000 1.835000 2.610000 2.005000 ;
        RECT 1.440000 2.005000 1.770000 2.465000 ;
        RECT 2.280000 0.265000 2.610000 0.735000 ;
        RECT 2.280000 1.495000 3.135000 1.665000 ;
        RECT 2.280000 1.665000 2.610000 1.835000 ;
        RECT 2.280000 2.005000 2.610000 2.465000 ;
        RECT 2.790000 0.905000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.595000 ;
      RECT 0.155000  1.495000 1.615000 1.665000 ;
      RECT 0.155000  1.665000 0.515000 2.465000 ;
      RECT 0.515000  0.290000 0.845000 0.825000 ;
      RECT 0.515000  0.825000 0.695000 1.495000 ;
      RECT 1.060000  0.085000 1.230000 0.825000 ;
      RECT 1.060000  1.835000 1.230000 2.635000 ;
      RECT 1.410000  1.075000 2.620000 1.245000 ;
      RECT 1.410000  1.245000 1.615000 1.495000 ;
      RECT 1.940000  0.085000 2.110000 0.565000 ;
      RECT 1.940000  2.175000 2.110000 2.635000 ;
      RECT 2.780000  0.085000 2.950000 0.565000 ;
      RECT 2.780000  1.835000 2.950000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_4
END LIBRARY

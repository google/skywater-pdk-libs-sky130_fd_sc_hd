* File: sky130_fd_sc_hd__ha_1.pex.spice
* Created: Thu Aug 27 14:21:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__HA_1%A_79_21# 1 2 7 9 12 14 17 20 22 23 24 28 30 31
c68 17 0 1.6846e-19 $X=0.655 $Y=1.16
r69 31 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.595 $Y=2.02
+ $X2=1.595 $Y2=2.19
r70 25 28 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=0.51
+ $X2=1.2 $Y2=0.51
r71 23 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=2.02
+ $X2=1.595 $Y2=2.02
r72 23 24 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.51 $Y=2.02
+ $X2=1.13 $Y2=2.02
r73 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.045 $Y=1.935
+ $X2=1.13 $Y2=2.02
r74 21 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=1.245
+ $X2=1.045 $Y2=1.16
r75 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.045 $Y=1.245
+ $X2=1.045 $Y2=1.935
r76 20 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=1.075
+ $X2=1.045 $Y2=1.16
r77 19 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.675
+ $X2=1.045 $Y2=0.51
r78 19 20 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.045 $Y=0.675
+ $X2=1.045 $Y2=1.075
r79 17 36 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.47 $Y2=1.16
r80 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.655
+ $Y=1.16 $X2=0.655 $Y2=1.16
r81 14 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=1.16
+ $X2=1.045 $Y2=1.16
r82 14 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.96 $Y=1.16
+ $X2=0.655 $Y2=1.16
r83 10 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r84 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r85 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r86 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
r87 2 34 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=2.065 $X2=1.595 $Y2=2.19
r88 1 28 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%A_250_199# 1 2 9 13 17 20 22 26 28 32 34 35 36
+ 37 38 42 44 50 54
c131 44 0 1.73601e-19 $X=3.085 $Y=0.8
c132 38 0 1.6846e-19 $X=1.385 $Y=1.06
r133 50 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.16
+ $X2=4.075 $Y2=1.325
r134 50 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.16
+ $X2=4.075 $Y2=0.995
r135 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.075
+ $Y=1.16 $X2=4.075 $Y2=1.16
r136 47 49 17.3597 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=3.997 $Y=0.8
+ $X2=3.997 $Y2=1.16
r137 44 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.085 $Y=0.8
+ $X2=3.085 $Y2=1.06
r138 42 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.385 $Y2=0.995
r139 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=1.16 $X2=1.385 $Y2=1.16
r140 38 41 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.385 $Y=1.06
+ $X2=1.385 $Y2=1.16
r141 36 49 9.27442 $w=2.53e-07 $l=1.99825e-07 $layer=LI1_cond $X=3.92 $Y=1.325
+ $X2=3.997 $Y2=1.16
r142 36 37 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.92 $Y=1.325
+ $X2=3.92 $Y2=1.785
r143 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.835 $Y=1.87
+ $X2=3.92 $Y2=1.785
r144 34 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.835 $Y=1.87
+ $X2=3.52 $Y2=1.87
r145 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.435 $Y=1.955
+ $X2=3.52 $Y2=1.87
r146 30 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.435 $Y=1.955
+ $X2=3.435 $Y2=2.19
r147 29 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=0.8
+ $X2=3.085 $Y2=0.8
r148 28 47 3.06467 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=3.835 $Y=0.8
+ $X2=3.997 $Y2=0.8
r149 28 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.835 $Y=0.8
+ $X2=3.17 $Y2=0.8
r150 24 44 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.715
+ $X2=3.085 $Y2=0.8
r151 24 26 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.085 $Y=0.715
+ $X2=3.085 $Y2=0.51
r152 23 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.47 $Y=1.06
+ $X2=1.385 $Y2=1.06
r153 22 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=1.06 $X2=3.085
+ $Y2=1.06
r154 22 23 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=3 $Y=1.06 $X2=1.47
+ $Y2=1.06
r155 20 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.13 $Y=1.985
+ $X2=4.13 $Y2=1.325
r156 17 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.56
+ $X2=4.13 $Y2=0.995
r157 13 52 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.41 $Y=0.445
+ $X2=1.41 $Y2=0.995
r158 7 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.16
r159 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=2.275
r160 2 32 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=2.065 $X2=3.435 $Y2=2.19
r161 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.085 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%B 3 7 10 13 15 17 20 22 23 24 31 37 38 46
c84 20 0 6.7589e-20 $X=3.295 $Y=0.81
c85 15 0 1.68655e-19 $X=3.295 $Y=0.735
r86 44 46 1.70033 $w=3.03e-07 $l=4.5e-08 $layer=LI1_cond $X=2.002 $Y=1.825
+ $X2=2.002 $Y2=1.87
r87 36 38 10.6716 $w=2.71e-07 $l=6e-08 $layer=POLY_cond $X=3 $Y=1.75 $X2=3.06
+ $Y2=1.75
r88 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=1.74
+ $X2=3 $Y2=1.74
r89 31 34 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=1.66 $X2=1.9
+ $Y2=1.825
r90 31 33 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=1.66 $X2=1.9
+ $Y2=1.495
r91 23 40 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.002 $Y=1.74
+ $X2=2.002 $Y2=1.655
r92 23 44 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.002 $Y=1.74
+ $X2=2.002 $Y2=1.825
r93 23 37 45.0626 $w=2.08e-07 $l=8.45e-07 $layer=LI1_cond $X=2.155 $Y=1.74 $X2=3
+ $Y2=1.74
r94 23 24 12.0912 $w=3.03e-07 $l=3.2e-07 $layer=LI1_cond $X=2.002 $Y=1.89
+ $X2=2.002 $Y2=2.21
r95 23 46 0.7557 $w=3.03e-07 $l=2e-08 $layer=LI1_cond $X=2.002 $Y=1.89 $X2=2.002
+ $Y2=1.87
r96 23 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.66 $X2=1.935 $Y2=1.66
r97 22 40 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=2.002 $Y=1.53
+ $X2=2.002 $Y2=1.655
r98 18 20 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.06 $Y=0.81
+ $X2=3.295 $Y2=0.81
r99 15 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.295 $Y=0.735
+ $X2=3.295 $Y2=0.81
r100 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.295 $Y=0.735
+ $X2=3.295 $Y2=0.445
r101 11 38 27.5683 $w=2.71e-07 $l=2.40312e-07 $layer=POLY_cond $X=3.215 $Y=1.925
+ $X2=3.06 $Y2=1.75
r102 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.215 $Y=1.925
+ $X2=3.215 $Y2=2.275
r103 10 38 16.5906 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.06 $Y=1.575
+ $X2=3.06 $Y2=1.75
r104 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.06 $Y=0.885
+ $X2=3.06 $Y2=0.81
r105 9 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.06 $Y=0.885
+ $X2=3.06 $Y2=1.575
r106 7 33 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.83 $Y=0.445
+ $X2=1.83 $Y2=1.495
r107 3 34 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.805 $Y=2.275
+ $X2=1.805 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%A 3 5 7 11 15 17 18 29
c81 17 0 6.7589e-20 $X=3.445 $Y=1.19
c82 15 0 5.82564e-20 $X=3.655 $Y=2.275
c83 5 0 4.94663e-21 $X=2.355 $Y=1.565
r84 26 29 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.48 $Y=1.32
+ $X2=3.655 $Y2=1.32
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.48
+ $Y=1.32 $X2=3.48 $Y2=1.32
r86 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5 $Y=1.4
+ $X2=2.5 $Y2=1.4
r87 18 27 4.09758 $w=2.23e-07 $l=8e-08 $layer=LI1_cond $X=3.472 $Y=1.4 $X2=3.472
+ $Y2=1.32
r88 18 24 45.8548 $w=2.08e-07 $l=8.6e-07 $layer=LI1_cond $X=3.36 $Y=1.4 $X2=2.5
+ $Y2=1.4
r89 17 27 6.65856 $w=2.23e-07 $l=1.3e-07 $layer=LI1_cond $X=3.472 $Y=1.19
+ $X2=3.472 $Y2=1.32
r90 13 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.485
+ $X2=3.655 $Y2=1.32
r91 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.655 $Y=1.485
+ $X2=3.655 $Y2=2.275
r92 9 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.155
+ $X2=3.655 $Y2=1.32
r93 9 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.655 $Y=1.155
+ $X2=3.655 $Y2=0.445
r94 5 23 38.7288 $w=3.45e-07 $l=1.87029e-07 $layer=POLY_cond $X=2.355 $Y=1.565
+ $X2=2.402 $Y2=1.4
r95 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.355 $Y=1.565
+ $X2=2.355 $Y2=2.275
r96 1 23 52.6998 $w=3.45e-07 $l=3.32423e-07 $layer=POLY_cond $X=2.25 $Y=1.135
+ $X2=2.402 $Y2=1.4
r97 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.25 $Y=1.135 $X2=2.25
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%SUM 1 2 7 8 9 10 11 12 23 30 36
r20 36 48 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.205 $Y=1.53
+ $X2=0.205 $Y2=1.565
r21 30 46 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.205 $Y=0.85
+ $X2=0.205 $Y2=0.825
r22 12 43 4.12815 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.33
r23 11 12 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=1.87
+ $X2=0.257 $Y2=2.21
r24 11 37 4.74738 $w=3.33e-07 $l=1.38e-07 $layer=LI1_cond $X=0.257 $Y=1.87
+ $X2=0.257 $Y2=1.732
r25 10 37 4.88498 $w=3.33e-07 $l=1.42e-07 $layer=LI1_cond $X=0.257 $Y=1.59
+ $X2=0.257 $Y2=1.732
r26 10 48 2.00123 $w=3.33e-07 $l=2.5e-08 $layer=LI1_cond $X=0.257 $Y=1.59
+ $X2=0.257 $Y2=1.565
r27 10 36 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.205 $Y=1.505
+ $X2=0.205 $Y2=1.53
r28 9 10 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.205 $Y=1.19
+ $X2=0.205 $Y2=1.505
r29 8 46 2.17324 $w=3.33e-07 $l=3e-08 $layer=LI1_cond $X=0.257 $Y=0.795
+ $X2=0.257 $Y2=0.825
r30 8 21 4.71298 $w=3.33e-07 $l=1.37e-07 $layer=LI1_cond $X=0.257 $Y=0.795
+ $X2=0.257 $Y2=0.658
r31 8 9 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.205 $Y=0.88
+ $X2=0.205 $Y2=1.19
r32 8 30 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=0.205 $Y=0.88 $X2=0.205
+ $Y2=0.85
r33 7 21 5.09139 $w=3.33e-07 $l=1.48e-07 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.658
r34 7 23 3.78414 $w=3.33e-07 $l=1.1e-07 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.4
r35 2 10 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
r36 2 43 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.33
r37 1 23 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%VPWR 1 2 3 12 16 18 30 37 38 42 48 52 58 60
r64 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 56 58 8.91451 $w=5.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.99 $Y=2.54
+ $X2=3.12 $Y2=2.54
r66 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 54 56 0.789863 $w=5.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.955 $Y=2.54
+ $X2=2.99 $Y2=2.54
r68 51 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 50 54 9.5912 $w=5.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.53 $Y=2.54
+ $X2=2.955 $Y2=2.54
r70 50 52 7.78613 $w=5.28e-07 $l=8e-08 $layer=LI1_cond $X=2.53 $Y=2.54 $X2=2.45
+ $Y2=2.54
r71 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 46 48 8.46316 $w=5.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.15 $Y=2.54
+ $X2=1.26 $Y2=2.54
r73 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 44 46 1.24121 $w=5.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.095 $Y=2.54
+ $X2=1.15 $Y2=2.54
r75 41 44 9.36552 $w=5.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.54
+ $X2=1.095 $Y2=2.54
r76 41 42 7.89897 $w=5.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.54
+ $X2=0.595 $Y2=2.54
r77 38 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r78 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r79 35 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=3.88 $Y2=2.72
r80 35 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=4.37 $Y2=2.72
r81 34 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r82 34 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 33 58 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.12 $Y2=2.72
r84 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 30 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.88 $Y2=2.72
r86 30 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.45 $Y2=2.72
r87 29 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r88 29 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 28 52 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.45 $Y2=2.72
r90 28 48 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.26 $Y2=2.72
r91 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r92 22 42 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.595 $Y2=2.72
r93 18 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 14 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.72
r96 14 16 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.29
r97 10 41 6.67551 $w=1.95e-07 $l=2.70934e-07 $layer=LI1_cond $X=0.692 $Y=2.275
+ $X2=0.68 $Y2=2.54
r98 10 12 33.8415 $w=1.93e-07 $l=5.95e-07 $layer=LI1_cond $X=0.692 $Y=2.275
+ $X2=0.692 $Y2=1.68
r99 3 16 600 $w=1.7e-07 $l=3.05573e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=2.065 $X2=3.92 $Y2=2.29
r100 2 54 300 $w=1.7e-07 $l=6.56125e-07 $layer=licon1_PDIFF $count=2 $X=2.43
+ $Y=2.065 $X2=2.955 $Y2=2.36
r101 1 44 600 $w=1.7e-07 $l=1.11664e-06 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=1.095 $Y2=2.36
r102 1 41 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.36
r103 1 12 300 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%COUT 1 2 11 12 13 14 15 27
c22 11 0 5.82564e-20 $X=4.34 $Y=1.65
r23 15 24 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=4.345 $Y=2.21
+ $X2=4.345 $Y2=2.33
r24 14 15 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=4.345 $Y=1.87
+ $X2=4.345 $Y2=2.21
r25 13 31 13.0555 $w=3.38e-07 $l=3.15e-07 $layer=LI1_cond $X=4.345 $Y=0.51
+ $X2=4.345 $Y2=0.825
r26 13 27 3.72849 $w=3.38e-07 $l=1.1e-07 $layer=LI1_cond $X=4.345 $Y=0.51
+ $X2=4.345 $Y2=0.4
r27 12 31 44.3636 $w=1.83e-07 $l=7.4e-07 $layer=LI1_cond $X=4.422 $Y=1.565
+ $X2=4.422 $Y2=0.825
r28 11 12 5.25957 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.345 $Y=1.65
+ $X2=4.345 $Y2=1.565
r29 9 14 4.57588 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=4.345 $Y=1.735
+ $X2=4.345 $Y2=1.87
r30 9 11 2.88111 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.345 $Y=1.735
+ $X2=4.345 $Y2=1.65
r31 2 24 400 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.485 $X2=4.34 $Y2=2.33
r32 2 11 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.485 $X2=4.34 $Y2=1.65
r33 1 27 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.205
+ $Y=0.235 $X2=4.34 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%VGND 1 2 3 12 16 20 22 24 29 34 44 45 48 51 54
r70 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r71 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r72 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r73 45 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r74 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r75 42 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=3.88
+ $Y2=0
r76 42 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.37
+ $Y2=0
r77 41 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r78 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r79 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r80 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r81 37 40 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r82 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r83 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r84 35 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.53
+ $Y2=0
r85 34 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.88
+ $Y2=0
r86 34 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.45
+ $Y2=0
r87 33 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r88 33 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r89 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r90 30 48 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.692
+ $Y2=0
r91 30 32 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=1.61
+ $Y2=0
r92 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r93 29 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.61
+ $Y2=0
r94 24 48 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.692
+ $Y2=0
r95 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r96 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r97 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r98 18 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0
r99 18 20 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0.38
r100 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r101 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.38
r102 10 48 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r103 10 12 16.7786 $w=1.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.38
r104 3 20 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.92 $Y2=0.38
r105 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.38
r106 1 12 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__HA_1%A_297_47# 1 2 9 11 12 15
r24 13 15 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.46 $Y=0.635
+ $X2=2.46 $Y2=0.51
r25 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=0.72
+ $X2=2.46 $Y2=0.635
r26 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.375 $Y=0.72
+ $X2=1.705 $Y2=0.72
r27 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=0.635
+ $X2=1.705 $Y2=0.72
r28 7 9 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.62 $Y=0.635
+ $X2=1.62 $Y2=0.51
r29 2 15 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.51
r30 1 9 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends


* File: sky130_fd_sc_hd__or3b_4.pxi.spice
* Created: Tue Sep  1 19:28:14 2020
* 
x_PM_SKY130_FD_SC_HD__OR3B_4%C_N N_C_N_M1013_g N_C_N_M1014_g C_N C_N
+ N_C_N_c_83_n PM_SKY130_FD_SC_HD__OR3B_4%C_N
x_PM_SKY130_FD_SC_HD__OR3B_4%A_176_21# N_A_176_21#_M1009_d N_A_176_21#_M1008_d
+ N_A_176_21#_M1001_d N_A_176_21#_c_109_n N_A_176_21#_M1002_g
+ N_A_176_21#_M1004_g N_A_176_21#_c_110_n N_A_176_21#_M1003_g
+ N_A_176_21#_M1007_g N_A_176_21#_c_111_n N_A_176_21#_M1005_g
+ N_A_176_21#_M1010_g N_A_176_21#_c_112_n N_A_176_21#_M1012_g
+ N_A_176_21#_M1015_g N_A_176_21#_c_113_n N_A_176_21#_c_114_n
+ N_A_176_21#_c_115_n N_A_176_21#_c_133_p N_A_176_21#_c_239_p
+ N_A_176_21#_c_124_n N_A_176_21#_c_116_n N_A_176_21#_c_117_n
+ N_A_176_21#_c_145_p N_A_176_21#_c_148_p N_A_176_21#_c_118_n
+ N_A_176_21#_c_119_n PM_SKY130_FD_SC_HD__OR3B_4%A_176_21#
x_PM_SKY130_FD_SC_HD__OR3B_4%A N_A_c_256_n N_A_M1009_g N_A_M1000_g N_A_c_260_n
+ N_A_c_257_n N_A_c_258_n A PM_SKY130_FD_SC_HD__OR3B_4%A
x_PM_SKY130_FD_SC_HD__OR3B_4%B N_B_M1006_g N_B_M1011_g B B N_B_c_303_n
+ N_B_c_304_n N_B_c_305_n PM_SKY130_FD_SC_HD__OR3B_4%B
x_PM_SKY130_FD_SC_HD__OR3B_4%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1014_s
+ N_A_27_47#_M1008_g N_A_27_47#_M1001_g N_A_27_47#_c_344_n N_A_27_47#_c_345_n
+ N_A_27_47#_c_346_n N_A_27_47#_c_363_n N_A_27_47#_c_347_n N_A_27_47#_c_373_n
+ N_A_27_47#_c_353_n N_A_27_47#_c_354_n N_A_27_47#_c_380_n N_A_27_47#_c_348_n
+ N_A_27_47#_c_349_n N_A_27_47#_c_350_n PM_SKY130_FD_SC_HD__OR3B_4%A_27_47#
x_PM_SKY130_FD_SC_HD__OR3B_4%VPWR N_VPWR_M1014_d N_VPWR_M1007_d N_VPWR_M1015_d
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n VPWR N_VPWR_c_446_n
+ N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_442_n N_VPWR_c_451_n
+ N_VPWR_c_452_n N_VPWR_c_453_n PM_SKY130_FD_SC_HD__OR3B_4%VPWR
x_PM_SKY130_FD_SC_HD__OR3B_4%X N_X_M1002_s N_X_M1005_s N_X_M1004_s N_X_M1010_s
+ N_X_c_508_n N_X_c_513_n N_X_c_509_n N_X_c_530_n N_X_c_510_n N_X_c_537_n
+ N_X_c_538_n X PM_SKY130_FD_SC_HD__OR3B_4%X
x_PM_SKY130_FD_SC_HD__OR3B_4%VGND N_VGND_M1013_d N_VGND_M1003_d N_VGND_M1012_d
+ N_VGND_M1006_d N_VGND_c_581_n N_VGND_c_582_n N_VGND_c_583_n N_VGND_c_584_n
+ N_VGND_c_585_n N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n
+ N_VGND_c_590_n VGND N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n VGND
+ PM_SKY130_FD_SC_HD__OR3B_4%VGND
cc_1 VNB N_C_N_M1013_g 0.0359089f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB C_N 0.00882738f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_83_n 0.0383384f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_176_21#_c_109_n 0.0162946f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_5 VNB N_A_176_21#_c_110_n 0.0157821f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_6 VNB N_A_176_21#_c_111_n 0.0157207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_176_21#_c_112_n 0.0152476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_176_21#_c_113_n 0.00227943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_176_21#_c_114_n 0.00130133f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_176_21#_c_115_n 0.00148375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_176_21#_c_116_n 0.0117914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_176_21#_c_117_n 0.0237879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_176_21#_c_118_n 0.0126408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_176_21#_c_119_n 0.0630913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_c_256_n 0.0161968f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_A_c_257_n 3.07343e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_17 VNB N_A_c_258_n 0.0221445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_c_303_n 0.0203489f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_19 VNB N_B_c_304_n 0.00332839f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_20 VNB N_B_c_305_n 0.0167656f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_21 VNB N_A_27_47#_c_344_n 0.0182298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_345_n 0.0039003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_346_n 0.00930805f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_24 VNB N_A_27_47#_c_347_n 0.006646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_348_n 0.00320906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_349_n 0.0224001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_350_n 0.0199081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_442_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_508_n 8.69458e-19 $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_30 VNB N_X_c_509_n 0.00353053f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_31 VNB N_X_c_510_n 0.0019307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_581_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_33 VNB N_VGND_c_582_n 0.00406558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_583_n 3.15634e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_584_n 3.95773e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_585_n 0.0187422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_586_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_587_n 0.0144207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_588_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_589_n 0.0111699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_590_n 0.00516067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_591_n 0.018223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_592_n 0.219992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_593_n 0.0218393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VPB N_C_N_M1014_g 0.049006f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.01
cc_46 VPB C_N 0.0160532f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_47 VPB N_C_N_c_83_n 0.0100411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_48 VPB N_A_176_21#_M1004_g 0.0202012f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_A_176_21#_M1007_g 0.0176242f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.53
cc_50 VPB N_A_176_21#_M1010_g 0.0176231f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_176_21#_M1015_g 0.0181714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_176_21#_c_124_n 0.0113342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_176_21#_c_117_n 0.0392226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_176_21#_c_119_n 0.0100546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_M1000_g 0.0169429f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.01
cc_56 VPB N_A_c_260_n 0.00283459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_c_257_n 0.00158529f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_58 VPB N_A_c_258_n 0.0046266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B_M1011_g 0.0179256f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.01
cc_60 VPB N_B_c_303_n 0.00468852f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_61 VPB N_B_c_304_n 0.00213983f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_62 VPB N_A_27_47#_M1001_g 0.0230655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_347_n 0.00552293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_353_n 0.00266045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_354_n 0.0187262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_348_n 0.00232434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_349_n 0.0057853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_443_n 0.00980242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_444_n 3.00801e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_445_n 3.94561e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_446_n 0.0172683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_447_n 0.0120084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_448_n 0.0118696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_449_n 0.041841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_442_n 0.0492078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_451_n 0.00565096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_452_n 0.00436419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_453_n 0.00449722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_X_c_508_n 8.69458e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_80 VPB X 0.00631179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 N_C_N_M1013_g N_A_176_21#_c_109_n 0.0187739f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_82 N_C_N_M1014_g N_A_176_21#_M1004_g 0.0187739f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_83 N_C_N_c_83_n N_A_176_21#_c_119_n 0.0187739f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_84 N_C_N_M1013_g N_A_27_47#_c_344_n 0.00239051f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_85 N_C_N_M1013_g N_A_27_47#_c_345_n 0.0170801f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_86 C_N N_A_27_47#_c_345_n 0.0060742f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_87 N_C_N_c_83_n N_A_27_47#_c_345_n 0.0012291f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_88 C_N N_A_27_47#_c_346_n 0.0227094f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_89 N_C_N_c_83_n N_A_27_47#_c_346_n 0.00599978f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_90 N_C_N_M1014_g N_A_27_47#_c_363_n 0.0151922f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_91 C_N N_A_27_47#_c_363_n 0.00445498f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_92 N_C_N_M1013_g N_A_27_47#_c_347_n 0.0130087f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_93 C_N N_A_27_47#_c_347_n 0.042517f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_94 C_N N_A_27_47#_c_354_n 0.0223722f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_95 N_C_N_c_83_n N_A_27_47#_c_354_n 8.87396e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_96 N_C_N_M1014_g N_VPWR_c_443_n 0.00394846f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_97 N_C_N_M1014_g N_VPWR_c_446_n 0.00378081f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_98 N_C_N_M1014_g N_VPWR_c_442_n 0.00502381f $X=0.47 $Y=2.01 $X2=0 $Y2=0
cc_99 N_C_N_M1013_g N_X_c_513_n 5.497e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_100 N_C_N_M1013_g N_VGND_c_581_n 0.00478935f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_101 N_C_N_M1013_g N_VGND_c_592_n 0.00718838f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_102 N_C_N_M1013_g N_VGND_c_593_n 0.00439206f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A_176_21#_c_112_n N_A_c_256_n 0.0240018f $X=2.215 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_176_21#_c_114_n N_A_c_256_n 0.00140826f $X=2.28 $Y=0.89 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_176_21#_c_115_n N_A_c_256_n 0.00207559f $X=2.28 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_106 N_A_176_21#_c_133_p N_A_c_256_n 0.0113009f $X=2.76 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_176_21#_M1015_g N_A_M1000_g 0.0421086f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_176_21#_M1015_g N_A_c_260_n 0.00188155f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_176_21#_c_133_p N_A_c_260_n 0.0038033f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_176_21#_M1015_g N_A_c_257_n 0.00171726f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_176_21#_c_113_n N_A_c_257_n 0.0137913f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_176_21#_c_115_n N_A_c_257_n 0.00571956f $X=2.28 $Y=1.075 $X2=0 $Y2=0
cc_113 N_A_176_21#_c_133_p N_A_c_257_n 0.0122714f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_176_21#_c_119_n N_A_c_257_n 8.25131e-19 $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_176_21#_c_113_n N_A_c_258_n 0.00109316f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_176_21#_c_115_n N_A_c_258_n 4.38315e-19 $X=2.28 $Y=1.075 $X2=0 $Y2=0
cc_117 N_A_176_21#_c_133_p N_A_c_258_n 7.47524e-19 $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_176_21#_c_145_p N_A_c_258_n 2.69871e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A_176_21#_c_119_n N_A_c_258_n 0.0210564f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_176_21#_c_124_n N_B_M1011_g 0.001139f $X=3.85 $Y=2.317 $X2=0 $Y2=0
cc_121 N_A_176_21#_c_148_p N_B_c_303_n 0.00227792f $X=3.66 $Y=0.715 $X2=0 $Y2=0
cc_122 N_A_176_21#_c_145_p N_B_c_304_n 0.00322337f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_176_21#_c_148_p N_B_c_304_n 0.0171667f $X=3.66 $Y=0.715 $X2=0 $Y2=0
cc_124 N_A_176_21#_c_148_p N_B_c_305_n 0.0116387f $X=3.66 $Y=0.715 $X2=0 $Y2=0
cc_125 N_A_176_21#_c_124_n N_A_27_47#_M1001_g 0.00744135f $X=3.85 $Y=2.317 $X2=0
+ $Y2=0
cc_126 N_A_176_21#_c_117_n N_A_27_47#_M1001_g 0.00854324f $X=3.952 $Y=2.21 $X2=0
+ $Y2=0
cc_127 N_A_176_21#_c_109_n N_A_27_47#_c_345_n 0.0013109f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_A_176_21#_c_109_n N_A_27_47#_c_347_n 0.00850451f $X=0.955 $Y=0.995
+ $X2=0 $Y2=0
cc_129 N_A_176_21#_M1004_g N_A_27_47#_c_373_n 0.0135875f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_176_21#_M1007_g N_A_27_47#_c_373_n 0.0116058f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_176_21#_M1010_g N_A_27_47#_c_373_n 0.0116058f $X=1.795 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_176_21#_M1015_g N_A_27_47#_c_373_n 0.0125f $X=2.215 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_176_21#_c_113_n N_A_27_47#_c_373_n 0.00340069f $X=2.195 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_176_21#_c_124_n N_A_27_47#_c_373_n 0.00660479f $X=3.85 $Y=2.317 $X2=0
+ $Y2=0
cc_135 N_A_176_21#_c_117_n N_A_27_47#_c_353_n 0.0215607f $X=3.952 $Y=2.21 $X2=0
+ $Y2=0
cc_136 N_A_176_21#_M1004_g N_A_27_47#_c_380_n 0.00162764f $X=0.955 $Y=1.985
+ $X2=0 $Y2=0
cc_137 N_A_176_21#_c_117_n N_A_27_47#_c_348_n 0.0249158f $X=3.952 $Y=2.21 $X2=0
+ $Y2=0
cc_138 N_A_176_21#_c_148_p N_A_27_47#_c_348_n 0.0181856f $X=3.66 $Y=0.715 $X2=0
+ $Y2=0
cc_139 N_A_176_21#_c_117_n N_A_27_47#_c_349_n 0.00756781f $X=3.952 $Y=2.21 $X2=0
+ $Y2=0
cc_140 N_A_176_21#_c_118_n N_A_27_47#_c_349_n 0.00233368f $X=3.952 $Y=0.715
+ $X2=0 $Y2=0
cc_141 N_A_176_21#_c_117_n N_A_27_47#_c_350_n 0.00550363f $X=3.952 $Y=2.21 $X2=0
+ $Y2=0
cc_142 N_A_176_21#_c_148_p N_A_27_47#_c_350_n 0.0133375f $X=3.66 $Y=0.715 $X2=0
+ $Y2=0
cc_143 N_A_176_21#_M1004_g N_VPWR_c_443_n 0.0100525f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_176_21#_M1007_g N_VPWR_c_443_n 0.00123638f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_176_21#_M1004_g N_VPWR_c_444_n 0.00123489f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_176_21#_M1007_g N_VPWR_c_444_n 0.00889313f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_176_21#_M1010_g N_VPWR_c_444_n 0.00885947f $X=1.795 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_176_21#_M1015_g N_VPWR_c_444_n 0.00123111f $X=2.215 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_176_21#_M1010_g N_VPWR_c_445_n 0.00124518f $X=1.795 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_176_21#_M1015_g N_VPWR_c_445_n 0.00912635f $X=2.215 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_176_21#_M1004_g N_VPWR_c_447_n 0.00344532f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_176_21#_M1007_g N_VPWR_c_447_n 0.00344532f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_176_21#_M1010_g N_VPWR_c_448_n 0.00344532f $X=1.795 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_176_21#_M1015_g N_VPWR_c_448_n 0.00330146f $X=2.215 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_176_21#_c_124_n N_VPWR_c_449_n 0.0270932f $X=3.85 $Y=2.317 $X2=0
+ $Y2=0
cc_156 N_A_176_21#_M1001_d N_VPWR_c_442_n 0.00211645f $X=3.61 $Y=1.485 $X2=0
+ $Y2=0
cc_157 N_A_176_21#_M1004_g N_VPWR_c_442_n 0.00407565f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_176_21#_M1007_g N_VPWR_c_442_n 0.00407565f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_176_21#_M1010_g N_VPWR_c_442_n 0.00407565f $X=1.795 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_176_21#_M1015_g N_VPWR_c_442_n 0.00392934f $X=2.215 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_176_21#_c_124_n N_VPWR_c_442_n 0.0192963f $X=3.85 $Y=2.317 $X2=0
+ $Y2=0
cc_162 N_A_176_21#_c_109_n N_X_c_508_n 0.00176417f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_176_21#_M1004_g N_X_c_508_n 0.00176417f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_176_21#_c_110_n N_X_c_508_n 0.00177623f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_176_21#_M1007_g N_X_c_508_n 0.00177623f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_176_21#_c_113_n N_X_c_508_n 0.0127974f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_176_21#_c_119_n N_X_c_508_n 0.0166904f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_176_21#_c_109_n N_X_c_513_n 0.00687212f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_176_21#_c_110_n N_X_c_513_n 0.00618135f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_176_21#_c_111_n N_X_c_513_n 5.19613e-19 $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_176_21#_c_110_n N_X_c_509_n 0.00845772f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_176_21#_c_111_n N_X_c_509_n 0.0109841f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_176_21#_c_112_n N_X_c_509_n 0.00119027f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_176_21#_c_113_n N_X_c_509_n 0.0501269f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_176_21#_c_114_n N_X_c_509_n 0.0130974f $X=2.28 $Y=0.89 $X2=0 $Y2=0
cc_176 N_A_176_21#_c_115_n N_X_c_509_n 0.00117611f $X=2.28 $Y=1.075 $X2=0 $Y2=0
cc_177 N_A_176_21#_c_119_n N_X_c_509_n 0.00388181f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_176_21#_c_111_n N_X_c_530_n 0.00333989f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_176_21#_c_112_n N_X_c_530_n 0.00194172f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_176_21#_c_114_n N_X_c_530_n 0.00525339f $X=2.28 $Y=0.89 $X2=0 $Y2=0
cc_181 N_A_176_21#_c_109_n N_X_c_510_n 0.00440045f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_176_21#_c_110_n N_X_c_510_n 0.0011047f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_176_21#_c_113_n N_X_c_510_n 0.00426971f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_176_21#_c_119_n N_X_c_510_n 0.00279996f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_176_21#_M1004_g N_X_c_537_n 0.00639858f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_176_21#_c_110_n N_X_c_538_n 5.20925e-19 $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_176_21#_c_111_n N_X_c_538_n 0.00346461f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_176_21#_c_113_n N_X_c_538_n 0.00198266f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_176_21#_c_119_n N_X_c_538_n 4.98263e-19 $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_176_21#_M1007_g X 0.0122249f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_176_21#_M1010_g X 0.0122249f $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_176_21#_M1015_g X 0.00698802f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_176_21#_c_113_n X 0.0690662f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_176_21#_c_119_n X 0.00715867f $X=2.215 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_176_21#_c_114_n N_VGND_M1012_d 0.00126113f $X=2.28 $Y=0.89 $X2=0
+ $Y2=0
cc_196 N_A_176_21#_c_133_p N_VGND_M1012_d 0.00300025f $X=2.76 $Y=0.74 $X2=0
+ $Y2=0
cc_197 N_A_176_21#_c_148_p N_VGND_M1006_d 0.0084162f $X=3.66 $Y=0.715 $X2=0
+ $Y2=0
cc_198 N_A_176_21#_c_109_n N_VGND_c_581_n 0.00434912f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_176_21#_c_110_n N_VGND_c_582_n 0.00268723f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_176_21#_c_111_n N_VGND_c_582_n 0.00137415f $X=1.795 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_176_21#_c_111_n N_VGND_c_583_n 4.79856e-19 $X=1.795 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_176_21#_c_112_n N_VGND_c_583_n 0.0070037f $X=2.215 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_176_21#_c_114_n N_VGND_c_583_n 0.00651354f $X=2.28 $Y=0.89 $X2=0
+ $Y2=0
cc_204 N_A_176_21#_c_133_p N_VGND_c_583_n 0.0099168f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_176_21#_c_148_p N_VGND_c_584_n 0.0206674f $X=3.66 $Y=0.715 $X2=0
+ $Y2=0
cc_206 N_A_176_21#_c_109_n N_VGND_c_585_n 0.00479157f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_176_21#_c_110_n N_VGND_c_585_n 0.00425617f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_176_21#_c_111_n N_VGND_c_587_n 0.0043257f $X=1.795 $Y=0.995 $X2=0
+ $Y2=0
cc_209 N_A_176_21#_c_112_n N_VGND_c_587_n 0.00402685f $X=2.215 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_176_21#_c_114_n N_VGND_c_587_n 9.65875e-19 $X=2.28 $Y=0.89 $X2=0
+ $Y2=0
cc_211 N_A_176_21#_c_133_p N_VGND_c_589_n 0.00232396f $X=2.76 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_176_21#_c_239_p N_VGND_c_589_n 0.00846569f $X=2.845 $Y=0.47 $X2=0
+ $Y2=0
cc_213 N_A_176_21#_c_148_p N_VGND_c_589_n 0.00232396f $X=3.66 $Y=0.715 $X2=0
+ $Y2=0
cc_214 N_A_176_21#_c_116_n N_VGND_c_591_n 0.0126179f $X=3.745 $Y=0.47 $X2=0
+ $Y2=0
cc_215 N_A_176_21#_c_148_p N_VGND_c_591_n 0.00232396f $X=3.66 $Y=0.715 $X2=0
+ $Y2=0
cc_216 N_A_176_21#_c_118_n N_VGND_c_591_n 0.00281072f $X=3.952 $Y=0.715 $X2=0
+ $Y2=0
cc_217 N_A_176_21#_M1009_d N_VGND_c_592_n 0.00256656f $X=2.71 $Y=0.235 $X2=0
+ $Y2=0
cc_218 N_A_176_21#_M1008_d N_VGND_c_592_n 0.00231589f $X=3.61 $Y=0.235 $X2=0
+ $Y2=0
cc_219 N_A_176_21#_c_109_n N_VGND_c_592_n 0.00770375f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_176_21#_c_110_n N_VGND_c_592_n 0.00573783f $X=1.375 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_176_21#_c_111_n N_VGND_c_592_n 0.00582201f $X=1.795 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_176_21#_c_112_n N_VGND_c_592_n 0.00579963f $X=2.215 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_176_21#_c_114_n N_VGND_c_592_n 0.00217608f $X=2.28 $Y=0.89 $X2=0
+ $Y2=0
cc_224 N_A_176_21#_c_133_p N_VGND_c_592_n 0.00495795f $X=2.76 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_176_21#_c_239_p N_VGND_c_592_n 0.00625722f $X=2.845 $Y=0.47 $X2=0
+ $Y2=0
cc_226 N_A_176_21#_c_116_n N_VGND_c_592_n 0.00927792f $X=3.745 $Y=0.47 $X2=0
+ $Y2=0
cc_227 N_A_176_21#_c_148_p N_VGND_c_592_n 0.00996249f $X=3.66 $Y=0.715 $X2=0
+ $Y2=0
cc_228 N_A_176_21#_c_118_n N_VGND_c_592_n 0.0041615f $X=3.952 $Y=0.715 $X2=0
+ $Y2=0
cc_229 N_A_M1000_g N_B_M1011_g 0.0628571f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_c_260_n N_B_M1011_g 3.36535e-19 $X=2.627 $Y=1.415 $X2=0 $Y2=0
cc_231 N_A_c_257_n N_B_M1011_g 2.29135e-19 $X=2.635 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_c_257_n N_B_c_303_n 3.21144e-19 $X=2.635 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_c_258_n N_B_c_303_n 0.0201765f $X=2.635 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_M1000_g N_B_c_304_n 0.00125605f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_c_260_n N_B_c_304_n 0.0142283f $X=2.627 $Y=1.415 $X2=0 $Y2=0
cc_236 N_A_c_257_n N_B_c_304_n 0.0320748f $X=2.635 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_c_258_n N_B_c_304_n 0.00199269f $X=2.635 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_c_256_n N_B_c_305_n 0.0243978f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_M1000_g N_A_27_47#_c_373_n 0.0114643f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_c_260_n N_A_27_47#_c_373_n 0.0183689f $X=2.627 $Y=1.415 $X2=0 $Y2=0
cc_241 N_A_c_258_n N_A_27_47#_c_373_n 7.32583e-19 $X=2.635 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_c_260_n N_VPWR_M1015_d 0.00294065f $X=2.627 $Y=1.415 $X2=0 $Y2=0
cc_243 N_A_M1000_g N_VPWR_c_445_n 0.0106753f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A_M1000_g N_VPWR_c_449_n 0.00330146f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_M1000_g N_VPWR_c_442_n 0.00395759f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A_M1000_g X 2.48221e-19 $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_c_260_n X 0.0224672f $X=2.627 $Y=1.415 $X2=0 $Y2=0
cc_248 N_A_c_256_n N_VGND_c_583_n 0.00716819f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_c_256_n N_VGND_c_584_n 6.25182e-19 $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_c_256_n N_VGND_c_589_n 0.00341689f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_256_n N_VGND_c_592_n 0.00405445f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B_M1011_g N_A_27_47#_M1001_g 0.049098f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_253 N_B_c_304_n N_A_27_47#_M1001_g 0.00118139f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B_M1011_g N_A_27_47#_c_373_n 0.0121815f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B_c_303_n N_A_27_47#_c_373_n 0.00145405f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B_c_304_n N_A_27_47#_c_373_n 0.0150515f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B_M1011_g N_A_27_47#_c_353_n 0.00452731f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B_c_303_n N_A_27_47#_c_348_n 0.00199358f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B_c_304_n N_A_27_47#_c_348_n 0.050953f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B_c_303_n N_A_27_47#_c_349_n 0.0202262f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B_c_304_n N_A_27_47#_c_349_n 3.34918e-19 $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_262 N_B_c_305_n N_A_27_47#_c_350_n 0.0203981f $X=3.115 $Y=0.995 $X2=0 $Y2=0
cc_263 N_B_M1011_g N_VPWR_c_445_n 0.00242481f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_264 N_B_M1011_g N_VPWR_c_449_n 0.00431606f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B_M1011_g N_VPWR_c_442_n 0.00618933f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_266 N_B_c_304_n A_542_297# 0.00218202f $X=3.115 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_267 N_B_c_304_n A_626_297# 0.00211207f $X=3.115 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_268 N_B_c_305_n N_VGND_c_583_n 6.21849e-19 $X=3.115 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B_c_305_n N_VGND_c_584_n 0.0074276f $X=3.115 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B_c_305_n N_VGND_c_589_n 0.00341689f $X=3.115 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B_c_305_n N_VGND_c_592_n 0.00405445f $X=3.115 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_347_n N_VPWR_M1014_d 0.00417312f $X=0.68 $Y=1.81 $X2=-0.19
+ $Y2=-0.24
cc_273 N_A_27_47#_c_373_n N_VPWR_M1014_d 0.00276232f $X=3.39 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_274 N_A_27_47#_c_380_n N_VPWR_M1014_d 0.0024773f $X=0.68 $Y=1.925 $X2=-0.19
+ $Y2=-0.24
cc_275 N_A_27_47#_c_373_n N_VPWR_M1007_d 0.00317505f $X=3.39 $Y=1.955 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_373_n N_VPWR_M1015_d 0.00437469f $X=3.39 $Y=1.955 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_373_n N_VPWR_c_443_n 0.0065098f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_380_n N_VPWR_c_443_n 0.0138837f $X=0.68 $Y=1.925 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_373_n N_VPWR_c_444_n 0.0161795f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_373_n N_VPWR_c_445_n 0.0169033f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_363_n N_VPWR_c_446_n 0.00272266f $X=0.595 $Y=1.925 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_354_n N_VPWR_c_446_n 0.00662803f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_373_n N_VPWR_c_447_n 0.00699808f $X=3.39 $Y=1.955 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_373_n N_VPWR_c_448_n 0.00692422f $X=3.39 $Y=1.955 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_M1001_g N_VPWR_c_449_n 0.00392252f $X=3.535 $Y=1.985 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_373_n N_VPWR_c_449_n 0.0127815f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_287 N_A_27_47#_M1001_g N_VPWR_c_442_n 0.0067573f $X=3.535 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_363_n N_VPWR_c_442_n 0.00572244f $X=0.595 $Y=1.925 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_373_n N_VPWR_c_442_n 0.0529157f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_354_n N_VPWR_c_442_n 0.00838075f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_380_n N_VPWR_c_442_n 7.87123e-19 $X=0.68 $Y=1.925 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_373_n N_X_M1004_s 0.00442708f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_373_n N_X_M1010_s 0.00442755f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_347_n N_X_c_508_n 0.0363015f $X=0.68 $Y=1.81 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_344_n N_X_c_513_n 0.00325423f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_345_n N_X_c_510_n 0.0148935f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_347_n N_X_c_537_n 0.0224924f $X=0.68 $Y=1.81 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_373_n N_X_c_537_n 0.00861686f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_299 N_A_27_47#_c_373_n X 0.06067f $X=3.39 $Y=1.955 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_373_n A_542_297# 0.00781724f $X=3.39 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_301 N_A_27_47#_c_373_n A_626_297# 0.0101698f $X=3.39 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_302 N_A_27_47#_c_353_n A_626_297# 0.00412914f $X=3.505 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_303 N_A_27_47#_c_345_n N_VGND_M1013_d 0.00308856f $X=0.595 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_304 N_A_27_47#_c_345_n N_VGND_c_581_n 0.0124847f $X=0.595 $Y=0.82 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_350_n N_VGND_c_584_n 0.0104844f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_350_n N_VGND_c_591_n 0.00341689f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_M1013_s N_VGND_c_592_n 0.00236396f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_344_n N_VGND_c_592_n 0.00973659f $X=0.26 $Y=0.455 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_345_n N_VGND_c_592_n 0.00709158f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_350_n N_VGND_c_592_n 0.00512785f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_344_n N_VGND_c_593_n 0.014595f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_345_n N_VGND_c_593_n 0.00385657f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_442_n N_X_M1004_s 0.00333025f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_c_442_n N_X_M1010_s 0.00333025f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_M1007_d X 0.00168902f $X=1.45 $Y=1.485 $X2=0 $Y2=0
cc_316 N_VPWR_c_442_n A_542_297# 0.00333025f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_317 N_VPWR_c_442_n A_626_297# 0.00406927f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_318 N_X_c_509_n N_VGND_M1003_d 0.00162006f $X=1.855 $Y=0.82 $X2=0 $Y2=0
cc_319 N_X_c_513_n N_VGND_c_581_n 0.0175677f $X=1.165 $Y=0.395 $X2=0 $Y2=0
cc_320 N_X_c_509_n N_VGND_c_582_n 0.0122414f $X=1.855 $Y=0.82 $X2=0 $Y2=0
cc_321 N_X_c_513_n N_VGND_c_585_n 0.0158178f $X=1.165 $Y=0.395 $X2=0 $Y2=0
cc_322 N_X_c_509_n N_VGND_c_585_n 0.00193763f $X=1.855 $Y=0.82 $X2=0 $Y2=0
cc_323 N_X_c_510_n N_VGND_c_585_n 9.39298e-19 $X=1.132 $Y=0.82 $X2=0 $Y2=0
cc_324 N_X_c_509_n N_VGND_c_587_n 0.00213422f $X=1.855 $Y=0.82 $X2=0 $Y2=0
cc_325 N_X_c_538_n N_VGND_c_587_n 0.013896f $X=2.005 $Y=0.42 $X2=0 $Y2=0
cc_326 N_X_M1002_s N_VGND_c_592_n 0.00216698f $X=1.03 $Y=0.235 $X2=0 $Y2=0
cc_327 N_X_M1005_s N_VGND_c_592_n 0.0038878f $X=1.87 $Y=0.235 $X2=0 $Y2=0
cc_328 N_X_c_513_n N_VGND_c_592_n 0.0120119f $X=1.165 $Y=0.395 $X2=0 $Y2=0
cc_329 N_X_c_509_n N_VGND_c_592_n 0.00857624f $X=1.855 $Y=0.82 $X2=0 $Y2=0
cc_330 N_X_c_510_n N_VGND_c_592_n 0.00148235f $X=1.132 $Y=0.82 $X2=0 $Y2=0
cc_331 N_X_c_538_n N_VGND_c_592_n 0.00878527f $X=2.005 $Y=0.42 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__fa_1.spice
* Created: Tue Sep  1 19:08:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__fa_1.pex.spice"
.subckt sky130_fd_sc_hd__fa_1  VNB VPB A B CIN COUT VPWR SUM VGND
* 
* VGND	VGND
* SUM	SUM
* VPWR	VPWR
* COUT	COUT
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_A_76_199#_M1024_g N_COUT_M1024_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12435 AS=0.169 PD=1.20888 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1020 A_208_47# N_A_M1020_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.42 AD=0.063
+ AS=0.0803495 PD=0.72 PS=0.781121 NRD=27.132 NRS=19.992 M=1 R=2.8 SA=75000.7
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1025 N_A_76_199#_M1025_d N_B_M1025_g A_208_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.063 PD=0.69 PS=0.72 NRD=0 NRS=27.132 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1023 N_A_382_47#_M1023_d N_CIN_M1023_g N_A_76_199#_M1025_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_382_47#_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_382_47#_M1000_d N_B_M1000_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_A_738_47#_M1026_d N_B_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_CIN_M1014_g N_A_738_47#_M1026_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1019 N_A_738_47#_M1019_d N_A_M1019_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.0567 PD=0.715 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_995_47#_M1007_d N_A_76_199#_M1007_g N_A_738_47#_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0693 AS=0.06195 PD=0.75 PS=0.715 NRD=15.708 NRS=5.712 M=1
+ R=2.8 SA=75001.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1002 A_1091_47# N_CIN_M1002_g N_A_995_47#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0693 PD=0.63 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1004 A_1163_47# N_B_M1004_g A_1091_47# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0441 PD=0.75 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8 SA=75002.3 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g A_1163_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0803495 AS=0.0693 PD=0.781121 PS=0.75 NRD=0 NRS=31.428 M=1 R=2.8
+ SA=75002.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_SUM_M1016_d N_A_995_47#_M1016_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12435 PD=1.82 PS=1.20888 NRD=0 NRS=12.912 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1017 N_VPWR_M1017_d N_A_76_199#_M1017_g N_COUT_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.208239 AS=0.26 PD=1.89437 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1011 A_208_413# N_A_M1011_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=0.42 AD=0.063
+ AS=0.0874606 PD=0.72 PS=0.795634 NRD=44.5417 NRS=32.8202 M=1 R=2.8 SA=75000.7
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1018 N_A_76_199#_M1018_d N_B_M1018_g A_208_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.063 PD=0.69 PS=0.72 NRD=0 NRS=44.5417 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_A_382_413#_M1012_d N_CIN_M1012_g N_A_76_199#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_A_382_413#_M1012_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_382_413#_M1005_d N_B_M1005_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_738_413#_M1022_d N_B_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_CIN_M1008_g N_A_738_413#_M1022_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_738_413#_M1003_d N_A_M1003_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06195 AS=0.0567 PD=0.715 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 N_A_995_47#_M1010_d N_A_76_199#_M1010_g N_A_738_413#_M1003_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0693 AS=0.06195 PD=0.75 PS=0.715 NRD=25.7873 NRS=9.3772 M=1
+ R=2.8 SA=75001.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1021 A_1091_413# N_CIN_M1021_g N_A_995_47#_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0693 PD=0.63 PS=0.75 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1027 A_1163_413# N_B_M1027_g A_1091_413# VPB PHIGHVT L=0.15 W=0.42 AD=0.0693
+ AS=0.0441 PD=0.75 PS=0.63 NRD=51.5943 NRS=23.443 M=1 R=2.8 SA=75002.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g A_1163_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0874606 AS=0.0693 PD=0.795634 PS=0.75 NRD=32.8202 NRS=51.5943 M=1 R=2.8
+ SA=75002.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_SUM_M1006_d N_A_995_47#_M1006_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.208239 PD=2.52 PS=1.89437 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=12.4227 P=18.69
c_175 VPB 0 1.32337e-19 $X=0.15 $Y=2.635
c_1263 A_208_413# 0 7.82359e-20 $X=1.04 $Y=2.065
*
.include "sky130_fd_sc_hd__fa_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_inputiso1p_1.pex.spice
* Created: Tue Sep  1 19:12:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_1%A 3 7 9 10 18
r28 17 18 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.615 $Y=1.16
+ $X2=0.675 $Y2=1.16
r29 14 17 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.415 $Y=1.16
+ $X2=0.615 $Y2=1.16
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.415
+ $Y=1.16 $X2=0.415 $Y2=1.16
r31 10 15 0.973895 $w=3.53e-07 $l=3e-08 $layer=LI1_cond $X=0.322 $Y=1.19
+ $X2=0.322 $Y2=1.16
r32 9 15 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.322 $Y=0.85
+ $X2=0.322 $Y2=1.16
r33 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.675 $Y=1.325
+ $X2=0.675 $Y2=1.16
r34 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.675 $Y=1.325
+ $X2=0.675 $Y2=1.695
r35 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=1.16
r36 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.615 $Y=0.995
+ $X2=0.615 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_1%SLEEP 3 7 9 10 14
r37 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.16
+ $X2=1.095 $Y2=1.325
r38 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.16
+ $X2=1.095 $Y2=0.995
r39 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.16 $X2=1.095 $Y2=1.16
r40 9 10 13.4814 $w=2.63e-07 $l=3.1e-07 $layer=LI1_cond $X=1.142 $Y=0.85
+ $X2=1.142 $Y2=1.16
r41 7 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.035 $Y=1.695
+ $X2=1.035 $Y2=1.325
r42 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.035 $Y=0.445
+ $X2=1.035 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_1%A_68_297# 1 2 9 12 15 16 17 20
+ 21 27 31
c54 20 0 9.5905e-20 $X=1.61 $Y=1.16
c55 15 0 1.0136e-19 $X=0.755 $Y=1.495
r56 27 29 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=0.43
+ $X2=0.81 $Y2=0.595
r57 21 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.61 $Y2=1.325
r58 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.61 $Y2=0.995
r59 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.16 $X2=1.61 $Y2=1.16
r60 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.61 $Y=1.495
+ $X2=1.61 $Y2=1.16
r61 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.58
+ $X2=1.61 $Y2=1.495
r62 16 17 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.525 $Y=1.58
+ $X2=0.84 $Y2=1.58
r63 15 17 5.63966 $w=2.89e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.755 $Y=1.495
+ $X2=0.84 $Y2=1.58
r64 15 24 12.2422 $w=2.89e-07 $l=3.66033e-07 $layer=LI1_cond $X=0.755 $Y=1.495
+ $X2=0.465 $Y2=1.667
r65 15 29 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=0.755 $Y=1.495
+ $X2=0.755 $Y2=0.595
r66 12 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.52 $Y=1.985
+ $X2=1.52 $Y2=1.325
r67 9 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.52 $Y=0.56 $X2=1.52
+ $Y2=0.995
r68 2 24 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.485 $X2=0.465 $Y2=1.66
r69 1 27 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.235 $X2=0.825 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_1%VPWR 1 6 8 10 17 18 21
r20 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r21 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r22 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r23 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.31 $Y2=2.72
r24 15 17 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=2.07 $Y2=2.72
r25 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=2.72
+ $X2=1.31 $Y2=2.72
r26 10 12 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.145 $Y=2.72
+ $X2=0.23 $Y2=2.72
r27 8 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r28 8 12 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r29 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=2.635 $X2=1.31
+ $Y2=2.72
r30 4 6 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=1.31 $Y=2.635
+ $X2=1.31 $Y2=1.92
r31 1 6 300 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.485 $X2=1.31 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_1%X 1 2 10 13 19
c25 2 0 9.5905e-20 $X=1.595 $Y=1.485
r26 19 20 2.56478 $w=5.33e-07 $l=2.5e-08 $layer=LI1_cond $X=1.912 $Y=1.87
+ $X2=1.912 $Y2=1.845
r27 13 23 2.23566 $w=5.33e-07 $l=1e-07 $layer=LI1_cond $X=1.912 $Y=1.9 $X2=1.912
+ $Y2=2
r28 13 19 0.670698 $w=5.33e-07 $l=3e-08 $layer=LI1_cond $X=1.912 $Y=1.9
+ $X2=1.912 $Y2=1.87
r29 13 20 1.09756 $w=3.13e-07 $l=3e-08 $layer=LI1_cond $X=2.022 $Y=1.815
+ $X2=2.022 $Y2=1.845
r30 11 13 36.2196 $w=3.13e-07 $l=9.9e-07 $layer=LI1_cond $X=2.022 $Y=0.825
+ $X2=2.022 $Y2=1.815
r31 10 11 4.21929 $w=3.15e-07 $l=2.85e-07 $layer=LI1_cond $X=2.022 $Y=0.54
+ $X2=2.022 $Y2=0.825
r32 8 10 6.12728 $w=5.68e-07 $l=2.92e-07 $layer=LI1_cond $X=1.73 $Y=0.54
+ $X2=2.022 $Y2=0.54
r33 2 23 300 $w=1.7e-07 $l=6.13148e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.485 $X2=1.81 $Y2=2
r34 1 8 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.595
+ $Y=0.235 $X2=1.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO1P_1%VGND 1 2 7 9 13 16 17 18 25 26
r30 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r31 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r32 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r33 20 29 3.81131 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.49 $Y=0 $X2=0.245
+ $Y2=0
r34 20 22 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=0.49 $Y=0 $X2=1.15
+ $Y2=0
r35 18 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r36 18 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r37 16 22 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.15
+ $Y2=0
r38 16 17 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.287
+ $Y2=0
r39 15 25 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=2.07
+ $Y2=0
r40 15 17 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.287
+ $Y2=0
r41 11 17 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.287 $Y=0.085
+ $X2=1.287 $Y2=0
r42 11 13 18.4927 $w=2.13e-07 $l=3.45e-07 $layer=LI1_cond $X=1.287 $Y=0.085
+ $X2=1.287 $Y2=0.43
r43 7 29 3.26684 $w=2.4e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.245 $Y2=0
r44 7 9 16.5664 $w=2.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.43
r45 2 13 182 $w=1.7e-07 $l=2.75772e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.235 $X2=1.305 $Y2=0.43
r46 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.28
+ $Y=0.235 $X2=0.405 $Y2=0.43
.ends


* File: sky130_fd_sc_hd__lpflow_decapkapwr_8.pex.spice
* Created: Thu Aug 27 14:24:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%VGND 1 9 10 11 12 21 33 36
r22 35 36 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r23 33 35 0.445255 $w=8.22e-07 $l=3e-08 $layer=LI1_cond $X=3.42 $Y=0.385
+ $X2=3.45 $Y2=0.385
r24 30 36 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=3.45
+ $Y2=0
r25 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r26 23 26 0.262178 $w=1.396e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.645
+ $X2=0.26 $Y2=0.645
r27 20 29 7.51576 $w=1.396e-06 $l=8.6e-07 $layer=LI1_cond $X=1.55 $Y=0.645
+ $X2=0.69 $Y2=0.645
r28 19 21 8.47369 $w=1.49e-06 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.87
+ $X2=1.715 $Y2=1.87
r29 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.29 $X2=1.55 $Y2=1.29
r30 16 29 1.1361 $w=1.396e-06 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=0.645
+ $X2=0.69 $Y2=0.645
r31 16 26 2.62178 $w=1.396e-06 $l=3e-07 $layer=LI1_cond $X=0.56 $Y=0.645
+ $X2=0.26 $Y2=0.645
r32 15 19 32.8283 $w=1.49e-06 $l=9.9e-07 $layer=POLY_cond $X=0.56 $Y=1.87
+ $X2=1.55 $Y2=1.87
r33 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.56
+ $Y=1.29 $X2=0.56 $Y2=1.29
r34 12 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r35 12 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r36 11 20 2.92381 $w=1.396e-06 $l=3.40147e-07 $layer=LI1_cond $X=1.735 $Y=0.385
+ $X2=1.55 $Y2=0.645
r37 10 33 4.05283 $w=9.4e-07 $l=2.95e-07 $layer=LI1_cond $X=3.125 $Y=0.385
+ $X2=3.42 $Y2=0.385
r38 10 11 18.0404 $w=9.38e-07 $l=1.39e-06 $layer=LI1_cond $X=3.125 $Y=0.385
+ $X2=1.735 $Y2=0.385
r39 9 21 5.33186 $w=1.13e-06 $l=1.25e-07 $layer=POLY_cond $X=1.84 $Y=2.05
+ $X2=1.715 $Y2=2.05
r40 1 33 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=3.285 $Y=0.235
+ $X2=3.42 $Y2=0.475
r41 1 26 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%KAPWR 1 9 12 18 20 31 36 37 39
+ 41
c25 37 0 7.9696e-20 $X=3.45 $Y=2.21
r26 39 41 0.0085136 $w=2.6e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=2.21
+ $X2=0.23 $Y2=2.21
r27 36 37 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=2.21
+ $X2=3.45 $Y2=2.21
r28 34 36 0.254167 $w=1.438e-06 $l=3e-08 $layer=LI1_cond $X=3.42 $Y=1.745
+ $X2=3.45 $Y2=1.745
r29 29 31 21.8141 $w=9.18e-07 $l=1.645e-06 $layer=LI1_cond $X=0.26 $Y=2.005
+ $X2=1.905 $Y2=2.005
r30 25 29 0.397826 $w=9.18e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=2.005
+ $X2=0.26 $Y2=2.005
r31 25 41 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=2.21
+ $X2=0.23 $Y2=2.21
r32 21 34 2.54167 $w=1.438e-06 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.745
+ $X2=3.42 $Y2=1.745
r33 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.11 $X2=3.12 $Y2=1.11
r34 17 21 8.72639 $w=1.438e-06 $l=1.03e-06 $layer=LI1_cond $X=2.09 $Y=1.745
+ $X2=3.12 $Y2=1.745
r35 17 31 3.1528 $w=1.438e-06 $l=1.85e-07 $layer=LI1_cond $X=2.09 $Y=1.745
+ $X2=1.905 $Y2=1.745
r36 16 20 45.2647 $w=1.17e-06 $l=1.03e-06 $layer=POLY_cond $X=2.09 $Y=0.69
+ $X2=3.12 $Y2=0.69
r37 16 18 12.167 $w=1.17e-06 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=0.69
+ $X2=1.925 $Y2=0.69
r38 16 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.11 $X2=2.09 $Y2=1.11
r39 12 39 0.0120192 $w=2.6e-07 $l=2.5e-08 $layer=MET1_cond $X=0.19 $Y=2.21
+ $X2=0.215 $Y2=2.21
r40 12 37 1.80091 $w=2.6e-07 $l=3.173e-06 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=3.45 $Y2=2.21
r41 12 41 0.0266759 $w=2.6e-07 $l=4.7e-08 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=0.23 $Y2=2.21
r42 9 18 5.05802 $w=8.1e-07 $l=8.5e-08 $layer=POLY_cond $X=1.84 $Y=0.51
+ $X2=1.925 $Y2=0.51
r43 1 34 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.615 $X2=3.42 $Y2=1.83
r44 1 29 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_8%VPWR 1 8 9
c10 8 0 7.9696e-20 $X=3.45 $Y=2.72
r11 8 9 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r12 4 8 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=3.45
+ $Y2=2.72
r13 1 9 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.45 $Y2=2.72
r14 1 4 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
.ends


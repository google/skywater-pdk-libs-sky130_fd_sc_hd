* File: sky130_fd_sc_hd__and4bb_4.pxi.spice
* Created: Thu Aug 27 14:09:17 2020
* 
x_PM_SKY130_FD_SC_HD__AND4BB_4%B_N N_B_N_M1017_g N_B_N_M1009_g B_N B_N B_N
+ N_B_N_c_104_n PM_SKY130_FD_SC_HD__AND4BB_4%B_N
x_PM_SKY130_FD_SC_HD__AND4BB_4%A_174_21# N_A_174_21#_M1018_d N_A_174_21#_M1016_d
+ N_A_174_21#_M1005_d N_A_174_21#_M1001_g N_A_174_21#_c_145_n
+ N_A_174_21#_M1000_g N_A_174_21#_M1003_g N_A_174_21#_c_146_n
+ N_A_174_21#_M1002_g N_A_174_21#_M1007_g N_A_174_21#_c_147_n
+ N_A_174_21#_M1011_g N_A_174_21#_M1019_g N_A_174_21#_c_148_n
+ N_A_174_21#_M1012_g N_A_174_21#_c_190_p N_A_174_21#_c_140_n
+ N_A_174_21#_c_141_n N_A_174_21#_c_159_p N_A_174_21#_c_244_p
+ N_A_174_21#_c_191_p N_A_174_21#_c_156_p N_A_174_21#_c_172_p
+ N_A_174_21#_c_142_n N_A_174_21#_c_173_p N_A_174_21#_c_143_n
+ N_A_174_21#_c_144_n PM_SKY130_FD_SC_HD__AND4BB_4%A_174_21#
x_PM_SKY130_FD_SC_HD__AND4BB_4%D N_D_M1004_g N_D_M1016_g D N_D_c_281_n
+ N_D_c_282_n PM_SKY130_FD_SC_HD__AND4BB_4%D
x_PM_SKY130_FD_SC_HD__AND4BB_4%C N_C_M1008_g N_C_M1010_g C C N_C_c_320_n
+ N_C_c_321_n PM_SKY130_FD_SC_HD__AND4BB_4%C
x_PM_SKY130_FD_SC_HD__AND4BB_4%A_27_47# N_A_27_47#_M1017_s N_A_27_47#_M1009_s
+ N_A_27_47#_M1013_g N_A_27_47#_M1005_g N_A_27_47#_c_354_n N_A_27_47#_c_362_n
+ N_A_27_47#_c_363_n N_A_27_47#_c_355_n N_A_27_47#_c_365_n N_A_27_47#_c_356_n
+ N_A_27_47#_c_366_n N_A_27_47#_c_357_n N_A_27_47#_c_358_n N_A_27_47#_c_359_n
+ PM_SKY130_FD_SC_HD__AND4BB_4%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4BB_4%A_832_21# N_A_832_21#_M1014_d N_A_832_21#_M1006_d
+ N_A_832_21#_c_445_n N_A_832_21#_M1018_g N_A_832_21#_M1015_g
+ N_A_832_21#_c_446_n N_A_832_21#_c_447_n N_A_832_21#_c_448_n
+ N_A_832_21#_c_449_n N_A_832_21#_c_450_n N_A_832_21#_c_455_n
+ N_A_832_21#_c_456_n N_A_832_21#_c_504_p N_A_832_21#_c_488_p
+ PM_SKY130_FD_SC_HD__AND4BB_4%A_832_21#
x_PM_SKY130_FD_SC_HD__AND4BB_4%A_N N_A_N_M1014_g N_A_N_M1006_g A_N A_N
+ N_A_N_c_511_n N_A_N_c_512_n PM_SKY130_FD_SC_HD__AND4BB_4%A_N
x_PM_SKY130_FD_SC_HD__AND4BB_4%VPWR N_VPWR_M1009_d N_VPWR_M1002_d N_VPWR_M1012_d
+ N_VPWR_M1010_d N_VPWR_M1015_d N_VPWR_c_535_n N_VPWR_c_536_n N_VPWR_c_537_n
+ N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_542_n
+ VPWR N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n
+ N_VPWR_c_534_n N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n
+ N_VPWR_c_552_n PM_SKY130_FD_SC_HD__AND4BB_4%VPWR
x_PM_SKY130_FD_SC_HD__AND4BB_4%X N_X_M1001_d N_X_M1007_d N_X_M1000_s N_X_M1011_s
+ N_X_c_660_p N_X_c_663_p N_X_c_634_n X X X N_X_c_630_n X X N_X_c_646_n
+ PM_SKY130_FD_SC_HD__AND4BB_4%X
x_PM_SKY130_FD_SC_HD__AND4BB_4%VGND N_VGND_M1017_d N_VGND_M1003_s N_VGND_M1019_s
+ N_VGND_M1014_s N_VGND_c_671_n N_VGND_c_672_n N_VGND_c_673_n N_VGND_c_674_n
+ N_VGND_c_675_n N_VGND_c_676_n VGND N_VGND_c_677_n N_VGND_c_678_n
+ N_VGND_c_679_n N_VGND_c_680_n N_VGND_c_681_n N_VGND_c_682_n N_VGND_c_683_n
+ N_VGND_c_684_n PM_SKY130_FD_SC_HD__AND4BB_4%VGND
cc_1 VNB N_B_N_M1017_g 0.0321427f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB B_N 0.00354643f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_3 VNB N_B_N_c_104_n 0.0231135f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_4 VNB N_A_174_21#_M1001_g 0.0173209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_174_21#_M1003_g 0.0172377f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.325
cc_6 VNB N_A_174_21#_M1007_g 0.0172667f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.53
cc_7 VNB N_A_174_21#_M1019_g 0.0183688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_174_21#_c_140_n 0.00276841f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_174_21#_c_141_n 4.44797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_174_21#_c_142_n 0.012601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_174_21#_c_143_n 0.00104297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_174_21#_c_144_n 0.0691048f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB D 0.00431502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_D_c_281_n 0.0203084f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_15 VNB N_D_c_282_n 0.0176898f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB C 0.00300637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_C_c_320_n 0.0261176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_C_c_321_n 0.0176357f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_19 VNB N_A_27_47#_c_354_n 0.033106f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_20 VNB N_A_27_47#_c_355_n 0.00721425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_356_n 0.0128993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_357_n 0.00103878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_358_n 0.0217269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_359_n 0.0182267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_832_21#_c_445_n 0.0210055f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_26 VNB N_A_832_21#_c_446_n 0.00918427f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_27 VNB N_A_832_21#_c_447_n 0.00427151f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.325
cc_28 VNB N_A_832_21#_c_448_n 0.067178f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.85
cc_29 VNB N_A_832_21#_c_449_n 0.0218622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_832_21#_c_450_n 0.00350079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_N_M1014_g 0.0431418f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_32 VNB N_A_N_c_511_n 0.0263794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_N_c_512_n 0.0153089f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_34 VNB N_VPWR_c_534_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB X 0.00134056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_671_n 0.00271064f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_37 VNB N_VGND_c_672_n 3.05427e-19 $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.325
cc_38 VNB N_VGND_c_673_n 0.00278678f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.16
cc_39 VNB N_VGND_c_674_n 0.00899889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_675_n 0.0588037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_676_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_677_n 0.0178546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_678_n 0.0112618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_679_n 0.0123863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_680_n 0.0206251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_681_n 0.311093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_682_n 0.00507198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_683_n 0.00436184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_684_n 0.00518879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_B_N_M1009_g 0.0549471f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_51 VPB B_N 0.00193391f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_52 VPB N_B_N_c_104_n 0.00473762f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_53 VPB N_A_174_21#_c_145_n 0.0162256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_174_21#_c_146_n 0.0157459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_174_21#_c_147_n 0.0157686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_174_21#_c_148_n 0.0166323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_174_21#_c_141_n 0.00328606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_174_21#_c_144_n 0.0203908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_D_M1016_g 0.0206086f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_60 VPB D 0.00194512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_D_c_281_n 0.00419043f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_62 VPB N_C_M1010_g 0.0213457f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_63 VPB C 0.00303377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_C_c_320_n 0.00727566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_M1005_g 0.0213394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_354_n 0.0290594f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_67 VPB N_A_27_47#_c_362_n 0.0147617f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_68 VPB N_A_27_47#_c_363_n 0.00204048f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.85
cc_69 VPB N_A_27_47#_c_355_n 0.00215394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_365_n 0.00363704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_366_n 0.0110158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_357_n 7.01922e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_358_n 0.00432329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_832_21#_M1015_g 0.0228461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_832_21#_c_446_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_76 VPB N_A_832_21#_c_447_n 0.014747f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.325
cc_77 VPB N_A_832_21#_c_448_n 0.0390084f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.85
cc_78 VPB N_A_832_21#_c_455_n 0.018053f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.16
cc_79 VPB N_A_832_21#_c_456_n 0.00263967f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.19
cc_80 VPB N_A_N_M1006_g 0.0730399f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_81 VPB N_A_N_c_511_n 0.00491122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_N_c_512_n 0.0163234f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_83 VPB N_VPWR_c_535_n 0.00215067f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=0.995
cc_84 VPB N_VPWR_c_536_n 3.11529e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_537_n 0.00271156f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.53
cc_86 VPB N_VPWR_c_538_n 0.00562936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_539_n 0.0113234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_540_n 0.00872784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_541_n 0.011815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_542_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_543_n 0.014294f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_544_n 0.0143676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_545_n 0.0204795f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_546_n 0.0187885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_534_n 0.0455327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_548_n 0.00507168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_549_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_550_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_551_n 0.0191102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_552_n 0.00874105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB X 0.00105123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 N_B_N_M1017_g N_A_174_21#_M1001_g 0.019386f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_103 B_N N_A_174_21#_M1001_g 0.00673925f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_104 N_B_N_c_104_n N_A_174_21#_M1001_g 0.0201431f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B_N_M1009_g N_A_174_21#_c_144_n 0.0350771f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_106 N_B_N_M1017_g N_A_27_47#_c_354_n 0.010442f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_107 N_B_N_M1009_g N_A_27_47#_c_354_n 0.0161302f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_108 B_N N_A_27_47#_c_354_n 0.0657471f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_109 N_B_N_c_104_n N_A_27_47#_c_354_n 0.00753785f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B_N_M1009_g N_A_27_47#_c_363_n 0.0147588f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_111 B_N N_A_27_47#_c_363_n 0.0192342f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_112 N_B_N_c_104_n N_A_27_47#_c_363_n 7.40595e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_113 B_N N_VPWR_M1009_d 0.00387935f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_114 N_B_N_M1009_g N_VPWR_c_535_n 0.00832549f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_115 N_B_N_M1009_g N_VPWR_c_543_n 0.00339367f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_116 N_B_N_M1009_g N_VPWR_c_534_n 0.00489827f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_117 N_B_N_M1017_g X 6.24427e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_118 B_N X 0.00435374f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_119 N_B_N_M1009_g N_X_c_630_n 4.75342e-19 $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_120 B_N N_X_c_630_n 0.0071243f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_121 B_N X 0.0542375f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_122 N_B_N_c_104_n X 2.84869e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_123 B_N N_VGND_M1017_d 0.00337458f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_124 N_B_N_M1017_g N_VGND_c_671_n 0.00310635f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_125 B_N N_VGND_c_671_n 0.0101817f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_126 N_B_N_c_104_n N_VGND_c_671_n 2.92234e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B_N_M1017_g N_VGND_c_677_n 0.00585385f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_128 N_B_N_M1017_g N_VGND_c_681_n 0.00810792f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_129 B_N N_VGND_c_681_n 0.00602577f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_130 N_A_174_21#_c_148_n N_D_M1016_g 0.0190428f $X=2.205 $Y=1.375 $X2=0 $Y2=0
cc_131 N_A_174_21#_c_156_p N_D_M1016_g 0.010347f $X=3.985 $Y=1.63 $X2=0 $Y2=0
cc_132 N_A_174_21#_c_140_n D 0.00576147f $X=2.415 $Y=1.075 $X2=0 $Y2=0
cc_133 N_A_174_21#_c_141_n D 0.00576147f $X=2.415 $Y=1.545 $X2=0 $Y2=0
cc_134 N_A_174_21#_c_159_p D 0.0150695f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_135 N_A_174_21#_c_156_p D 0.022188f $X=3.985 $Y=1.63 $X2=0 $Y2=0
cc_136 N_A_174_21#_c_142_n D 0.00443117f $X=4.255 $Y=0.385 $X2=0 $Y2=0
cc_137 N_A_174_21#_c_143_n D 0.0139777f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_174_21#_c_144_n D 2.68365e-19 $X=2.205 $Y=1.2 $X2=0 $Y2=0
cc_139 N_A_174_21#_c_141_n N_D_c_281_n 0.00545094f $X=2.415 $Y=1.545 $X2=0 $Y2=0
cc_140 N_A_174_21#_c_159_p N_D_c_281_n 0.00252445f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_141 N_A_174_21#_c_156_p N_D_c_281_n 0.00245882f $X=3.985 $Y=1.63 $X2=0 $Y2=0
cc_142 N_A_174_21#_c_143_n N_D_c_281_n 0.00113172f $X=2.415 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_174_21#_c_144_n N_D_c_281_n 0.0356623f $X=2.205 $Y=1.2 $X2=0 $Y2=0
cc_144 N_A_174_21#_M1019_g N_D_c_282_n 0.0177362f $X=2.205 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A_174_21#_c_140_n N_D_c_282_n 0.00522591f $X=2.415 $Y=1.075 $X2=0 $Y2=0
cc_146 N_A_174_21#_c_159_p N_D_c_282_n 0.0126868f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_147 N_A_174_21#_c_172_p N_D_c_282_n 0.00368086f $X=2.855 $Y=0.615 $X2=0 $Y2=0
cc_148 N_A_174_21#_c_173_p N_D_c_282_n 0.00422018f $X=2.94 $Y=0.385 $X2=0 $Y2=0
cc_149 N_A_174_21#_c_156_p N_C_M1010_g 0.013565f $X=3.985 $Y=1.63 $X2=0 $Y2=0
cc_150 N_A_174_21#_c_159_p C 0.00153582f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_151 N_A_174_21#_c_156_p C 0.0171891f $X=3.985 $Y=1.63 $X2=0 $Y2=0
cc_152 N_A_174_21#_c_142_n C 0.0114881f $X=4.255 $Y=0.385 $X2=0 $Y2=0
cc_153 N_A_174_21#_c_156_p N_C_c_320_n 0.00125861f $X=3.985 $Y=1.63 $X2=0 $Y2=0
cc_154 N_A_174_21#_c_142_n N_C_c_320_n 7.39795e-19 $X=4.255 $Y=0.385 $X2=0 $Y2=0
cc_155 N_A_174_21#_c_159_p N_C_c_321_n 0.00407095f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_156 N_A_174_21#_c_172_p N_C_c_321_n 0.00303963f $X=2.855 $Y=0.615 $X2=0 $Y2=0
cc_157 N_A_174_21#_c_142_n N_C_c_321_n 0.0152586f $X=4.255 $Y=0.385 $X2=0 $Y2=0
cc_158 N_A_174_21#_c_156_p N_A_27_47#_M1005_g 0.0110208f $X=3.985 $Y=1.63 $X2=0
+ $Y2=0
cc_159 N_A_174_21#_M1016_d N_A_27_47#_c_363_n 0.00616873f $X=2.78 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_174_21#_M1005_d N_A_27_47#_c_363_n 0.00615835f $X=3.83 $Y=1.485 $X2=0
+ $Y2=0
cc_161 N_A_174_21#_c_145_n N_A_27_47#_c_363_n 0.0148185f $X=0.945 $Y=1.375 $X2=0
+ $Y2=0
cc_162 N_A_174_21#_c_146_n N_A_27_47#_c_363_n 0.0116333f $X=1.365 $Y=1.375 $X2=0
+ $Y2=0
cc_163 N_A_174_21#_c_147_n N_A_27_47#_c_363_n 0.0116333f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_164 N_A_174_21#_c_148_n N_A_27_47#_c_363_n 0.0137059f $X=2.205 $Y=1.375 $X2=0
+ $Y2=0
cc_165 N_A_174_21#_c_190_p N_A_27_47#_c_363_n 0.00311226f $X=2.33 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_174_21#_c_191_p N_A_27_47#_c_363_n 0.0117088f $X=2.5 $Y=1.63 $X2=0
+ $Y2=0
cc_167 N_A_174_21#_c_156_p N_A_27_47#_c_363_n 0.0788813f $X=3.985 $Y=1.63 $X2=0
+ $Y2=0
cc_168 N_A_174_21#_c_144_n N_A_27_47#_c_363_n 5.68379e-19 $X=2.205 $Y=1.2 $X2=0
+ $Y2=0
cc_169 N_A_174_21#_c_156_p N_A_27_47#_c_355_n 0.0137593f $X=3.985 $Y=1.63 $X2=0
+ $Y2=0
cc_170 N_A_174_21#_c_142_n N_A_27_47#_c_355_n 0.00960477f $X=4.255 $Y=0.385
+ $X2=0 $Y2=0
cc_171 N_A_174_21#_c_156_p N_A_27_47#_c_357_n 0.00822672f $X=3.985 $Y=1.63 $X2=0
+ $Y2=0
cc_172 N_A_174_21#_c_142_n N_A_27_47#_c_357_n 0.00403727f $X=4.255 $Y=0.385
+ $X2=0 $Y2=0
cc_173 N_A_174_21#_c_156_p N_A_27_47#_c_358_n 0.00143746f $X=3.985 $Y=1.63 $X2=0
+ $Y2=0
cc_174 N_A_174_21#_c_142_n N_A_27_47#_c_358_n 0.00151018f $X=4.255 $Y=0.385
+ $X2=0 $Y2=0
cc_175 N_A_174_21#_c_142_n N_A_27_47#_c_359_n 0.0154295f $X=4.255 $Y=0.385 $X2=0
+ $Y2=0
cc_176 N_A_174_21#_c_142_n N_A_832_21#_c_445_n 0.0198002f $X=4.255 $Y=0.385
+ $X2=0 $Y2=0
cc_177 N_A_174_21#_c_142_n N_A_832_21#_c_448_n 0.00919115f $X=4.255 $Y=0.385
+ $X2=0 $Y2=0
cc_178 N_A_174_21#_c_142_n N_A_832_21#_c_450_n 0.00851485f $X=4.255 $Y=0.385
+ $X2=0 $Y2=0
cc_179 N_A_174_21#_c_141_n N_VPWR_M1012_d 0.00102719f $X=2.415 $Y=1.545 $X2=0
+ $Y2=0
cc_180 N_A_174_21#_c_191_p N_VPWR_M1012_d 0.00296279f $X=2.5 $Y=1.63 $X2=0 $Y2=0
cc_181 N_A_174_21#_c_156_p N_VPWR_M1012_d 0.00356965f $X=3.985 $Y=1.63 $X2=0
+ $Y2=0
cc_182 N_A_174_21#_c_156_p N_VPWR_M1010_d 0.00938792f $X=3.985 $Y=1.63 $X2=0
+ $Y2=0
cc_183 N_A_174_21#_c_145_n N_VPWR_c_535_n 0.0016047f $X=0.945 $Y=1.375 $X2=0
+ $Y2=0
cc_184 N_A_174_21#_c_145_n N_VPWR_c_536_n 0.00114039f $X=0.945 $Y=1.375 $X2=0
+ $Y2=0
cc_185 N_A_174_21#_c_146_n N_VPWR_c_536_n 0.00842528f $X=1.365 $Y=1.375 $X2=0
+ $Y2=0
cc_186 N_A_174_21#_c_147_n N_VPWR_c_536_n 0.00810864f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_187 N_A_174_21#_c_148_n N_VPWR_c_536_n 0.00110281f $X=2.205 $Y=1.375 $X2=0
+ $Y2=0
cc_188 N_A_174_21#_c_147_n N_VPWR_c_537_n 0.00110281f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_189 N_A_174_21#_c_148_n N_VPWR_c_537_n 0.00815407f $X=2.205 $Y=1.375 $X2=0
+ $Y2=0
cc_190 N_A_174_21#_c_147_n N_VPWR_c_541_n 0.00339367f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_191 N_A_174_21#_c_148_n N_VPWR_c_541_n 0.00339367f $X=2.205 $Y=1.375 $X2=0
+ $Y2=0
cc_192 N_A_174_21#_c_145_n N_VPWR_c_544_n 0.00425094f $X=0.945 $Y=1.375 $X2=0
+ $Y2=0
cc_193 N_A_174_21#_c_146_n N_VPWR_c_544_n 0.00339367f $X=1.365 $Y=1.375 $X2=0
+ $Y2=0
cc_194 N_A_174_21#_M1016_d N_VPWR_c_534_n 0.00385378f $X=2.78 $Y=1.485 $X2=0
+ $Y2=0
cc_195 N_A_174_21#_M1005_d N_VPWR_c_534_n 0.00385378f $X=3.83 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_A_174_21#_c_145_n N_VPWR_c_534_n 0.00580516f $X=0.945 $Y=1.375 $X2=0
+ $Y2=0
cc_197 N_A_174_21#_c_146_n N_VPWR_c_534_n 0.00398704f $X=1.365 $Y=1.375 $X2=0
+ $Y2=0
cc_198 N_A_174_21#_c_147_n N_VPWR_c_534_n 0.00398704f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_199 N_A_174_21#_c_148_n N_VPWR_c_534_n 0.00398704f $X=2.205 $Y=1.375 $X2=0
+ $Y2=0
cc_200 N_A_174_21#_M1003_g N_X_c_634_n 0.015219f $X=1.365 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_174_21#_M1007_g N_X_c_634_n 0.0115365f $X=1.785 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A_174_21#_c_190_p N_X_c_634_n 0.0300956f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_174_21#_c_144_n N_X_c_634_n 0.00417342f $X=2.205 $Y=1.2 $X2=0 $Y2=0
cc_204 N_A_174_21#_M1001_g X 0.00673409f $X=0.945 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A_174_21#_c_145_n N_X_c_630_n 0.00391178f $X=0.945 $Y=1.375 $X2=0 $Y2=0
cc_206 N_A_174_21#_M1001_g X 0.00437659f $X=0.945 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_174_21#_c_145_n X 0.00309782f $X=0.945 $Y=1.375 $X2=0 $Y2=0
cc_208 N_A_174_21#_M1003_g X 0.00392198f $X=1.365 $Y=0.56 $X2=0 $Y2=0
cc_209 N_A_174_21#_c_146_n X 0.0028656f $X=1.365 $Y=1.375 $X2=0 $Y2=0
cc_210 N_A_174_21#_c_190_p X 0.0132531f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_174_21#_c_144_n X 0.0266213f $X=2.205 $Y=1.2 $X2=0 $Y2=0
cc_212 N_A_174_21#_c_146_n N_X_c_646_n 0.0123431f $X=1.365 $Y=1.375 $X2=0 $Y2=0
cc_213 N_A_174_21#_c_147_n N_X_c_646_n 0.00929518f $X=1.785 $Y=1.375 $X2=0 $Y2=0
cc_214 N_A_174_21#_c_148_n N_X_c_646_n 0.00274959f $X=2.205 $Y=1.375 $X2=0 $Y2=0
cc_215 N_A_174_21#_c_190_p N_X_c_646_n 0.0280758f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_174_21#_c_144_n N_X_c_646_n 0.00434986f $X=2.205 $Y=1.2 $X2=0 $Y2=0
cc_217 N_A_174_21#_c_140_n N_VGND_M1019_s 0.00148984f $X=2.415 $Y=1.075 $X2=0
+ $Y2=0
cc_218 N_A_174_21#_c_159_p N_VGND_M1019_s 0.00348067f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_219 N_A_174_21#_c_244_p N_VGND_M1019_s 0.00272918f $X=2.5 $Y=0.7 $X2=0 $Y2=0
cc_220 N_A_174_21#_M1001_g N_VGND_c_671_n 0.00769236f $X=0.945 $Y=0.56 $X2=0
+ $Y2=0
cc_221 N_A_174_21#_M1003_g N_VGND_c_671_n 5.10275e-19 $X=1.365 $Y=0.56 $X2=0
+ $Y2=0
cc_222 N_A_174_21#_M1001_g N_VGND_c_672_n 5.10275e-19 $X=0.945 $Y=0.56 $X2=0
+ $Y2=0
cc_223 N_A_174_21#_M1003_g N_VGND_c_672_n 0.00670862f $X=1.365 $Y=0.56 $X2=0
+ $Y2=0
cc_224 N_A_174_21#_M1007_g N_VGND_c_672_n 0.00675643f $X=1.785 $Y=0.56 $X2=0
+ $Y2=0
cc_225 N_A_174_21#_M1019_g N_VGND_c_672_n 5.18673e-19 $X=2.205 $Y=0.56 $X2=0
+ $Y2=0
cc_226 N_A_174_21#_M1007_g N_VGND_c_673_n 4.92041e-19 $X=1.785 $Y=0.56 $X2=0
+ $Y2=0
cc_227 N_A_174_21#_M1019_g N_VGND_c_673_n 0.00565488f $X=2.205 $Y=0.56 $X2=0
+ $Y2=0
cc_228 N_A_174_21#_c_190_p N_VGND_c_673_n 7.71914e-19 $X=2.33 $Y=1.16 $X2=0
+ $Y2=0
cc_229 N_A_174_21#_c_159_p N_VGND_c_673_n 0.00550144f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_230 N_A_174_21#_c_244_p N_VGND_c_673_n 0.0136474f $X=2.5 $Y=0.7 $X2=0 $Y2=0
cc_231 N_A_174_21#_c_144_n N_VGND_c_673_n 2.89755e-19 $X=2.205 $Y=1.2 $X2=0
+ $Y2=0
cc_232 N_A_174_21#_c_142_n N_VGND_c_674_n 0.00814718f $X=4.255 $Y=0.385 $X2=0
+ $Y2=0
cc_233 N_A_174_21#_c_159_p N_VGND_c_675_n 0.00269343f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_234 N_A_174_21#_c_142_n N_VGND_c_675_n 0.075401f $X=4.255 $Y=0.385 $X2=0
+ $Y2=0
cc_235 N_A_174_21#_c_173_p N_VGND_c_675_n 0.00759604f $X=2.94 $Y=0.385 $X2=0
+ $Y2=0
cc_236 N_A_174_21#_M1001_g N_VGND_c_678_n 0.00403236f $X=0.945 $Y=0.56 $X2=0
+ $Y2=0
cc_237 N_A_174_21#_M1003_g N_VGND_c_678_n 0.00341112f $X=1.365 $Y=0.56 $X2=0
+ $Y2=0
cc_238 N_A_174_21#_M1007_g N_VGND_c_679_n 0.00341112f $X=1.785 $Y=0.56 $X2=0
+ $Y2=0
cc_239 N_A_174_21#_M1019_g N_VGND_c_679_n 0.00544582f $X=2.205 $Y=0.56 $X2=0
+ $Y2=0
cc_240 N_A_174_21#_M1018_d N_VGND_c_681_n 0.00212021f $X=4.31 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_A_174_21#_M1001_g N_VGND_c_681_n 0.00596417f $X=0.945 $Y=0.56 $X2=0
+ $Y2=0
cc_242 N_A_174_21#_M1003_g N_VGND_c_681_n 0.00397316f $X=1.365 $Y=0.56 $X2=0
+ $Y2=0
cc_243 N_A_174_21#_M1007_g N_VGND_c_681_n 0.00397316f $X=1.785 $Y=0.56 $X2=0
+ $Y2=0
cc_244 N_A_174_21#_M1019_g N_VGND_c_681_n 0.00912034f $X=2.205 $Y=0.56 $X2=0
+ $Y2=0
cc_245 N_A_174_21#_c_159_p N_VGND_c_681_n 0.00459547f $X=2.77 $Y=0.7 $X2=0 $Y2=0
cc_246 N_A_174_21#_c_244_p N_VGND_c_681_n 8.89004e-19 $X=2.5 $Y=0.7 $X2=0 $Y2=0
cc_247 N_A_174_21#_c_142_n N_VGND_c_681_n 0.0586418f $X=4.255 $Y=0.385 $X2=0
+ $Y2=0
cc_248 N_A_174_21#_c_173_p N_VGND_c_681_n 0.00628982f $X=2.94 $Y=0.385 $X2=0
+ $Y2=0
cc_249 N_A_174_21#_c_159_p A_556_47# 0.00330744f $X=2.77 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_250 N_A_174_21#_c_172_p A_556_47# 0.00165856f $X=2.855 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_251 N_A_174_21#_c_142_n A_556_47# 0.00323394f $X=4.255 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_252 N_A_174_21#_c_173_p A_556_47# 0.00109783f $X=2.94 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_174_21#_c_142_n A_652_47# 0.00954505f $X=4.255 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_254 N_A_174_21#_c_142_n A_766_47# 0.00906169f $X=4.255 $Y=0.385 $X2=-0.19
+ $Y2=-0.24
cc_255 N_D_M1016_g N_C_M1010_g 0.0373813f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_256 D C 0.0262737f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_257 N_D_c_281_n C 2.39128e-19 $X=2.765 $Y=1.16 $X2=0 $Y2=0
cc_258 N_D_c_282_n C 9.98121e-19 $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_259 D N_C_c_320_n 0.0025442f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_260 N_D_c_281_n N_C_c_320_n 0.0204721f $X=2.765 $Y=1.16 $X2=0 $Y2=0
cc_261 N_D_c_282_n N_C_c_321_n 0.0316565f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_262 N_D_M1016_g N_A_27_47#_c_363_n 0.0126173f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_263 N_D_M1016_g N_VPWR_c_537_n 0.00417809f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_264 N_D_M1016_g N_VPWR_c_545_n 0.00425094f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_265 N_D_M1016_g N_VPWR_c_534_n 0.00614772f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_266 N_D_c_282_n N_VGND_c_673_n 0.00311379f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_267 N_D_c_282_n N_VGND_c_675_n 0.00418433f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_268 N_D_c_282_n N_VGND_c_681_n 0.00596249f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_269 N_C_M1010_g N_A_27_47#_M1005_g 0.0338739f $X=3.185 $Y=1.985 $X2=0 $Y2=0
cc_270 N_C_M1010_g N_A_27_47#_c_363_n 0.012933f $X=3.185 $Y=1.985 $X2=0 $Y2=0
cc_271 C N_A_27_47#_c_357_n 0.0231705f $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_272 N_C_c_320_n N_A_27_47#_c_357_n 3.32159e-19 $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_273 N_C_c_320_n N_A_27_47#_c_358_n 0.0202449f $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_274 C N_A_27_47#_c_359_n 0.00811617f $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_275 N_C_c_321_n N_A_27_47#_c_359_n 0.0261739f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_276 N_C_M1010_g N_VPWR_c_538_n 0.00941682f $X=3.185 $Y=1.985 $X2=0 $Y2=0
cc_277 N_C_M1010_g N_VPWR_c_545_n 0.00425094f $X=3.185 $Y=1.985 $X2=0 $Y2=0
cc_278 N_C_M1010_g N_VPWR_c_534_n 0.00634388f $X=3.185 $Y=1.985 $X2=0 $Y2=0
cc_279 N_C_c_321_n N_VGND_c_675_n 0.00367119f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_280 N_C_c_321_n N_VGND_c_681_n 0.00582183f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_281 C A_652_47# 0.00500756f $X=3.37 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_282 N_A_27_47#_c_359_n N_A_832_21#_c_445_n 0.0346039f $X=3.815 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_M1005_g N_A_832_21#_M1015_g 0.0366942f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_363_n N_A_832_21#_M1015_g 0.015032f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_365_n N_A_832_21#_M1015_g 0.0151211f $X=4.405 $Y=1.915 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_355_n N_A_832_21#_c_446_n 0.0132138f $X=4.32 $Y=1.24 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_357_n N_A_832_21#_c_446_n 0.00119722f $X=3.815 $Y=1.16 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_358_n N_A_832_21#_c_446_n 0.0224341f $X=3.815 $Y=1.16 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_355_n N_A_832_21#_c_447_n 0.00569154f $X=4.32 $Y=1.24 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_365_n N_A_832_21#_c_447_n 0.021623f $X=4.405 $Y=1.915 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_355_n N_A_832_21#_c_448_n 0.0138054f $X=4.32 $Y=1.24 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_363_n N_A_832_21#_c_456_n 0.00759698f $X=4.32 $Y=2 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_363_n N_VPWR_M1009_d 0.00553685f $X=4.32 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_294 N_A_27_47#_c_363_n N_VPWR_M1002_d 0.00327016f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_363_n N_VPWR_M1012_d 0.005014f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_363_n N_VPWR_M1010_d 0.00710632f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_363_n N_VPWR_M1015_d 0.00437261f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_365_n N_VPWR_M1015_d 0.00897148f $X=4.405 $Y=1.915 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_363_n N_VPWR_c_535_n 0.0181288f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_363_n N_VPWR_c_536_n 0.0159625f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_363_n N_VPWR_c_537_n 0.0200362f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_302 N_A_27_47#_M1005_g N_VPWR_c_538_n 0.00327828f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_363_n N_VPWR_c_538_n 0.0222787f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_363_n N_VPWR_c_540_n 0.0102692f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_363_n N_VPWR_c_541_n 0.0077537f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_362_n N_VPWR_c_543_n 0.0179169f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_363_n N_VPWR_c_543_n 0.00244309f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_363_n N_VPWR_c_544_n 0.00848923f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_309 N_A_27_47#_c_363_n N_VPWR_c_545_n 0.0110602f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_310 N_A_27_47#_M1009_s N_VPWR_c_534_n 0.00226392f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_M1005_g N_VPWR_c_534_n 0.00616215f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_362_n N_VPWR_c_534_n 0.00991829f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_363_n N_VPWR_c_534_n 0.0767149f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_314 N_A_27_47#_M1005_g N_VPWR_c_551_n 0.00425094f $X=3.755 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_363_n N_VPWR_c_551_n 0.010089f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_363_n N_X_M1000_s 0.004392f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_363_n N_X_M1011_s 0.00439557f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_318 N_A_27_47#_c_363_n N_X_c_630_n 0.0151802f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_319 N_A_27_47#_c_363_n N_X_c_646_n 0.0396402f $X=4.32 $Y=2 $X2=0 $Y2=0
cc_320 N_A_27_47#_c_359_n N_VGND_c_675_n 0.00367119f $X=3.815 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_356_n N_VGND_c_677_n 0.0177247f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_322 N_A_27_47#_M1017_s N_VGND_c_681_n 0.00382897f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_356_n N_VGND_c_681_n 0.00987844f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_324 N_A_27_47#_c_359_n N_VGND_c_681_n 0.00582183f $X=3.815 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_A_832_21#_c_447_n N_A_N_M1014_g 0.00495664f $X=5.035 $Y=1.16 $X2=0
+ $Y2=0
cc_326 N_A_832_21#_c_449_n N_A_N_M1014_g 0.0164119f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A_832_21#_c_447_n N_A_N_M1006_g 0.0138718f $X=5.035 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_832_21#_c_455_n N_A_N_M1006_g 0.0167965f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_329 N_A_832_21#_c_447_n N_A_N_c_511_n 9.97711e-19 $X=5.035 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A_832_21#_c_448_n N_A_N_c_511_n 0.0210419f $X=5.035 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_832_21#_c_449_n N_A_N_c_511_n 8.93472e-19 $X=5.635 $Y=0.74 $X2=0
+ $Y2=0
cc_332 N_A_832_21#_c_455_n N_A_N_c_511_n 4.7524e-19 $X=5.635 $Y=2 $X2=0 $Y2=0
cc_333 N_A_832_21#_c_447_n N_A_N_c_512_n 0.0254402f $X=5.035 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_832_21#_c_448_n N_A_N_c_512_n 0.00131484f $X=5.035 $Y=1.16 $X2=0
+ $Y2=0
cc_335 N_A_832_21#_c_449_n N_A_N_c_512_n 0.026727f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A_832_21#_c_455_n N_A_N_c_512_n 0.0182316f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_337 N_A_832_21#_c_455_n N_VPWR_M1015_d 0.00283287f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_338 N_A_832_21#_c_456_n N_VPWR_M1015_d 0.00230774f $X=5.12 $Y=2 $X2=0 $Y2=0
cc_339 N_A_832_21#_c_456_n N_VPWR_c_539_n 0.0142055f $X=5.12 $Y=2 $X2=0 $Y2=0
cc_340 N_A_832_21#_M1015_g N_VPWR_c_540_n 0.00923307f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_832_21#_c_455_n N_VPWR_c_546_n 0.00363176f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_342 N_A_832_21#_c_488_p N_VPWR_c_546_n 0.01143f $X=5.72 $Y=2.3 $X2=0 $Y2=0
cc_343 N_A_832_21#_M1006_d N_VPWR_c_534_n 0.00368727f $X=5.585 $Y=2.065 $X2=0
+ $Y2=0
cc_344 N_A_832_21#_M1015_g N_VPWR_c_534_n 0.00730283f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_345 N_A_832_21#_c_455_n N_VPWR_c_534_n 0.00782241f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_346 N_A_832_21#_c_456_n N_VPWR_c_534_n 8.5692e-19 $X=5.12 $Y=2 $X2=0 $Y2=0
cc_347 N_A_832_21#_c_488_p N_VPWR_c_534_n 0.00643448f $X=5.72 $Y=2.3 $X2=0 $Y2=0
cc_348 N_A_832_21#_M1015_g N_VPWR_c_551_n 0.00425094f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_832_21#_c_455_n N_VPWR_c_552_n 0.0189398f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_350 N_A_832_21#_c_450_n N_VGND_M1014_s 0.00117425f $X=5.12 $Y=0.74 $X2=0
+ $Y2=0
cc_351 N_A_832_21#_c_445_n N_VGND_c_674_n 0.00229482f $X=4.235 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A_832_21#_c_448_n N_VGND_c_674_n 7.23671e-19 $X=5.035 $Y=1.16 $X2=0
+ $Y2=0
cc_353 N_A_832_21#_c_449_n N_VGND_c_674_n 0.0129893f $X=5.635 $Y=0.74 $X2=0
+ $Y2=0
cc_354 N_A_832_21#_c_450_n N_VGND_c_674_n 0.0111742f $X=5.12 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A_832_21#_c_445_n N_VGND_c_675_n 0.00368502f $X=4.235 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_832_21#_c_450_n N_VGND_c_675_n 4.7797e-19 $X=5.12 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A_832_21#_c_449_n N_VGND_c_680_n 0.005481f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A_832_21#_c_504_p N_VGND_c_680_n 0.011459f $X=5.72 $Y=0.42 $X2=0 $Y2=0
cc_359 N_A_832_21#_M1014_d N_VGND_c_681_n 0.00370147f $X=5.585 $Y=0.235 $X2=0
+ $Y2=0
cc_360 N_A_832_21#_c_445_n N_VGND_c_681_n 0.006734f $X=4.235 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_832_21#_c_449_n N_VGND_c_681_n 0.00927486f $X=5.635 $Y=0.74 $X2=0
+ $Y2=0
cc_362 N_A_832_21#_c_450_n N_VGND_c_681_n 0.00152708f $X=5.12 $Y=0.74 $X2=0
+ $Y2=0
cc_363 N_A_832_21#_c_504_p N_VGND_c_681_n 0.00644035f $X=5.72 $Y=0.42 $X2=0
+ $Y2=0
cc_364 N_A_N_M1006_g N_VPWR_c_546_n 0.00425094f $X=5.51 $Y=2.275 $X2=0 $Y2=0
cc_365 N_A_N_M1006_g N_VPWR_c_534_n 0.00807745f $X=5.51 $Y=2.275 $X2=0 $Y2=0
cc_366 N_A_N_M1006_g N_VPWR_c_552_n 0.0106802f $X=5.51 $Y=2.275 $X2=0 $Y2=0
cc_367 N_A_N_M1014_g N_VGND_c_674_n 0.00943588f $X=5.51 $Y=0.445 $X2=0 $Y2=0
cc_368 N_A_N_M1014_g N_VGND_c_680_n 0.00428022f $X=5.51 $Y=0.445 $X2=0 $Y2=0
cc_369 N_A_N_M1014_g N_VGND_c_681_n 0.00821349f $X=5.51 $Y=0.445 $X2=0 $Y2=0
cc_370 N_VPWR_c_534_n N_X_M1000_s 0.00315309f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_371 N_VPWR_c_534_n N_X_M1011_s 0.00315309f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_M1002_d N_X_c_646_n 0.0036439f $X=1.44 $Y=1.485 $X2=0 $Y2=0
cc_373 N_X_c_634_n N_VGND_M1003_s 0.0033771f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_374 N_X_c_634_n N_VGND_c_672_n 0.0152323f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_375 N_X_c_660_p N_VGND_c_678_n 0.0113958f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_376 N_X_c_634_n N_VGND_c_678_n 0.00235782f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_377 X N_VGND_c_678_n 0.00151341f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_378 N_X_c_663_p N_VGND_c_679_n 0.0112485f $X=1.995 $Y=0.42 $X2=0 $Y2=0
cc_379 N_X_c_634_n N_VGND_c_679_n 0.00235782f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_380 N_X_M1001_d N_VGND_c_681_n 0.00251404f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_381 N_X_M1007_d N_VGND_c_681_n 0.00406917f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_382 N_X_c_660_p N_VGND_c_681_n 0.00646998f $X=1.155 $Y=0.42 $X2=0 $Y2=0
cc_383 N_X_c_663_p N_VGND_c_681_n 0.0064389f $X=1.995 $Y=0.42 $X2=0 $Y2=0
cc_384 N_X_c_634_n N_VGND_c_681_n 0.00972604f $X=1.91 $Y=0.735 $X2=0 $Y2=0
cc_385 X N_VGND_c_681_n 0.00292428f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_386 N_VGND_c_681_n A_556_47# 0.00268492f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_387 N_VGND_c_681_n A_652_47# 0.00342801f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_388 N_VGND_c_681_n A_766_47# 0.00268551f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24

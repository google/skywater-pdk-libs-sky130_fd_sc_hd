* File: sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2.spice.pex
* Created: Thu Aug 27 14:26:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%VGND 1 2 3 4 5 6 7 8
+ 37 51 55 59 63 67 71 75 79 90 93 96 99 102 104 105 130 140 147 162
c149 75 0 7.6696e-20 $X=5 $Y=0.42
r150 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=5.44
+ $X2=6.21 $Y2=5.44
r151 158 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=5.44
+ $X2=4.83 $Y2=5.44
r152 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r153 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=5.44
+ $X2=0.23 $Y2=5.44
r154 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r155 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r156 144 162 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=5.44
+ $X2=6.21 $Y2=5.44
r157 144 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=5.44
+ $X2=4.83 $Y2=5.44
r158 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=5.44
+ $X2=5.75 $Y2=5.44
r159 141 158 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.955 $Y=5.44
+ $X2=4.7 $Y2=5.44
r160 141 143 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.955 $Y=5.44
+ $X2=5.75 $Y2=5.44
r161 140 161 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=6.065 $Y=5.44
+ $X2=6.252 $Y2=5.44
r162 140 143 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.065 $Y=5.44
+ $X2=5.75 $Y2=5.44
r163 139 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r164 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r165 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r166 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r167 133 159 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=5.44
+ $X2=4.83 $Y2=5.44
r168 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=5.44
+ $X2=4.37 $Y2=5.44
r169 130 158 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.445 $Y=5.44
+ $X2=4.7 $Y2=5.44
r170 130 132 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.445 $Y=5.44
+ $X2=4.37 $Y2=5.44
r171 129 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r172 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r173 126 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=5.44
+ $X2=4.37 $Y2=5.44
r174 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=5.44
+ $X2=3.45 $Y2=5.44
r175 123 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r176 123 156 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r177 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r178 120 155 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0
+ $X2=2.185 $Y2=0
r179 120 122 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.99
+ $Y2=0
r180 119 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=5.44
+ $X2=3.45 $Y2=5.44
r181 118 119 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=5.44
+ $X2=2.53 $Y2=5.44
r182 116 119 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=5.44
+ $X2=2.53 $Y2=5.44
r183 115 118 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=5.44
+ $X2=2.53 $Y2=5.44
r184 115 116 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=5.44
+ $X2=0.69 $Y2=5.44
r185 113 152 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=5.44
+ $X2=0.187 $Y2=5.44
r186 113 115 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=5.44
+ $X2=0.69 $Y2=5.44
r187 112 156 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r188 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r189 109 149 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r190 109 111 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.69 $Y2=0
r191 108 155 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=0
+ $X2=2.185 $Y2=0
r192 108 111 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=2.02 $Y=0
+ $X2=0.69 $Y2=0
r193 105 112 0.0554856 $w=4.8e-07 $l=1.95e-07 $layer=MET1_cond $X=0.495 $Y=0
+ $X2=0.69 $Y2=0
r194 105 150 0.0754035 $w=4.8e-07 $l=2.65e-07 $layer=MET1_cond $X=0.495 $Y=0
+ $X2=0.23 $Y2=0
r195 104 116 0.0825171 $w=4.8e-07 $l=2.9e-07 $layer=MET1_cond $X=0.4 $Y=5.44
+ $X2=0.69 $Y2=5.44
r196 104 153 0.0483721 $w=4.8e-07 $l=1.7e-07 $layer=MET1_cond $X=0.4 $Y=5.44
+ $X2=0.23 $Y2=5.44
r197 102 138 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.75 $Y2=0
r198 102 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.99 $Y2=0
r199 101 146 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=6.155 $Y=0
+ $X2=6.21 $Y2=0
r200 101 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=0
+ $X2=5.99 $Y2=0
r201 99 135 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.83
+ $Y2=0
r202 99 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r203 98 138 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.75 $Y2=0
r204 98 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r205 96 128 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=0
+ $X2=3.91 $Y2=0
r206 96 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.14
+ $Y2=0
r207 95 135 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.305 $Y=0
+ $X2=4.83 $Y2=0
r208 95 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.14
+ $Y2=0
r209 93 125 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=5.44
+ $X2=3.45 $Y2=5.44
r210 93 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.575 $Y=5.44
+ $X2=3.67 $Y2=5.44
r211 92 132 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.765 $Y=5.44
+ $X2=4.37 $Y2=5.44
r212 92 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.765 $Y=5.44
+ $X2=3.67 $Y2=5.44
r213 90 122 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=0
+ $X2=2.99 $Y2=0
r214 90 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.28
+ $Y2=0
r215 89 128 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.91 $Y2=0
r216 89 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.28
+ $Y2=0
r217 87 118 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.645 $Y=5.44
+ $X2=2.53 $Y2=5.44
r218 87 88 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.645 $Y=5.44
+ $X2=2.775 $Y2=5.44
r219 86 125 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.905 $Y=5.44
+ $X2=3.45 $Y2=5.44
r220 86 88 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.905 $Y=5.44
+ $X2=2.775 $Y2=5.44
r221 81 161 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.21 $Y=5.355
+ $X2=6.252 $Y2=5.44
r222 77 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0
r223 77 79 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0.42
r224 73 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r225 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.42
r226 69 158 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=5.355
+ $X2=4.7 $Y2=5.44
r227 69 71 14.5406 $w=5.08e-07 $l=6.2e-07 $layer=LI1_cond $X=4.7 $Y=5.355
+ $X2=4.7 $Y2=4.735
r228 65 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r229 65 67 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.42
r230 61 94 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=5.355
+ $X2=3.67 $Y2=5.44
r231 61 63 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=3.67 $Y=5.355
+ $X2=3.67 $Y2=4.735
r232 57 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0
r233 57 59 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0.42
r234 53 88 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=5.355
+ $X2=2.775 $Y2=5.44
r235 53 55 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=2.775 $Y=5.355
+ $X2=2.775 $Y2=4.7
r236 49 155 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0
r237 49 51 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0.62
r238 44 152 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=5.355
+ $X2=0.187 $Y2=5.44
r239 39 149 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.187 $Y2=0
r240 37 81 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=6.21 $Y=4.8
+ $X2=6.21 $Y2=5.355
r241 37 44 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=0.23 $Y=4.8
+ $X2=0.23 $Y2=5.355
r242 37 39 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=0.23 $Y=0.64
+ $X2=0.23 $Y2=0.085
r243 8 79 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.85
+ $Y=0.235 $X2=5.99 $Y2=0.42
r244 7 75 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=0.235 $X2=5 $Y2=0.42
r245 6 71 45.5 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=4 $X=4.39
+ $Y=4.555 $X2=4.87 $Y2=4.735
r246 5 67 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.235 $X2=4.14 $Y2=0.42
r247 4 63 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.53 $Y=4.555
+ $X2=3.67 $Y2=4.735
r248 3 59 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.135
+ $Y=0.235 $X2=3.28 $Y2=0.42
r249 2 55 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.685
+ $Y=4.555 $X2=2.81 $Y2=4.7
r250 1 51 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.41 $X2=2.245 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%VPB 7 8 11 15 17 20 23
+ 28 34
r85 20 34 0.00371286 $w=1.4e-07 $l=3e-09 $layer=MET1_cond $X=0.557 $Y=3.57
+ $X2=0.56 $Y2=3.57
r86 18 28 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=6.21 $Y=3.57 $X2=6.21
+ $Y2=3.29
r87 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.155 $Y=3.57
+ $X2=6.155 $Y2=3.57
r88 15 34 6.74504 $w=1.4e-07 $l=5.45e-06 $layer=MET1_cond $X=6.01 $Y=3.57
+ $X2=0.56 $Y2=3.57
r89 15 17 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.01 $Y=3.57
+ $X2=6.155 $Y2=3.57
r90 14 23 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=0.23 $Y=3.57 $X2=0.23
+ $Y2=3.29
r91 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.225 $Y=3.57
+ $X2=0.225 $Y2=3.57
r92 11 20 0.231435 $w=1.4e-07 $l=1.87e-07 $layer=MET1_cond $X=0.37 $Y=3.57
+ $X2=0.557 $Y2=3.57
r93 11 13 0.0980892 $w=2.27e-07 $l=1.45e-07 $layer=MET1_cond $X=0.37 $Y=3.57
+ $X2=0.225 $Y2=3.57
r94 8 28 91 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=6.125 $Y=3.04 $X2=6.21 $Y2=3.29
r95 7 23 91 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=0.145 $Y=3.04 $X2=0.23 $Y2=3.29
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%LOWLVPWR 1 7 11 16 17
+ 20 25 26 30 32 34
c58 25 0 2.86228e-19 $X=2.225 $Y=2.2
r59 30 32 1.10767 $w=1.4e-07 $l=8.95e-07 $layer=MET1_cond $X=1.36 $Y=2.21
+ $X2=0.465 $Y2=2.21
r60 26 34 2.07418 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.2
+ $X2=2.06 $Y2=2.2
r61 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.225 $Y=2.2
+ $X2=2.225 $Y2=2.2
r62 23 34 23.6891 $w=2.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.505 $Y=2.2
+ $X2=2.06 $Y2=2.2
r63 22 25 0.461955 $w=2.3e-07 $l=7.2e-07 $layer=MET1_cond $X=1.505 $Y=2.2
+ $X2=2.225 $Y2=2.2
r64 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.505 $Y=2.2
+ $X2=1.505 $Y2=2.2
r65 20 30 0.0864037 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=1.475 $Y=2.2
+ $X2=1.36 $Y2=2.2
r66 20 22 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=1.475 $Y=2.2
+ $X2=1.505 $Y2=2.2
r67 16 17 17.048 $w=7.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.435 $Y=3.49
+ $X2=2.435 $Y2=2.66
r68 13 26 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.225 $Y=2.335
+ $X2=2.225 $Y2=2.2
r69 13 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.225 $Y=2.335
+ $X2=2.225 $Y2=2.66
r70 9 26 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=2.2
r71 9 11 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=1.79
r72 7 16 91 $w=1.7e-07 $l=6.45697e-07 $layer=licon1_NTAP_notbjt $count=2 $X=2.1
+ $Y=3.27 $X2=2.645 $Y2=3.49
r73 1 11 300 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_PDIFF $count=2 $X=2.1
+ $Y=1.485 $X2=2.225 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%A_505_297# 1 2 7 9 10
+ 12 13 14 15 17 18 20 22 28 31 35 36 39 40
c84 40 0 1.64106e-19 $X=3.225 $Y=3.84
c85 39 0 1.09489e-19 $X=3.225 $Y=3.84
r86 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=3.84 $X2=3.225 $Y2=3.84
r87 37 39 51.3361 $w=3.28e-07 $l=1.47e-06 $layer=LI1_cond $X=3.225 $Y=2.37
+ $X2=3.225 $Y2=3.84
r88 35 37 7.03987 $w=2.4e-07 $l=2.16852e-07 $layer=LI1_cond $X=3.06 $Y=2.25
+ $X2=3.225 $Y2=2.37
r89 35 36 12.4848 $w=2.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.06 $Y=2.25 $X2=2.8
+ $Y2=2.25
r90 31 34 56.1816 $w=2.38e-07 $l=1.17e-06 $layer=LI1_cond $X=2.68 $Y=0.62
+ $X2=2.68 $Y2=1.79
r91 29 36 6.81649 $w=2.4e-07 $l=1.69706e-07 $layer=LI1_cond $X=2.68 $Y=2.13
+ $X2=2.8 $Y2=2.25
r92 29 34 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.68 $Y=2.13
+ $X2=2.68 $Y2=1.79
r93 26 40 80.7859 $w=3.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.235 $Y=4.33
+ $X2=3.235 $Y2=3.84
r94 26 27 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.235 $Y=4.405
+ $X2=3.455 $Y2=4.405
r95 23 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.025 $Y=4.405
+ $X2=3.235 $Y2=4.405
r96 20 22 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.315 $Y=4.48
+ $X2=4.315 $Y2=4.88
r97 19 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.96 $Y=4.405
+ $X2=3.885 $Y2=4.405
r98 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.24 $Y=4.405
+ $X2=4.315 $Y2=4.48
r99 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.24 $Y=4.405
+ $X2=3.96 $Y2=4.405
r100 15 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.885 $Y=4.48
+ $X2=3.885 $Y2=4.405
r101 15 17 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.885 $Y=4.48
+ $X2=3.885 $Y2=4.88
r102 14 27 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.53 $Y=4.405
+ $X2=3.455 $Y2=4.405
r103 13 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.81 $Y=4.405
+ $X2=3.885 $Y2=4.405
r104 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.81 $Y=4.405
+ $X2=3.53 $Y2=4.405
r105 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.455 $Y=4.48
+ $X2=3.455 $Y2=4.405
r106 10 12 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.455 $Y=4.48
+ $X2=3.455 $Y2=4.88
r107 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.025 $Y=4.48
+ $X2=3.025 $Y2=4.405
r108 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.025 $Y=4.48 $X2=3.025
+ $Y2=4.88
r109 2 34 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=2.525
+ $Y=1.485 $X2=2.675 $Y2=1.79
r110 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.41 $X2=2.675 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%A_714_47# 1 2 3 10 11
+ 14 19 22 23 24 28 29 30 31 34 38 45
c103 28 0 1.64375e-19 $X=4.105 $Y=2.07
c104 14 0 7.6696e-20 $X=4.78 $Y=1.955
c105 11 0 1.09489e-19 $X=4.27 $Y=2.58
c106 10 0 1.90316e-19 $X=4.705 $Y=2.58
r107 43 45 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.765 $Y=2.49
+ $X2=4.105 $Y2=2.49
r108 40 42 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=3.71 $Y=0.855
+ $X2=4.105 $Y2=0.855
r109 36 38 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=4.57 $Y=0.73
+ $X2=4.57 $Y2=0.42
r110 32 34 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.555 $Y=3.47
+ $X2=4.555 $Y2=3.235
r111 31 42 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.855
+ $X2=4.105 $Y2=0.855
r112 30 36 6.98266 $w=2.5e-07 $l=1.65831e-07 $layer=LI1_cond $X=4.475 $Y=0.855
+ $X2=4.57 $Y2=0.73
r113 30 31 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.475 $Y=0.855
+ $X2=4.19 $Y2=0.855
r114 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.105
+ $Y=2.07 $X2=4.105 $Y2=2.07
r115 26 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=2.405
+ $X2=4.105 $Y2=2.49
r116 26 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.105 $Y=2.405
+ $X2=4.105 $Y2=2.07
r117 25 42 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.105 $Y=0.98
+ $X2=4.105 $Y2=0.855
r118 25 28 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.105 $Y=0.98
+ $X2=4.105 $Y2=2.07
r119 23 32 9.70995 $w=1.99e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.39 $Y=3.555
+ $X2=4.555 $Y2=3.47
r120 23 24 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.39 $Y=3.555
+ $X2=3.85 $Y2=3.555
r121 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=3.47
+ $X2=3.85 $Y2=3.555
r122 21 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=2.575
+ $X2=3.765 $Y2=2.49
r123 21 22 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.765 $Y=2.575
+ $X2=3.765 $Y2=3.47
r124 17 40 2.34666 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.71 $Y=0.73
+ $X2=3.71 $Y2=0.855
r125 17 19 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=3.71 $Y=0.73
+ $X2=3.71 $Y2=0.42
r126 16 29 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=4.105 $Y=2.505
+ $X2=4.105 $Y2=2.07
r127 12 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.78 $Y=2.505
+ $X2=4.78 $Y2=1.955
r128 11 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.27 $Y=2.58
+ $X2=4.105 $Y2=2.505
r129 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.705 $Y=2.58
+ $X2=4.78 $Y2=2.505
r130 10 11 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=2.58
+ $X2=4.27 $Y2=2.58
r131 3 34 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=3.09 $X2=4.555 $Y2=3.235
r132 2 38 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.43
+ $Y=0.235 $X2=4.57 $Y2=0.42
r133 1 19 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.57
+ $Y=0.235 $X2=3.71 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%A 3 5 7 8 12 14 15 18
+ 20 24 26 30 32 33 34 35 39
c71 15 0 1.64375e-19 $X=3.63 $Y=1.145
r72 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.25 $X2=3.125 $Y2=1.25
r73 35 39 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=3.13 $Y=1.425
+ $X2=3.13 $Y2=1.25
r74 28 30 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.785 $Y=1.07
+ $X2=4.785 $Y2=0.56
r75 27 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.43 $Y=1.145
+ $X2=4.355 $Y2=1.145
r76 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.71 $Y=1.145
+ $X2=4.785 $Y2=1.07
r77 26 27 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.71 $Y=1.145
+ $X2=4.43 $Y2=1.145
r78 22 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.355 $Y=1.07
+ $X2=4.355 $Y2=1.145
r79 22 24 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.355 $Y=1.07
+ $X2=4.355 $Y2=0.56
r80 21 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4 $Y=1.145 $X2=3.925
+ $Y2=1.145
r81 20 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.28 $Y=1.145
+ $X2=4.355 $Y2=1.145
r82 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.28 $Y=1.145 $X2=4
+ $Y2=1.145
r83 16 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=1.07
+ $X2=3.925 $Y2=1.145
r84 16 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.925 $Y=1.07
+ $X2=3.925 $Y2=0.56
r85 14 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.85 $Y=1.145
+ $X2=3.925 $Y2=1.145
r86 14 15 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.85 $Y=1.145
+ $X2=3.63 $Y2=1.145
r87 10 15 33.8325 $w=2.41e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.63 $Y2=1.145
r88 10 38 74 $w=2.41e-07 $l=4.75857e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.125 $Y2=1.312
r89 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.495 $Y2=0.56
r90 9 32 4.83878 $w=1.55e-07 $l=9.38083e-08 $layer=POLY_cond $X=2.535 $Y=1.147
+ $X2=2.455 $Y2=1.117
r91 8 38 39.1212 $w=2.41e-07 $l=2.33345e-07 $layer=POLY_cond $X=2.96 $Y=1.147
+ $X2=3.125 $Y2=1.312
r92 8 9 203.325 $w=1.55e-07 $l=4.25e-07 $layer=POLY_cond $X=2.96 $Y=1.147
+ $X2=2.535 $Y2=1.147
r93 5 32 20.9729 $w=1.5e-07 $l=1.09471e-07 $layer=POLY_cond $X=2.46 $Y=1.01
+ $X2=2.455 $Y2=1.117
r94 5 7 125.32 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.46 $Y=1.01 $X2=2.46
+ $Y2=0.62
r95 1 32 20.9729 $w=1.5e-07 $l=1.10472e-07 $layer=POLY_cond $X=2.45 $Y=1.225
+ $X2=2.455 $Y2=1.117
r96 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.45 $Y=1.225 $X2=2.45
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%A_620_911# 1 2 3 10 11
+ 12 17 18 20 24 29 31 32 34 38 40 41 44 48 49 53 56 57 60 62 63
c126 60 0 1.02426e-19 $X=4.555 $Y=1.79
c127 44 0 7.14482e-20 $X=4.1 $Y=4.735
c128 38 0 9.26578e-20 $X=3.24 $Y=4.735
c129 31 0 8.23968e-20 $X=4.78 $Y=2.94
c130 24 0 9.10198e-20 $X=5.085 $Y=4.88
c131 18 0 1.25592e-19 $X=5.16 $Y=2.94
c132 11 0 1.76914e-21 $X=4.27 $Y=2.94
c133 10 0 7.64702e-20 $X=4.705 $Y=2.94
r134 58 60 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.555 $Y=2.745
+ $X2=4.555 $Y2=1.79
r135 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.47 $Y=2.83
+ $X2=4.555 $Y2=2.745
r136 56 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.47 $Y=2.83
+ $X2=4.19 $Y2=2.83
r137 54 63 10.0555 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.105 $Y=4.045
+ $X2=4.105 $Y2=3.97
r138 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=3.975 $X2=4.105 $Y2=3.975
r139 51 62 3.70735 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.105 $Y=4.155
+ $X2=3.935 $Y2=4.155
r140 51 53 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.105 $Y=4.155
+ $X2=4.105 $Y2=3.975
r141 49 63 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=4.105 $Y=3.135
+ $X2=4.105 $Y2=3.97
r142 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=3.135 $X2=4.105 $Y2=3.135
r143 46 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=2.915
+ $X2=4.19 $Y2=2.83
r144 46 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.105 $Y=2.915
+ $X2=4.105 $Y2=3.135
r145 42 62 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=4.1 $Y=4.325
+ $X2=3.935 $Y2=4.155
r146 42 44 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.1 $Y=4.325
+ $X2=4.1 $Y2=4.735
r147 40 62 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=4.24
+ $X2=3.935 $Y2=4.155
r148 40 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.935 $Y=4.24
+ $X2=3.405 $Y2=4.24
r149 36 41 17.4739 $w=1.11e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.24 $Y=4.325
+ $X2=3.405 $Y2=4.24
r150 36 38 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.24 $Y=4.325
+ $X2=3.24 $Y2=4.735
r151 33 34 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.085 $Y=4.045
+ $X2=5.235 $Y2=4.045
r152 30 49 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=4.105 $Y=3.015
+ $X2=4.105 $Y2=3.135
r153 27 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.235 $Y=3.97
+ $X2=5.235 $Y2=4.045
r154 27 29 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.235 $Y=3.97
+ $X2=5.235 $Y2=3.485
r155 26 29 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.235 $Y=3.015
+ $X2=5.235 $Y2=3.485
r156 22 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.085 $Y=4.12
+ $X2=5.085 $Y2=4.045
r157 22 24 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.085 $Y=4.12
+ $X2=5.085 $Y2=4.88
r158 21 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=4.045
+ $X2=4.78 $Y2=4.045
r159 20 33 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.01 $Y=4.045
+ $X2=5.085 $Y2=4.045
r160 20 21 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.01 $Y=4.045
+ $X2=4.855 $Y2=4.045
r161 19 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=2.94
+ $X2=4.78 $Y2=2.94
r162 18 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.16 $Y=2.94
+ $X2=5.235 $Y2=3.015
r163 18 19 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=5.16 $Y=2.94
+ $X2=4.855 $Y2=2.94
r164 15 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=3.97
+ $X2=4.78 $Y2=4.045
r165 15 17 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.78 $Y=3.97
+ $X2=4.78 $Y2=3.485
r166 14 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=3.015
+ $X2=4.78 $Y2=2.94
r167 14 17 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.78 $Y=3.015 $X2=4.78
+ $Y2=3.485
r168 13 54 22.122 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=4.045
+ $X2=4.105 $Y2=4.045
r169 12 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=4.045
+ $X2=4.78 $Y2=4.045
r170 12 13 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=4.045
+ $X2=4.27 $Y2=4.045
r171 11 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.27 $Y=2.94
+ $X2=4.105 $Y2=3.015
r172 10 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=2.94
+ $X2=4.78 $Y2=2.94
r173 10 11 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=2.94
+ $X2=4.27 $Y2=2.94
r174 3 60 300 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.56 $X2=4.555 $Y2=1.79
r175 2 44 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.96 $Y=4.555
+ $X2=4.1 $Y2=4.735
r176 1 38 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.1 $Y=4.555
+ $X2=3.24 $Y2=4.735
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%A_1032_911# 1 2 9 11
+ 13 14 18 23 24 25 28 32 35 38
c69 28 0 9.10198e-20 $X=5.455 $Y=3.235
c70 11 0 1.02426e-19 $X=5.255 $Y=1.41
r71 35 37 12.4159 $w=4.52e-07 $l=4.6e-07 $layer=LI1_cond $X=5.45 $Y=4.24
+ $X2=5.45 $Y2=4.7
r72 33 38 19.468 $w=3.59e-07 $l=1.45e-07 $layer=POLY_cond $X=5.92 $Y=4.195
+ $X2=5.775 $Y2=4.195
r73 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.92
+ $Y=4.21 $X2=5.92 $Y2=4.21
r74 30 35 4.69682 $w=2.3e-07 $l=3.15e-07 $layer=LI1_cond $X=5.765 $Y=4.24
+ $X2=5.45 $Y2=4.24
r75 30 32 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.765 $Y=4.24
+ $X2=5.92 $Y2=4.24
r76 26 35 7.30083 $w=4.52e-07 $l=1.17473e-07 $layer=LI1_cond $X=5.455 $Y=4.125
+ $X2=5.45 $Y2=4.24
r77 26 28 51.9522 $w=1.88e-07 $l=8.9e-07 $layer=LI1_cond $X=5.455 $Y=4.125
+ $X2=5.455 $Y2=3.235
r78 21 38 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.775 $Y=4.015
+ $X2=5.775 $Y2=4.195
r79 21 23 1040.91 $w=1.5e-07 $l=2.03e-06 $layer=POLY_cond $X=5.775 $Y=4.015
+ $X2=5.775 $Y2=1.985
r80 20 25 36.6911 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=5.775 $Y=1.41
+ $X2=5.775 $Y2=1.247
r81 20 23 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.775 $Y=1.41
+ $X2=5.775 $Y2=1.985
r82 16 25 36.6911 $w=1.5e-07 $l=1.62e-07 $layer=POLY_cond $X=5.775 $Y=1.085
+ $X2=5.775 $Y2=1.247
r83 16 18 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.775 $Y=1.085
+ $X2=5.775 $Y2=0.56
r84 15 24 4.85217 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=5.33 $Y=1.247
+ $X2=5.255 $Y2=1.247
r85 14 25 4.85217 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=5.7 $Y=1.247
+ $X2=5.775 $Y2=1.247
r86 14 15 65.694 $w=3.25e-07 $l=3.7e-07 $layer=POLY_cond $X=5.7 $Y=1.247
+ $X2=5.33 $Y2=1.247
r87 11 24 36.6911 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=5.255 $Y=1.41
+ $X2=5.255 $Y2=1.247
r88 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.255 $Y=1.41
+ $X2=5.255 $Y2=1.985
r89 7 24 36.6911 $w=1.5e-07 $l=1.62e-07 $layer=POLY_cond $X=5.255 $Y=1.085
+ $X2=5.255 $Y2=1.247
r90 7 9 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.255 $Y=1.085
+ $X2=5.255 $Y2=0.56
r91 2 28 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.31
+ $Y=3.09 $X2=5.455 $Y2=3.235
r92 1 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.16
+ $Y=4.555 $X2=5.3 $Y2=4.7
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%VPWR 1 2 3 12 16 20 23
+ 25 26 27 34 41 42 49
c86 23 0 1.90316e-19 $X=5.005 $Y=2.72
r87 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r88 39 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r89 39 49 0.611765 $w=4.8e-07 $l=2.15e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.6 $Y2=2.72
r90 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r91 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r92 31 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 30 34 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 27 49 0.13658 $w=4.8e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=2.72 $X2=3.6
+ $Y2=2.72
r96 27 35 0.429658 $w=4.8e-07 $l=1.51e-06 $layer=MET1_cond $X=3.12 $Y=2.72
+ $X2=1.61 $Y2=2.72
r97 25 38 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=5.75 $Y2=2.72
r98 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=5.99 $Y2=2.72
r99 24 41 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=6.21 $Y2=2.72
r100 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=2.72
+ $X2=5.99 $Y2=2.72
r101 22 38 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=5.75 $Y2=2.72
r102 22 23 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=5.005 $Y2=2.72
r103 18 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=2.635
+ $X2=5.99 $Y2=2.72
r104 18 20 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.99 $Y=2.635
+ $X2=5.99 $Y2=1.79
r105 14 23 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.805
+ $X2=5.005 $Y2=2.72
r106 14 16 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.005 $Y=2.805
+ $X2=5.005 $Y2=3.235
r107 10 23 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.635
+ $X2=5.005 $Y2=2.72
r108 10 12 42.3398 $w=2.28e-07 $l=8.45e-07 $layer=LI1_cond $X=5.005 $Y=2.635
+ $X2=5.005 $Y2=1.79
r109 3 20 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=5.85
+ $Y=1.485 $X2=5.99 $Y2=1.79
r110 2 12 300 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.56 $X2=5.005 $Y2=1.79
r111 1 16 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=3.09 $X2=5.005 $Y2=3.235
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_ISOWELL_TAP_2%X 1 2 9 11 12 18
r23 18 26 3.14303 $w=2.73e-07 $l=7.5e-08 $layer=LI1_cond $X=5.497 $Y=1.055
+ $X2=5.497 $Y2=0.98
r24 12 23 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=5.497 $Y=1.425
+ $X2=5.497 $Y2=1.79
r25 11 26 0.293093 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=5.485 $Y=0.975
+ $X2=5.485 $Y2=0.98
r26 11 12 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=5.497 $Y=1.06
+ $X2=5.497 $Y2=1.425
r27 11 18 0.209535 $w=2.73e-07 $l=5e-09 $layer=LI1_cond $X=5.497 $Y=1.06
+ $X2=5.497 $Y2=1.055
r28 7 11 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=5.485 $Y=0.83
+ $X2=5.485 $Y2=0.975
r29 7 9 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=5.485 $Y=0.83
+ $X2=5.485 $Y2=0.42
r30 2 23 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=5.33
+ $Y=1.485 $X2=5.47 $Y2=1.79
r31 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.33
+ $Y=0.235 $X2=5.47 $Y2=0.42
.ends


* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_4.pex.spice
* Created: Thu Aug 27 14:23:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%A 3 7 9 10 14
c37 14 0 2.23144e-19 $X=0.51 $Y=1.16
r38 14 17 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.495 $Y2=1.325
r39 14 16 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.495 $Y2=0.995
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r41 10 15 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.6 $Y=1.19 $X2=0.6
+ $Y2=1.16
r42 9 15 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.6 $Y=0.85 $X2=0.6
+ $Y2=1.16
r43 7 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r44 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%A_27_47# 1 2 9 13 17 21 25 29
+ 33 37 40 43 45 48 49 54 60 62 71
c114 49 0 1.51549e-19 $X=1.115 $Y=1.16
c115 48 0 2.75502e-19 $X=1.03 $Y=1.495
c116 25 0 1.24224e-19 $X=1.815 $Y=1.985
r117 71 72 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=2.245 $Y=1.157
+ $X2=2.25 $Y2=1.157
r118 68 69 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=1.815 $Y=1.157
+ $X2=1.82 $Y2=1.157
r119 67 68 74.7628 $w=2.74e-07 $l=4.25e-07 $layer=POLY_cond $X=1.39 $Y=1.157
+ $X2=1.815 $Y2=1.157
r120 66 67 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=1.385 $Y=1.157
+ $X2=1.39 $Y2=1.157
r121 63 64 0.879562 $w=2.74e-07 $l=5e-09 $layer=POLY_cond $X=0.955 $Y=1.157
+ $X2=0.96 $Y2=1.157
r122 57 60 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r123 55 71 57.1715 $w=2.74e-07 $l=3.25e-07 $layer=POLY_cond $X=1.92 $Y=1.157
+ $X2=2.245 $Y2=1.157
r124 55 69 17.5912 $w=2.74e-07 $l=1e-07 $layer=POLY_cond $X=1.92 $Y=1.157
+ $X2=1.82 $Y2=1.157
r125 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r126 52 66 25.5073 $w=2.74e-07 $l=1.45e-07 $layer=POLY_cond $X=1.24 $Y=1.157
+ $X2=1.385 $Y2=1.157
r127 52 64 49.2555 $w=2.74e-07 $l=2.8e-07 $layer=POLY_cond $X=1.24 $Y=1.157
+ $X2=0.96 $Y2=1.157
r128 51 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.24 $Y=1.16
+ $X2=1.92 $Y2=1.16
r129 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.24
+ $Y=1.16 $X2=1.24 $Y2=1.16
r130 49 51 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.115 $Y=1.16
+ $X2=1.24 $Y2=1.16
r131 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.03 $Y=1.245
+ $X2=1.115 $Y2=1.16
r132 47 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.03 $Y=1.245
+ $X2=1.03 $Y2=1.495
r133 46 62 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.355 $Y=1.58
+ $X2=0.22 $Y2=1.58
r134 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.945 $Y=1.58
+ $X2=1.03 $Y2=1.495
r135 45 46 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.945 $Y=1.58
+ $X2=0.355 $Y2=1.58
r136 41 62 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=1.58
r137 41 43 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=1.69
r138 40 62 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.17 $Y=1.495
+ $X2=0.22 $Y2=1.58
r139 39 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r140 39 40 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.495
r141 35 72 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=2.25 $Y=1.02
+ $X2=2.25 $Y2=1.157
r142 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.25 $Y=1.02
+ $X2=2.25 $Y2=0.445
r143 31 71 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=2.245 $Y=1.295
+ $X2=2.245 $Y2=1.157
r144 31 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.245 $Y=1.295
+ $X2=2.245 $Y2=1.985
r145 27 69 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=1.82 $Y=1.02
+ $X2=1.82 $Y2=1.157
r146 27 29 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.82 $Y=1.02
+ $X2=1.82 $Y2=0.445
r147 23 68 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=1.815 $Y=1.295
+ $X2=1.815 $Y2=1.157
r148 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.815 $Y=1.295
+ $X2=1.815 $Y2=1.985
r149 19 67 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=1.39 $Y=1.02
+ $X2=1.39 $Y2=1.157
r150 19 21 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.39 $Y=1.02
+ $X2=1.39 $Y2=0.445
r151 15 66 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=1.385 $Y=1.295
+ $X2=1.385 $Y2=1.157
r152 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.385 $Y=1.295
+ $X2=1.385 $Y2=1.985
r153 11 64 16.847 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=0.96 $Y=1.02
+ $X2=0.96 $Y2=1.157
r154 11 13 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.96 $Y=1.02
+ $X2=0.96 $Y2=0.445
r155 7 63 16.847 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=0.955 $Y=1.295
+ $X2=0.955 $Y2=1.157
r156 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.955 $Y=1.295
+ $X2=0.955 $Y2=1.985
r157 2 43 300 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.69
r158 1 60 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%KAPWR 1 2 3 12 18 19 22 23 24
+ 28 31 40 47
r56 28 47 0.00230263 $w=2e-07 $l=3e-09 $layer=MET1_cond $X=0.242 $Y=2.24
+ $X2=0.245 $Y2=2.24
r57 27 40 11.3222 $w=2.83e-07 $l=2.8e-07 $layer=LI1_cond $X=2.477 $Y=2.21
+ $X2=2.477 $Y2=1.93
r58 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.46 $Y=2.21
+ $X2=2.46 $Y2=2.21
r59 21 24 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.58 $Y=2.21
+ $X2=1.725 $Y2=2.21
r60 21 23 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=1.58 $Y=2.21
+ $X2=1.435 $Y2=2.21
r61 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.58 $Y=2.225
+ $X2=1.58 $Y2=2.225
r62 19 23 0.456689 $w=2e-07 $l=5.95e-07 $layer=MET1_cond $X=0.84 $Y=2.24
+ $X2=1.435 $Y2=2.24
r63 18 47 0.234101 $w=2e-07 $l=3.05e-07 $layer=MET1_cond $X=0.55 $Y=2.24
+ $X2=0.245 $Y2=2.24
r64 17 31 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.69 $Y=2.21
+ $X2=0.69 $Y2=2
r65 16 19 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.695 $Y=2.21
+ $X2=0.84 $Y2=2.21
r66 16 18 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.695 $Y=2.21
+ $X2=0.55 $Y2=2.21
r67 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=2.21
+ $X2=0.695 $Y2=2.21
r68 12 26 0.0784173 $w=2.46e-07 $l=1.59295e-07 $layer=MET1_cond $X=2.315 $Y=2.24
+ $X2=2.46 $Y2=2.21
r69 12 24 0.452852 $w=2e-07 $l=5.9e-07 $layer=MET1_cond $X=2.315 $Y=2.24
+ $X2=1.725 $Y2=2.24
r70 3 40 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.485 $X2=2.46 $Y2=1.93
r71 2 22 600 $w=1.7e-07 $l=9.02289e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.485 $X2=1.6 $Y2=2.32
r72 1 31 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%X 1 2 3 4 15 19 21 22 23 24 27
+ 34 35 36 37 47
c85 24 0 1.24224e-19 $X=1.39 $Y=1.857
c86 3 0 1.06215e-19 $X=1.03 $Y=1.485
r87 37 47 6.40246 $w=4.03e-07 $l=2.25e-07 $layer=LI1_cond $X=2.457 $Y=1.19
+ $X2=2.457 $Y2=1.415
r88 36 46 4.76257 $w=1.68e-07 $l=7.3e-08 $layer=LI1_cond $X=2.53 $Y=0.82
+ $X2=2.457 $Y2=0.82
r89 36 37 7.68295 $w=4.03e-07 $l=2.7e-07 $layer=LI1_cond $X=2.457 $Y=0.92
+ $X2=2.457 $Y2=1.19
r90 36 46 0.426831 $w=4.03e-07 $l=1.5e-08 $layer=LI1_cond $X=2.457 $Y=0.92
+ $X2=2.457 $Y2=0.905
r91 35 47 25.2481 $w=1.68e-07 $l=3.87e-07 $layer=LI1_cond $X=2.07 $Y=1.5
+ $X2=2.457 $Y2=1.5
r92 35 43 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.07 $Y=1.5
+ $X2=2.035 $Y2=1.5
r93 35 43 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=2.035 $Y=1.6
+ $X2=2.035 $Y2=1.585
r94 32 35 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=2.035 $Y=1.75
+ $X2=2.035 $Y2=1.6
r95 32 34 4.62773 $w=2.45e-07 $l=1.07e-07 $layer=LI1_cond $X=2.035 $Y=1.75
+ $X2=2.035 $Y2=1.857
r96 25 46 27.5316 $w=1.68e-07 $l=4.22e-07 $layer=LI1_cond $X=2.035 $Y=0.82
+ $X2=2.457 $Y2=0.82
r97 25 27 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=2.035 $Y=0.735
+ $X2=2.035 $Y2=0.51
r98 23 34 1.81688 $w=2.15e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=1.857
+ $X2=2.035 $Y2=1.857
r99 23 24 27.605 $w=2.13e-07 $l=5.15e-07 $layer=LI1_cond $X=1.905 $Y=1.857
+ $X2=1.39 $Y2=1.857
r100 21 25 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=0.82
+ $X2=2.035 $Y2=0.82
r101 21 22 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.905 $Y=0.82
+ $X2=1.305 $Y2=0.82
r102 17 24 13.9799 $w=2.15e-07 $l=2.54804e-07 $layer=LI1_cond $X=1.145 $Y=1.877
+ $X2=1.39 $Y2=1.857
r103 17 19 7.68295 $w=2.38e-07 $l=1.6e-07 $layer=LI1_cond $X=1.145 $Y=2.005
+ $X2=1.145 $Y2=2.165
r104 13 22 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.157 $Y=0.735
+ $X2=1.305 $Y2=0.82
r105 13 15 8.78982 $w=2.93e-07 $l=2.25e-07 $layer=LI1_cond $X=1.157 $Y=0.735
+ $X2=1.157 $Y2=0.51
r106 4 35 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.485 $X2=2.03 $Y2=1.62
r107 4 34 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=1.485 $X2=2.03 $Y2=1.96
r108 3 19 600 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.17 $Y2=2.165
r109 2 27 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.035 $Y2=0.51
r110 1 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.175 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%VGND 1 2 3 12 16 18 20 22 24 29
+ 34 40 43 47
r45 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r46 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r47 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r49 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r50 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r51 35 43 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.602
+ $Y2=0
r52 35 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=2.07
+ $Y2=0
r53 34 46 4.22854 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.547
+ $Y2=0
r54 34 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.07
+ $Y2=0
r55 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r56 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r57 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 30 40 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.692
+ $Y2=0
r59 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.15
+ $Y2=0
r60 29 43 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.602
+ $Y2=0
r61 29 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.15
+ $Y2=0
r62 24 40 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.692
+ $Y2=0
r63 24 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.23
+ $Y2=0
r64 22 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r65 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 18 46 3.13151 $w=2.8e-07 $l=1.15521e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.547 $Y2=0
r67 18 20 12.965 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.4
r68 14 43 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0
r69 14 16 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0.4
r70 10 40 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r71 10 12 13.2007 $w=2.73e-07 $l=3.15e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.4
r72 3 20 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.465 $Y2=0.4
r73 2 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.235 $X2=1.605 $Y2=0.4
r74 1 12 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%VPWR 1 8 9
r38 8 9 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72 $X2=2.53
+ $Y2=2.72
r39 4 8 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r40 1 9 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r41 1 4 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends


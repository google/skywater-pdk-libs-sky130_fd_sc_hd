* File: sky130_fd_sc_hd__nand2_2.pex.spice
* Created: Tue Sep  1 19:15:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND2_2%B 1 3 6 8 10 13 15 16 24
c45 16 0 1.81089e-19 $X=0.695 $Y=1.19
c46 8 0 9.09144e-20 $X=0.89 $Y=0.995
r47 22 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.68 $Y=1.16
+ $X2=0.89 $Y2=1.16
r48 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.68 $Y2=1.16
r49 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=1.16 $X2=0.68 $Y2=1.16
r50 15 16 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.235 $Y=1.2
+ $X2=0.68 $Y2=1.2
r51 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r52 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r53 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r54 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r55 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r56 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r57 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_2%A 1 3 6 8 10 13 15 16 24
c45 24 0 1.81089e-19 $X=1.73 $Y=1.16
c46 1 0 5.77853e-20 $X=1.31 $Y=0.995
r47 22 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.73 $Y2=1.16
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r49 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r50 16 23 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.2
+ $X2=1.52 $Y2=1.2
r51 15 23 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.2
+ $X2=1.52 $Y2=1.2
r52 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r54 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r56 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_2%VPWR 1 2 3 10 12 18 20 22 25 26 27 33 42
c35 3 0 1.4808e-19 $X=1.805 $Y=1.485
r36 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r39 33 41 3.96354 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=2.077 $Y2=2.72
r40 33 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r41 32 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 29 38 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r44 29 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 27 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 27 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r47 25 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72 $X2=1.1
+ $Y2=2.72
r49 24 35 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72 $X2=1.1
+ $Y2=2.72
r51 20 41 3.21368 $w=2.55e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.982 $Y=2.635
+ $X2=2.077 $Y2=2.72
r52 20 22 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=1.982 $Y=2.635
+ $X2=1.982 $Y2=2
r53 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r54 16 18 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r55 12 15 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r56 10 38 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r57 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r58 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r59 2 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r60 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r61 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_2%Y 1 2 3 10 12 14 16 22 24 29 30 31 32 38 39
c53 30 0 1.4808e-19 $X=2.075 $Y=0.85
c54 16 0 9.09144e-20 $X=1.935 $Y=0.78
r55 32 39 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=1.58
+ $X2=2.075 $Y2=1.495
r56 32 39 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.075 $Y=1.47
+ $X2=2.075 $Y2=1.495
r57 31 32 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=2.075 $Y=1.19
+ $X2=2.075 $Y2=1.47
r58 30 38 3.22874 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.78
+ $X2=2.075 $Y2=0.905
r59 30 31 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=2.075 $Y=0.92
+ $X2=2.075 $Y2=1.19
r60 30 38 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.075 $Y=0.92
+ $X2=2.075 $Y2=0.905
r61 25 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.58
+ $X2=1.52 $Y2=1.58
r62 24 32 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.935 $Y=1.58
+ $X2=2.075 $Y2=1.58
r63 24 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.935 $Y=1.58
+ $X2=1.685 $Y2=1.58
r64 20 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=1.58
r65 20 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=1.665
+ $X2=1.52 $Y2=2.34
r66 16 30 3.61619 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=1.935 $Y=0.78
+ $X2=2.075 $Y2=0.78
r67 16 18 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=1.935 $Y=0.78
+ $X2=1.52 $Y2=0.78
r68 15 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.58
+ $X2=0.68 $Y2=1.58
r69 14 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.58
+ $X2=1.52 $Y2=1.58
r70 14 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.58
+ $X2=0.845 $Y2=1.58
r71 10 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.665 $X2=0.68
+ $Y2=1.58
r72 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r73 3 29 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r74 3 22 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r75 2 27 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r76 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r77 1 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_2%A_27_47# 1 2 3 12 14 15 16 17 25 26
c42 25 0 5.77853e-20 $X=1.94 $Y=0.38
r43 25 26 8.37661 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0.37
+ $X2=1.775 $Y2=0.37
r44 19 21 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.185 $Y=0.36
+ $X2=1.06 $Y2=0.36
r45 19 26 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=1.185 $Y=0.36
+ $X2=1.775 $Y2=0.36
r46 17 23 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.715
+ $X2=1.06 $Y2=0.8
r47 16 21 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.06 $Y=0.465
+ $X2=1.06 $Y2=0.36
r48 16 17 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.06 $Y=0.465
+ $X2=1.06 $Y2=0.715
r49 14 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.935 $Y=0.8
+ $X2=1.06 $Y2=0.8
r50 14 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.8
+ $X2=0.425 $Y2=0.8
r51 10 15 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.425 $Y2=0.8
r52 10 12 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.38
r53 3 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r54 2 23 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.72
r55 2 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r56 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2_2%VGND 1 6 8 10 17 18 21
r32 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r33 18 22 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=0.69
+ $Y2=0
r34 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r35 15 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r36 15 17 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=0.765 $Y=0 $X2=2.07
+ $Y2=0
r37 10 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r38 10 12 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r39 8 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r40 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r41 4 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r42 4 6 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0.38
r43 1 6 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__dfsbp_2.spice.pex
* Created: Thu Aug 27 14:15:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFSBP_2%CLK 4 5 7 8 10 13 17 19 20 24 26
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r47 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.265 $Y=1.19
+ $X2=0.265 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_27_47# 1 2 9 13 15 17 20 24 28 31 35 36 37
+ 40 42 46 47 50 51 52 54 55 59 61 62 63 64 73 78 85 86 92 93 96
c273 92 0 3.28258e-19 $X=5.155 $Y=1.74
c274 86 0 3.30612e-20 $X=2.765 $Y=1.74
c275 85 0 2.53448e-20 $X=2.765 $Y=1.74
c276 73 0 1.81067e-19 $X=5.29 $Y=1.87
c277 63 0 1.39518e-19 $X=5.145 $Y=1.87
c278 61 0 1.01003e-19 $X=2.385 $Y=1.87
c279 52 0 3.16972e-20 $X=5.07 $Y=0.81
c280 51 0 1.753e-19 $X=5.82 $Y=0.81
c281 47 0 9.52104e-20 $X=2.435 $Y=0.87
c282 46 0 1.76471e-19 $X=2.435 $Y=0.87
c283 40 0 1.81794e-19 $X=0.725 $Y=1.795
c284 37 0 3.29888e-20 $X=0.61 $Y=1.88
c285 24 0 7.27138e-20 $X=5.065 $Y=2.275
r286 93 104 6.31985 $w=3.08e-07 $l=1.7e-07 $layer=LI1_cond $X=5.155 $Y=1.81
+ $X2=4.985 $Y2=1.81
r287 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.74 $X2=5.155 $Y2=1.74
r288 89 92 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.065 $Y=1.74
+ $X2=5.155 $Y2=1.74
r289 85 88 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.765 $Y=1.74
+ $X2=2.765 $Y2=1.875
r290 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.74 $X2=2.765 $Y2=1.74
r291 73 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r292 71 86 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.765 $Y2=1.765
r293 71 99 2.12292 $w=3.78e-07 $l=7e-08 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.46 $Y2=1.765
r294 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=1.87
r295 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=1.87
+ $X2=0.73 $Y2=1.87
r296 64 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.87
+ $X2=2.53 $Y2=1.87
r297 63 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r298 63 64 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=2.675 $Y2=1.87
r299 62 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=1.87
+ $X2=0.73 $Y2=1.87
r300 61 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=2.53 $Y2=1.87
r301 61 62 1.86881 $w=1.4e-07 $l=1.51e-06 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=0.875 $Y2=1.87
r302 59 96 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.985 $Y=0.93
+ $X2=5.985 $Y2=0.765
r303 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=0.93 $X2=5.985 $Y2=0.93
r304 55 58 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.985 $Y=0.81
+ $X2=5.985 $Y2=0.93
r305 51 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.985 $Y2=0.81
r306 51 52 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.07 $Y2=0.81
r307 50 104 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.985 $Y=1.655
+ $X2=4.985 $Y2=1.81
r308 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.985 $Y=0.895
+ $X2=5.07 $Y2=0.81
r309 49 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.985 $Y=0.895
+ $X2=4.985 $Y2=1.655
r310 47 80 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.435 $Y=0.87
+ $X2=2.305 $Y2=0.87
r311 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=0.87 $X2=2.435 $Y2=0.87
r312 44 99 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=1.765
r313 44 46 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=0.87
r314 43 78 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r315 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r316 40 67 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r317 40 42 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r318 39 42 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r319 38 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r320 37 67 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r321 37 38 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r322 35 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r323 35 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r324 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r325 29 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r326 28 96 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.045 $Y=0.445
+ $X2=6.045 $Y2=0.765
r327 22 89 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=1.74
r328 22 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=2.275
r329 20 88 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.875
r330 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r331 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r332 11 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r333 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r334 7 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r335 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r336 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r337 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%D 3 7 9 10 14 15
c39 14 0 1.34441e-19 $X=1.855 $Y=1.17
c40 7 0 1.76471e-19 $X=1.83 $Y=2.065
r41 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.335
r42 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.005
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.17 $X2=1.855 $Y2=1.17
r44 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.53
r45 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.17
r46 7 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.83 $Y=2.065
+ $X2=1.83 $Y2=1.335
r47 3 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.83 $Y=0.555
+ $X2=1.83 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_193_47# 1 2 9 11 12 15 18 21 23 25 28 29
+ 30 32 33 34 41 42 45 46 53 58
c196 46 0 4.72633e-20 $X=5.33 $Y=1.19
c197 45 0 2.56901e-19 $X=5.33 $Y=1.19
c198 41 0 3.30612e-20 $X=2.99 $Y=0.85
c199 34 0 2.53448e-20 $X=3.135 $Y=1.19
c200 33 0 1.51904e-19 $X=5.185 $Y=1.19
c201 32 0 9.52104e-20 $X=3.027 $Y=1.12
c202 25 0 1.67681e-19 $X=5.605 $Y=2.275
c203 23 0 1.753e-19 $X=5.605 $Y=1.455
c204 9 0 4.43992e-20 $X=2.315 $Y=2.275
r205 53 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=1.095
r206 53 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=0.765
r207 46 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.335
+ $Y=1.26 $X2=5.335 $Y2=1.26
r208 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.33 $Y=1.19
+ $X2=5.33 $Y2=1.19
r209 42 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=0.93 $X2=2.915 $Y2=0.93
r210 41 43 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.965
r211 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.85
r212 37 62 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.96
r213 37 58 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.51
r214 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0.85
+ $X2=1.15 $Y2=0.85
r215 33 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.19
+ $X2=5.33 $Y2=1.19
r216 33 34 2.53712 $w=1.4e-07 $l=2.05e-06 $layer=MET1_cond $X=5.185 $Y=1.19
+ $X2=3.135 $Y2=1.19
r217 32 34 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.135 $Y2=1.19
r218 32 43 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.027 $Y2=0.965
r219 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=0.85
+ $X2=1.15 $Y2=0.85
r220 29 41 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=2.99 $Y2=0.85
r221 29 30 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=1.295 $Y2=0.85
r222 28 49 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=5.47 $Y=1.26
+ $X2=5.335 $Y2=1.26
r223 23 28 52.102 $w=1.88e-07 $l=2.09464e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.575 $Y2=1.26
r224 23 25 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.605 $Y2=2.275
r225 19 28 36.719 $w=1.88e-07 $l=1.39911e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.575 $Y2=1.26
r226 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.565 $Y2=0.445
r227 18 56 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.855 $Y=1.245
+ $X2=2.855 $Y2=1.095
r228 15 55 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.855 $Y=0.415
+ $X2=2.855 $Y2=0.765
r229 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.855 $Y2=1.245
r230 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.39 $Y2=1.32
r231 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.39 $Y2=1.32
r232 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.315 $Y2=2.275
r233 2 62 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r234 1 58 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_652_21# 1 2 9 13 15 19 21 25 28 30 31 35
+ 38
c115 38 0 1.32054e-19 $X=4.625 $Y=0.895
c116 35 0 2.11834e-19 $X=4.075 $Y=1.96
c117 28 0 3.22473e-19 $X=4.625 $Y=1.835
c118 21 0 1.87283e-19 $X=4.54 $Y=1.96
r119 36 38 6.44012 $w=3.38e-07 $l=1.9e-07 $layer=LI1_cond $X=4.435 $Y=0.895
+ $X2=4.625 $Y2=0.895
r120 31 42 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.905
r121 31 41 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.575
r122 30 33 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=3.485 $Y=1.74
+ $X2=3.485 $Y2=1.96
r123 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.74 $X2=3.445 $Y2=1.74
r124 27 38 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=0.895
r125 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=1.835
r126 23 36 2.53954 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.895
r127 23 25 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.46
r128 22 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.96
+ $X2=4.075 $Y2=1.96
r129 21 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.625 $Y2=1.835
r130 21 22 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.16 $Y2=1.96
r131 17 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=1.96
r132 17 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=2.21
r133 16 33 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.61 $Y=1.96
+ $X2=3.485 $Y2=1.96
r134 15 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=4.075 $Y2=1.96
r135 15 16 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=3.61 $Y2=1.96
r136 13 42 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.335 $Y=2.275
+ $X2=3.335 $Y2=1.905
r137 9 41 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.335 $Y=0.445
+ $X2=3.335 $Y2=1.575
r138 2 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.065 $X2=4.075 $Y2=2.21
r139 1 25 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.235 $X2=4.475 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%SET_B 1 3 7 11 17 19 20 24 26 27 29 30 36 37
c135 37 0 1.72331e-19 $X=7.13 $Y=0.85
c136 29 0 2.95874e-19 $X=6.985 $Y=0.85
c137 26 0 1.49785e-19 $X=6.99 $Y=0.9
c138 19 0 1.94282e-20 $X=6.895 $Y=1.535
c139 1 0 9.39349e-20 $X=3.865 $Y=1.145
r140 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0.85
+ $X2=7.13 $Y2=0.85
r141 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=0.85
+ $X2=3.91 $Y2=0.85
r142 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=7.13 $Y2=0.85
r143 29 30 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=4.055 $Y2=0.85
r144 27 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=0.98 $X2=3.775 $Y2=0.98
r145 27 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0.85
+ $X2=3.91 $Y2=0.85
r146 26 37 5.97563 $w=2.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.99 $Y=0.87
+ $X2=7.13 $Y2=0.87
r147 24 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=0.98
+ $X2=6.825 $Y2=1.145
r148 24 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=0.98
+ $X2=6.825 $Y2=0.815
r149 23 26 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=0.9
+ $X2=6.99 $Y2=0.9
r150 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.825
+ $Y=0.98 $X2=6.825 $Y2=0.98
r151 19 20 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=6.895 $Y=1.535
+ $X2=6.895 $Y2=1.685
r152 19 44 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.885 $Y=1.535
+ $X2=6.885 $Y2=1.145
r153 17 20 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.905 $Y=2.275
+ $X2=6.905 $Y2=1.685
r154 11 43 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.765 $Y=0.445
+ $X2=6.765 $Y2=0.815
r155 5 40 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.81 $Y2=0.98
r156 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.905 $Y2=0.445
r157 1 40 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.81 $Y2=0.98
r158 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.865 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_476_47# 1 2 7 9 11 14 16 20 22 24 25 26 30
+ 35 37 38 43 44 53
c157 53 0 1.95729e-19 $X=4.705 $Y=1.4
c158 43 0 4.43992e-20 $X=3.44 $Y=1.3
c159 26 0 1.01003e-19 $X=3.02 $Y=2.335
c160 22 0 3.81194e-20 $X=5.205 $Y=0.735
c161 16 0 1.15925e-19 $X=5.13 $Y=0.825
c162 7 0 3.16972e-20 $X=4.265 $Y=0.735
r163 48 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.705 $Y2=1.4
r164 48 50 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.265 $Y2=1.4
r165 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.285
+ $Y=1.4 $X2=4.285 $Y2=1.4
r166 44 47 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.245 $Y=1.32
+ $X2=4.245 $Y2=1.4
r167 42 43 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=1.3
+ $X2=3.44 $Y2=1.3
r168 40 42 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=3.105 $Y=1.3
+ $X2=3.355 $Y2=1.3
r169 38 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=4.245 $Y2=1.32
r170 38 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=3.44 $Y2=1.32
r171 37 42 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.355 $Y=1.195
+ $X2=3.355 $Y2=1.3
r172 36 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.355 $Y=0.465
+ $X2=3.355 $Y2=1.195
r173 34 40 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=1.3
r174 34 35 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=2.25
r175 30 36 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=3.355 $Y2=0.465
r176 30 32 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=2.59 $Y2=0.365
r177 26 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=3.105 $Y2=2.25
r178 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=2.525 $Y2=2.335
r179 22 24 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.205 $Y=0.735
+ $X2=5.205 $Y2=0.445
r180 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=1.4
r181 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=2.275
r182 17 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.34 $Y=0.825
+ $X2=4.265 $Y2=0.825
r183 16 22 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=5.205 $Y2=0.735
r184 16 17 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=4.34 $Y2=0.825
r185 12 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=1.4
r186 12 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=2.275
r187 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.235
+ $X2=4.265 $Y2=1.4
r188 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=0.825
r189 10 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=1.235
r190 7 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.825
r191 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.445
r192 2 28 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.065 $X2=2.525 $Y2=2.335
r193 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.59 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_1178_261# 1 2 8 11 15 19 24 28 31 35 38 39
c76 38 0 1.67681e-19 $X=7.51 $Y=1.67
c77 31 0 1.94282e-20 $X=7.735 $Y=1.575
c78 19 0 6.59327e-20 $X=6.405 $Y=1.38
r79 37 39 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.735 $Y2=1.67
r80 37 38 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.51 $Y2=1.67
r81 33 35 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.595 $Y=0.515
+ $X2=7.735 $Y2=0.515
r82 31 39 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=7.735 $Y=1.575
+ $X2=7.735 $Y2=1.67
r83 30 35 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.735 $Y=0.68
+ $X2=7.735 $Y2=0.515
r84 30 31 52.244 $w=1.88e-07 $l=8.95e-07 $layer=LI1_cond $X=7.735 $Y=0.68
+ $X2=7.735 $Y2=1.575
r85 26 37 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.67
r86 26 28 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.87
r87 24 42 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=6.06 $Y=1.66
+ $X2=6.06 $Y2=1.825
r88 23 38 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=6.095 $Y=1.66
+ $X2=7.51 $Y2=1.66
r89 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.095
+ $Y=1.66 $X2=6.095 $Y2=1.66
r90 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=1.38
r91 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=0.445
r92 11 42 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.965 $Y=2.275
+ $X2=5.965 $Y2=1.825
r93 8 24 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=6.06 $Y=1.655 $X2=6.06
+ $Y2=1.66
r94 7 19 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.06 $Y=1.38
+ $X2=6.405 $Y2=1.38
r95 7 8 33.9437 $w=3.4e-07 $l=2e-07 $layer=POLY_cond $X=6.06 $Y=1.455 $X2=6.06
+ $Y2=1.655
r96 2 28 300 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=2 $X=7.46
+ $Y=1.645 $X2=7.595 $Y2=1.87
r97 1 33 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_1028_413# 1 2 3 12 16 18 19 22 26 30 34 36
+ 37 40 44 48 49 54 55 59 60 61 64 69 71 74 76 78
c191 74 0 9.39049e-20 $X=6.405 $Y=1.32
c192 54 0 7.27138e-20 $X=5.675 $Y=1.915
c193 49 0 1.39518e-19 $X=5.59 $Y=2.29
c194 40 0 1.2453e-19 $X=9.685 $Y=0.56
r195 77 81 10.5355 $w=3.66e-07 $l=8e-08 $layer=POLY_cond $X=7.305 $Y=1.225
+ $X2=7.385 $Y2=1.225
r196 76 78 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=1.29
+ $X2=7.14 $Y2=1.29
r197 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.305
+ $Y=1.26 $X2=7.305 $Y2=1.26
r198 67 69 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=2.085
+ $X2=6.66 $Y2=2.21
r199 66 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=6.405 $Y2=1.32
r200 66 78 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=7.14 $Y2=1.32
r201 64 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.235
+ $X2=6.405 $Y2=1.32
r202 63 64 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.405 $Y=0.475
+ $X2=6.405 $Y2=1.235
r203 62 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2 $X2=5.675
+ $Y2=2
r204 61 67 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=6.54 $Y=2
+ $X2=6.66 $Y2=2.085
r205 61 62 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.54 $Y=2 $X2=5.76
+ $Y2=2
r206 59 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=6.405 $Y2=1.32
r207 59 60 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=5.76 $Y2=1.32
r208 55 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=6.405 $Y2=0.475
r209 55 57 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=5.805 $Y2=0.39
r210 54 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=1.915
+ $X2=5.675 $Y2=2
r211 53 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.675 $Y=1.405
+ $X2=5.76 $Y2=1.32
r212 53 54 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.675 $Y=1.405
+ $X2=5.675 $Y2=1.915
r213 49 71 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.675 $Y=2.29
+ $X2=5.675 $Y2=2
r214 49 51 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=5.59 $Y=2.29
+ $X2=5.275 $Y2=2.29
r215 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.325 $Y=1.16
+ $X2=8.745 $Y2=1.16
r216 42 48 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.685 $Y=1.295
+ $X2=9.685 $Y2=1.16
r217 42 44 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.685 $Y=1.295
+ $X2=9.685 $Y2=1.985
r218 38 48 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.685 $Y=1.025
+ $X2=9.685 $Y2=1.16
r219 38 40 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.685 $Y=1.025
+ $X2=9.685 $Y2=0.56
r220 37 47 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=8.82 $Y=1.16
+ $X2=8.745 $Y2=1.16
r221 36 48 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=9.61 $Y=1.16
+ $X2=9.685 $Y2=1.16
r222 36 37 175.517 $w=2.7e-07 $l=7.9e-07 $layer=POLY_cond $X=9.61 $Y=1.16
+ $X2=8.82 $Y2=1.16
r223 32 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.745 $Y=1.295
+ $X2=8.745 $Y2=1.16
r224 32 34 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.745 $Y=1.295
+ $X2=8.745 $Y2=1.985
r225 28 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.745 $Y=1.025
+ $X2=8.745 $Y2=1.16
r226 28 30 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.745 $Y=1.025
+ $X2=8.745 $Y2=0.56
r227 24 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.325 $Y=1.295
+ $X2=8.325 $Y2=1.16
r228 24 26 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.325 $Y=1.295
+ $X2=8.325 $Y2=1.985
r229 20 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.325 $Y=1.025
+ $X2=8.325 $Y2=1.16
r230 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.325 $Y=1.025
+ $X2=8.325 $Y2=0.56
r231 19 81 13.2898 $w=3.66e-07 $l=1.0247e-07 $layer=POLY_cond $X=7.46 $Y=1.16
+ $X2=7.385 $Y2=1.225
r232 18 46 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=8.25 $Y=1.16
+ $X2=8.325 $Y2=1.16
r233 18 19 175.517 $w=2.7e-07 $l=7.9e-07 $layer=POLY_cond $X=8.25 $Y=1.16
+ $X2=7.46 $Y2=1.16
r234 14 81 23.7042 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.385 $Y=1.425
+ $X2=7.385 $Y2=1.225
r235 14 16 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.385 $Y=1.425
+ $X2=7.385 $Y2=2.065
r236 10 81 23.7042 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.385 $Y=1.025
+ $X2=7.385 $Y2=1.225
r237 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.385 $Y=1.025
+ $X2=7.385 $Y2=0.505
r238 3 69 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=2.065 $X2=6.695 $Y2=2.21
r239 2 51 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=2.065 $X2=5.275 $Y2=2.33
r240 1 57 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=5.64
+ $Y=0.235 $X2=5.805 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_1870_47# 1 2 7 9 12 14 16 19 23 27 33 36
+ 39
c71 39 0 1.91378e-19 $X=10.525 $Y=1.16
r72 34 39 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=10.105 $Y=1.16
+ $X2=10.525 $Y2=1.16
r73 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.105
+ $Y=1.16 $X2=10.105 $Y2=1.16
r74 31 36 0.881669 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.64 $Y=1.16
+ $X2=9.475 $Y2=1.16
r75 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.64 $Y=1.16
+ $X2=10.105 $Y2=1.16
r76 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.475 $Y=1.66
+ $X2=9.475 $Y2=2.34
r77 25 36 5.74456 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=1.325
+ $X2=9.475 $Y2=1.16
r78 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.475 $Y=1.325
+ $X2=9.475 $Y2=1.66
r79 21 36 5.74456 $w=2.9e-07 $l=1.83916e-07 $layer=LI1_cond $X=9.435 $Y=0.995
+ $X2=9.475 $Y2=1.16
r80 21 23 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=9.435 $Y=0.995
+ $X2=9.435 $Y2=0.51
r81 17 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.525 $Y=1.325
+ $X2=10.525 $Y2=1.16
r82 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.525 $Y=1.325
+ $X2=10.525 $Y2=1.985
r83 14 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.525 $Y=0.995
+ $X2=10.525 $Y2=1.16
r84 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.525 $Y=0.995
+ $X2=10.525 $Y2=0.56
r85 10 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.105 $Y=1.325
+ $X2=10.105 $Y2=1.16
r86 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.105 $Y=1.325
+ $X2=10.105 $Y2=1.985
r87 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.105 $Y=0.995
+ $X2=10.105 $Y2=1.16
r88 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.105 $Y=0.995
+ $X2=10.105 $Y2=0.56
r89 2 29 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=9.35
+ $Y=1.485 $X2=9.475 $Y2=2.34
r90 2 27 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=9.35
+ $Y=1.485 $X2=9.475 $Y2=1.66
r91 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=9.35
+ $Y=0.235 $X2=9.475 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 39 43 47 49
+ 53 59 63 67 71 73 75 77 79 85 90 95 103 108 113 119 122 125 132 135 142 145
+ 148 151 155
c196 155 0 1.81794e-19 $X=10.81 $Y=2.72
c197 67 0 1.91378e-19 $X=9.895 $Y=1.66
c198 10 0 3.98522e-20 $X=10.6 $Y=1.485
c199 1 0 3.29888e-20 $X=0.545 $Y=1.815
r200 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r201 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r202 149 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r203 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r204 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r205 143 146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r206 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r207 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r208 135 138 10.6812 $w=4.08e-07 $l=3.8e-07 $layer=LI1_cond $X=6.135 $Y=2.34
+ $X2=6.135 $Y2=2.72
r209 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r210 129 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r211 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r212 125 128 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.62 $Y=2.34
+ $X2=3.62 $Y2=2.72
r213 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r214 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r215 117 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r216 117 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.89 $Y2=2.72
r217 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r218 114 151 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.98 $Y=2.72
+ $X2=9.895 $Y2=2.72
r219 114 116 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.98 $Y=2.72
+ $X2=10.35 $Y2=2.72
r220 113 154 4.12062 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=10.65 $Y=2.72
+ $X2=10.845 $Y2=2.72
r221 113 116 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.65 $Y=2.72
+ $X2=10.35 $Y2=2.72
r222 112 149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r223 112 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r224 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r225 109 145 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.2 $Y=2.72 $X2=8.11
+ $Y2=2.72
r226 109 111 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.2 $Y=2.72
+ $X2=8.51 $Y2=2.72
r227 108 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.87 $Y=2.72
+ $X2=8.995 $Y2=2.72
r228 108 111 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.87 $Y=2.72
+ $X2=8.51 $Y2=2.72
r229 107 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r230 107 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r231 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r232 104 138 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.135 $Y2=2.72
r233 104 106 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.67 $Y2=2.72
r234 103 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=7.175 $Y2=2.72
r235 103 106 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=6.67 $Y2=2.72
r236 102 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r237 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r238 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r239 99 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r240 98 101 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r241 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r242 96 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.495 $Y2=2.72
r243 96 98 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.83 $Y2=2.72
r244 95 138 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.93 $Y=2.72
+ $X2=6.135 $Y2=2.72
r245 95 101 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.93 $Y=2.72
+ $X2=5.75 $Y2=2.72
r246 94 129 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r247 94 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r248 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r249 91 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r250 91 93 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r251 90 128 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=3.62 $Y2=2.72
r252 90 93 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=2.07 $Y2=2.72
r253 89 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r254 89 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r255 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r256 86 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r257 86 88 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r258 85 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r259 85 88 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r260 79 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r261 77 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r262 75 79 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r263 75 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r264 71 154 3.12744 $w=2.65e-07 $l=1.12161e-07 $layer=LI1_cond $X=10.782
+ $Y=2.635 $X2=10.845 $Y2=2.72
r265 71 73 27.6151 $w=2.63e-07 $l=6.35e-07 $layer=LI1_cond $X=10.782 $Y=2.635
+ $X2=10.782 $Y2=2
r266 67 70 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.895 $Y=1.66
+ $X2=9.895 $Y2=2.34
r267 65 151 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.895 $Y=2.635
+ $X2=9.895 $Y2=2.72
r268 65 70 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.895 $Y=2.635
+ $X2=9.895 $Y2=2.34
r269 64 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.12 $Y=2.72
+ $X2=8.995 $Y2=2.72
r270 63 151 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=2.72
+ $X2=9.895 $Y2=2.72
r271 63 64 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.81 $Y=2.72
+ $X2=9.12 $Y2=2.72
r272 59 62 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=8.995 $Y=1.66
+ $X2=8.995 $Y2=2.34
r273 57 148 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.995 $Y=2.635
+ $X2=8.995 $Y2=2.72
r274 57 62 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.995 $Y=2.635
+ $X2=8.995 $Y2=2.34
r275 53 56 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=8.11 $Y=1.66
+ $X2=8.11 $Y2=2.34
r276 51 145 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=2.635
+ $X2=8.11 $Y2=2.72
r277 51 56 18.1768 $w=1.78e-07 $l=2.95e-07 $layer=LI1_cond $X=8.11 $Y=2.635
+ $X2=8.11 $Y2=2.34
r278 50 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.175 $Y2=2.72
r279 49 145 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.02 $Y=2.72 $X2=8.11
+ $Y2=2.72
r280 49 50 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.02 $Y=2.72
+ $X2=7.34 $Y2=2.72
r281 45 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.72
r282 45 47 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.21
r283 41 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.72
r284 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.34
r285 40 128 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.81 $Y=2.72
+ $X2=3.62 $Y2=2.72
r286 39 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=4.495 $Y2=2.72
r287 39 40 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=3.81 $Y2=2.72
r288 35 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r289 35 37 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.22
r290 31 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r291 31 33 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r292 10 73 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=10.6
+ $Y=1.485 $X2=10.735 $Y2=2
r293 9 70 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.76
+ $Y=1.485 $X2=9.895 $Y2=2.34
r294 9 67 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.76
+ $Y=1.485 $X2=9.895 $Y2=1.66
r295 8 62 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.82
+ $Y=1.485 $X2=8.955 $Y2=2.34
r296 8 59 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.82
+ $Y=1.485 $X2=8.955 $Y2=1.66
r297 7 56 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=1.485 $X2=8.115 $Y2=2.34
r298 7 53 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=1.485 $X2=8.115 $Y2=1.66
r299 6 47 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=2.065 $X2=7.175 $Y2=2.21
r300 5 135 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.04
+ $Y=2.065 $X2=6.175 $Y2=2.34
r301 4 43 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.065 $X2=4.495 $Y2=2.34
r302 3 125 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.065 $X2=3.595 $Y2=2.34
r303 2 37 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.645 $X2=1.62 $Y2=2.22
r304 1 33 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%A_381_47# 1 2 8 9 10 11 12 15 20
c59 20 0 1.34441e-19 $X=2.04 $Y=1.96
r60 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r61 11 20 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.88
r62 11 12 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.6 $Y2=1.88
r63 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r64 9 10 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=1.6 $Y2=0.73
r65 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.795
+ $X2=1.6 $Y2=1.88
r66 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.6 $Y2=0.73
r67 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.515 $Y2=1.795
r68 2 20 300 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.645 $X2=2.04 $Y2=1.96
r69 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%Q_N 1 2 7 8 9 10 11 12 20
r19 12 37 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.535 $Y=2.21
+ $X2=8.535 $Y2=2.34
r20 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=1.87
+ $X2=8.535 $Y2=2.21
r21 11 31 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8.535 $Y=1.87
+ $X2=8.535 $Y2=1.66
r22 10 31 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.535 $Y=1.53
+ $X2=8.535 $Y2=1.66
r23 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=1.19
+ $X2=8.535 $Y2=1.53
r24 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=0.85
+ $X2=8.535 $Y2=1.19
r25 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.535 $Y=0.51
+ $X2=8.535 $Y2=0.85
r26 7 20 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=8.535 $Y=0.51
+ $X2=8.535 $Y2=0.4
r27 2 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.4
+ $Y=1.485 $X2=8.535 $Y2=2.34
r28 2 31 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.4
+ $Y=1.485 $X2=8.535 $Y2=1.66
r29 1 20 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.4
+ $Y=0.235 $X2=8.535 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%Q 1 2 10 13 15 16 17 18
c32 18 0 3.37075e-19 $X=10.81 $Y=1.19
r33 17 32 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.315 $Y=2.21
+ $X2=10.315 $Y2=2.34
r34 16 17 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.315 $Y=1.87
+ $X2=10.315 $Y2=2.21
r35 14 18 7.43508 $w=5.53e-07 $l=3.45e-07 $layer=LI1_cond $X=10.637 $Y=0.845
+ $X2=10.637 $Y2=1.19
r36 13 15 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=10.355 $Y=0.72
+ $X2=10.355 $Y2=0.51
r37 13 14 2.28979 $w=6.66e-07 $l=3.38783e-07 $layer=LI1_cond $X=10.355 $Y=0.72
+ $X2=10.637 $Y2=0.845
r38 12 16 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=10.315 $Y=1.665
+ $X2=10.315 $Y2=1.87
r39 11 18 6.57304 $w=5.53e-07 $l=3.05e-07 $layer=LI1_cond $X=10.637 $Y=1.495
+ $X2=10.637 $Y2=1.19
r40 10 12 4.02047 $w=7.63e-07 $l=5e-09 $layer=LI1_cond $X=10.532 $Y=1.66
+ $X2=10.532 $Y2=1.665
r41 10 11 3.50193 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=10.532 $Y=1.66
+ $X2=10.532 $Y2=1.495
r42 2 32 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=10.18
+ $Y=1.485 $X2=10.315 $Y2=2.34
r43 2 10 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=10.18
+ $Y=1.485 $X2=10.315 $Y2=1.66
r44 1 15 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=10.18
+ $Y=0.235 $X2=10.315 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DFSBP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 44 48 52
+ 56 58 60 62 64 66 72 77 85 95 100 105 111 114 117 120 125 131 133 136 139 143
c182 143 0 1.99443e-19 $X=10.81 $Y=0
c183 125 0 1.49785e-19 $X=6.67 $Y=0.24
c184 9 0 1.72693e-19 $X=10.6 $Y=0.235
r185 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r186 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r187 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r188 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r189 130 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r190 129 131 11.126 $w=6.48e-07 $l=2e-07 $layer=LI1_cond $X=7.13 $Y=0.24
+ $X2=7.33 $Y2=0.24
r191 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r192 127 129 1.01207 $w=6.48e-07 $l=5.5e-08 $layer=LI1_cond $X=7.075 $Y=0.24
+ $X2=7.13 $Y2=0.24
r193 124 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r194 123 127 7.45249 $w=6.48e-07 $l=4.05e-07 $layer=LI1_cond $X=6.67 $Y=0.24
+ $X2=7.075 $Y2=0.24
r195 123 125 7.44573 $w=6.48e-07 $l=4.45988e-08 $layer=LI1_cond $X=6.67 $Y=0.24
+ $X2=6.67 $Y2=0.24
r196 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r197 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r198 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r199 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r200 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r201 109 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r202 109 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=9.89 $Y2=0
r203 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r204 106 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.06 $Y=0
+ $X2=9.895 $Y2=0
r205 106 108 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.06 $Y=0
+ $X2=10.35 $Y2=0
r206 105 142 4.12062 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=10.65 $Y=0
+ $X2=10.845 $Y2=0
r207 105 108 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.65 $Y=0
+ $X2=10.35 $Y2=0
r208 104 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r209 104 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.97 $Y2=0
r210 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r211 101 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.12 $Y=0
+ $X2=8.995 $Y2=0
r212 101 103 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.12 $Y=0
+ $X2=9.43 $Y2=0
r213 100 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.73 $Y=0
+ $X2=9.895 $Y2=0
r214 100 103 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.73 $Y=0 $X2=9.43
+ $Y2=0
r215 99 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r216 99 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r217 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r218 96 133 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.2 $Y=0 $X2=8.11
+ $Y2=0
r219 96 98 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.2 $Y=0 $X2=8.51
+ $Y2=0
r220 95 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.87 $Y=0
+ $X2=8.995 $Y2=0
r221 95 98 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.87 $Y=0 $X2=8.51
+ $Y2=0
r222 94 124 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r223 94 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r224 93 125 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r225 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r226 91 120 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.91
+ $Y2=0
r227 91 93 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.29
+ $Y2=0
r228 89 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r229 89 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r230 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r231 86 117 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.02 $Y=0
+ $X2=3.815 $Y2=0
r232 86 88 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.37
+ $Y2=0
r233 85 120 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.91
+ $Y2=0
r234 85 88 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.37
+ $Y2=0
r235 84 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r236 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r237 81 84 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r238 81 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r239 80 83 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r240 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r241 78 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.62 $Y2=0
r242 78 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r243 77 117 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.61 $Y=0
+ $X2=3.815 $Y2=0
r244 77 83 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.45
+ $Y2=0
r245 76 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r246 76 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r247 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r248 73 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r249 73 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r250 72 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.62 $Y2=0
r251 72 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r252 66 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r253 64 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r254 62 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r255 62 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r256 58 142 3.12744 $w=2.65e-07 $l=1.12161e-07 $layer=LI1_cond $X=10.782
+ $Y=0.085 $X2=10.845 $Y2=0
r257 58 60 13.0465 $w=2.63e-07 $l=3e-07 $layer=LI1_cond $X=10.782 $Y=0.085
+ $X2=10.782 $Y2=0.385
r258 54 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.895 $Y=0.085
+ $X2=9.895 $Y2=0
r259 54 56 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.895 $Y=0.085
+ $X2=9.895 $Y2=0.38
r260 50 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.995 $Y=0.085
+ $X2=8.995 $Y2=0
r261 50 52 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=8.995 $Y=0.085
+ $X2=8.995 $Y2=0.4
r262 46 133 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=0.085
+ $X2=8.11 $Y2=0
r263 46 48 19.4091 $w=1.78e-07 $l=3.15e-07 $layer=LI1_cond $X=8.11 $Y=0.085
+ $X2=8.11 $Y2=0.4
r264 44 133 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.02 $Y=0 $X2=8.11
+ $Y2=0
r265 44 131 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.02 $Y=0 $X2=7.33
+ $Y2=0
r266 40 120 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=0.085
+ $X2=4.91 $Y2=0
r267 40 42 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=4.91 $Y=0.085
+ $X2=4.91 $Y2=0.38
r268 36 117 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r269 36 38 7.7298 $w=4.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.36
r270 32 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r271 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.38
r272 28 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r273 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r274 9 60 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=10.6
+ $Y=0.235 $X2=10.735 $Y2=0.385
r275 8 56 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=9.76
+ $Y=0.235 $X2=9.895 $Y2=0.38
r276 7 52 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=8.82
+ $Y=0.235 $X2=8.955 $Y2=0.4
r277 6 48 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=7.99
+ $Y=0.235 $X2=8.115 $Y2=0.4
r278 5 127 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=6.84
+ $Y=0.235 $X2=7.075 $Y2=0.48
r279 4 42 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=4.995 $Y2=0.38
r280 3 38 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.235 $X2=3.695 $Y2=0.36
r281 2 34 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r282 1 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


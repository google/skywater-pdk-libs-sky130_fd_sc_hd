* File: sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1.pex.spice
* Created: Tue Sep  1 19:13:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VGND 1 2 3 4 5 6 7
+ 38 52 56 60 64 68 72 76 92 95 98 101 104 107 109 110 135 151 154
c139 76 0 7.6696e-20 $X=5 $Y=0.475
r140 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=5.44
+ $X2=4.83 $Y2=5.44
r141 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r142 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=5.44
+ $X2=0.23 $Y2=5.44
r143 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r144 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=5.44
+ $X2=6.21 $Y2=5.44
r145 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r146 148 154 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=5.44
+ $X2=6.21 $Y2=5.44
r147 148 166 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=5.44
+ $X2=4.83 $Y2=5.44
r148 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=5.44
+ $X2=5.75 $Y2=5.44
r149 145 165 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.955 $Y=5.44
+ $X2=4.7 $Y2=5.44
r150 145 147 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.955 $Y=5.44
+ $X2=5.75 $Y2=5.44
r151 144 151 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r152 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r153 141 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r154 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r155 138 166 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=5.44
+ $X2=4.83 $Y2=5.44
r156 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=5.44
+ $X2=4.37 $Y2=5.44
r157 135 165 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.445 $Y=5.44
+ $X2=4.7 $Y2=5.44
r158 135 137 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.445 $Y=5.44
+ $X2=4.37 $Y2=5.44
r159 134 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r160 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r161 131 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=5.44
+ $X2=4.37 $Y2=5.44
r162 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=5.44
+ $X2=3.45 $Y2=5.44
r163 128 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r164 128 163 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r165 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r166 125 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0
+ $X2=2.185 $Y2=0
r167 125 127 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.99
+ $Y2=0
r168 124 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=5.44
+ $X2=3.45 $Y2=5.44
r169 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=5.44
+ $X2=2.53 $Y2=5.44
r170 121 124 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=5.44
+ $X2=2.53 $Y2=5.44
r171 120 123 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=5.44
+ $X2=2.53 $Y2=5.44
r172 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=5.44
+ $X2=0.69 $Y2=5.44
r173 118 159 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=5.44
+ $X2=0.187 $Y2=5.44
r174 118 120 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=5.44
+ $X2=0.69 $Y2=5.44
r175 117 163 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r176 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r177 114 156 4.42505 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r178 114 116 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.69 $Y2=0
r179 113 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=0
+ $X2=2.185 $Y2=0
r180 113 116 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=2.02 $Y=0
+ $X2=0.69 $Y2=0
r181 110 117 0.0554856 $w=4.8e-07 $l=1.95e-07 $layer=MET1_cond $X=0.495 $Y=0
+ $X2=0.69 $Y2=0
r182 110 157 0.0754035 $w=4.8e-07 $l=2.65e-07 $layer=MET1_cond $X=0.495 $Y=0
+ $X2=0.23 $Y2=0
r183 109 121 0.0825171 $w=4.8e-07 $l=2.9e-07 $layer=MET1_cond $X=0.4 $Y=5.44
+ $X2=0.69 $Y2=5.44
r184 109 160 0.0483721 $w=4.8e-07 $l=1.7e-07 $layer=MET1_cond $X=0.4 $Y=5.44
+ $X2=0.23 $Y2=5.44
r185 107 147 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.865 $Y=5.44
+ $X2=5.75 $Y2=5.44
r186 107 108 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.865 $Y=5.44
+ $X2=6.01 $Y2=5.44
r187 106 153 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=6.155 $Y=5.44
+ $X2=6.21 $Y2=5.44
r188 106 108 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.155 $Y=5.44
+ $X2=6.01 $Y2=5.44
r189 104 143 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.865 $Y=0
+ $X2=5.75 $Y2=0
r190 104 105 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.865 $Y=0
+ $X2=6.01 $Y2=0
r191 103 150 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=6.155 $Y=0
+ $X2=6.21 $Y2=0
r192 103 105 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.155 $Y=0
+ $X2=6.01 $Y2=0
r193 101 140 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.83 $Y2=0
r194 101 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r195 100 143 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.75 $Y2=0
r196 100 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r197 98 133 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=0
+ $X2=3.91 $Y2=0
r198 98 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.14
+ $Y2=0
r199 97 140 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.305 $Y=0
+ $X2=4.83 $Y2=0
r200 97 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.14
+ $Y2=0
r201 95 130 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=5.44
+ $X2=3.45 $Y2=5.44
r202 95 96 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.575 $Y=5.44
+ $X2=3.67 $Y2=5.44
r203 94 137 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.765 $Y=5.44
+ $X2=4.37 $Y2=5.44
r204 94 96 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.765 $Y=5.44
+ $X2=3.67 $Y2=5.44
r205 92 127 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=0
+ $X2=2.99 $Y2=0
r206 92 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.28
+ $Y2=0
r207 91 133 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.91 $Y2=0
r208 91 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.28
+ $Y2=0
r209 89 123 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.645 $Y=5.44
+ $X2=2.53 $Y2=5.44
r210 89 90 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.645 $Y=5.44
+ $X2=2.775 $Y2=5.44
r211 88 130 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.905 $Y=5.44
+ $X2=3.45 $Y2=5.44
r212 88 90 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.905 $Y=5.44
+ $X2=2.775 $Y2=5.44
r213 83 108 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=5.355
+ $X2=6.01 $Y2=5.44
r214 78 105 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=0.085
+ $X2=6.01 $Y2=0
r215 74 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r216 74 76 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.475
r217 70 165 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=5.355
+ $X2=4.7 $Y2=5.44
r218 70 72 14.5406 $w=5.08e-07 $l=6.2e-07 $layer=LI1_cond $X=4.7 $Y=5.355
+ $X2=4.7 $Y2=4.735
r219 66 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r220 66 68 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.475
r221 62 96 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=5.355
+ $X2=3.67 $Y2=5.44
r222 62 64 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=3.67 $Y=5.355
+ $X2=3.67 $Y2=4.735
r223 58 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0
r224 58 60 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0.475
r225 54 90 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=5.355
+ $X2=2.775 $Y2=5.44
r226 54 56 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=2.775 $Y=5.355
+ $X2=2.775 $Y2=4.7
r227 50 162 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0
r228 50 52 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0.62
r229 45 159 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=5.355
+ $X2=0.187 $Y2=5.44
r230 40 156 3.0128 $w=2.9e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.187 $Y2=0
r231 38 83 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=6.01 $Y=4.8
+ $X2=6.01 $Y2=5.355
r232 38 78 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=6.01 $Y=0.64
+ $X2=6.01 $Y2=0.085
r233 38 45 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=0.23 $Y=4.8
+ $X2=0.23 $Y2=5.355
r234 38 40 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=0.23 $Y=0.64
+ $X2=0.23 $Y2=0.085
r235 7 76 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=0.29 $X2=5 $Y2=0.475
r236 6 72 45.5 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=4 $X=4.39
+ $Y=4.555 $X2=4.87 $Y2=4.735
r237 5 68 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.29 $X2=4.14 $Y2=0.475
r238 4 64 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.53 $Y=4.555
+ $X2=3.67 $Y2=4.735
r239 3 60 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.135
+ $Y=0.29 $X2=3.28 $Y2=0.475
r240 2 56 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.685
+ $Y=4.555 $X2=2.81 $Y2=4.7
r241 1 52 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.41 $X2=2.245 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPB 7 8 11 15 19 22
+ 27 33
r79 19 33 0.00371286 $w=1.4e-07 $l=3e-09 $layer=MET1_cond $X=0.557 $Y=3.57
+ $X2=0.56 $Y2=3.57
r80 18 27 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=6.01 $Y=3.57 $X2=6.01
+ $Y2=3.29
r81 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.015 $Y=3.57
+ $X2=6.015 $Y2=3.57
r82 15 33 6.57177 $w=1.4e-07 $l=5.31e-06 $layer=MET1_cond $X=5.87 $Y=3.57
+ $X2=0.56 $Y2=3.57
r83 15 17 0.0980892 $w=2.27e-07 $l=1.45e-07 $layer=MET1_cond $X=5.87 $Y=3.57
+ $X2=6.015 $Y2=3.57
r84 14 22 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=0.23 $Y=3.57 $X2=0.23
+ $Y2=3.29
r85 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.225 $Y=3.57
+ $X2=0.225 $Y2=3.57
r86 11 19 0.231435 $w=1.4e-07 $l=1.87e-07 $layer=MET1_cond $X=0.37 $Y=3.57
+ $X2=0.557 $Y2=3.57
r87 11 13 0.0980892 $w=2.27e-07 $l=1.45e-07 $layer=MET1_cond $X=0.37 $Y=3.57
+ $X2=0.225 $Y2=3.57
r88 8 27 91 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=5.925 $Y=3.04 $X2=6.01 $Y2=3.29
r89 7 22 91 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=0.145 $Y=3.04 $X2=0.23 $Y2=3.29
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPWRIN 1 7 11 16 17
+ 20 25 26 30 32 34
c55 25 0 2.85357e-19 $X=2.225 $Y=2.2
r56 30 32 1.10767 $w=1.4e-07 $l=8.95e-07 $layer=MET1_cond $X=1.36 $Y=2.21
+ $X2=0.465 $Y2=2.21
r57 26 34 2.07418 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.2
+ $X2=2.06 $Y2=2.2
r58 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.225 $Y=2.2
+ $X2=2.225 $Y2=2.2
r59 23 34 23.6891 $w=2.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.505 $Y=2.2
+ $X2=2.06 $Y2=2.2
r60 22 25 0.461955 $w=2.3e-07 $l=7.2e-07 $layer=MET1_cond $X=1.505 $Y=2.2
+ $X2=2.225 $Y2=2.2
r61 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.505 $Y=2.2
+ $X2=1.505 $Y2=2.2
r62 20 30 0.0864037 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=1.475 $Y=2.2
+ $X2=1.36 $Y2=2.2
r63 20 22 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=1.475 $Y=2.2
+ $X2=1.505 $Y2=2.2
r64 16 17 17.048 $w=7.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.435 $Y=3.49
+ $X2=2.435 $Y2=2.66
r65 13 26 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.225 $Y=2.335
+ $X2=2.225 $Y2=2.2
r66 13 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.225 $Y=2.335
+ $X2=2.225 $Y2=2.66
r67 9 26 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=2.2
r68 9 11 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=1.79
r69 7 16 91 $w=1.7e-07 $l=6.45697e-07 $layer=licon1_NTAP_notbjt $count=2 $X=2.1
+ $Y=3.27 $X2=2.645 $Y2=3.49
r70 1 11 300 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_PDIFF $count=2 $X=2.1
+ $Y=1.485 $X2=2.225 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_505_297# 1 2 7 9
+ 10 12 13 14 15 17 18 20 22 28 31 35 36 39 40
c84 40 0 1.64106e-19 $X=3.225 $Y=3.84
c85 39 0 1.09489e-19 $X=3.225 $Y=3.84
r86 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=3.84 $X2=3.225 $Y2=3.84
r87 37 39 51.3361 $w=3.28e-07 $l=1.47e-06 $layer=LI1_cond $X=3.225 $Y=2.37
+ $X2=3.225 $Y2=3.84
r88 35 37 7.03987 $w=2.4e-07 $l=2.16852e-07 $layer=LI1_cond $X=3.06 $Y=2.25
+ $X2=3.225 $Y2=2.37
r89 35 36 12.4848 $w=2.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.06 $Y=2.25 $X2=2.8
+ $Y2=2.25
r90 31 34 56.1816 $w=2.38e-07 $l=1.17e-06 $layer=LI1_cond $X=2.68 $Y=0.62
+ $X2=2.68 $Y2=1.79
r91 29 36 6.81649 $w=2.4e-07 $l=1.69706e-07 $layer=LI1_cond $X=2.68 $Y=2.13
+ $X2=2.8 $Y2=2.25
r92 29 34 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.68 $Y=2.13
+ $X2=2.68 $Y2=1.79
r93 26 40 80.7859 $w=3.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.235 $Y=4.33
+ $X2=3.235 $Y2=3.84
r94 26 27 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.235 $Y=4.405
+ $X2=3.455 $Y2=4.405
r95 23 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.025 $Y=4.405
+ $X2=3.235 $Y2=4.405
r96 20 22 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.315 $Y=4.48
+ $X2=4.315 $Y2=4.88
r97 19 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.96 $Y=4.405
+ $X2=3.885 $Y2=4.405
r98 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.24 $Y=4.405
+ $X2=4.315 $Y2=4.48
r99 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.24 $Y=4.405
+ $X2=3.96 $Y2=4.405
r100 15 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.885 $Y=4.48
+ $X2=3.885 $Y2=4.405
r101 15 17 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.885 $Y=4.48
+ $X2=3.885 $Y2=4.88
r102 14 27 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.53 $Y=4.405
+ $X2=3.455 $Y2=4.405
r103 13 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.81 $Y=4.405
+ $X2=3.885 $Y2=4.405
r104 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.81 $Y=4.405
+ $X2=3.53 $Y2=4.405
r105 10 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.455 $Y=4.48
+ $X2=3.455 $Y2=4.405
r106 10 12 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.455 $Y=4.48
+ $X2=3.455 $Y2=4.88
r107 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.025 $Y=4.48
+ $X2=3.025 $Y2=4.405
r108 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.025 $Y=4.48 $X2=3.025
+ $Y2=4.88
r109 2 34 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=2.525
+ $Y=1.485 $X2=2.675 $Y2=1.79
r110 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.41 $X2=2.675 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_714_58# 1 2 3 10
+ 11 14 19 22 23 24 28 29 30 31 34 36 38 46
c104 28 0 1.64375e-19 $X=4.105 $Y=2.07
c105 14 0 7.6696e-20 $X=4.78 $Y=1.955
c106 11 0 1.09489e-19 $X=4.27 $Y=2.58
c107 10 0 1.83233e-19 $X=4.705 $Y=2.58
r108 44 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.765 $Y=2.49
+ $X2=4.105 $Y2=2.49
r109 42 43 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=3.71 $Y=0.855
+ $X2=4.105 $Y2=0.855
r110 36 49 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.57 $Y=0.73
+ $X2=4.57 $Y2=0.855
r111 36 38 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=4.57 $Y=0.73
+ $X2=4.57 $Y2=0.475
r112 32 34 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.555 $Y=3.47
+ $X2=4.555 $Y2=3.235
r113 31 43 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.855
+ $X2=4.105 $Y2=0.855
r114 30 49 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.475 $Y=0.855
+ $X2=4.57 $Y2=0.855
r115 30 31 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.475 $Y=0.855
+ $X2=4.19 $Y2=0.855
r116 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.105
+ $Y=2.07 $X2=4.105 $Y2=2.07
r117 26 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=2.405
+ $X2=4.105 $Y2=2.49
r118 26 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.105 $Y=2.405
+ $X2=4.105 $Y2=2.07
r119 25 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.105 $Y=0.98
+ $X2=4.105 $Y2=0.855
r120 25 28 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.105 $Y=0.98
+ $X2=4.105 $Y2=2.07
r121 23 32 9.70995 $w=1.99e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.39 $Y=3.555
+ $X2=4.555 $Y2=3.47
r122 23 24 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.39 $Y=3.555
+ $X2=3.85 $Y2=3.555
r123 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=3.47
+ $X2=3.85 $Y2=3.555
r124 21 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=2.575
+ $X2=3.765 $Y2=2.49
r125 21 22 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.765 $Y=2.575
+ $X2=3.765 $Y2=3.47
r126 17 42 2.34666 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.71 $Y=0.73
+ $X2=3.71 $Y2=0.855
r127 17 19 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=3.71 $Y=0.73
+ $X2=3.71 $Y2=0.475
r128 16 29 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=4.105 $Y=2.505
+ $X2=4.105 $Y2=2.07
r129 12 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.78 $Y=2.505
+ $X2=4.78 $Y2=1.955
r130 11 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.27 $Y=2.58
+ $X2=4.105 $Y2=2.505
r131 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.705 $Y=2.58
+ $X2=4.78 $Y2=2.505
r132 10 11 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=2.58
+ $X2=4.27 $Y2=2.58
r133 3 34 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=3.09 $X2=4.555 $Y2=3.235
r134 2 49 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.29 $X2=4.57 $Y2=0.815
r135 2 38 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.29 $X2=4.57 $Y2=0.475
r136 1 42 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.29 $X2=3.71 $Y2=0.815
r137 1 19 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.29 $X2=3.71 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A 3 5 7 8 12 14 15
+ 18 20 24 26 30 32 33 34 35 39
c71 15 0 1.64375e-19 $X=3.63 $Y=1.145
r72 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.25 $X2=3.125 $Y2=1.25
r73 35 39 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=3.13 $Y=1.425
+ $X2=3.13 $Y2=1.25
r74 28 30 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.785 $Y=1.07
+ $X2=4.785 $Y2=0.615
r75 27 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.43 $Y=1.145
+ $X2=4.355 $Y2=1.145
r76 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.71 $Y=1.145
+ $X2=4.785 $Y2=1.07
r77 26 27 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.71 $Y=1.145
+ $X2=4.43 $Y2=1.145
r78 22 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.355 $Y=1.07
+ $X2=4.355 $Y2=1.145
r79 22 24 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.355 $Y=1.07
+ $X2=4.355 $Y2=0.615
r80 21 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4 $Y=1.145 $X2=3.925
+ $Y2=1.145
r81 20 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.28 $Y=1.145
+ $X2=4.355 $Y2=1.145
r82 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.28 $Y=1.145 $X2=4
+ $Y2=1.145
r83 16 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=1.07
+ $X2=3.925 $Y2=1.145
r84 16 18 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.925 $Y=1.07
+ $X2=3.925 $Y2=0.615
r85 14 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.85 $Y=1.145
+ $X2=3.925 $Y2=1.145
r86 14 15 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.85 $Y=1.145
+ $X2=3.63 $Y2=1.145
r87 10 15 33.8325 $w=2.41e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.63 $Y2=1.145
r88 10 38 74 $w=2.41e-07 $l=4.75857e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.125 $Y2=1.312
r89 10 12 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.495 $Y=1.07
+ $X2=3.495 $Y2=0.615
r90 9 32 4.83878 $w=1.55e-07 $l=9.38083e-08 $layer=POLY_cond $X=2.535 $Y=1.147
+ $X2=2.455 $Y2=1.117
r91 8 38 39.1212 $w=2.41e-07 $l=2.33345e-07 $layer=POLY_cond $X=2.96 $Y=1.147
+ $X2=3.125 $Y2=1.312
r92 8 9 203.325 $w=1.55e-07 $l=4.25e-07 $layer=POLY_cond $X=2.96 $Y=1.147
+ $X2=2.535 $Y2=1.147
r93 5 32 20.9729 $w=1.5e-07 $l=1.09471e-07 $layer=POLY_cond $X=2.46 $Y=1.01
+ $X2=2.455 $Y2=1.117
r94 5 7 125.32 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.46 $Y=1.01 $X2=2.46
+ $Y2=0.62
r95 1 32 20.9729 $w=1.5e-07 $l=1.10472e-07 $layer=POLY_cond $X=2.45 $Y=1.225
+ $X2=2.455 $Y2=1.117
r96 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.45 $Y=1.225 $X2=2.45
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_620_911# 1 2 3 10
+ 11 12 17 18 20 24 29 31 32 34 38 40 41 44 48 49 53 56 57 60 62 63
c126 60 0 1.08173e-19 $X=4.555 $Y=1.79
c127 44 0 7.14482e-20 $X=4.1 $Y=4.735
c128 38 0 9.26578e-20 $X=3.24 $Y=4.735
c129 31 0 8.23968e-20 $X=4.78 $Y=2.94
c130 24 0 9.10198e-20 $X=5.085 $Y=4.88
c131 18 0 1.24721e-19 $X=5.16 $Y=2.94
c132 11 0 1.76914e-21 $X=4.27 $Y=2.94
c133 10 0 7.64702e-20 $X=4.705 $Y=2.94
r134 58 60 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.555 $Y=2.745
+ $X2=4.555 $Y2=1.79
r135 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.47 $Y=2.83
+ $X2=4.555 $Y2=2.745
r136 56 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.47 $Y=2.83
+ $X2=4.19 $Y2=2.83
r137 54 63 10.0555 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.105 $Y=4.045
+ $X2=4.105 $Y2=3.97
r138 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=3.975 $X2=4.105 $Y2=3.975
r139 51 62 3.70735 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.105 $Y=4.155
+ $X2=3.935 $Y2=4.155
r140 51 53 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.105 $Y=4.155
+ $X2=4.105 $Y2=3.975
r141 49 63 146.009 $w=3.3e-07 $l=8.35e-07 $layer=POLY_cond $X=4.105 $Y=3.135
+ $X2=4.105 $Y2=3.97
r142 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=3.135 $X2=4.105 $Y2=3.135
r143 46 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=2.915
+ $X2=4.19 $Y2=2.83
r144 46 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.105 $Y=2.915
+ $X2=4.105 $Y2=3.135
r145 42 62 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=4.1 $Y=4.325
+ $X2=3.935 $Y2=4.155
r146 42 44 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.1 $Y=4.325
+ $X2=4.1 $Y2=4.735
r147 40 62 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=4.24
+ $X2=3.935 $Y2=4.155
r148 40 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.935 $Y=4.24
+ $X2=3.405 $Y2=4.24
r149 36 41 17.4739 $w=1.11e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.24 $Y=4.325
+ $X2=3.405 $Y2=4.24
r150 36 38 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.24 $Y=4.325
+ $X2=3.24 $Y2=4.735
r151 33 34 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.085 $Y=4.045
+ $X2=5.235 $Y2=4.045
r152 30 49 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=4.105 $Y=3.015
+ $X2=4.105 $Y2=3.135
r153 27 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.235 $Y=3.97
+ $X2=5.235 $Y2=4.045
r154 27 29 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.235 $Y=3.97
+ $X2=5.235 $Y2=3.485
r155 26 29 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.235 $Y=3.015
+ $X2=5.235 $Y2=3.485
r156 22 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.085 $Y=4.12
+ $X2=5.085 $Y2=4.045
r157 22 24 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.085 $Y=4.12
+ $X2=5.085 $Y2=4.88
r158 21 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=4.045
+ $X2=4.78 $Y2=4.045
r159 20 33 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.01 $Y=4.045
+ $X2=5.085 $Y2=4.045
r160 20 21 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.01 $Y=4.045
+ $X2=4.855 $Y2=4.045
r161 19 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=2.94
+ $X2=4.78 $Y2=2.94
r162 18 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.16 $Y=2.94
+ $X2=5.235 $Y2=3.015
r163 18 19 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=5.16 $Y=2.94
+ $X2=4.855 $Y2=2.94
r164 15 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=3.97
+ $X2=4.78 $Y2=4.045
r165 15 17 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.78 $Y=3.97
+ $X2=4.78 $Y2=3.485
r166 14 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=3.015
+ $X2=4.78 $Y2=2.94
r167 14 17 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.78 $Y=3.015 $X2=4.78
+ $Y2=3.485
r168 13 54 22.122 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=4.045
+ $X2=4.105 $Y2=4.045
r169 12 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=4.045
+ $X2=4.78 $Y2=4.045
r170 12 13 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=4.045
+ $X2=4.27 $Y2=4.045
r171 11 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.27 $Y=2.94
+ $X2=4.105 $Y2=3.015
r172 10 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=2.94
+ $X2=4.78 $Y2=2.94
r173 10 11 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.705 $Y=2.94
+ $X2=4.27 $Y2=2.94
r174 3 60 300 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.56 $X2=4.555 $Y2=1.79
r175 2 44 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.96 $Y=4.555
+ $X2=4.1 $Y2=4.735
r176 1 38 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=3.1 $Y=4.555
+ $X2=3.24 $Y2=4.735
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%A_1028_32# 1 2 7 9
+ 13 14 15 17 19 21 23 26 30 33 36
c68 26 0 9.10198e-20 $X=5.455 $Y=3.235
c69 15 0 1.08173e-19 $X=5.305 $Y=2.58
r70 33 35 12.4159 $w=4.52e-07 $l=4.6e-07 $layer=LI1_cond $X=5.45 $Y=4.24
+ $X2=5.45 $Y2=4.7
r71 31 36 19.468 $w=3.59e-07 $l=1.45e-07 $layer=POLY_cond $X=5.92 $Y=4.195
+ $X2=5.775 $Y2=4.195
r72 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.92
+ $Y=4.21 $X2=5.92 $Y2=4.21
r73 28 33 4.69682 $w=2.3e-07 $l=3.15e-07 $layer=LI1_cond $X=5.765 $Y=4.24
+ $X2=5.45 $Y2=4.24
r74 28 30 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.765 $Y=4.24
+ $X2=5.92 $Y2=4.24
r75 24 33 7.30083 $w=4.52e-07 $l=1.17473e-07 $layer=LI1_cond $X=5.455 $Y=4.125
+ $X2=5.45 $Y2=4.24
r76 24 26 51.9522 $w=1.88e-07 $l=8.9e-07 $layer=LI1_cond $X=5.455 $Y=4.125
+ $X2=5.455 $Y2=3.235
r77 21 22 56.6142 $w=4.64e-07 $l=5.45e-07 $layer=POLY_cond $X=5.23 $Y=1.25
+ $X2=5.775 $Y2=1.25
r78 20 21 1.55819 $w=4.64e-07 $l=1.5e-08 $layer=POLY_cond $X=5.215 $Y=1.25
+ $X2=5.23 $Y2=1.25
r79 19 36 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.775 $Y=4.015
+ $X2=5.775 $Y2=4.195
r80 18 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.775 $Y=2.655
+ $X2=5.775 $Y2=2.58
r81 18 19 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=5.775 $Y=2.655
+ $X2=5.775 $Y2=4.015
r82 17 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.775 $Y=2.505
+ $X2=5.775 $Y2=2.58
r83 16 22 29.5305 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.775 $Y=1.485
+ $X2=5.775 $Y2=1.25
r84 16 17 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=5.775 $Y=1.485
+ $X2=5.775 $Y2=2.505
r85 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.7 $Y=2.58
+ $X2=5.775 $Y2=2.58
r86 14 15 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.7 $Y=2.58
+ $X2=5.305 $Y2=2.58
r87 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.23 $Y=2.505
+ $X2=5.305 $Y2=2.58
r88 11 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.23 $Y=2.505
+ $X2=5.23 $Y2=1.955
r89 10 21 29.5305 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.23 $Y=1.485
+ $X2=5.23 $Y2=1.25
r90 10 13 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.23 $Y=1.485 $X2=5.23
+ $Y2=1.955
r91 7 20 29.5305 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.215 $Y=1.015
+ $X2=5.215 $Y2=1.25
r92 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.215 $Y=1.015 $X2=5.215
+ $Y2=0.615
r93 2 26 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.31
+ $Y=3.09 $X2=5.455 $Y2=3.235
r94 1 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.16
+ $Y=4.555 $X2=5.3 $Y2=4.7
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%VPWR 1 2 9 13 16 17
+ 24 31 32 39
c81 16 0 1.83233e-19 $X=5.005 $Y=2.72
r82 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r83 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r84 29 39 0.480875 $w=4.8e-07 $l=1.69e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=3.6 $Y2=2.72
r85 28 31 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r86 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r87 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r88 21 25 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r89 20 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r90 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r91 17 39 0.13658 $w=4.8e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=2.72 $X2=3.6
+ $Y2=2.72
r92 17 25 0.429658 $w=4.8e-07 $l=1.51e-06 $layer=MET1_cond $X=3.12 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 15 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=5.29 $Y2=2.72
r94 15 16 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.12 $Y=2.72
+ $X2=5.005 $Y2=2.72
r95 11 16 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.805
+ $X2=5.005 $Y2=2.72
r96 11 13 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.005 $Y=2.805
+ $X2=5.005 $Y2=3.235
r97 7 16 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.635
+ $X2=5.005 $Y2=2.72
r98 7 9 42.3398 $w=2.28e-07 $l=8.45e-07 $layer=LI1_cond $X=5.005 $Y=2.635
+ $X2=5.005 $Y2=1.79
r99 2 13 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=3.09 $X2=5.005 $Y2=3.235
r100 1 9 300 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.56 $X2=5.005 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_LSBUF_LH_HL_ISOWELL_TAP_1%X 1 2 9 11 12 18
r21 18 26 3.14303 $w=2.73e-07 $l=7.5e-08 $layer=LI1_cond $X=5.497 $Y=1.055
+ $X2=5.497 $Y2=0.98
r22 12 23 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=5.497 $Y=1.425
+ $X2=5.497 $Y2=1.79
r23 11 26 0.293093 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=5.485 $Y=0.975
+ $X2=5.485 $Y2=0.98
r24 11 12 15.2961 $w=2.73e-07 $l=3.65e-07 $layer=LI1_cond $X=5.497 $Y=1.06
+ $X2=5.497 $Y2=1.425
r25 11 18 0.209535 $w=2.73e-07 $l=5e-09 $layer=LI1_cond $X=5.497 $Y=1.06
+ $X2=5.497 $Y2=1.055
r26 7 11 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=5.485 $Y=0.83
+ $X2=5.485 $Y2=0.975
r27 7 9 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=5.485 $Y=0.83
+ $X2=5.485 $Y2=0.475
r28 2 23 300 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=2 $X=5.305
+ $Y=1.56 $X2=5.455 $Y2=1.79
r29 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.29
+ $Y=0.29 $X2=5.43 $Y2=0.475
.ends


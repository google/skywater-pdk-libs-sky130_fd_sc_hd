* File: sky130_fd_sc_hd__o221ai_2.pex.spice
* Created: Tue Sep  1 19:22:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O221AI_2%C1 1 3 6 8 10 13 15 22
r41 21 22 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.475 $Y=1.16
+ $X2=0.895 $Y2=1.16
r42 18 21 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.16
+ $X2=0.475 $Y2=1.16
r43 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r44 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.325
+ $X2=0.895 $Y2=1.16
r45 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.895 $Y=1.325
+ $X2=0.895 $Y2=1.985
r46 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=0.995
+ $X2=0.895 $Y2=1.16
r47 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.895 $Y=0.995
+ $X2=0.895 $Y2=0.56
r48 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.16
r49 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.985
r50 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%B1 1 3 6 8 10 13 15 19 20 22 25 26 27
r82 24 26 10.5432 $w=5.38e-07 $l=2e-07 $layer=LI1_cond $X=1.835 $Y=1.345
+ $X2=2.035 $Y2=1.345
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=1.16 $X2=1.835 $Y2=1.16
r84 22 27 13.622 $w=5.38e-07 $l=6.15e-07 $layer=LI1_cond $X=1.765 $Y=1.345
+ $X2=1.15 $Y2=1.345
r85 22 24 1.55047 $w=5.38e-07 $l=7e-08 $layer=LI1_cond $X=1.765 $Y=1.345
+ $X2=1.835 $Y2=1.345
r86 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=1.16 $X2=3.095 $Y2=1.16
r87 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.095 $Y=1.445
+ $X2=3.095 $Y2=1.16
r88 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.93 $Y=1.53
+ $X2=3.095 $Y2=1.445
r89 15 26 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.93 $Y=1.53
+ $X2=2.035 $Y2=1.53
r90 11 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=1.325
+ $X2=3.095 $Y2=1.16
r91 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.095 $Y=1.325
+ $X2=3.095 $Y2=1.985
r92 8 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=0.995
+ $X2=3.095 $Y2=1.16
r93 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.095 $Y=0.995
+ $X2=3.095 $Y2=0.56
r94 4 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.325
+ $X2=1.835 $Y2=1.16
r95 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.835 $Y=1.325
+ $X2=1.835 $Y2=1.985
r96 1 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=0.995
+ $X2=1.835 $Y2=1.16
r97 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.835 $Y=0.995
+ $X2=1.835 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%B2 1 3 6 8 10 13 15 22
r41 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.465 $Y=1.16
+ $X2=2.675 $Y2=1.16
r42 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.255 $Y=1.16
+ $X2=2.465 $Y2=1.16
r43 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.465
+ $Y=1.16 $X2=2.465 $Y2=1.16
r44 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.325
+ $X2=2.675 $Y2=1.16
r45 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.675 $Y=1.325
+ $X2=2.675 $Y2=1.985
r46 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=0.995
+ $X2=2.675 $Y2=1.16
r47 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.675 $Y=0.995
+ $X2=2.675 $Y2=0.56
r48 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.325
+ $X2=2.255 $Y2=1.16
r49 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.255 $Y=1.325
+ $X2=2.255 $Y2=1.985
r50 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.995
+ $X2=2.255 $Y2=1.16
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.255 $Y=0.995
+ $X2=2.255 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%A1 1 3 6 8 10 13 17 18 20 21 23 24 25 29 33
c86 29 0 1.25382e-19 $X=4.855 $Y=1.16
c87 1 0 9.81989e-20 $X=3.595 $Y=0.995
r88 30 33 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=4.855 $Y=1.175
+ $X2=5.29 $Y2=1.175
r89 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.855
+ $Y=1.16 $X2=4.855 $Y2=1.16
r90 25 33 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=5.31 $Y=1.175 $X2=5.29
+ $Y2=1.175
r91 24 30 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=4.815 $Y=1.175
+ $X2=4.855 $Y2=1.175
r92 22 24 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.73 $Y=1.275
+ $X2=4.815 $Y2=1.175
r93 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.73 $Y=1.275
+ $X2=4.73 $Y2=1.445
r94 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.645 $Y=1.53
+ $X2=4.73 $Y2=1.445
r95 20 21 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.645 $Y=1.53
+ $X2=3.76 $Y2=1.53
r96 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.595
+ $Y=1.16 $X2=3.595 $Y2=1.16
r97 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.595 $Y=1.445
+ $X2=3.76 $Y2=1.53
r98 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.595 $Y=1.445
+ $X2=3.595 $Y2=1.16
r99 11 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.325
+ $X2=4.855 $Y2=1.16
r100 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.855 $Y=1.325
+ $X2=4.855 $Y2=1.985
r101 8 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=0.995
+ $X2=4.855 $Y2=1.16
r102 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.855 $Y=0.995
+ $X2=4.855 $Y2=0.56
r103 4 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.325
+ $X2=3.595 $Y2=1.16
r104 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.595 $Y=1.325
+ $X2=3.595 $Y2=1.985
r105 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=0.995
+ $X2=3.595 $Y2=1.16
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.595 $Y=0.995
+ $X2=3.595 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%A2 1 3 6 8 10 13 15 22
r48 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.225 $Y=1.16
+ $X2=4.435 $Y2=1.16
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.225
+ $Y=1.16 $X2=4.225 $Y2=1.16
r50 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.015 $Y=1.16
+ $X2=4.225 $Y2=1.16
r51 15 21 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=1.175
+ $X2=4.225 $Y2=1.175
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=1.325
+ $X2=4.435 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.435 $Y=1.325
+ $X2=4.435 $Y2=1.985
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=0.995
+ $X2=4.435 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.435 $Y=0.995
+ $X2=4.435 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.015 $Y=1.325
+ $X2=4.015 $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.015 $Y=0.995
+ $X2=4.015 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%VPWR 1 2 3 4 13 15 21 25 30 31 32 39 52 53
+ 61 64 66
r73 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r74 63 64 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=1.625 $Y=2.465
+ $X2=1.75 $Y2=2.465
r75 59 63 0.263841 $w=6.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.61 $Y=2.465
+ $X2=1.625 $Y2=2.465
r76 59 61 18.8554 $w=6.78e-07 $l=6.3e-07 $layer=LI1_cond $X=1.61 $Y=2.465
+ $X2=0.98 $Y2=2.465
r77 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r78 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 50 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r80 50 67 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r82 47 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=2.72
+ $X2=3.345 $Y2=2.72
r83 47 49 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=3.51 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 46 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r86 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r87 43 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r88 42 45 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r89 42 64 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72 $X2=1.75
+ $Y2=2.72
r90 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r91 39 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=2.72
+ $X2=3.345 $Y2=2.72
r92 39 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.18 $Y=2.72
+ $X2=2.99 $Y2=2.72
r93 38 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 37 61 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=0.98 $Y2=2.72
r95 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 35 56 3.97976 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=0.195 $Y2=2.72
r97 35 37 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=2.72 $X2=0.69
+ $Y2=2.72
r98 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r99 32 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r100 30 49 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.985 $Y=2.72
+ $X2=4.83 $Y2=2.72
r101 30 31 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.985 $Y=2.72
+ $X2=5.087 $Y2=2.72
r102 29 52 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.19 $Y=2.72 $X2=5.29
+ $Y2=2.72
r103 29 31 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=5.19 $Y=2.72
+ $X2=5.087 $Y2=2.72
r104 25 28 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.087 $Y=1.62
+ $X2=5.087 $Y2=2.3
r105 23 31 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.087 $Y=2.635
+ $X2=5.087 $Y2=2.72
r106 23 28 18.1242 $w=2.03e-07 $l=3.35e-07 $layer=LI1_cond $X=5.087 $Y=2.635
+ $X2=5.087 $Y2=2.3
r107 19 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=2.635
+ $X2=3.345 $Y2=2.72
r108 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.345 $Y=2.635
+ $X2=3.345 $Y2=2.3
r109 15 18 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.265 $Y=1.65
+ $X2=0.265 $Y2=2.33
r110 13 56 3.1634 $w=2.5e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.195 $Y2=2.72
r111 13 18 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.33
r112 4 28 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=1.485 $X2=5.07 $Y2=2.3
r113 4 25 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=1.485 $X2=5.07 $Y2=1.62
r114 3 21 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.17
+ $Y=1.485 $X2=3.305 $Y2=2.3
r115 2 63 300 $w=1.7e-07 $l=1.09455e-06 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=1.485 $X2=1.625 $Y2=2.3
r116 1 18 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=2.33
r117 1 15 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%Y 1 2 3 4 13 16 19 23 26 29 31 32 33 38 43
r65 38 41 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.225 $Y=1.87
+ $X2=4.225 $Y2=1.96
r66 33 43 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.34 $Y=1.87
+ $X2=1.63 $Y2=1.87
r67 32 36 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.465 $Y=1.87
+ $X2=2.465 $Y2=1.96
r68 32 33 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.465 $Y=1.87
+ $X2=2.34 $Y2=1.87
r69 30 43 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.85 $Y=1.87
+ $X2=1.63 $Y2=1.87
r70 30 31 3.05049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.85 $Y=1.87
+ $X2=0.705 $Y2=1.87
r71 28 29 27.2823 $w=2.43e-07 $l=5.8e-07 $layer=LI1_cond $X=0.727 $Y=0.865
+ $X2=0.727 $Y2=1.445
r72 26 28 5.50333 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.685 $Y=0.73
+ $X2=0.685 $Y2=0.865
r73 24 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.59 $Y=1.87
+ $X2=2.465 $Y2=1.87
r74 23 38 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.1 $Y=1.87
+ $X2=4.225 $Y2=1.87
r75 23 24 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=4.1 $Y=1.87
+ $X2=2.59 $Y2=1.87
r76 17 31 3.46198 $w=2.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=0.685 $Y=1.955
+ $X2=0.705 $Y2=1.87
r77 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.685 $Y=1.955
+ $X2=0.685 $Y2=1.96
r78 14 31 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.785
+ $X2=0.705 $Y2=1.87
r79 14 16 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=1.785
+ $X2=0.705 $Y2=1.62
r80 13 29 6.07313 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=0.705 $Y=1.59
+ $X2=0.705 $Y2=1.445
r81 13 16 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=0.705 $Y=1.59
+ $X2=0.705 $Y2=1.62
r82 4 41 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=1.485 $X2=4.225 $Y2=1.96
r83 3 36 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.485 $X2=2.465 $Y2=1.96
r84 2 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.685 $Y2=1.96
r85 2 16 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.685 $Y2=1.62
r86 1 26 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.685 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%A_382_297# 1 2 7 10 15
r21 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.885 $Y=2.3 $X2=2.885
+ $Y2=2.38
r22 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.045 $Y=2.3 $X2=2.045
+ $Y2=2.38
r23 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.17 $Y=2.38
+ $X2=2.045 $Y2=2.38
r24 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.76 $Y=2.38
+ $X2=2.885 $Y2=2.38
r25 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.76 $Y=2.38 $X2=2.17
+ $Y2=2.38
r26 2 15 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.75
+ $Y=1.485 $X2=2.885 $Y2=2.3
r27 1 10 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.485 $X2=2.045 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%A_734_297# 1 2 7 11 14
c17 11 0 1.25382e-19 $X=4.645 $Y=1.96
r18 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.805 $Y=2.3 $X2=3.805
+ $Y2=2.38
r19 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.645 $Y=2.295
+ $X2=4.645 $Y2=1.96
r20 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.93 $Y=2.38
+ $X2=3.805 $Y2=2.38
r21 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.52 $Y=2.38
+ $X2=4.645 $Y2=2.295
r22 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.52 $Y=2.38 $X2=3.93
+ $Y2=2.38
r23 2 11 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.51
+ $Y=1.485 $X2=4.645 $Y2=1.96
r24 1 14 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=1.485 $X2=3.805 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%A_28_47# 1 2 3 4 13 15 17 19 20 25
c49 25 0 6.89549e-20 $X=2.885 $Y=0.73
r50 23 25 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=2.045 $Y=0.775
+ $X2=2.885 $Y2=0.775
r51 21 32 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=1.27 $Y=0.775
+ $X2=1.145 $Y2=0.775
r52 21 23 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=1.27 $Y=0.775
+ $X2=2.045 $Y2=0.775
r53 20 32 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=1.145 $Y=0.645
+ $X2=1.145 $Y2=0.775
r54 19 30 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.145 $Y=0.475
+ $X2=1.145 $Y2=0.365
r55 19 20 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.145 $Y=0.475
+ $X2=1.145 $Y2=0.645
r56 18 28 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=0.35 $Y=0.365
+ $X2=0.225 $Y2=0.365
r57 17 30 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.02 $Y=0.365
+ $X2=1.145 $Y2=0.365
r58 17 18 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=1.02 $Y=0.365
+ $X2=0.35 $Y2=0.365
r59 13 28 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.225 $Y=0.475
+ $X2=0.225 $Y2=0.365
r60 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=0.475
+ $X2=0.225 $Y2=0.73
r61 4 25 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.75
+ $Y=0.235 $X2=2.885 $Y2=0.73
r62 3 23 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.235 $X2=2.045 $Y2=0.73
r63 2 32 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.235 $X2=1.105 $Y2=0.73
r64 2 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.235 $X2=1.105 $Y2=0.39
r65 1 28 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.39
r66 1 15 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%A_300_47# 1 2 3 4 5 16 22 25 26 27 30 32 36
+ 40
c73 40 0 2.9244e-20 $X=4.225 $Y=0.815
r74 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.065 $Y=0.725
+ $X2=5.065 $Y2=0.39
r75 33 40 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=0.815
+ $X2=4.225 $Y2=0.815
r76 32 34 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.9 $Y=0.815
+ $X2=5.065 $Y2=0.725
r77 32 33 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.9 $Y=0.815
+ $X2=4.39 $Y2=0.815
r78 28 40 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.225 $Y=0.725
+ $X2=4.225 $Y2=0.815
r79 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.225 $Y=0.725
+ $X2=4.225 $Y2=0.39
r80 26 40 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.06 $Y=0.82
+ $X2=4.225 $Y2=0.815
r81 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.06 $Y=0.82
+ $X2=3.55 $Y2=0.82
r82 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.385 $Y=0.735
+ $X2=3.55 $Y2=0.82
r83 23 25 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.385 $Y=0.735
+ $X2=3.385 $Y2=0.73
r84 22 39 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.385 $Y=0.475
+ $X2=3.385 $Y2=0.365
r85 22 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.385 $Y=0.475
+ $X2=3.385 $Y2=0.73
r86 18 21 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=1.625 $Y=0.365
+ $X2=2.465 $Y2=0.365
r87 16 39 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=0.365
+ $X2=3.385 $Y2=0.365
r88 16 21 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=3.22 $Y=0.365
+ $X2=2.465 $Y2=0.365
r89 5 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.93
+ $Y=0.235 $X2=5.065 $Y2=0.39
r90 4 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.09
+ $Y=0.235 $X2=4.225 $Y2=0.39
r91 3 39 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.35 $Y2=0.39
r92 3 25 182 $w=1.7e-07 $l=5.78035e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.35 $Y2=0.73
r93 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.235 $X2=2.465 $Y2=0.39
r94 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.235 $X2=1.625 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_2%VGND 1 2 9 13 16 17 19 20 21 34 35
r68 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r69 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r70 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r71 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r72 28 29 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r73 24 28 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=3.45
+ $Y2=0
r74 21 29 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=3.45
+ $Y2=0
r75 21 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 19 31 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.37
+ $Y2=0
r77 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.645
+ $Y2=0
r78 18 34 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=5.29
+ $Y2=0
r79 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.645
+ $Y2=0
r80 16 28 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.45
+ $Y2=0
r81 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.805
+ $Y2=0
r82 15 31 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.37
+ $Y2=0
r83 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.805
+ $Y2=0
r84 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=0.085
+ $X2=4.645 $Y2=0
r85 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.645 $Y=0.085
+ $X2=4.645 $Y2=0.39
r86 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0
r87 7 9 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0.39
r88 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.51
+ $Y=0.235 $X2=4.645 $Y2=0.39
r89 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.235 $X2=3.805 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__clkinv_8.spice.pex
* Created: Thu Aug 27 14:12:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKINV_8%A 1 3 4 6 7 9 12 14 16 19 21 23 26 28 30 33
+ 35 37 40 42 44 47 49 51 54 56 58 61 63 65 66 68 69 70 71 72 73 74 75 76 77 112
+ 113
r168 111 113 36.7542 $w=5.75e-07 $l=3.95e-07 $layer=POLY_cond $X=4.7 $Y=1.097
+ $X2=5.095 $Y2=1.097
r169 111 112 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=4.7
+ $Y=1.16 $X2=4.7 $Y2=1.16
r170 109 111 2.32622 $w=5.75e-07 $l=2.5e-08 $layer=POLY_cond $X=4.675 $Y=1.097
+ $X2=4.7 $Y2=1.097
r171 92 93 39.5457 $w=5.75e-07 $l=4.25e-07 $layer=POLY_cond $X=0.89 $Y=1.097
+ $X2=1.315 $Y2=1.097
r172 90 92 25.1231 $w=5.75e-07 $l=2.7e-07 $layer=POLY_cond $X=0.62 $Y=1.097
+ $X2=0.89 $Y2=1.097
r173 87 90 13.9573 $w=5.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.47 $Y=1.097
+ $X2=0.62 $Y2=1.097
r174 77 112 14.688 $w=2.53e-07 $l=3.25e-07 $layer=LI1_cond $X=4.375 $Y=1.162
+ $X2=4.7 $Y2=1.162
r175 76 77 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=3.915 $Y=1.162
+ $X2=4.375 $Y2=1.162
r176 75 76 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=3.455 $Y=1.162
+ $X2=3.915 $Y2=1.162
r177 74 75 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=2.995 $Y=1.162
+ $X2=3.455 $Y2=1.162
r178 73 74 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.162
+ $X2=2.995 $Y2=1.162
r179 72 73 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=2.075 $Y=1.162
+ $X2=2.535 $Y2=1.162
r180 71 72 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=1.615 $Y=1.162
+ $X2=2.075 $Y2=1.162
r181 70 71 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=1.155 $Y=1.162
+ $X2=1.615 $Y2=1.162
r182 69 70 24.1787 $w=2.53e-07 $l=5.35e-07 $layer=LI1_cond $X=0.62 $Y=1.162
+ $X2=1.155 $Y2=1.162
r183 69 90 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r184 66 113 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=5.095 $Y=1.385
+ $X2=5.095 $Y2=1.097
r185 66 68 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.095 $Y=1.385
+ $X2=5.095 $Y2=1.985
r186 63 109 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=4.675 $Y=1.385
+ $X2=4.675 $Y2=1.097
r187 63 65 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.675 $Y=1.385
+ $X2=4.675 $Y2=1.985
r188 59 109 23.2622 $w=5.75e-07 $l=2.5e-07 $layer=POLY_cond $X=4.425 $Y=1.097
+ $X2=4.675 $Y2=1.097
r189 59 107 15.8183 $w=5.75e-07 $l=1.7e-07 $layer=POLY_cond $X=4.425 $Y=1.097
+ $X2=4.255 $Y2=1.097
r190 59 61 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=4.425 $Y=0.81
+ $X2=4.425 $Y2=0.445
r191 56 107 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=4.255 $Y=1.385
+ $X2=4.255 $Y2=1.097
r192 56 58 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.255 $Y=1.385
+ $X2=4.255 $Y2=1.985
r193 52 107 24.1926 $w=5.75e-07 $l=2.6e-07 $layer=POLY_cond $X=3.995 $Y=1.097
+ $X2=4.255 $Y2=1.097
r194 52 105 14.8878 $w=5.75e-07 $l=1.6e-07 $layer=POLY_cond $X=3.995 $Y=1.097
+ $X2=3.835 $Y2=1.097
r195 52 54 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.995 $Y=0.81
+ $X2=3.995 $Y2=0.445
r196 49 105 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=3.835 $Y=1.385
+ $X2=3.835 $Y2=1.097
r197 49 51 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.835 $Y=1.385
+ $X2=3.835 $Y2=1.985
r198 45 105 25.1231 $w=5.75e-07 $l=2.7e-07 $layer=POLY_cond $X=3.565 $Y=1.097
+ $X2=3.835 $Y2=1.097
r199 45 103 13.9573 $w=5.75e-07 $l=1.5e-07 $layer=POLY_cond $X=3.565 $Y=1.097
+ $X2=3.415 $Y2=1.097
r200 45 47 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.565 $Y=0.81
+ $X2=3.565 $Y2=0.445
r201 42 103 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=3.415 $Y=1.385
+ $X2=3.415 $Y2=1.097
r202 42 44 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.415 $Y=1.385
+ $X2=3.415 $Y2=1.985
r203 38 103 26.0536 $w=5.75e-07 $l=2.8e-07 $layer=POLY_cond $X=3.135 $Y=1.097
+ $X2=3.415 $Y2=1.097
r204 38 101 13.0268 $w=5.75e-07 $l=1.4e-07 $layer=POLY_cond $X=3.135 $Y=1.097
+ $X2=2.995 $Y2=1.097
r205 38 40 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.135 $Y=0.81
+ $X2=3.135 $Y2=0.445
r206 35 101 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.995 $Y=1.385
+ $X2=2.995 $Y2=1.097
r207 35 37 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.995 $Y=1.385
+ $X2=2.995 $Y2=1.985
r208 31 101 26.9841 $w=5.75e-07 $l=2.9e-07 $layer=POLY_cond $X=2.705 $Y=1.097
+ $X2=2.995 $Y2=1.097
r209 31 99 12.0963 $w=5.75e-07 $l=1.3e-07 $layer=POLY_cond $X=2.705 $Y=1.097
+ $X2=2.575 $Y2=1.097
r210 31 33 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.705 $Y=0.81
+ $X2=2.705 $Y2=0.445
r211 28 99 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.575 $Y=1.385
+ $X2=2.575 $Y2=1.097
r212 28 30 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.575 $Y=1.385
+ $X2=2.575 $Y2=1.985
r213 24 99 27.9146 $w=5.75e-07 $l=3e-07 $layer=POLY_cond $X=2.275 $Y=1.097
+ $X2=2.575 $Y2=1.097
r214 24 97 11.1658 $w=5.75e-07 $l=1.2e-07 $layer=POLY_cond $X=2.275 $Y=1.097
+ $X2=2.155 $Y2=1.097
r215 24 26 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.275 $Y=0.81
+ $X2=2.275 $Y2=0.445
r216 21 97 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=2.155 $Y=1.385
+ $X2=2.155 $Y2=1.097
r217 21 23 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.155 $Y=1.385
+ $X2=2.155 $Y2=1.985
r218 17 97 28.8451 $w=5.75e-07 $l=3.1e-07 $layer=POLY_cond $X=1.845 $Y=1.097
+ $X2=2.155 $Y2=1.097
r219 17 95 10.2353 $w=5.75e-07 $l=1.1e-07 $layer=POLY_cond $X=1.845 $Y=1.097
+ $X2=1.735 $Y2=1.097
r220 17 19 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.845 $Y=0.81
+ $X2=1.845 $Y2=0.445
r221 14 95 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.097
r222 14 16 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.985
r223 10 95 29.7756 $w=5.75e-07 $l=3.2e-07 $layer=POLY_cond $X=1.415 $Y=1.097
+ $X2=1.735 $Y2=1.097
r224 10 93 9.30486 $w=5.75e-07 $l=1e-07 $layer=POLY_cond $X=1.415 $Y=1.097
+ $X2=1.315 $Y2=1.097
r225 10 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.415 $Y=0.81
+ $X2=1.415 $Y2=0.445
r226 7 93 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=1.315 $Y=1.385
+ $X2=1.315 $Y2=1.097
r227 7 9 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.315 $Y=1.385 $X2=1.315
+ $Y2=1.985
r228 4 92 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=0.89 $Y=1.385
+ $X2=0.89 $Y2=1.097
r229 4 6 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.89 $Y=1.385 $X2=0.89
+ $Y2=1.985
r230 1 87 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=0.47 $Y=1.385
+ $X2=0.47 $Y2=1.097
r231 1 3 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.47 $Y=1.385 $X2=0.47
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_8%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 42 46
+ 50 53 54 56 57 58 59 60 62 77 84 85 91 94 97
r93 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r94 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r95 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r96 85 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r97 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r98 82 97 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.43 $Y=2.72
+ $X2=5.302 $Y2=2.72
r99 82 84 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.43 $Y=2.72 $X2=5.75
+ $Y2=2.72
r100 81 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r101 81 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r102 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r103 78 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=4.47 $Y2=2.72
r104 78 80 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=4.83 $Y2=2.72
r105 77 97 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=5.175 $Y=2.72
+ $X2=5.302 $Y2=2.72
r106 77 80 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.175 $Y=2.72
+ $X2=4.83 $Y2=2.72
r107 76 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r108 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r109 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r110 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r111 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 70 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r113 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 67 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.105 $Y2=2.72
r115 67 69 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.61 $Y2=2.72
r116 66 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 63 88 4.06843 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r119 63 65 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 62 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=1.105 $Y2=2.72
r121 62 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 60 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 60 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 58 75 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.495 $Y=2.72
+ $X2=3.45 $Y2=2.72
r125 58 59 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.495 $Y=2.72
+ $X2=3.622 $Y2=2.72
r126 56 72 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.665 $Y=2.72
+ $X2=2.53 $Y2=2.72
r127 56 57 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=2.665 $Y=2.72
+ $X2=2.787 $Y2=2.72
r128 55 75 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 55 57 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=2.91 $Y=2.72
+ $X2=2.787 $Y2=2.72
r130 53 69 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.61 $Y2=2.72
r131 53 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.945 $Y2=2.72
r132 52 72 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=2.53 $Y2=2.72
r133 52 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=1.945 $Y2=2.72
r134 48 97 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.302 $Y=2.635
+ $X2=5.302 $Y2=2.72
r135 48 50 30.2799 $w=2.53e-07 $l=6.7e-07 $layer=LI1_cond $X=5.302 $Y=2.635
+ $X2=5.302 $Y2=1.965
r136 44 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.47 $Y=2.635
+ $X2=4.47 $Y2=2.72
r137 44 46 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=4.47 $Y=2.635
+ $X2=4.47 $Y2=1.965
r138 43 59 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=3.75 $Y=2.72
+ $X2=3.622 $Y2=2.72
r139 42 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.345 $Y=2.72
+ $X2=4.47 $Y2=2.72
r140 42 43 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.345 $Y=2.72
+ $X2=3.75 $Y2=2.72
r141 38 59 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.622 $Y=2.635
+ $X2=3.622 $Y2=2.72
r142 38 40 30.2799 $w=2.53e-07 $l=6.7e-07 $layer=LI1_cond $X=3.622 $Y=2.635
+ $X2=3.622 $Y2=1.965
r143 34 57 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.787 $Y=2.635
+ $X2=2.787 $Y2=2.72
r144 34 36 31.5158 $w=2.43e-07 $l=6.7e-07 $layer=LI1_cond $X=2.787 $Y=2.635
+ $X2=2.787 $Y2=1.965
r145 30 54 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=2.635
+ $X2=1.945 $Y2=2.72
r146 30 32 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=1.945 $Y=2.635
+ $X2=1.945 $Y2=1.965
r147 26 91 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=2.635
+ $X2=1.105 $Y2=2.72
r148 26 28 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=2.635
+ $X2=1.105 $Y2=1.965
r149 22 88 3.14379 $w=2.6e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.197 $Y2=2.72
r150 22 24 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=1.965
r151 7 50 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=5.17
+ $Y=1.485 $X2=5.305 $Y2=1.965
r152 6 46 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=4.33
+ $Y=1.485 $X2=4.465 $Y2=1.965
r153 5 40 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=3.49
+ $Y=1.485 $X2=3.625 $Y2=1.965
r154 4 36 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=2.65
+ $Y=1.485 $X2=2.785 $Y2=1.965
r155 3 32 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=1.81
+ $Y=1.485 $X2=1.945 $Y2=1.965
r156 2 28 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.105 $Y2=1.965
r157 1 24 300 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_8%Y 1 2 3 4 5 6 7 8 9 10 32 33 34 35 36 39 41
+ 45 49 51 53 57 61 63 65 69 73 75 77 81 85 87 89 93 95 96 97 98 99 100 101 102
+ 103 104 105 106 112 113
r171 106 113 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.295 $Y=1.545
+ $X2=5.305 $Y2=1.545
r172 106 113 0.341465 $w=2.68e-07 $l=8e-09 $layer=LI1_cond $X=5.305 $Y=1.452
+ $X2=5.305 $Y2=1.46
r173 105 106 11.183 $w=2.68e-07 $l=2.62e-07 $layer=LI1_cond $X=5.305 $Y=1.19
+ $X2=5.305 $Y2=1.452
r174 104 112 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.305 $Y=0.78
+ $X2=5.305 $Y2=0.865
r175 104 105 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.305 $Y=0.9
+ $X2=5.305 $Y2=1.19
r176 104 112 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.305 $Y=0.9
+ $X2=5.305 $Y2=0.865
r177 91 106 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.885 $Y=1.545
+ $X2=5.295 $Y2=1.545
r178 91 93 9.60369 $w=2.38e-07 $l=2e-07 $layer=LI1_cond $X=4.885 $Y=1.63
+ $X2=4.885 $Y2=1.83
r179 90 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.305 $Y=0.78
+ $X2=4.21 $Y2=0.78
r180 89 104 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.17 $Y=0.78
+ $X2=5.305 $Y2=0.78
r181 89 90 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=5.17 $Y=0.78
+ $X2=4.305 $Y2=0.78
r182 88 102 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.175 $Y=1.545
+ $X2=4.047 $Y2=1.545
r183 87 91 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.765 $Y=1.545
+ $X2=4.885 $Y2=1.545
r184 87 88 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.765 $Y=1.545
+ $X2=4.175 $Y2=1.545
r185 83 103 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.21 $Y=0.695
+ $X2=4.21 $Y2=0.78
r186 83 85 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=4.21 $Y=0.695
+ $X2=4.21 $Y2=0.445
r187 79 102 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.047 $Y=1.63
+ $X2=4.047 $Y2=1.545
r188 79 81 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=4.047 $Y=1.63
+ $X2=4.047 $Y2=1.83
r189 78 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.445 $Y=0.78
+ $X2=3.35 $Y2=0.78
r190 77 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.115 $Y=0.78
+ $X2=4.21 $Y2=0.78
r191 77 78 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.115 $Y=0.78
+ $X2=3.445 $Y2=0.78
r192 76 100 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.325 $Y=1.545
+ $X2=3.202 $Y2=1.545
r193 75 102 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.92 $Y=1.545
+ $X2=4.047 $Y2=1.545
r194 75 76 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.92 $Y=1.545
+ $X2=3.325 $Y2=1.545
r195 71 101 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.695
+ $X2=3.35 $Y2=0.78
r196 71 73 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.35 $Y=0.695
+ $X2=3.35 $Y2=0.445
r197 67 100 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.202 $Y=1.63
+ $X2=3.202 $Y2=1.545
r198 67 69 9.4077 $w=2.43e-07 $l=2e-07 $layer=LI1_cond $X=3.202 $Y=1.63
+ $X2=3.202 $Y2=1.83
r199 66 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.585 $Y=0.78
+ $X2=2.49 $Y2=0.78
r200 65 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.255 $Y=0.78
+ $X2=3.35 $Y2=0.78
r201 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.255 $Y=0.78
+ $X2=2.585 $Y2=0.78
r202 64 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.495 $Y=1.545
+ $X2=2.37 $Y2=1.545
r203 63 100 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=3.08 $Y=1.545
+ $X2=3.202 $Y2=1.545
r204 63 64 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.08 $Y=1.545
+ $X2=2.495 $Y2=1.545
r205 59 99 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.695
+ $X2=2.49 $Y2=0.78
r206 59 61 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=2.49 $Y=0.695
+ $X2=2.49 $Y2=0.445
r207 55 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=1.63
+ $X2=2.37 $Y2=1.545
r208 55 57 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=2.37 $Y=1.63 $X2=2.37
+ $Y2=1.83
r209 54 97 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=0.78
+ $X2=1.63 $Y2=0.78
r210 53 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.395 $Y=0.78
+ $X2=2.49 $Y2=0.78
r211 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.395 $Y=0.78
+ $X2=1.725 $Y2=0.78
r212 52 96 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.645 $Y=1.545
+ $X2=1.525 $Y2=1.545
r213 51 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=1.545
+ $X2=2.37 $Y2=1.545
r214 51 52 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.245 $Y=1.545
+ $X2=1.645 $Y2=1.545
r215 47 97 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.695
+ $X2=1.63 $Y2=0.78
r216 47 49 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.63 $Y=0.695
+ $X2=1.63 $Y2=0.445
r217 43 96 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=1.63
+ $X2=1.525 $Y2=1.545
r218 43 45 9.60369 $w=2.38e-07 $l=2e-07 $layer=LI1_cond $X=1.525 $Y=1.63
+ $X2=1.525 $Y2=1.83
r219 42 95 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.805 $Y=1.545
+ $X2=0.685 $Y2=1.545
r220 41 96 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.405 $Y=1.545
+ $X2=1.525 $Y2=1.545
r221 41 42 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.405 $Y=1.545
+ $X2=0.805 $Y2=1.545
r222 37 95 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=1.63
+ $X2=0.685 $Y2=1.545
r223 37 39 14.4055 $w=2.38e-07 $l=3e-07 $layer=LI1_cond $X=0.685 $Y=1.63
+ $X2=0.685 $Y2=1.93
r224 35 95 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.565 $Y=1.545
+ $X2=0.685 $Y2=1.545
r225 35 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.565 $Y=1.545
+ $X2=0.285 $Y2=1.545
r226 33 97 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.535 $Y=0.78
+ $X2=1.63 $Y2=0.78
r227 33 34 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.535 $Y=0.78
+ $X2=0.285 $Y2=0.78
r228 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.46
+ $X2=0.285 $Y2=1.545
r229 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.285 $Y2=0.78
r230 31 32 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.2 $Y2=1.46
r231 10 93 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=4.75
+ $Y=1.485 $X2=4.885 $Y2=1.83
r232 9 81 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=3.91
+ $Y=1.485 $X2=4.045 $Y2=1.83
r233 8 69 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=3.07
+ $Y=1.485 $X2=3.205 $Y2=1.83
r234 7 57 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=2.23
+ $Y=1.485 $X2=2.365 $Y2=1.83
r235 6 45 300 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_PDIFF $count=2 $X=1.39
+ $Y=1.485 $X2=1.525 $Y2=1.83
r236 5 39 300 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.93
r237 4 85 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.07
+ $Y=0.235 $X2=4.21 $Y2=0.445
r238 3 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.21
+ $Y=0.235 $X2=3.35 $Y2=0.445
r239 2 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.49 $Y2=0.445
r240 1 49 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.235 $X2=1.63 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_8%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 42 44 49 54 70 71 74 77 80 83
r90 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r91 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r92 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r93 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r94 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r95 67 70 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r96 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r97 65 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r98 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r99 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r100 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r101 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r102 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=2.92
+ $Y2=0
r103 59 61 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0
+ $X2=3.45 $Y2=0
r104 58 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r105 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r106 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r107 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.06
+ $Y2=0
r108 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.53 $Y2=0
r109 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.92
+ $Y2=0
r110 54 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.755 $Y=0
+ $X2=2.53 $Y2=0
r111 53 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r112 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r113 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r114 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r115 50 52 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r116 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.06
+ $Y2=0
r117 49 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=1.61 $Y2=0
r118 47 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r119 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r120 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r121 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r122 42 47 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r123 42 83 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r124 40 64 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r125 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.64
+ $Y2=0
r126 39 67 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.83
+ $Y2=0
r127 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.64
+ $Y2=0
r128 37 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0
+ $X2=3.45 $Y2=0
r129 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.78
+ $Y2=0
r130 36 64 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.945 $Y=0
+ $X2=4.37 $Y2=0
r131 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=3.78
+ $Y2=0
r132 32 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r133 32 34 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.39
r134 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0
r135 28 30 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.78 $Y=0.085
+ $X2=3.78 $Y2=0.39
r136 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0
r137 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0.39
r138 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.06 $Y2=0
r139 20 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.06 $Y2=0.39
r140 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r141 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r142 5 34 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.5
+ $Y=0.235 $X2=4.64 $Y2=0.39
r143 4 30 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.64
+ $Y=0.235 $X2=3.78 $Y2=0.39
r144 3 26 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.235 $X2=2.92 $Y2=0.39
r145 2 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.235 $X2=2.06 $Y2=0.39
r146 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__a21boi_1.pxi.spice
* Created: Thu Aug 27 14:00:30 2020
* 
x_PM_SKY130_FD_SC_HD__A21BOI_1%B1_N N_B1_N_c_56_n N_B1_N_c_57_n N_B1_N_c_60_n
+ N_B1_N_M1001_g N_B1_N_c_58_n N_B1_N_M1007_g N_B1_N_c_61_n B1_N B1_N
+ N_B1_N_c_59_n PM_SKY130_FD_SC_HD__A21BOI_1%B1_N
x_PM_SKY130_FD_SC_HD__A21BOI_1%A_27_413# N_A_27_413#_M1007_s N_A_27_413#_M1001_s
+ N_A_27_413#_c_92_n N_A_27_413#_M1002_g N_A_27_413#_c_100_n N_A_27_413#_M1006_g
+ N_A_27_413#_c_94_n N_A_27_413#_c_102_n N_A_27_413#_c_95_n N_A_27_413#_c_103_n
+ N_A_27_413#_c_104_n N_A_27_413#_c_96_n N_A_27_413#_c_97_n N_A_27_413#_c_98_n
+ PM_SKY130_FD_SC_HD__A21BOI_1%A_27_413#
x_PM_SKY130_FD_SC_HD__A21BOI_1%A1 N_A1_M1003_g N_A1_M1004_g A1 A1 A1
+ N_A1_c_161_n N_A1_c_162_n PM_SKY130_FD_SC_HD__A21BOI_1%A1
x_PM_SKY130_FD_SC_HD__A21BOI_1%A2 N_A2_c_197_n N_A2_M1005_g N_A2_M1000_g A2
+ N_A2_c_199_n PM_SKY130_FD_SC_HD__A21BOI_1%A2
x_PM_SKY130_FD_SC_HD__A21BOI_1%VPWR N_VPWR_M1001_d N_VPWR_M1004_d N_VPWR_c_222_n
+ N_VPWR_c_223_n VPWR N_VPWR_c_224_n N_VPWR_c_225_n N_VPWR_c_226_n
+ N_VPWR_c_221_n N_VPWR_c_228_n N_VPWR_c_229_n PM_SKY130_FD_SC_HD__A21BOI_1%VPWR
x_PM_SKY130_FD_SC_HD__A21BOI_1%Y N_Y_M1002_d N_Y_M1006_s N_Y_c_262_n Y Y Y Y Y
+ N_Y_c_263_n PM_SKY130_FD_SC_HD__A21BOI_1%Y
x_PM_SKY130_FD_SC_HD__A21BOI_1%A_300_297# N_A_300_297#_M1006_d
+ N_A_300_297#_M1000_d N_A_300_297#_c_307_n N_A_300_297#_c_298_n
+ N_A_300_297#_c_301_n N_A_300_297#_c_311_n
+ PM_SKY130_FD_SC_HD__A21BOI_1%A_300_297#
x_PM_SKY130_FD_SC_HD__A21BOI_1%VGND N_VGND_M1007_d N_VGND_M1005_d N_VGND_c_314_n
+ N_VGND_c_315_n N_VGND_c_316_n VGND N_VGND_c_317_n N_VGND_c_318_n
+ N_VGND_c_319_n N_VGND_c_320_n PM_SKY130_FD_SC_HD__A21BOI_1%VGND
cc_1 VNB N_B1_N_c_56_n 0.0311339f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0.83
cc_2 VNB N_B1_N_c_57_n 0.022461f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=0.83
cc_3 VNB N_B1_N_c_58_n 0.0200728f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=0.755
cc_4 VNB N_B1_N_c_59_n 0.0398605f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_5 VNB N_A_27_413#_c_92_n 0.0149112f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=0.445
cc_6 VNB N_A_27_413#_M1002_g 0.0308142f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.815
cc_7 VNB N_A_27_413#_c_94_n 0.0102035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_413#_c_95_n 0.00272003f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.53
cc_9 VNB N_A_27_413#_c_96_n 0.019694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_413#_c_97_n 0.00577707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_413#_c_98_n 0.00845379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A1 0.00230204f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=0.445
cc_13 VNB A1 0.00235155f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.89
cc_14 VNB N_A1_c_161_n 0.0223996f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_15 VNB N_A1_c_162_n 0.0178888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_197_n 0.0214152f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0.83
cc_17 VNB A2 0.011534f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=0.445
cc_18 VNB N_A2_c_199_n 0.0343496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_221_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_262_n 0.00346252f $X=-0.19 $Y=-0.24 $X2=0.765 $Y2=0.445
cc_21 VNB N_Y_c_263_n 0.00579612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_314_n 0.00506742f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=0.905
cc_23 VNB N_VGND_c_315_n 0.0106846f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.815
cc_24 VNB N_VGND_c_316_n 0.0259694f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.89
cc_25 VNB N_VGND_c_317_n 0.0280913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_318_n 0.0306256f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.16
cc_27 VNB N_VGND_c_319_n 0.00442399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_320_n 0.16743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_B1_N_c_60_n 0.0221502f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.965
cc_30 VPB N_B1_N_c_61_n 0.0333525f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.89
cc_31 VPB N_B1_N_c_59_n 0.0498291f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_32 VPB N_A_27_413#_c_92_n 0.0114465f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=0.445
cc_33 VPB N_A_27_413#_c_100_n 0.018805f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.89
cc_34 VPB N_A_27_413#_c_94_n 0.00628762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_413#_c_102_n 0.0155042f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_36 VPB N_A_27_413#_c_103_n 0.0153722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_413#_c_104_n 0.00648879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_413#_c_98_n 0.0246952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A1_M1004_g 0.0189127f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=0.755
cc_40 VPB A1 0.00268428f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.89
cc_41 VPB N_A1_c_161_n 0.00438486f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_42 VPB N_A2_M1000_g 0.0258474f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=0.755
cc_43 VPB A2 0.00562721f $X=-0.19 $Y=1.305 $X2=0.765 $Y2=0.445
cc_44 VPB N_A2_c_199_n 0.00949519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_222_n 0.00565992f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=0.905
cc_46 VPB N_VPWR_c_223_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.89
cc_47 VPB N_VPWR_c_224_n 0.0148038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_225_n 0.0275422f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_49 VPB N_VPWR_c_226_n 0.0162531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_221_n 0.0536141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_228_n 0.00510306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_229_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB Y 0.0106006f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.89
cc_54 VPB N_Y_c_263_n 0.00223038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_B1_N_c_58_n N_A_27_413#_M1002_g 0.0151603f $X=0.765 $Y=0.755 $X2=0 $Y2=0
cc_56 N_B1_N_c_60_n N_A_27_413#_c_102_n 9.97451e-19 $X=0.475 $Y=1.965 $X2=0
+ $Y2=0
cc_57 N_B1_N_c_61_n N_A_27_413#_c_102_n 0.0017983f $X=0.475 $Y=1.89 $X2=0 $Y2=0
cc_58 N_B1_N_c_56_n N_A_27_413#_c_95_n 0.00244253f $X=0.69 $Y=0.83 $X2=0 $Y2=0
cc_59 N_B1_N_c_60_n N_A_27_413#_c_103_n 0.00759264f $X=0.475 $Y=1.965 $X2=0
+ $Y2=0
cc_60 N_B1_N_c_61_n N_A_27_413#_c_103_n 0.0241801f $X=0.475 $Y=1.89 $X2=0 $Y2=0
cc_61 B1_N N_A_27_413#_c_103_n 0.0167934f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_62 N_B1_N_c_61_n N_A_27_413#_c_104_n 0.00299548f $X=0.475 $Y=1.89 $X2=0 $Y2=0
cc_63 N_B1_N_c_57_n N_A_27_413#_c_96_n 0.00669307f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_64 N_B1_N_c_58_n N_A_27_413#_c_96_n 0.00752819f $X=0.765 $Y=0.755 $X2=0 $Y2=0
cc_65 N_B1_N_c_56_n N_A_27_413#_c_97_n 0.018432f $X=0.69 $Y=0.83 $X2=0 $Y2=0
cc_66 N_B1_N_c_58_n N_A_27_413#_c_97_n 0.00115613f $X=0.765 $Y=0.755 $X2=0 $Y2=0
cc_67 B1_N N_A_27_413#_c_97_n 0.0505851f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_68 N_B1_N_c_59_n N_A_27_413#_c_97_n 0.0174827f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_69 N_B1_N_c_56_n N_A_27_413#_c_98_n 0.0116751f $X=0.69 $Y=0.83 $X2=0 $Y2=0
cc_70 B1_N N_A_27_413#_c_98_n 4.32293e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_71 N_B1_N_c_59_n N_A_27_413#_c_98_n 0.0258101f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B1_N_c_60_n N_VPWR_c_222_n 0.0104774f $X=0.475 $Y=1.965 $X2=0 $Y2=0
cc_73 N_B1_N_c_60_n N_VPWR_c_224_n 0.00358332f $X=0.475 $Y=1.965 $X2=0 $Y2=0
cc_74 N_B1_N_c_61_n N_VPWR_c_224_n 2.91333e-19 $X=0.475 $Y=1.89 $X2=0 $Y2=0
cc_75 N_B1_N_c_60_n N_VPWR_c_221_n 0.00520749f $X=0.475 $Y=1.965 $X2=0 $Y2=0
cc_76 N_B1_N_c_60_n Y 0.00381331f $X=0.475 $Y=1.965 $X2=0 $Y2=0
cc_77 N_B1_N_c_61_n Y 8.75976e-19 $X=0.475 $Y=1.89 $X2=0 $Y2=0
cc_78 N_B1_N_c_58_n N_VGND_c_314_n 0.00818075f $X=0.765 $Y=0.755 $X2=0 $Y2=0
cc_79 N_B1_N_c_56_n N_VGND_c_317_n 3.9459e-19 $X=0.69 $Y=0.83 $X2=0 $Y2=0
cc_80 N_B1_N_c_57_n N_VGND_c_317_n 0.00533101f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_81 N_B1_N_c_58_n N_VGND_c_317_n 0.00504158f $X=0.765 $Y=0.755 $X2=0 $Y2=0
cc_82 N_B1_N_c_57_n N_VGND_c_320_n 0.00698293f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_83 N_B1_N_c_58_n N_VGND_c_320_n 0.0101627f $X=0.765 $Y=0.755 $X2=0 $Y2=0
cc_84 N_A_27_413#_c_94_n N_A1_M1004_g 0.0249305f $X=1.425 $Y=1.285 $X2=0 $Y2=0
cc_85 N_A_27_413#_M1002_g N_A1_c_161_n 0.00480829f $X=1.255 $Y=0.56 $X2=0 $Y2=0
cc_86 N_A_27_413#_c_94_n N_A1_c_161_n 0.00812765f $X=1.425 $Y=1.285 $X2=0 $Y2=0
cc_87 N_A_27_413#_M1002_g N_A1_c_162_n 0.0176506f $X=1.255 $Y=0.56 $X2=0 $Y2=0
cc_88 N_A_27_413#_c_100_n N_VPWR_c_222_n 0.00247375f $X=1.425 $Y=1.385 $X2=0
+ $Y2=0
cc_89 N_A_27_413#_c_103_n N_VPWR_c_222_n 0.0222414f $X=0.685 $Y=1.845 $X2=0
+ $Y2=0
cc_90 N_A_27_413#_c_100_n N_VPWR_c_223_n 0.00125731f $X=1.425 $Y=1.385 $X2=0
+ $Y2=0
cc_91 N_A_27_413#_c_102_n N_VPWR_c_224_n 0.0143731f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_92 N_A_27_413#_c_103_n N_VPWR_c_224_n 0.00267771f $X=0.685 $Y=1.845 $X2=0
+ $Y2=0
cc_93 N_A_27_413#_c_100_n N_VPWR_c_225_n 0.00549284f $X=1.425 $Y=1.385 $X2=0
+ $Y2=0
cc_94 N_A_27_413#_M1001_s N_VPWR_c_221_n 0.00234906f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_95 N_A_27_413#_c_100_n N_VPWR_c_221_n 0.0111873f $X=1.425 $Y=1.385 $X2=0
+ $Y2=0
cc_96 N_A_27_413#_c_102_n N_VPWR_c_221_n 0.00964021f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_97 N_A_27_413#_c_103_n N_VPWR_c_221_n 0.00556583f $X=0.685 $Y=1.845 $X2=0
+ $Y2=0
cc_98 N_A_27_413#_M1002_g N_Y_c_262_n 0.00683614f $X=1.255 $Y=0.56 $X2=0 $Y2=0
cc_99 N_A_27_413#_c_94_n N_Y_c_262_n 8.81115e-19 $X=1.425 $Y=1.285 $X2=0 $Y2=0
cc_100 N_A_27_413#_c_97_n N_Y_c_262_n 0.00544819f $X=0.685 $Y=1.165 $X2=0 $Y2=0
cc_101 N_A_27_413#_c_92_n Y 0.00473069f $X=1.18 $Y=1.285 $X2=0 $Y2=0
cc_102 N_A_27_413#_c_100_n Y 0.0135562f $X=1.425 $Y=1.385 $X2=0 $Y2=0
cc_103 N_A_27_413#_c_94_n Y 0.00399746f $X=1.425 $Y=1.285 $X2=0 $Y2=0
cc_104 N_A_27_413#_c_103_n Y 0.0161894f $X=0.685 $Y=1.845 $X2=0 $Y2=0
cc_105 N_A_27_413#_c_104_n Y 0.0373268f $X=0.72 $Y=1.44 $X2=0 $Y2=0
cc_106 N_A_27_413#_c_98_n Y 0.00191906f $X=0.72 $Y=1.285 $X2=0 $Y2=0
cc_107 N_A_27_413#_c_92_n N_Y_c_263_n 0.00707405f $X=1.18 $Y=1.285 $X2=0 $Y2=0
cc_108 N_A_27_413#_M1002_g N_Y_c_263_n 0.0130213f $X=1.255 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_27_413#_c_94_n N_Y_c_263_n 0.0149341f $X=1.425 $Y=1.285 $X2=0 $Y2=0
cc_110 N_A_27_413#_c_95_n N_Y_c_263_n 0.0129833f $X=0.685 $Y=1.335 $X2=0 $Y2=0
cc_111 N_A_27_413#_c_97_n N_Y_c_263_n 0.00674892f $X=0.685 $Y=1.165 $X2=0 $Y2=0
cc_112 N_A_27_413#_c_92_n N_VGND_c_314_n 0.00493063f $X=1.18 $Y=1.285 $X2=0
+ $Y2=0
cc_113 N_A_27_413#_M1002_g N_VGND_c_314_n 0.00301887f $X=1.255 $Y=0.56 $X2=0
+ $Y2=0
cc_114 N_A_27_413#_c_96_n N_VGND_c_314_n 0.0433487f $X=0.55 $Y=0.45 $X2=0 $Y2=0
cc_115 N_A_27_413#_c_96_n N_VGND_c_317_n 0.0227625f $X=0.55 $Y=0.45 $X2=0 $Y2=0
cc_116 N_A_27_413#_M1002_g N_VGND_c_318_n 0.00585385f $X=1.255 $Y=0.56 $X2=0
+ $Y2=0
cc_117 N_A_27_413#_M1007_s N_VGND_c_320_n 0.00214551f $X=0.425 $Y=0.235 $X2=0
+ $Y2=0
cc_118 N_A_27_413#_M1002_g N_VGND_c_320_n 0.0111439f $X=1.255 $Y=0.56 $X2=0
+ $Y2=0
cc_119 N_A_27_413#_c_96_n N_VGND_c_320_n 0.0141679f $X=0.55 $Y=0.45 $X2=0 $Y2=0
cc_120 A1 N_A2_c_197_n 0.00493426f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_121 N_A1_c_162_n N_A2_c_197_n 0.0339945f $X=1.855 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A1_M1004_g N_A2_M1000_g 0.0289648f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_123 A1 A2 0.025159f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A1_c_161_n A2 2.4762e-19 $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_125 A1 N_A2_c_199_n 0.00266155f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_126 N_A1_c_161_n N_A2_c_199_n 0.0207062f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A1_M1004_g N_VPWR_c_223_n 0.0112076f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A1_M1004_g N_VPWR_c_225_n 0.00486043f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A1_M1004_g N_VPWR_c_221_n 0.00825064f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_130 A1 N_Y_c_262_n 0.00700653f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_131 A1 N_Y_c_262_n 0.00369411f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A1_c_161_n N_Y_c_262_n 4.20116e-19 $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A1_c_162_n N_Y_c_262_n 0.00185288f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A1_M1004_g Y 0.00123204f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_135 A1 N_Y_c_263_n 0.0240875f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A1_c_161_n N_Y_c_263_n 0.00209538f $X=1.855 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A1_M1004_g N_A_300_297#_c_298_n 0.01509f $X=1.855 $Y=1.985 $X2=0 $Y2=0
cc_138 A1 N_A_300_297#_c_298_n 0.0262092f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A1_c_161_n N_A_300_297#_c_298_n 2.71876e-19 $X=1.855 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A1_c_161_n N_A_300_297#_c_301_n 3.64332e-19 $X=1.855 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A1_c_162_n N_VGND_c_316_n 0.00161536f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_142 A1 N_VGND_c_318_n 0.00738499f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_143 N_A1_c_162_n N_VGND_c_318_n 0.00585385f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_144 A1 N_VGND_c_320_n 0.00747148f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_145 N_A1_c_162_n N_VGND_c_320_n 0.0112692f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_146 A1 A_384_47# 0.00611095f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_147 N_A2_M1000_g N_VPWR_c_223_n 0.0122778f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A2_M1000_g N_VPWR_c_226_n 0.00486043f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A2_M1000_g N_VPWR_c_221_n 0.00915791f $X=2.285 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A2_M1000_g N_A_300_297#_c_298_n 0.0213106f $X=2.285 $Y=1.985 $X2=0
+ $Y2=0
cc_151 A2 N_A_300_297#_c_298_n 0.0170232f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A2_c_199_n N_A_300_297#_c_298_n 0.00126208f $X=2.485 $Y=1.16 $X2=0
+ $Y2=0
cc_153 N_A2_c_197_n N_VGND_c_316_n 0.0140185f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_154 A2 N_VGND_c_316_n 0.0206827f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A2_c_199_n N_VGND_c_316_n 0.00611831f $X=2.485 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A2_c_197_n N_VGND_c_318_n 0.00486043f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A2_c_197_n N_VGND_c_320_n 0.0083285f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_158 N_VPWR_c_221_n N_Y_M1006_s 0.00213747f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_159 N_VPWR_c_222_n Y 0.0177105f $X=0.69 $Y=2.34 $X2=0 $Y2=0
cc_160 N_VPWR_c_225_n Y 0.0197891f $X=1.905 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_221_n Y 0.0123896f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_162 N_VPWR_c_221_n N_A_300_297#_M1006_d 0.00535906f $X=2.53 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_163 N_VPWR_c_221_n N_A_300_297#_M1000_d 0.00546898f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_225_n N_A_300_297#_c_307_n 0.0117061f $X=1.905 $Y=2.72 $X2=0
+ $Y2=0
cc_165 N_VPWR_c_221_n N_A_300_297#_c_307_n 0.00720598f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_166 N_VPWR_M1004_d N_A_300_297#_c_298_n 0.00360453f $X=1.93 $Y=1.485 $X2=0
+ $Y2=0
cc_167 N_VPWR_c_223_n N_A_300_297#_c_298_n 0.0165341f $X=2.07 $Y=2.02 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_226_n N_A_300_297#_c_311_n 0.0110687f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_221_n N_A_300_297#_c_311_n 0.006434f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_170 N_Y_c_263_n N_A_300_297#_c_301_n 0.00237414f $X=1.457 $Y=1.195 $X2=0
+ $Y2=0
cc_171 N_Y_c_263_n N_VGND_c_314_n 0.00766771f $X=1.457 $Y=1.195 $X2=0 $Y2=0
cc_172 Y N_VGND_c_318_n 0.0248017f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_173 N_Y_M1002_d N_VGND_c_320_n 0.00396852f $X=1.33 $Y=0.235 $X2=0 $Y2=0
cc_174 Y N_VGND_c_320_n 0.0163582f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_175 N_VGND_c_320_n A_384_47# 0.00485956f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__einvn_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645000 0.995000 7.800000 1.285000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.345000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.870000 0.620000 8.195000 0.825000 ;
        RECT 4.870000 1.455000 8.195000 1.625000 ;
        RECT 4.870000 1.625000 5.200000 2.125000 ;
        RECT 5.710000 1.625000 6.040000 2.125000 ;
        RECT 6.550000 1.625000 6.880000 2.125000 ;
        RECT 7.390000 1.625000 7.720000 2.125000 ;
        RECT 7.970000 0.825000 8.195000 1.455000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.280000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.485000 ;
        RECT 1.455000  0.085000 1.785000 0.485000 ;
        RECT 2.295000  0.085000 2.625000 0.485000 ;
        RECT 3.135000  0.085000 3.465000 0.485000 ;
        RECT 3.975000  0.085000 4.315000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.280000 2.805000 ;
        RECT 0.515000 1.835000 0.845000 2.635000 ;
        RECT 1.410000 1.835000 1.740000 2.635000 ;
        RECT 2.250000 1.835000 2.580000 2.635000 ;
        RECT 3.090000 1.835000 3.420000 2.635000 ;
        RECT 3.930000 1.835000 4.280000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 0.345000 0.655000 ;
      RECT 0.090000 0.655000 0.845000 0.825000 ;
      RECT 0.090000 1.495000 0.845000 1.665000 ;
      RECT 0.090000 1.665000 0.345000 2.465000 ;
      RECT 0.515000 0.825000 0.845000 0.995000 ;
      RECT 0.515000 0.995000 4.475000 1.325000 ;
      RECT 0.515000 1.325000 0.845000 1.495000 ;
      RECT 1.015000 0.255000 1.285000 0.655000 ;
      RECT 1.015000 0.655000 4.700000 0.825000 ;
      RECT 1.015000 1.495000 4.700000 1.665000 ;
      RECT 1.015000 1.665000 1.240000 2.465000 ;
      RECT 1.910000 1.665000 2.080000 2.465000 ;
      RECT 1.955000 0.255000 2.125000 0.655000 ;
      RECT 2.750000 1.665000 2.920000 2.465000 ;
      RECT 2.795000 0.255000 2.965000 0.655000 ;
      RECT 3.590000 1.665000 3.760000 2.465000 ;
      RECT 3.635000 0.255000 3.805000 0.655000 ;
      RECT 4.450000 1.665000 4.700000 2.295000 ;
      RECT 4.450000 2.295000 8.195000 2.465000 ;
      RECT 4.485000 0.255000 8.195000 0.450000 ;
      RECT 4.485000 0.450000 4.700000 0.655000 ;
      RECT 5.370000 1.795000 5.540000 2.295000 ;
      RECT 6.210000 1.795000 6.380000 2.295000 ;
      RECT 7.050000 1.795000 7.220000 2.295000 ;
      RECT 7.890000 1.795000 8.195000 2.295000 ;
  END
END sky130_fd_sc_hd__einvn_8

* File: sky130_fd_sc_hd__o311ai_1.spice
* Created: Thu Aug 27 14:39:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o311ai_1.spice.pex"
.subckt sky130_fd_sc_hd__o311ai_1  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_A_138_47#_M1006_d N_A1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_138_47#_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1003 N_A_138_47#_M1003_d N_A3_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.08775 PD=1.26 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1008 A_458_47# N_B1_M1008_g N_A_138_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.19825 PD=0.86 PS=1.26 NRD=9.228 NRS=61.836 M=1 R=4.33333
+ SA=75001.8 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g A_458_47# VNB NSHORT L=0.15 W=0.65 AD=0.182
+ AS=0.06825 PD=1.86 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.2 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1009 A_138_297# N_A1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.28 PD=1.27 PS=2.56 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002.2
+ A=0.15 P=2.3 MULT=1
MM1002 A_222_297# N_A2_M1002_g A_138_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A3_M1001_g A_222_297# VPB PHIGHVT L=0.15 W=1 AD=0.225
+ AS=0.135 PD=1.45 PS=1.27 NRD=16.7253 NRS=15.7403 M=1 R=6.66667 SA=75001
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=1 AD=0.185
+ AS=0.225 PD=1.37 PS=1.45 NRD=8.8453 NRS=16.7253 M=1 R=6.66667 SA=75001.6
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1005_d N_C1_M1005_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1 AD=0.31
+ AS=0.185 PD=2.62 PS=1.37 NRD=4.9053 NRS=8.8453 M=1 R=6.66667 SA=75002.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__o311ai_1.spice.SKY130_FD_SC_HD__O311AI_1.pxi"
*
.ends
*
*

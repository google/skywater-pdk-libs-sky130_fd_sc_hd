* NGSPICE file created from sky130_fd_sc_hd__o211ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=1.025e+12p pd=6.05e+06u as=6.55e+11p ps=5.31e+06u
M1001 Y A2 a_110_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1002 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.535e+11p pd=2.08e+06u as=4.2575e+11p ps=3.91e+06u
M1003 a_110_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_326_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=0p ps=0u
M1007 Y C1 a_326_47# VNB nshort w=650000u l=150000u
+  ad=3.9325e+11p pd=2.51e+06u as=0p ps=0u
.ends


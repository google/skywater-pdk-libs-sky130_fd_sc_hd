* File: sky130_fd_sc_hd__a31o_1.spice
* Created: Tue Sep  1 18:55:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a31o_1.pex.spice"
.subckt sky130_fd_sc_hd__a31o_1  VNB VPB A3 A2 A1 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_80_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.112125 AS=0.17225 PD=0.995 PS=1.83 NRD=12.912 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1004 A_209_47# N_A3_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.112125 PD=0.97 PS=0.995 NRD=19.38 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1001 A_303_47# N_A2_M1001_g A_209_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.104 PD=0.98 PS=0.97 NRD=20.304 NRS=19.38 M=1 R=4.33333 SA=75001.2
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_80_21#_M1006_d N_A1_M1006_g A_303_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0.912 NRS=20.304 M=1 R=4.33333
+ SA=75001.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_B1_M1007_g N_A_80_21#_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.208 AS=0.10725 PD=1.94 PS=0.98 NRD=4.608 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_80_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1725 AS=0.265 PD=1.345 PS=2.53 NRD=5.91 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1008 N_A_209_297#_M1008_d N_A3_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.1725 PD=1.32 PS=1.345 NRD=2.9353 NRS=6.8753 M=1 R=6.66667
+ SA=75000.7 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_209_297#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.16 PD=1.33 PS=1.32 NRD=4.9053 NRS=4.9053 M=1 R=6.66667
+ SA=75001.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_209_297#_M1000_d N_A1_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.165 PD=1.33 PS=1.33 NRD=4.9053 NRS=4.9053 M=1 R=6.66667
+ SA=75001.6 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_A_80_21#_M1009_d N_B1_M1009_g N_A_209_297#_M1000_d VPB PHIGHVT L=0.15
+ W=1 AD=0.32 AS=0.165 PD=2.64 PS=1.33 NRD=10.8153 NRS=4.9053 M=1 R=6.66667
+ SA=75002.1 SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_59 VPB 0 1.20212e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__a31o_1.pxi.spice"
*
.ends
*
*

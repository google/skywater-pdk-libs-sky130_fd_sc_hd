* File: sky130_fd_sc_hd__xor2_1.pxi.spice
* Created: Tue Sep  1 19:33:21 2020
* 
x_PM_SKY130_FD_SC_HD__XOR2_1%B N_B_c_59_n N_B_M1005_g N_B_M1009_g N_B_c_60_n
+ N_B_M1003_g N_B_M1002_g N_B_c_61_n N_B_c_62_n N_B_c_63_n N_B_c_70_n B
+ N_B_c_64_n N_B_c_65_n B PM_SKY130_FD_SC_HD__XOR2_1%B
x_PM_SKY130_FD_SC_HD__XOR2_1%A N_A_c_143_n N_A_M1008_g N_A_M1006_g N_A_c_144_n
+ N_A_M1000_g N_A_M1004_g A N_A_c_146_n PM_SKY130_FD_SC_HD__XOR2_1%A
x_PM_SKY130_FD_SC_HD__XOR2_1%A_35_297# N_A_35_297#_M1005_d N_A_35_297#_M1009_s
+ N_A_35_297#_c_187_n N_A_35_297#_M1001_g N_A_35_297#_M1007_g
+ N_A_35_297#_c_188_n N_A_35_297#_c_189_n N_A_35_297#_c_196_n
+ N_A_35_297#_c_197_n N_A_35_297#_c_206_n N_A_35_297#_c_190_n
+ N_A_35_297#_c_262_p N_A_35_297#_c_209_n N_A_35_297#_c_191_n
+ N_A_35_297#_c_192_n N_A_35_297#_c_222_n PM_SKY130_FD_SC_HD__XOR2_1%A_35_297#
x_PM_SKY130_FD_SC_HD__XOR2_1%VPWR N_VPWR_M1006_d N_VPWR_M1002_d N_VPWR_c_277_n
+ N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n
+ VPWR N_VPWR_c_283_n N_VPWR_c_276_n PM_SKY130_FD_SC_HD__XOR2_1%VPWR
x_PM_SKY130_FD_SC_HD__XOR2_1%A_285_297# N_A_285_297#_M1004_d
+ N_A_285_297#_M1007_s N_A_285_297#_c_318_n N_A_285_297#_c_325_n
+ N_A_285_297#_c_319_n PM_SKY130_FD_SC_HD__XOR2_1%A_285_297#
x_PM_SKY130_FD_SC_HD__XOR2_1%X N_X_M1003_d N_X_M1007_d N_X_c_348_n N_X_c_345_n X
+ PM_SKY130_FD_SC_HD__XOR2_1%X
x_PM_SKY130_FD_SC_HD__XOR2_1%VGND N_VGND_M1005_s N_VGND_M1008_d N_VGND_M1001_d
+ N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n
+ VGND N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n
+ PM_SKY130_FD_SC_HD__XOR2_1%VGND
cc_1 VNB N_B_c_59_n 0.0186432f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_2 VNB N_B_c_60_n 0.01967f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=0.995
cc_3 VNB N_B_c_61_n 6.73802e-19 $X=-0.19 $Y=-0.24 $X2=1.645 $Y2=1.445
cc_4 VNB N_B_c_62_n 0.00380468f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_5 VNB N_B_c_63_n 0.0195056f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_6 VNB N_B_c_64_n 0.0224001f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_7 VNB N_B_c_65_n 0.00321074f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_8 VNB N_A_c_143_n 0.0160202f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_9 VNB N_A_c_144_n 0.0160211f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=0.995
cc_10 VNB A 0.00152291f $X=-0.19 $Y=-0.24 $X2=1.645 $Y2=1.245
cc_11 VNB N_A_c_146_n 0.0300352f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_35_297#_c_187_n 0.025013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_35_297#_c_188_n 0.0341732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_35_297#_c_189_n 0.0233289f $X=-0.19 $Y=-0.24 $X2=1.645 $Y2=1.245
cc_15 VNB N_A_35_297#_c_190_n 0.00850627f $X=-0.19 $Y=-0.24 $X2=1.56 $Y2=1.53
cc_16 VNB N_A_35_297#_c_191_n 0.00421405f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=1.53
cc_17 VNB N_A_35_297#_c_192_n 0.0220236f $X=-0.19 $Y=-0.24 $X2=0.722 $Y2=1.53
cc_18 VNB N_VPWR_c_276_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0.722 $Y2=1.53
cc_19 VNB N_X_c_345_n 8.44928e-19 $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.985
cc_20 VNB N_VGND_c_378_n 0.0113652f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=0.56
cc_21 VNB N_VGND_c_379_n 0.0122648f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.985
cc_22 VNB N_VGND_c_380_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.645 $Y2=1.445
cc_23 VNB N_VGND_c_381_n 0.0104904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_382_n 0.0361949f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_25 VNB N_VGND_c_383_n 0.0112517f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_26 VNB N_VGND_c_384_n 0.0381509f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_27 VNB N_VGND_c_385_n 0.00436214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_386_n 0.180198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_B_M1009_g 0.0223541f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.985
cc_30 VPB N_B_M1002_g 0.0228143f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_31 VPB N_B_c_61_n 0.00130531f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.445
cc_32 VPB N_B_c_63_n 0.00460655f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_33 VPB N_B_c_70_n 0.00721195f $X=-0.19 $Y=1.305 $X2=1.56 $Y2=1.53
cc_34 VPB B 3.66229e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_35 VPB N_B_c_64_n 0.00472672f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_36 VPB N_B_c_65_n 0.00251016f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_37 VPB N_A_M1006_g 0.0183378f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.985
cc_38 VPB N_A_M1004_g 0.0183338f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_39 VPB N_A_c_146_n 0.00400357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_35_297#_M1007_g 0.0282319f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_41 VPB N_A_35_297#_c_188_n 0.0157226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_35_297#_c_189_n 0.00202895f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.245
cc_43 VPB N_A_35_297#_c_196_n 0.00782983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_35_297#_c_197_n 0.0207996f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_45 VPB N_A_35_297#_c_191_n 0.00342144f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.53
cc_46 VPB N_A_35_297#_c_192_n 0.0195818f $X=-0.19 $Y=1.305 $X2=0.722 $Y2=1.53
cc_47 VPB N_VPWR_c_277_n 0.00415222f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.56
cc_48 VPB N_VPWR_c_278_n 0.00416524f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_49 VPB N_VPWR_c_279_n 0.0320302f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.445
cc_50 VPB N_VPWR_c_280_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.16
cc_51 VPB N_VPWR_c_281_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_52 VPB N_VPWR_c_282_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_53 VPB N_VPWR_c_283_n 0.032149f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.53
cc_54 VPB N_VPWR_c_276_n 0.046844f $X=-0.19 $Y=1.305 $X2=0.722 $Y2=1.53
cc_55 VPB N_A_285_297#_c_318_n 0.00419921f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.56
cc_56 VPB N_A_285_297#_c_319_n 0.00995644f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.445
cc_57 VPB N_X_c_345_n 9.56278e-19 $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_58 VPB X 0.0527968f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_59 N_B_c_59_n N_A_c_143_n 0.0242458f $X=0.51 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_60 N_B_M1009_g N_A_M1006_g 0.0583861f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_61 N_B_c_70_n N_A_M1006_g 0.0149047f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_62 N_B_c_60_n N_A_c_144_n 0.0430295f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_63 N_B_M1002_g N_A_M1004_g 0.0272174f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_64 N_B_c_70_n N_A_M1004_g 0.0144798f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_65 N_B_c_61_n A 0.00227864f $X=1.645 $Y=1.445 $X2=0 $Y2=0
cc_66 N_B_c_62_n A 0.0140779f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B_c_70_n A 0.0388786f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_68 N_B_c_64_n A 6.73416e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_69 N_B_c_65_n A 0.016854f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_70 N_B_c_61_n N_A_c_146_n 0.00384105f $X=1.645 $Y=1.445 $X2=0 $Y2=0
cc_71 N_B_c_62_n N_A_c_146_n 0.00110046f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B_c_63_n N_A_c_146_n 0.0221254f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_73 N_B_c_70_n N_A_c_146_n 0.00214031f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_74 N_B_c_64_n N_A_c_146_n 0.0214761f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B_c_65_n N_A_c_146_n 0.00607121f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B_c_62_n N_A_35_297#_c_188_n 5.50196e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B_c_63_n N_A_35_297#_c_188_n 0.0209943f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B_M1009_g N_A_35_297#_c_196_n 0.00438682f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_79 B N_A_35_297#_c_196_n 0.00243774f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_80 N_B_c_64_n N_A_35_297#_c_196_n 8.13752e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B_M1009_g N_A_35_297#_c_197_n 0.00937391f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_82 N_B_c_59_n N_A_35_297#_c_206_n 0.0125738f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B_c_64_n N_A_35_297#_c_206_n 0.00108358f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B_c_65_n N_A_35_297#_c_206_n 0.0137887f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_85 N_B_c_60_n N_A_35_297#_c_209_n 0.0128444f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B_c_62_n N_A_35_297#_c_209_n 0.0165152f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B_c_63_n N_A_35_297#_c_209_n 0.00244591f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B_c_70_n N_A_35_297#_c_209_n 0.0044708f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_89 N_B_c_60_n N_A_35_297#_c_191_n 0.00544572f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B_c_61_n N_A_35_297#_c_191_n 0.00325552f $X=1.645 $Y=1.445 $X2=0 $Y2=0
cc_91 N_B_c_62_n N_A_35_297#_c_191_n 0.0138117f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_92 N_B_c_63_n N_A_35_297#_c_191_n 0.00276653f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B_c_59_n N_A_35_297#_c_192_n 0.00572387f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B_M1009_g N_A_35_297#_c_192_n 0.00776159f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_95 B N_A_35_297#_c_192_n 0.00807294f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_96 N_B_c_64_n N_A_35_297#_c_192_n 0.00753248f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_c_65_n N_A_35_297#_c_192_n 0.0334999f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_98 N_B_c_70_n N_A_35_297#_c_222_n 0.00412186f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_99 N_B_c_65_n N_A_35_297#_c_222_n 0.00268565f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B_c_70_n A_117_297# 0.00484576f $X=1.56 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_101 B A_117_297# 0.00120458f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_102 N_B_c_70_n N_VPWR_M1006_d 0.00165831f $X=1.56 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_103 N_B_c_70_n N_VPWR_c_277_n 0.0126919f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_104 N_B_M1002_g N_VPWR_c_278_n 0.00316354f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B_M1009_g N_VPWR_c_279_n 0.00541359f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B_M1002_g N_VPWR_c_281_n 0.00541359f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B_M1009_g N_VPWR_c_276_n 0.0107189f $X=0.51 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B_M1002_g N_VPWR_c_276_n 0.00714876f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_109 N_B_c_70_n N_A_285_297#_M1004_d 0.00165495f $X=1.56 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_110 N_B_M1002_g N_A_285_297#_c_318_n 0.0114405f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_111 N_B_c_62_n N_A_285_297#_c_318_n 0.00483807f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B_c_63_n N_A_285_297#_c_318_n 9.05168e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B_c_70_n N_A_285_297#_c_318_n 2.89797e-19 $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_114 N_B_M1002_g N_A_285_297#_c_325_n 0.00812439f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B_c_70_n N_A_285_297#_c_325_n 0.0176705f $X=1.56 $Y=1.53 $X2=0 $Y2=0
cc_116 N_B_M1002_g N_A_285_297#_c_319_n 0.00326978f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B_c_60_n N_X_c_348_n 0.00683228f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B_c_60_n N_X_c_345_n 0.0030103f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B_M1002_g N_X_c_345_n 8.1591e-19 $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B_M1002_g X 0.00409202f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B_c_59_n N_VGND_c_379_n 0.0084203f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_59_n N_VGND_c_380_n 6.98115e-19 $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_60_n N_VGND_c_380_n 0.00188705f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_59_n N_VGND_c_383_n 0.00341689f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B_c_60_n N_VGND_c_384_n 0.00379767f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B_c_59_n N_VGND_c_386_n 0.00405445f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_60_n N_VGND_c_386_n 0.00671337f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_M1006_g N_A_35_297#_c_196_n 0.0020618f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_c_143_n N_A_35_297#_c_209_n 0.0114901f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_144_n N_A_35_297#_c_209_n 0.0123413f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_131 A N_A_35_297#_c_209_n 0.0249659f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A_c_146_n N_A_35_297#_c_209_n 0.00210097f $X=1.35 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_M1006_g N_VPWR_c_277_n 0.00268723f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_M1004_g N_VPWR_c_277_n 0.00146448f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1006_g N_VPWR_c_279_n 0.00585385f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1004_g N_VPWR_c_281_n 0.00541359f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_M1006_g N_VPWR_c_276_n 0.0106412f $X=0.93 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_M1004_g N_VPWR_c_276_n 0.00952874f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_M1004_g N_A_285_297#_c_325_n 0.00773497f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_c_144_n N_X_c_348_n 5.95155e-19 $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_c_143_n N_VGND_c_379_n 6.98115e-19 $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_143_n N_VGND_c_380_n 0.0073188f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_c_144_n N_VGND_c_380_n 0.00929354f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_143_n N_VGND_c_383_n 0.00341689f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_144_n N_VGND_c_384_n 0.00341689f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_143_n N_VGND_c_386_n 0.00405445f $X=0.93 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_144_n N_VGND_c_386_n 0.00405445f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_35_297#_M1007_g N_VPWR_c_278_n 0.00230662f $X=2.71 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_35_297#_c_197_n N_VPWR_c_279_n 0.0246229f $X=0.3 $Y=2 $X2=0 $Y2=0
cc_150 N_A_35_297#_M1007_g N_VPWR_c_283_n 0.00585385f $X=2.71 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_35_297#_M1009_s N_VPWR_c_276_n 0.00209319f $X=0.175 $Y=1.485 $X2=0
+ $Y2=0
cc_152 N_A_35_297#_M1007_g N_VPWR_c_276_n 0.0129764f $X=2.71 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_35_297#_c_197_n N_VPWR_c_276_n 0.0143524f $X=0.3 $Y=2 $X2=0 $Y2=0
cc_154 N_A_35_297#_c_188_n N_A_285_297#_c_318_n 6.67948e-19 $X=2.615 $Y=1.16
+ $X2=0 $Y2=0
cc_155 N_A_35_297#_c_191_n N_A_285_297#_c_318_n 0.00487667f $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_156 N_A_35_297#_c_188_n N_A_285_297#_c_319_n 0.00624889f $X=2.615 $Y=1.16
+ $X2=0 $Y2=0
cc_157 N_A_35_297#_c_191_n N_A_285_297#_c_319_n 0.00417041f $X=2.25 $Y=1.16
+ $X2=0 $Y2=0
cc_158 N_A_35_297#_c_209_n N_X_M1003_d 0.0156228f $X=2.105 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_35_297#_c_191_n N_X_M1003_d 0.00127987f $X=2.25 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_35_297#_c_187_n N_X_c_348_n 0.00288241f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_35_297#_c_188_n N_X_c_348_n 0.00522174f $X=2.615 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_35_297#_c_209_n N_X_c_348_n 0.0397607f $X=2.105 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_35_297#_c_187_n N_X_c_345_n 0.0154416f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_35_297#_M1007_g N_X_c_345_n 0.00240415f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_35_297#_c_188_n N_X_c_345_n 0.0118816f $X=2.615 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_35_297#_c_189_n N_X_c_345_n 0.0145988f $X=2.615 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_35_297#_c_209_n N_X_c_345_n 0.0138308f $X=2.105 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_35_297#_c_191_n N_X_c_345_n 0.0357973f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_35_297#_M1007_g X 0.0191917f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_35_297#_c_188_n X 0.00130054f $X=2.615 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_35_297#_c_206_n N_VGND_M1005_s 0.00582184f $X=0.635 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_172 N_A_35_297#_c_190_n N_VGND_M1005_s 0.00162259f $X=0.255 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_173 N_A_35_297#_c_192_n N_VGND_M1005_s 9.20807e-19 $X=0.275 $Y=1.785
+ $X2=-0.19 $Y2=-0.24
cc_174 N_A_35_297#_c_209_n N_VGND_M1008_d 0.00335176f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_35_297#_c_190_n N_VGND_c_378_n 9.77208e-19 $X=0.255 $Y=0.74 $X2=0
+ $Y2=0
cc_176 N_A_35_297#_c_206_n N_VGND_c_379_n 0.0108815f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_35_297#_c_190_n N_VGND_c_379_n 0.00971556f $X=0.255 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_35_297#_c_209_n N_VGND_c_380_n 0.0152567f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_35_297#_c_187_n N_VGND_c_382_n 0.00843132f $X=2.69 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_35_297#_c_206_n N_VGND_c_383_n 0.00232396f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_181 N_A_35_297#_c_262_p N_VGND_c_383_n 0.00735006f $X=0.72 $Y=0.5 $X2=0 $Y2=0
cc_182 N_A_35_297#_c_209_n N_VGND_c_383_n 0.00232396f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_35_297#_c_187_n N_VGND_c_384_n 0.00499198f $X=2.69 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_35_297#_c_209_n N_VGND_c_384_n 0.0059291f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_A_35_297#_M1005_d N_VGND_c_386_n 0.0025909f $X=0.585 $Y=0.235 $X2=0
+ $Y2=0
cc_186 N_A_35_297#_c_187_n N_VGND_c_386_n 0.0107744f $X=2.69 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_35_297#_c_206_n N_VGND_c_386_n 0.00506455f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_188 N_A_35_297#_c_190_n N_VGND_c_386_n 0.0021233f $X=0.255 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_35_297#_c_262_p N_VGND_c_386_n 0.00613703f $X=0.72 $Y=0.5 $X2=0 $Y2=0
cc_190 N_A_35_297#_c_209_n N_VGND_c_386_n 0.0171406f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_35_297#_c_209_n A_285_47# 0.00529999f $X=2.105 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_192 A_117_297# N_VPWR_c_276_n 0.0115413f $X=0.585 $Y=1.485 $X2=0.722 $Y2=1.53
cc_193 N_VPWR_c_276_n N_A_285_297#_M1004_d 0.00215201f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_194 N_VPWR_c_276_n N_A_285_297#_M1007_s 0.00209319f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_195 N_VPWR_M1002_d N_A_285_297#_c_318_n 0.0102575f $X=1.845 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_278_n N_A_285_297#_c_318_n 0.0128043f $X=1.98 $Y=2.29 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_276_n N_A_285_297#_c_318_n 0.0121493f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_281_n N_A_285_297#_c_325_n 0.0189039f $X=1.895 $Y=2.72 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_276_n N_A_285_297#_c_325_n 0.0122217f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_278_n N_A_285_297#_c_319_n 0.0269205f $X=1.98 $Y=2.29 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_283_n N_A_285_297#_c_319_n 0.0262277f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_276_n N_A_285_297#_c_319_n 0.0153277f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_276_n N_X_M1007_d 0.00346258f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_204 N_VPWR_c_283_n X 0.0215235f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_205 N_VPWR_c_276_n X 0.0122467f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_206 N_A_285_297#_M1007_s X 0.00193056f $X=2.375 $Y=1.485 $X2=0 $Y2=0
cc_207 N_A_285_297#_c_319_n X 0.00446318f $X=2.5 $Y=1.95 $X2=0 $Y2=0
cc_208 N_X_c_348_n N_VGND_c_380_n 0.00615876f $X=2.505 $Y=0.4 $X2=0 $Y2=0
cc_209 N_X_c_348_n N_VGND_c_382_n 0.0138777f $X=2.505 $Y=0.4 $X2=0 $Y2=0
cc_210 N_X_c_345_n N_VGND_c_382_n 0.0318709f $X=2.59 $Y=1.365 $X2=0 $Y2=0
cc_211 X N_VGND_c_382_n 0.0124789f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_212 N_X_c_348_n N_VGND_c_384_n 0.0417462f $X=2.505 $Y=0.4 $X2=0 $Y2=0
cc_213 N_X_M1003_d N_VGND_c_386_n 0.00636643f $X=1.845 $Y=0.235 $X2=0 $Y2=0
cc_214 N_X_c_348_n N_VGND_c_386_n 0.0334945f $X=2.505 $Y=0.4 $X2=0 $Y2=0
cc_215 N_VGND_c_386_n A_285_47# 0.00323135f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* NGSPICE file created from sky130_fd_sc_hd__nor3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
M1000 Y B VGND VNB nshort w=650000u l=150000u
+  ad=3.965e+11p pd=3.82e+06u as=3.76e+11p ps=3.81e+06u
M1001 a_91_199# C_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=2.915e+11p ps=2.67e+06u
M1002 a_245_297# B a_161_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u
M1003 a_161_297# a_91_199# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1004 a_91_199# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1005 VPWR A a_245_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_91_199# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__and4b_2.pex.spice
* Created: Thu Aug 27 14:08:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4B_2%A_N 3 7 9 10 11 19
r30 16 19 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r31 10 11 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.16
+ $X2=0.235 $Y2=1.53
r32 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r33 9 10 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.235 $Y=0.85
+ $X2=0.235 $Y2=1.16
r34 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r35 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.275
r36 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r37 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%A_27_413# 1 2 7 9 11 13 15 18 20 21 23 25 27
+ 33
r65 34 36 79.2176 $w=2.16e-07 $l=3.55e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=0.805
r66 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r67 30 33 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=1.16
+ $X2=0.89 $Y2=1.16
r68 27 29 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=0.42 $X2=0.7
+ $Y2=0.585
r69 24 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.325
+ $X2=0.72 $Y2=1.16
r70 24 25 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.72 $Y=1.325
+ $X2=0.72 $Y2=1.83
r71 23 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=0.995
+ $X2=0.72 $Y2=1.16
r72 23 29 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.72 $Y=0.995
+ $X2=0.72 $Y2=0.585
r73 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.635 $Y=1.915
+ $X2=0.72 $Y2=1.83
r74 20 21 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.635 $Y=1.915
+ $X2=0.345 $Y2=1.915
r75 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=2
+ $X2=0.345 $Y2=1.915
r76 16 18 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.26 $Y=2 $X2=0.26
+ $Y2=2.3
r77 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.41 $Y=0.73 $X2=1.41
+ $Y2=0.445
r78 12 36 11.3495 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.025 $Y=0.805
+ $X2=0.89 $Y2=0.805
r79 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=0.805
+ $X2=1.41 $Y2=0.73
r80 11 12 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.335 $Y=0.805
+ $X2=1.025 $Y2=0.805
r81 7 34 41.3672 $w=2.16e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r82 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=2.275
r83 2 18 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r84 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%B 3 7 12 13 14 15 16 17 23
r44 16 17 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=1.635 $Y=1.19
+ $X2=1.635 $Y2=1.53
r45 16 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.24 $X2=1.66 $Y2=1.24
r46 15 16 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=1.635 $Y=0.85
+ $X2=1.635 $Y2=1.19
r47 14 15 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=1.635 $Y=0.51
+ $X2=1.635 $Y2=0.85
r48 12 23 49.9064 $w=3.7e-07 $l=3.2e-07 $layer=POLY_cond $X=1.62 $Y=1.56
+ $X2=1.62 $Y2=1.24
r49 12 13 49.8761 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=1.62 $Y=1.56
+ $X2=1.62 $Y2=1.745
r50 10 23 44.4176 $w=3.7e-07 $l=1.5e-07 $layer=POLY_cond $X=1.64 $Y=1.09
+ $X2=1.64 $Y2=1.24
r51 7 10 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=1.77 $Y=0.445
+ $X2=1.77 $Y2=1.09
r52 3 13 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.51 $Y=2.275
+ $X2=1.51 $Y2=1.745
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%C 3 7 9 10 11 12 18
r39 18 21 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.16 $X2=2.2
+ $Y2=1.325
r40 18 20 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.16 $X2=2.2
+ $Y2=0.995
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.16 $X2=2.19 $Y2=1.16
r42 11 12 12.4391 $w=3.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.117 $Y=1.19
+ $X2=2.117 $Y2=1.53
r43 11 19 1.09756 $w=3.13e-07 $l=3e-08 $layer=LI1_cond $X=2.117 $Y=1.19
+ $X2=2.117 $Y2=1.16
r44 10 19 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=2.117 $Y=0.85
+ $X2=2.117 $Y2=1.16
r45 9 10 12.4391 $w=3.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.117 $Y=0.51
+ $X2=2.117 $Y2=0.85
r46 7 21 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.27 $Y=2.275
+ $X2=2.27 $Y2=1.325
r47 3 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.27 $Y=0.445
+ $X2=2.27 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%D 3 7 9 10 11 16
c44 16 0 6.00848e-20 $X=2.69 $Y=1.16
r45 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=1.325
r46 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=0.995
r47 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.16 $X2=2.69 $Y2=1.16
r48 10 11 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.61 $Y=1.19
+ $X2=2.61 $Y2=1.53
r49 10 17 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=2.61 $Y=1.19 $X2=2.61
+ $Y2=1.16
r50 9 17 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.61 $Y=0.85 $X2=2.61
+ $Y2=1.16
r51 7 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.325
r52 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.715 $Y=0.445
+ $X2=2.715 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%A_193_413# 1 2 3 10 12 15 17 19 22 26 30 34
+ 36 39 40 41 44 47 53 59
r112 58 59 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=3.215 $Y=1.16
+ $X2=3.67 $Y2=1.16
r113 54 58 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.17 $Y=1.16
+ $X2=3.215 $Y2=1.16
r114 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.16 $X2=3.17 $Y2=1.16
r115 50 53 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.08 $Y=1.16 $X2=3.17
+ $Y2=1.16
r116 47 49 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.525 $Y=1.88
+ $X2=2.525 $Y2=2
r117 44 46 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=0.42
+ $X2=1.205 $Y2=0.585
r118 41 46 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=1.23 $Y=1.66
+ $X2=1.23 $Y2=0.585
r119 40 42 5.41145 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2
+ $X2=1.165 $Y2=2.085
r120 40 41 15.2072 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=2
+ $X2=1.165 $Y2=1.66
r121 38 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=1.325
+ $X2=3.08 $Y2=1.16
r122 38 39 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.08 $Y=1.325
+ $X2=3.08 $Y2=1.795
r123 37 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.88
+ $X2=2.525 $Y2=1.88
r124 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=1.88
+ $X2=3.08 $Y2=1.795
r125 36 37 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.995 $Y=1.88
+ $X2=2.61 $Y2=1.88
r126 32 49 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=2.085
+ $X2=2.525 $Y2=2
r127 32 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.525 $Y=2.085
+ $X2=2.525 $Y2=2.3
r128 31 40 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.315 $Y=2 $X2=1.165
+ $Y2=2
r129 30 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=2 $X2=2.525
+ $Y2=2
r130 30 31 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=2.44 $Y=2
+ $X2=1.315 $Y2=2
r131 26 42 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.1 $Y=2.3 $X2=1.1
+ $Y2=2.085
r132 20 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r133 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.985
r134 17 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=1.16
r135 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=0.56
r136 13 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.325
+ $X2=3.215 $Y2=1.16
r137 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.215 $Y=1.325
+ $X2=3.215 $Y2=1.985
r138 10 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=0.995
+ $X2=3.215 $Y2=1.16
r139 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.215 $Y=0.995
+ $X2=3.215 $Y2=0.56
r140 3 34 600 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=2.065 $X2=2.525 $Y2=2.3
r141 2 26 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=2.065 $X2=1.1 $Y2=2.3
r142 1 44 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%VPWR 1 2 3 4 15 21 23 25 27 29 34 39 45 50
+ 56 58 62
r71 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r72 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 54 56 9.61451 $w=5.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.07 $Y=2.53
+ $X2=2.225 $Y2=2.53
r74 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r75 52 54 0.217469 $w=5.48e-07 $l=1e-08 $layer=LI1_cond $X=2.06 $Y=2.53 $X2=2.07
+ $Y2=2.53
r76 49 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r77 48 52 9.7861 $w=5.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.61 $Y=2.53 $X2=2.06
+ $Y2=2.53
r78 48 50 7.43982 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=1.61 $Y=2.53
+ $X2=1.555 $Y2=2.53
r79 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r80 46 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 43 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r83 43 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r84 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 40 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=3.005 $Y2=2.72
r86 40 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.17 $Y=2.72
+ $X2=3.45 $Y2=2.72
r87 39 61 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.927 $Y2=2.72
r88 39 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 38 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r90 38 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r91 37 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.225 $Y2=2.72
r92 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r93 34 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=2.72
+ $X2=3.005 $Y2=2.72
r94 34 37 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.84 $Y=2.72
+ $X2=2.53 $Y2=2.72
r95 29 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r96 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 27 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r98 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r99 23 61 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.882 $Y=2.635
+ $X2=3.927 $Y2=2.72
r100 23 25 21.8448 $w=3.33e-07 $l=6.35e-07 $layer=LI1_cond $X=3.882 $Y=2.635
+ $X2=3.882 $Y2=2
r101 19 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=2.635
+ $X2=3.005 $Y2=2.72
r102 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.005 $Y=2.635
+ $X2=3.005 $Y2=2.34
r103 18 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r104 18 50 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.555 $Y2=2.72
r105 13 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r106 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r107 4 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=2
r108 3 21 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.065 $X2=3.005 $Y2=2.34
r109 2 52 300 $w=1.7e-07 $l=5.96867e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=2.065 $X2=2.06 $Y2=2.34
r110 1 15 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%X 1 2 7 8 9 10 11 12 23 38 44
c34 38 0 6.00848e-20 $X=3.905 $Y=0.85
r35 44 49 0.0949269 $w=6.28e-07 $l=5e-09 $layer=LI1_cond $X=3.74 $Y=1.53
+ $X2=3.74 $Y2=1.535
r36 38 47 0.474634 $w=6.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.74 $Y=0.85
+ $X2=3.74 $Y2=0.825
r37 12 50 9.62535 $w=7.13e-07 $l=1.7e-07 $layer=LI1_cond $X=3.697 $Y=1.575
+ $X2=3.697 $Y2=1.745
r38 12 49 0.868241 $w=7.13e-07 $l=4e-08 $layer=LI1_cond $X=3.697 $Y=1.575
+ $X2=3.697 $Y2=1.535
r39 12 44 0.759415 $w=6.28e-07 $l=4e-08 $layer=LI1_cond $X=3.74 $Y=1.49 $X2=3.74
+ $Y2=1.53
r40 11 12 5.69561 $w=6.28e-07 $l=3e-07 $layer=LI1_cond $X=3.74 $Y=1.19 $X2=3.74
+ $Y2=1.49
r41 10 47 1.00031 $w=7.93e-07 $l=3e-08 $layer=LI1_cond $X=3.657 $Y=0.795
+ $X2=3.657 $Y2=0.825
r42 10 46 7.53242 $w=7.93e-07 $l=1.55e-07 $layer=LI1_cond $X=3.657 $Y=0.795
+ $X2=3.657 $Y2=0.64
r43 10 11 5.88547 $w=6.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.74 $Y=0.88
+ $X2=3.74 $Y2=1.19
r44 10 38 0.569561 $w=6.28e-07 $l=3e-08 $layer=LI1_cond $X=3.74 $Y=0.88 $X2=3.74
+ $Y2=0.85
r45 9 31 13.5255 $w=2.03e-07 $l=2.5e-07 $layer=LI1_cond $X=3.442 $Y=2.21
+ $X2=3.442 $Y2=1.96
r46 8 31 4.86918 $w=2.03e-07 $l=9e-08 $layer=LI1_cond $X=3.442 $Y=1.87 $X2=3.442
+ $Y2=1.96
r47 8 50 6.76275 $w=2.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.442 $Y=1.87
+ $X2=3.442 $Y2=1.745
r48 7 46 5.25676 $w=2.83e-07 $l=1.3e-07 $layer=LI1_cond $X=3.402 $Y=0.51
+ $X2=3.402 $Y2=0.64
r49 7 23 3.63929 $w=2.83e-07 $l=9e-08 $layer=LI1_cond $X=3.402 $Y=0.51 $X2=3.402
+ $Y2=0.42
r50 2 31 300 $w=1.7e-07 $l=5.53512e-07 $layer=licon1_PDIFF $count=2 $X=3.29
+ $Y=1.485 $X2=3.46 $Y2=1.96
r51 1 23 182 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.235 $X2=3.46 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_2%VGND 1 2 3 10 12 16 18 20 22 24 32 41 45
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r63 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r64 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r65 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r66 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r67 33 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=2.925
+ $Y2=0
r68 33 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=3.45
+ $Y2=0
r69 32 44 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.927
+ $Y2=0
r70 32 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.45
+ $Y2=0
r71 31 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r72 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r73 28 31 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r74 27 30 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r75 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r76 25 38 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r77 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r78 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.925
+ $Y2=0
r79 24 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.53
+ $Y2=0
r80 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r81 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r82 18 44 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.882 $Y=0.085
+ $X2=3.927 $Y2=0
r83 18 20 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=3.882 $Y=0.085
+ $X2=3.882 $Y2=0.38
r84 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.085
+ $X2=2.925 $Y2=0
r85 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.925 $Y=0.085
+ $X2=2.925 $Y2=0.38
r86 10 38 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r87 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r88 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.38
r89 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.235 $X2=2.925 $Y2=0.38
r90 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


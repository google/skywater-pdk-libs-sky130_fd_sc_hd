* File: sky130_fd_sc_hd__o221a_2.pxi.spice
* Created: Thu Aug 27 14:36:55 2020
* 
x_PM_SKY130_FD_SC_HD__O221A_2%C1 N_C1_c_76_n N_C1_M1006_g N_C1_M1011_g
+ N_C1_c_77_n N_C1_c_78_n C1 C1 PM_SKY130_FD_SC_HD__O221A_2%C1
x_PM_SKY130_FD_SC_HD__O221A_2%B1 N_B1_c_108_n N_B1_M1003_g N_B1_M1005_g B1
+ N_B1_c_110_n PM_SKY130_FD_SC_HD__O221A_2%B1
x_PM_SKY130_FD_SC_HD__O221A_2%B2 N_B2_M1007_g N_B2_M1009_g B2 B2 N_B2_c_148_n
+ N_B2_c_149_n PM_SKY130_FD_SC_HD__O221A_2%B2
x_PM_SKY130_FD_SC_HD__O221A_2%A2 N_A2_M1001_g N_A2_M1010_g A2 A2 N_A2_c_189_n
+ N_A2_c_190_n N_A2_c_191_n PM_SKY130_FD_SC_HD__O221A_2%A2
x_PM_SKY130_FD_SC_HD__O221A_2%A1 N_A1_M1012_g N_A1_c_226_n N_A1_M1013_g A1
+ N_A1_c_228_n PM_SKY130_FD_SC_HD__O221A_2%A1
x_PM_SKY130_FD_SC_HD__O221A_2%A_38_47# N_A_38_47#_M1006_s N_A_38_47#_M1011_s
+ N_A_38_47#_M1009_d N_A_38_47#_c_261_n N_A_38_47#_M1004_g N_A_38_47#_M1000_g
+ N_A_38_47#_c_262_n N_A_38_47#_M1008_g N_A_38_47#_M1002_g N_A_38_47#_c_263_n
+ N_A_38_47#_c_276_n N_A_38_47#_c_264_n N_A_38_47#_c_270_n N_A_38_47#_c_282_n
+ N_A_38_47#_c_305_n N_A_38_47#_c_298_n N_A_38_47#_c_312_n N_A_38_47#_c_271_n
+ N_A_38_47#_c_272_n N_A_38_47#_c_273_n N_A_38_47#_c_265_n N_A_38_47#_c_274_n
+ N_A_38_47#_c_299_n N_A_38_47#_c_329_n N_A_38_47#_c_266_n
+ PM_SKY130_FD_SC_HD__O221A_2%A_38_47#
x_PM_SKY130_FD_SC_HD__O221A_2%VPWR N_VPWR_M1011_d N_VPWR_M1012_d N_VPWR_M1002_d
+ N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n
+ N_VPWR_c_403_n VPWR N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n
+ N_VPWR_c_397_n VPWR PM_SKY130_FD_SC_HD__O221A_2%VPWR
x_PM_SKY130_FD_SC_HD__O221A_2%X N_X_M1004_d N_X_M1000_s N_X_c_471_n N_X_c_473_n
+ N_X_c_477_n N_X_c_478_n N_X_c_466_n X N_X_c_469_n X
+ PM_SKY130_FD_SC_HD__O221A_2%X
x_PM_SKY130_FD_SC_HD__O221A_2%A_141_47# N_A_141_47#_M1006_d N_A_141_47#_M1007_d
+ N_A_141_47#_c_507_n PM_SKY130_FD_SC_HD__O221A_2%A_141_47#
x_PM_SKY130_FD_SC_HD__O221A_2%A_225_47# N_A_225_47#_M1003_d N_A_225_47#_M1001_d
+ N_A_225_47#_c_523_n N_A_225_47#_c_536_n N_A_225_47#_c_524_n
+ PM_SKY130_FD_SC_HD__O221A_2%A_225_47#
x_PM_SKY130_FD_SC_HD__O221A_2%VGND N_VGND_M1001_s N_VGND_M1013_d N_VGND_M1008_s
+ N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n
+ N_VGND_c_564_n N_VGND_c_565_n VGND N_VGND_c_566_n N_VGND_c_567_n
+ N_VGND_c_568_n VGND PM_SKY130_FD_SC_HD__O221A_2%VGND
cc_1 VNB N_C1_c_76_n 0.0183705f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.975
cc_2 VNB N_C1_c_77_n 0.0360749f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_3 VNB N_C1_c_78_n 0.00863986f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.15
cc_4 VNB C1 0.013421f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_5 VNB N_B1_c_108_n 0.0163468f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.975
cc_6 VNB B1 0.00399303f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_7 VNB N_B1_c_110_n 0.0199953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB B2 0.00163232f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_9 VNB N_B2_c_148_n 0.0276719f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_10 VNB N_B2_c_149_n 0.0217056f $X=-0.19 $Y=-0.24 $X2=0.205 $Y2=1.15
cc_11 VNB A2 5.11253e-19 $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.15
cc_12 VNB N_A2_c_189_n 0.0279389f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_13 VNB N_A2_c_190_n 0.00297345f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_14 VNB N_A2_c_191_n 0.0217006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_c_226_n 0.0163355f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.985
cc_16 VNB A1 0.00561882f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_17 VNB N_A1_c_228_n 0.0208016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_38_47#_c_261_n 0.0161247f $X=-0.19 $Y=-0.24 $X2=0.12 $Y2=1.105
cc_19 VNB N_A_38_47#_c_262_n 0.0191379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_38_47#_c_263_n 0.0146062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_38_47#_c_264_n 0.00644512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_38_47#_c_265_n 0.00694881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_38_47#_c_266_n 0.0335883f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_397_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_466_n 0.0114835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0219853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_141_47#_c_507_n 0.00264592f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_225_47#_c_523_n 0.0191936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_225_47#_c_524_n 0.00464057f $X=-0.19 $Y=-0.24 $X2=0.205 $Y2=1.15
cc_30 VNB N_VGND_c_559_n 0.00416643f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.15
cc_31 VNB N_VGND_c_560_n 0.0176326f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_32 VNB N_VGND_c_561_n 0.00571887f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.15
cc_33 VNB N_VGND_c_562_n 0.0106982f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_563_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_564_n 0.0543564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_565_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_566_n 0.0175996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_567_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_568_n 0.225167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_C1_M1011_g 0.0230215f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.985
cc_41 VPB N_C1_c_77_n 0.015268f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.15
cc_42 VPB N_C1_c_78_n 5.21542e-19 $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.15
cc_43 VPB C1 0.00218988f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_44 VPB N_B1_M1005_g 0.0187261f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.985
cc_45 VPB N_B1_c_110_n 0.0041626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_B2_M1009_g 0.0228028f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.985
cc_47 VPB B2 0.00136064f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.15
cc_48 VPB N_B2_c_148_n 0.00766493f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_A2_M1010_g 0.0212875f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.985
cc_50 VPB A2 0.00270944f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.15
cc_51 VPB N_A2_c_189_n 0.00788918f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_52 VPB N_A1_M1012_g 0.0182919f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=0.56
cc_53 VPB N_A1_c_228_n 0.00419406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_38_47#_M1000_g 0.018603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_38_47#_M1002_g 0.0209096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_38_47#_c_264_n 0.00557645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_38_47#_c_270_n 0.00920323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_38_47#_c_271_n 0.00513631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_38_47#_c_272_n 0.00218372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_38_47#_c_273_n 9.75527e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_38_47#_c_274_n 0.00158837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_38_47#_c_266_n 0.00488293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_398_n 0.00506753f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.15
cc_64 VPB N_VPWR_c_399_n 0.00202949f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.15
cc_65 VPB N_VPWR_c_400_n 0.0101786f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.15
cc_66 VPB N_VPWR_c_401_n 0.0137183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_402_n 0.0227999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_403_n 0.00458712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_404_n 0.0461856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_405_n 0.0144994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_406_n 0.00495714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_397_n 0.0491867f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB X 0.0250492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_X_c_469_n 0.00765661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 N_C1_c_76_n N_B1_c_108_n 0.0252809f $X=0.63 $Y=0.975 $X2=-0.19 $Y2=-0.24
cc_76 N_C1_M1011_g N_B1_M1005_g 0.022634f $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_77 N_C1_c_78_n B1 6.39292e-19 $X=0.63 $Y=1.15 $X2=0 $Y2=0
cc_78 N_C1_c_78_n N_B1_c_110_n 0.0210676f $X=0.63 $Y=1.15 $X2=0 $Y2=0
cc_79 N_C1_M1011_g N_A_38_47#_c_276_n 0.00977645f $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_80 N_C1_c_76_n N_A_38_47#_c_264_n 0.00571024f $X=0.63 $Y=0.975 $X2=0 $Y2=0
cc_81 N_C1_M1011_g N_A_38_47#_c_264_n 0.00381586f $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_82 N_C1_c_77_n N_A_38_47#_c_264_n 0.00577431f $X=0.555 $Y=1.15 $X2=0 $Y2=0
cc_83 N_C1_c_78_n N_A_38_47#_c_264_n 0.00545906f $X=0.63 $Y=1.15 $X2=0 $Y2=0
cc_84 C1 N_A_38_47#_c_264_n 0.0215078f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_85 N_C1_M1011_g N_A_38_47#_c_282_n 4.863e-19 $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_86 N_C1_c_76_n N_A_38_47#_c_265_n 0.0100253f $X=0.63 $Y=0.975 $X2=0 $Y2=0
cc_87 N_C1_c_77_n N_A_38_47#_c_265_n 0.0107449f $X=0.555 $Y=1.15 $X2=0 $Y2=0
cc_88 C1 N_A_38_47#_c_265_n 0.0130074f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_89 N_C1_M1011_g N_A_38_47#_c_274_n 0.0131927f $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_90 N_C1_c_77_n N_A_38_47#_c_274_n 0.010045f $X=0.555 $Y=1.15 $X2=0 $Y2=0
cc_91 C1 N_A_38_47#_c_274_n 0.00787756f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_92 N_C1_M1011_g N_VPWR_c_398_n 0.00290109f $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_93 N_C1_M1011_g N_VPWR_c_402_n 0.0054895f $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_94 N_C1_M1011_g N_VPWR_c_397_n 0.010918f $X=0.63 $Y=1.985 $X2=0 $Y2=0
cc_95 N_C1_c_76_n N_A_141_47#_c_507_n 0.00273074f $X=0.63 $Y=0.975 $X2=0 $Y2=0
cc_96 N_C1_c_76_n N_A_225_47#_c_524_n 2.76854e-19 $X=0.63 $Y=0.975 $X2=0 $Y2=0
cc_97 N_C1_c_76_n N_VGND_c_564_n 0.00411332f $X=0.63 $Y=0.975 $X2=0 $Y2=0
cc_98 N_C1_c_76_n N_VGND_c_568_n 0.0068433f $X=0.63 $Y=0.975 $X2=0 $Y2=0
cc_99 N_B1_M1005_g N_B2_M1009_g 0.0712986f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_100 B1 B2 0.0159956f $X=1.04 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B1_c_110_n B2 2.23755e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B1_M1005_g B2 2.21525e-19 $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_c_110_n B2 9.1141e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_104 B1 N_B2_c_148_n 0.00114659f $X=1.04 $Y=1.105 $X2=0 $Y2=0
cc_105 N_B1_c_110_n N_B2_c_148_n 0.0216372f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B1_c_108_n N_B2_c_149_n 0.0270258f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_M1005_g N_A_38_47#_c_276_n 6.30547e-19 $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B1_c_108_n N_A_38_47#_c_264_n 0.0020136f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B1_M1005_g N_A_38_47#_c_264_n 0.00210546f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_110 B1 N_A_38_47#_c_264_n 0.0158213f $X=1.04 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B1_c_110_n N_A_38_47#_c_264_n 0.00311953f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B1_M1005_g N_A_38_47#_c_270_n 0.0151833f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_113 B1 N_A_38_47#_c_270_n 0.0256593f $X=1.04 $Y=1.105 $X2=0 $Y2=0
cc_114 N_B1_c_110_n N_A_38_47#_c_270_n 0.00312275f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B1_M1005_g N_A_38_47#_c_282_n 0.00477737f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B1_M1005_g N_A_38_47#_c_298_n 0.00398406f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B1_M1005_g N_A_38_47#_c_299_n 0.0011746f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_118 N_B1_M1005_g N_VPWR_c_398_n 0.00290109f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B1_M1005_g N_VPWR_c_404_n 0.00559613f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B1_M1005_g N_VPWR_c_397_n 0.00986947f $X=1.11 $Y=1.985 $X2=0 $Y2=0
cc_121 N_B1_c_108_n N_A_141_47#_c_507_n 0.00937225f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_122 B1 N_A_141_47#_c_507_n 0.00426882f $X=1.04 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B1_c_110_n N_A_141_47#_c_507_n 8.43661e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_124 N_B1_c_108_n N_A_225_47#_c_524_n 0.00531066f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_125 B1 N_A_225_47#_c_524_n 0.0108737f $X=1.04 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B1_c_110_n N_A_225_47#_c_524_n 0.00175264f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B1_c_108_n N_VGND_c_564_n 0.00366111f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_c_108_n N_VGND_c_568_n 0.00529554f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B2_M1009_g A2 0.00168105f $X=1.485 $Y=1.985 $X2=0 $Y2=0
cc_130 B2 A2 0.0311571f $X=1.5 $Y=1.445 $X2=0 $Y2=0
cc_131 B2 N_A2_c_189_n 5.92437e-19 $X=1.5 $Y=1.105 $X2=0 $Y2=0
cc_132 N_B2_c_148_n N_A2_c_189_n 0.012064f $X=1.625 $Y=1.16 $X2=0 $Y2=0
cc_133 B2 N_A2_c_190_n 0.0167105f $X=1.5 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B2_c_148_n N_A2_c_190_n 7.88278e-19 $X=1.625 $Y=1.16 $X2=0 $Y2=0
cc_135 B2 N_A_38_47#_M1009_d 0.00468574f $X=1.5 $Y=1.445 $X2=0 $Y2=0
cc_136 N_B2_M1009_g N_A_38_47#_c_270_n 0.00156496f $X=1.485 $Y=1.985 $X2=0 $Y2=0
cc_137 B2 N_A_38_47#_c_270_n 0.0184838f $X=1.5 $Y=1.445 $X2=0 $Y2=0
cc_138 N_B2_M1009_g N_A_38_47#_c_282_n 0.0039954f $X=1.485 $Y=1.985 $X2=0 $Y2=0
cc_139 B2 N_A_38_47#_c_282_n 0.00252222f $X=1.5 $Y=1.445 $X2=0 $Y2=0
cc_140 N_B2_M1009_g N_A_38_47#_c_305_n 0.0102565f $X=1.485 $Y=1.985 $X2=0 $Y2=0
cc_141 B2 N_A_38_47#_c_305_n 0.00229244f $X=1.5 $Y=1.105 $X2=0 $Y2=0
cc_142 B2 N_A_38_47#_c_305_n 0.00367469f $X=1.5 $Y=1.445 $X2=0 $Y2=0
cc_143 N_B2_M1009_g N_A_38_47#_c_299_n 0.00734847f $X=1.485 $Y=1.985 $X2=0 $Y2=0
cc_144 B2 N_A_38_47#_c_299_n 0.0160501f $X=1.5 $Y=1.445 $X2=0 $Y2=0
cc_145 N_B2_c_148_n N_A_38_47#_c_299_n 6.25866e-19 $X=1.625 $Y=1.16 $X2=0 $Y2=0
cc_146 N_B2_M1009_g N_VPWR_c_404_n 0.00426014f $X=1.485 $Y=1.985 $X2=0 $Y2=0
cc_147 N_B2_M1009_g N_VPWR_c_397_n 0.00712214f $X=1.485 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B2_c_149_n N_A_141_47#_c_507_n 0.00816386f $X=1.577 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_B2_c_148_n N_A_225_47#_c_523_n 0.00536062f $X=1.625 $Y=1.16 $X2=0 $Y2=0
cc_150 N_B2_c_149_n N_A_225_47#_c_523_n 0.00751382f $X=1.577 $Y=0.995 $X2=0
+ $Y2=0
cc_151 B2 N_A_225_47#_c_524_n 0.0298732f $X=1.5 $Y=1.105 $X2=0 $Y2=0
cc_152 N_B2_c_149_n N_A_225_47#_c_524_n 0.00794375f $X=1.577 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_B2_c_149_n N_VGND_c_559_n 0.00241512f $X=1.577 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B2_c_149_n N_VGND_c_564_n 0.00366111f $X=1.577 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B2_c_149_n N_VGND_c_568_n 0.0065944f $X=1.577 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_M1010_g N_A1_M1012_g 0.049724f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A2_c_191_n N_A1_c_226_n 0.0124239f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A2_c_189_n A1 0.0012719f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_c_190_n A1 0.0174852f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A2_c_189_n N_A1_c_228_n 0.049724f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A2_c_190_n N_A1_c_228_n 2.22082e-19 $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_162 A2 N_A_38_47#_M1009_d 0.008584f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_163 N_A2_M1010_g N_A_38_47#_c_312_n 0.00910191f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A2_M1010_g N_A_38_47#_c_272_n 0.0041103f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_165 A2 N_A_38_47#_c_272_n 0.00835836f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_166 N_A2_c_190_n N_A_38_47#_c_272_n 7.63998e-19 $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A2_M1010_g N_A_38_47#_c_299_n 0.0100982f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_168 A2 N_A_38_47#_c_299_n 0.0255756f $X=1.98 $Y=1.445 $X2=0 $Y2=0
cc_169 N_A2_c_189_n N_A_38_47#_c_299_n 5.89807e-19 $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A2_c_190_n N_A_38_47#_c_299_n 0.00362757f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A2_M1010_g N_VPWR_c_399_n 0.00271246f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A2_M1010_g N_VPWR_c_404_n 0.00430753f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A2_M1010_g N_VPWR_c_397_n 0.00711996f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A2_c_189_n N_A_225_47#_c_523_n 0.00542239f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A2_c_190_n N_A_225_47#_c_523_n 0.0353147f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A2_c_191_n N_A_225_47#_c_523_n 0.0119689f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A2_c_191_n N_A_225_47#_c_536_n 0.011223f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A2_c_191_n N_VGND_c_559_n 0.00316354f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A2_c_191_n N_VGND_c_560_n 0.00425021f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_191_n N_VGND_c_568_n 0.00709f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_226_n N_A_38_47#_c_261_n 0.012217f $X=2.83 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_M1012_g N_A_38_47#_M1000_g 0.0216984f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A1_M1012_g N_A_38_47#_c_312_n 0.00426825f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A1_M1012_g N_A_38_47#_c_271_n 0.0133047f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_185 A1 N_A_38_47#_c_271_n 0.0320618f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_186 N_A1_c_228_n N_A_38_47#_c_271_n 0.00306699f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A1_M1012_g N_A_38_47#_c_273_n 6.83246e-19 $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A1_c_228_n N_A_38_47#_c_273_n 2.39937e-19 $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A1_M1012_g N_A_38_47#_c_299_n 0.00117263f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_190 A1 N_A_38_47#_c_329_n 0.0170082f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_191 A1 N_A_38_47#_c_266_n 0.00148661f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_192 N_A1_c_228_n N_A_38_47#_c_266_n 0.0224924f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A1_M1012_g N_VPWR_c_399_n 0.0170007f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A1_M1012_g N_VPWR_c_404_n 0.00388479f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A1_M1012_g N_VPWR_c_397_n 0.00660209f $X=2.77 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A1_c_226_n N_A_225_47#_c_523_n 0.00240112f $X=2.83 $Y=0.995 $X2=0 $Y2=0
cc_197 A1 N_A_225_47#_c_523_n 0.0122986f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_198 N_A1_c_228_n N_A_225_47#_c_523_n 0.00179264f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A1_c_226_n N_A_225_47#_c_536_n 0.00509815f $X=2.83 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A1_c_226_n N_VGND_c_560_n 0.00541964f $X=2.83 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A1_c_226_n N_VGND_c_561_n 0.00159991f $X=2.83 $Y=0.995 $X2=0 $Y2=0
cc_202 A1 N_VGND_c_561_n 0.0101626f $X=2.9 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A1_c_228_n N_VGND_c_561_n 2.31083e-19 $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A1_c_226_n N_VGND_c_568_n 0.00955661f $X=2.83 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_38_47#_c_270_n N_VPWR_M1011_d 0.00237235f $X=1.16 $Y=1.557 $X2=-0.19
+ $Y2=-0.24
cc_206 N_A_38_47#_c_271_n N_VPWR_M1012_d 0.00229612f $X=3.245 $Y=1.54 $X2=0
+ $Y2=0
cc_207 N_A_38_47#_c_270_n N_VPWR_c_398_n 0.0171618f $X=1.16 $Y=1.557 $X2=0 $Y2=0
cc_208 N_A_38_47#_M1000_g N_VPWR_c_399_n 0.00154076f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_38_47#_c_312_n N_VPWR_c_399_n 0.00587059f $X=2.54 $Y=1.875 $X2=0
+ $Y2=0
cc_210 N_A_38_47#_c_271_n N_VPWR_c_399_n 0.0212639f $X=3.245 $Y=1.54 $X2=0 $Y2=0
cc_211 N_A_38_47#_c_299_n N_VPWR_c_399_n 0.0140384f $X=2.2 $Y=1.96 $X2=0 $Y2=0
cc_212 N_A_38_47#_M1000_g N_VPWR_c_401_n 4.806e-19 $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_38_47#_M1002_g N_VPWR_c_401_n 0.00836929f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_38_47#_c_276_n N_VPWR_c_402_n 0.0209953f $X=0.415 $Y=2.3 $X2=0 $Y2=0
cc_215 N_A_38_47#_c_305_n N_VPWR_c_404_n 0.00294965f $X=1.55 $Y=1.96 $X2=0 $Y2=0
cc_216 N_A_38_47#_c_298_n N_VPWR_c_404_n 0.00245917f $X=1.33 $Y=1.96 $X2=0 $Y2=0
cc_217 N_A_38_47#_c_299_n N_VPWR_c_404_n 0.0541324f $X=2.2 $Y=1.96 $X2=0 $Y2=0
cc_218 N_A_38_47#_M1000_g N_VPWR_c_405_n 0.00541359f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_38_47#_M1002_g N_VPWR_c_405_n 0.00343969f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_38_47#_M1011_s N_VPWR_c_397_n 0.00335509f $X=0.23 $Y=1.485 $X2=0
+ $Y2=0
cc_221 N_A_38_47#_M1009_d N_VPWR_c_397_n 0.00639913f $X=1.56 $Y=1.485 $X2=0
+ $Y2=0
cc_222 N_A_38_47#_M1000_g N_VPWR_c_397_n 0.00966934f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_38_47#_M1002_g N_VPWR_c_397_n 0.0040221f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_38_47#_c_276_n N_VPWR_c_397_n 0.0124444f $X=0.415 $Y=2.3 $X2=0 $Y2=0
cc_225 N_A_38_47#_c_305_n N_VPWR_c_397_n 0.005334f $X=1.55 $Y=1.96 $X2=0 $Y2=0
cc_226 N_A_38_47#_c_298_n N_VPWR_c_397_n 0.00480871f $X=1.33 $Y=1.96 $X2=0 $Y2=0
cc_227 N_A_38_47#_c_299_n N_VPWR_c_397_n 0.0371063f $X=2.2 $Y=1.96 $X2=0 $Y2=0
cc_228 N_A_38_47#_c_270_n A_237_297# 0.00157343f $X=1.16 $Y=1.557 $X2=-0.19
+ $Y2=-0.24
cc_229 N_A_38_47#_c_282_n A_237_297# 0.00214842f $X=1.245 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_230 N_A_38_47#_c_305_n A_237_297# 0.00124064f $X=1.55 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_231 N_A_38_47#_c_298_n A_237_297# 0.00167595f $X=1.33 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_232 N_A_38_47#_c_312_n A_497_297# 0.00250865f $X=2.54 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_233 N_A_38_47#_c_271_n A_497_297# 4.57867e-19 $X=3.245 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_234 N_A_38_47#_c_299_n A_497_297# 0.00302312f $X=2.2 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_235 N_A_38_47#_c_271_n N_X_M1000_s 0.00202435f $X=3.245 $Y=1.54 $X2=0 $Y2=0
cc_236 N_A_38_47#_c_261_n N_X_c_471_n 0.00524267f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_38_47#_c_262_n N_X_c_471_n 0.0110762f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_38_47#_M1000_g N_X_c_473_n 0.00229286f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A_38_47#_c_271_n N_X_c_473_n 0.00382129f $X=3.245 $Y=1.54 $X2=0 $Y2=0
cc_240 N_A_38_47#_c_329_n N_X_c_473_n 0.00377116f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_38_47#_c_266_n N_X_c_473_n 0.00162837f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_38_47#_M1000_g N_X_c_477_n 0.00465162f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_38_47#_M1002_g N_X_c_478_n 0.0121245f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A_38_47#_c_261_n N_X_c_466_n 0.00254326f $X=3.25 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_38_47#_c_262_n N_X_c_466_n 0.0158689f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_38_47#_c_329_n N_X_c_466_n 0.0202299f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_38_47#_c_266_n N_X_c_466_n 0.00221825f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_38_47#_c_262_n X 0.0282469f $X=3.67 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_38_47#_c_271_n X 0.00548357f $X=3.245 $Y=1.54 $X2=0 $Y2=0
cc_250 N_A_38_47#_c_273_n X 0.00827294f $X=3.33 $Y=1.455 $X2=0 $Y2=0
cc_251 N_A_38_47#_c_329_n X 0.016457f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A_38_47#_M1002_g N_X_c_469_n 0.00340695f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_38_47#_c_265_n N_A_141_47#_c_507_n 0.00221744f $X=0.63 $Y=0.72 $X2=0
+ $Y2=0
cc_254 N_A_38_47#_c_271_n N_A_225_47#_c_523_n 3.54336e-19 $X=3.245 $Y=1.54 $X2=0
+ $Y2=0
cc_255 N_A_38_47#_c_272_n N_A_225_47#_c_523_n 0.00631957f $X=2.625 $Y=1.54 $X2=0
+ $Y2=0
cc_256 N_A_38_47#_c_264_n N_A_225_47#_c_524_n 0.00262277f $X=0.63 $Y=1.445 $X2=0
+ $Y2=0
cc_257 N_A_38_47#_c_270_n N_A_225_47#_c_524_n 0.00385463f $X=1.16 $Y=1.557 $X2=0
+ $Y2=0
cc_258 N_A_38_47#_c_261_n N_VGND_c_561_n 0.00161689f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_38_47#_c_271_n N_VGND_c_561_n 0.00182844f $X=3.245 $Y=1.54 $X2=0
+ $Y2=0
cc_260 N_A_38_47#_c_262_n N_VGND_c_563_n 0.00316354f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_261 N_A_38_47#_c_263_n N_VGND_c_564_n 0.0221115f $X=0.335 $Y=0.36 $X2=0 $Y2=0
cc_262 N_A_38_47#_c_265_n N_VGND_c_564_n 0.00244804f $X=0.63 $Y=0.72 $X2=0 $Y2=0
cc_263 N_A_38_47#_c_261_n N_VGND_c_566_n 0.00540789f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_38_47#_c_262_n N_VGND_c_566_n 0.00423846f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_38_47#_M1006_s N_VGND_c_568_n 0.00316631f $X=0.19 $Y=0.235 $X2=0
+ $Y2=0
cc_266 N_A_38_47#_c_261_n N_VGND_c_568_n 0.00948307f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A_38_47#_c_262_n N_VGND_c_568_n 0.00670547f $X=3.67 $Y=0.995 $X2=0
+ $Y2=0
cc_268 N_A_38_47#_c_263_n N_VGND_c_568_n 0.0124438f $X=0.335 $Y=0.36 $X2=0 $Y2=0
cc_269 N_A_38_47#_c_265_n N_VGND_c_568_n 0.00437724f $X=0.63 $Y=0.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_397_n A_237_297# 0.00275653f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_271 N_VPWR_c_397_n A_497_297# 0.00470663f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_272 N_VPWR_c_397_n N_X_M1000_s 0.00235129f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_273 N_VPWR_c_405_n N_X_c_477_n 0.015017f $X=3.715 $Y=2.72 $X2=0 $Y2=0
cc_274 N_VPWR_c_397_n N_X_c_477_n 0.00931087f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_275 N_VPWR_c_401_n N_X_c_478_n 0.00202396f $X=3.88 $Y=2.3 $X2=0 $Y2=0
cc_276 N_VPWR_c_405_n N_X_c_478_n 0.00221836f $X=3.715 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_397_n N_X_c_478_n 0.00415554f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_M1002_d X 0.00316886f $X=3.745 $Y=1.485 $X2=0 $Y2=0
cc_279 N_VPWR_M1002_d N_X_c_469_n 0.00293827f $X=3.745 $Y=1.485 $X2=0 $Y2=0
cc_280 N_VPWR_c_401_n N_X_c_469_n 0.0216603f $X=3.88 $Y=2.3 $X2=0 $Y2=0
cc_281 N_VPWR_c_397_n N_X_c_469_n 0.0014493f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_282 N_X_c_466_n N_VGND_M1008_s 0.00311706f $X=3.9 $Y=0.905 $X2=0 $Y2=0
cc_283 N_X_c_466_n N_VGND_c_561_n 0.00775692f $X=3.9 $Y=0.905 $X2=0 $Y2=0
cc_284 N_X_c_466_n N_VGND_c_562_n 0.00131872f $X=3.9 $Y=0.905 $X2=0 $Y2=0
cc_285 N_X_c_466_n N_VGND_c_563_n 0.0127122f $X=3.9 $Y=0.905 $X2=0 $Y2=0
cc_286 N_X_c_471_n N_VGND_c_566_n 0.0174129f $X=3.46 $Y=0.39 $X2=0 $Y2=0
cc_287 N_X_c_466_n N_VGND_c_566_n 0.00196939f $X=3.9 $Y=0.905 $X2=0 $Y2=0
cc_288 N_X_M1004_d N_VGND_c_568_n 0.00215535f $X=3.325 $Y=0.235 $X2=0 $Y2=0
cc_289 N_X_c_471_n N_VGND_c_568_n 0.0120402f $X=3.46 $Y=0.39 $X2=0 $Y2=0
cc_290 N_X_c_466_n N_VGND_c_568_n 0.00689009f $X=3.9 $Y=0.905 $X2=0 $Y2=0
cc_291 N_A_141_47#_c_507_n N_A_225_47#_M1003_d 0.00326577f $X=1.68 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_292 N_A_141_47#_M1007_d N_A_225_47#_c_523_n 0.0032442f $X=1.545 $Y=0.235
+ $X2=0 $Y2=0
cc_293 N_A_141_47#_c_507_n N_A_225_47#_c_523_n 0.0151035f $X=1.68 $Y=0.38 $X2=0
+ $Y2=0
cc_294 N_A_141_47#_c_507_n N_A_225_47#_c_524_n 0.0177578f $X=1.68 $Y=0.38 $X2=0
+ $Y2=0
cc_295 N_A_141_47#_c_507_n N_VGND_c_559_n 0.0102966f $X=1.68 $Y=0.38 $X2=0 $Y2=0
cc_296 N_A_141_47#_c_507_n N_VGND_c_564_n 0.0530818f $X=1.68 $Y=0.38 $X2=0 $Y2=0
cc_297 N_A_141_47#_M1006_d N_VGND_c_568_n 0.00216803f $X=0.705 $Y=0.235 $X2=0
+ $Y2=0
cc_298 N_A_141_47#_M1007_d N_VGND_c_568_n 0.00211652f $X=1.545 $Y=0.235 $X2=0
+ $Y2=0
cc_299 N_A_141_47#_c_507_n N_VGND_c_568_n 0.0413007f $X=1.68 $Y=0.38 $X2=0 $Y2=0
cc_300 N_A_225_47#_c_523_n N_VGND_M1001_s 0.00315719f $X=2.455 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_301 N_A_225_47#_c_523_n N_VGND_c_559_n 0.012101f $X=2.455 $Y=0.82 $X2=0 $Y2=0
cc_302 N_A_225_47#_c_523_n N_VGND_c_560_n 0.00193763f $X=2.455 $Y=0.82 $X2=0
+ $Y2=0
cc_303 N_A_225_47#_c_536_n N_VGND_c_560_n 0.0171957f $X=2.62 $Y=0.39 $X2=0 $Y2=0
cc_304 N_A_225_47#_c_523_n N_VGND_c_561_n 0.00787895f $X=2.455 $Y=0.82 $X2=0
+ $Y2=0
cc_305 N_A_225_47#_c_523_n N_VGND_c_564_n 0.00384963f $X=2.455 $Y=0.82 $X2=0
+ $Y2=0
cc_306 N_A_225_47#_M1003_d N_VGND_c_568_n 0.00219239f $X=1.125 $Y=0.235 $X2=0
+ $Y2=0
cc_307 N_A_225_47#_M1001_d N_VGND_c_568_n 0.00215764f $X=2.485 $Y=0.235 $X2=0
+ $Y2=0
cc_308 N_A_225_47#_c_523_n N_VGND_c_568_n 0.0122492f $X=2.455 $Y=0.82 $X2=0
+ $Y2=0
cc_309 N_A_225_47#_c_536_n N_VGND_c_568_n 0.0121066f $X=2.62 $Y=0.39 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dfxtp_4.spice
* Created: Tue Sep  1 19:04:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dfxtp_4.pex.spice"
.subckt sky130_fd_sc_hd__dfxtp_4  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_CLK_M1024_g N_A_27_47#_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_193_47#_M1014_d N_A_27_47#_M1014_g N_VGND_M1024_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_381_47#_M1001_d N_D_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.1092 PD=0.802308 PS=1.36 NRD=2.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1022 N_A_475_413#_M1022_d N_A_27_47#_M1022_g N_A_381_47#_M1001_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0594 AS=0.0609231 PD=0.69 PS=0.687692 NRD=14.988 NRS=11.664
+ M=1 R=2.4 SA=75000.7 SB=75003.4 A=0.054 P=1.02 MULT=1
MM1026 A_572_47# N_A_193_47#_M1026_g N_A_475_413#_M1022_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0634154 AS=0.0594 PD=0.701538 PS=0.69 NRD=40.38 NRS=1.656 M=1
+ R=2.4 SA=75001.1 SB=75002.9 A=0.054 P=1.02 MULT=1
MM1009 N_VGND_M1009_d N_A_634_183#_M1009_g A_572_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.118313 AS=0.0739846 PD=0.966792 PS=0.818462 NRD=47.136 NRS=34.608 M=1
+ R=2.8 SA=75001.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1016 N_A_634_183#_M1016_d N_A_475_413#_M1016_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.126592 AS=0.180287 PD=1.2736 PS=1.47321 NRD=4.68 NRS=25.308
+ M=1 R=4.26667 SA=75001.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1003 N_A_891_413#_M1003_d N_A_193_47#_M1003_g N_A_634_183#_M1016_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0657 AS=0.071208 PD=0.725 PS=0.7164 NRD=26.664 NRS=16.656
+ M=1 R=2.4 SA=75002.9 SB=75001.2 A=0.054 P=1.02 MULT=1
MM1027 A_1020_47# N_A_27_47#_M1027_g N_A_891_413#_M1003_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0657 PD=0.687692 PS=0.725 NRD=38.076 NRS=1.656 M=1
+ R=2.4 SA=75003.4 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1008 N_VGND_M1008_d N_A_1062_300#_M1008_g A_1020_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0710769 PD=1.41 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75003.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_891_413#_M1017_g N_A_1062_300#_M1017_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.105625 AS=0.169 PD=0.975 PS=1.82 NRD=5.532 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75002 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1017_d N_A_1062_300#_M1004_g N_Q_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.08775 PD=0.975 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_1062_300#_M1005_g N_Q_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.08775 PD=0.935 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1005_d N_A_1062_300#_M1010_g N_Q_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.092625 AS=0.08775 PD=0.935 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1029 N_VGND_M1029_d N_A_1062_300#_M1029_g N_Q_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.08775 PD=1.87 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_CLK_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_381_47#_M1018_d N_D_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.1092 PD=0.74 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.8 A=0.063 P=1.14 MULT=1
MM1012 N_A_475_413#_M1012_d N_A_193_47#_M1012_g N_A_381_47#_M1018_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06615 AS=0.0672 PD=0.735 PS=0.74 NRD=9.3772 NRS=21.0987 M=1
+ R=2.8 SA=75000.7 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1006 A_568_413# N_A_27_47#_M1006_g N_A_475_413#_M1012_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0693 AS=0.06615 PD=0.75 PS=0.735 NRD=51.5943 NRS=7.0329 M=1 R=2.8
+ SA=75001.1 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1028 N_VPWR_M1028_d N_A_634_183#_M1028_g A_568_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.128423 AS=0.0693 PD=0.904615 PS=0.75 NRD=111.384 NRS=51.5943 M=1 R=2.8
+ SA=75001.6 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1002 N_A_634_183#_M1002_d N_A_475_413#_M1002_g N_VPWR_M1028_d VPB PHIGHVT
+ L=0.15 W=0.75 AD=0.140385 AS=0.229327 PD=1.37821 PS=1.61538 NRD=0 NRS=0 M=1
+ R=5 SA=75001.4 SB=75001 A=0.1125 P=1.8 MULT=1
MM1019 N_A_891_413#_M1019_d N_A_27_47#_M1019_g N_A_634_183#_M1002_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.0786154 PD=0.69 PS=0.771795 NRD=0 NRS=23.443 M=1
+ R=2.8 SA=75002.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 A_975_413# N_A_193_47#_M1013_g N_A_891_413#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09135 AS=0.0567 PD=0.855 PS=0.69 NRD=76.2193 NRS=0 M=1 R=2.8
+ SA=75003.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_1062_300#_M1020_g A_975_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1218 AS=0.09135 PD=1.42 PS=0.855 NRD=0 NRS=76.2193 M=1 R=2.8 SA=75003.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_891_413#_M1023_g N_A_1062_300#_M1023_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.1625 AS=0.28 PD=1.325 PS=2.56 NRD=5.8903 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75002 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1023_d N_A_1062_300#_M1007_g N_Q_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1625 AS=0.135 PD=1.325 PS=1.27 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_1062_300#_M1015_g N_Q_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1425 AS=0.135 PD=1.285 PS=1.27 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1015_d N_A_1062_300#_M1021_g N_Q_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1425 AS=0.135 PD=1.285 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1025 N_VPWR_M1025_d N_A_1062_300#_M1025_g N_Q_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX30_noxref VNB VPB NWDIODE A=14.6376 P=21.45
c_178 VPB 0 1.42307e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dfxtp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a2111oi_0.spice
* Created: Thu Aug 27 13:58:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2111oi_0.spice.pex"
.subckt sky130_fd_sc_hd__a2111oi_0  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1008 N_Y_M1008_d N_D1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.126 PD=0.7 PS=1.44 NRD=0 NRS=9.996 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_C1_M1002_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=8.568 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=11.424 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_427_47# N_A1_M1003_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g A_427_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 A_169_369# N_D1_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1888 PD=0.85 PS=1.87 NRD=15.3857 NRS=9.2196 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1006 A_241_369# N_C1_M1006_g A_169_369# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0672 PD=0.85 PS=0.85 NRD=15.3857 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_313_369#_M1001_d N_B1_M1001_g A_241_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.9
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_313_369#_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1216 AS=0.0896 PD=1.02 PS=0.92 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_313_369#_M1005_d N_A2_M1005_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1952 AS=0.1216 PD=1.89 PS=1.02 NRD=12.2928 NRS=9.2196 M=1
+ R=4.26667 SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__a2111oi_0.spice.SKY130_FD_SC_HD__A2111OI_0.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a222oi_1.spice
* Created: Tue Sep  1 18:53:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a222oi_1.pex.spice"
.subckt sky130_fd_sc_hd__a222oi_1  VNB VPB C1 C2 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C2	C2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1011 A_109_47# N_C1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.64 AD=0.0672
+ AS=0.1664 PD=0.85 PS=1.8 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2 SB=75002.9
+ A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_C2_M1004_g A_109_47# VNB NSHORT L=0.15 W=0.64 AD=0.2912
+ AS=0.0672 PD=1.55 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75000.5 SB=75002.6
+ A=0.096 P=1.58 MULT=1
MM1003 A_393_47# N_B2_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.64 AD=0.0672
+ AS=0.2912 PD=0.85 PS=1.55 NRD=9.372 NRS=55.308 M=1 R=4.26667 SA=75001.6
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g A_393_47# VNB NSHORT L=0.15 W=0.64 AD=0.1056
+ AS=0.0672 PD=0.97 PS=0.85 NRD=2.808 NRS=9.372 M=1 R=4.26667 SA=75002
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 A_561_47# N_A1_M1006_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.64 AD=0.1056
+ AS=0.1056 PD=0.97 PS=0.97 NRD=20.616 NRS=6.552 M=1 R=4.26667 SA=75002.4
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g A_561_47# VNB NSHORT L=0.15 W=0.64 AD=0.1664
+ AS=0.1056 PD=1.8 PS=0.97 NRD=0 NRS=20.616 M=1 R=4.26667 SA=75002.9 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1009 N_A_109_297#_M1009_d N_C1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_C2_M1001_g N_A_109_297#_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1008 N_A_109_297#_M1008_d N_B2_M1008_g N_A_311_297#_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1007 N_A_311_297#_M1007_d N_B1_M1007_g N_A_109_297#_M1008_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_311_297#_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1000 N_A_311_297#_M1000_d N_A2_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.165 PD=2.52 PS=1.33 NRD=0 NRS=10.8153 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__a222oi_1.pxi.spice"
*
.ends
*
*

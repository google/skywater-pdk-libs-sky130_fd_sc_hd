* File: sky130_fd_sc_hd__bufinv_8.spice.pex
* Created: Thu Aug 27 14:10:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUFINV_8%A 1 3 6 8 14
r24 11 14 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r25 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r26 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r27 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r28 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r29 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_8%A_109_47# 1 2 9 13 17 21 25 29 33 37 40 45
+ 48 50 51 52 57
c94 45 0 1.44067e-19 $X=1.96 $Y=1.16
c95 29 0 1.25206e-19 $X=2.25 $Y=1.985
c96 25 0 1.25206e-19 $X=2.25 $Y=0.56
r97 53 55 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.41 $Y=1.16 $X2=1.83
+ $Y2=1.16
r98 50 51 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.63
+ $X2=0.68 $Y2=1.545
r99 46 57 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=1.96 $Y=1.16
+ $X2=2.25 $Y2=1.16
r100 46 55 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=1.96 $Y=1.16
+ $X2=1.83 $Y2=1.16
r101 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.96
+ $Y=1.16 $X2=1.96 $Y2=1.16
r102 43 52 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=1.175
+ $X2=0.76 $Y2=1.175
r103 43 45 61.8318 $w=1.98e-07 $l=1.115e-06 $layer=LI1_cond $X=0.845 $Y=1.175
+ $X2=1.96 $Y2=1.175
r104 41 52 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.76 $Y=1.275 $X2=0.76
+ $Y2=1.175
r105 41 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.76 $Y=1.275
+ $X2=0.76 $Y2=1.545
r106 40 52 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.76 $Y=1.075 $X2=0.76
+ $Y2=1.175
r107 40 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.76 $Y=1.075
+ $X2=0.76 $Y2=0.905
r108 35 50 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.68 $Y=1.71 $X2=0.68
+ $Y2=1.63
r109 35 37 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=0.68 $Y=1.71 $X2=0.68
+ $Y2=2.31
r110 31 48 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=0.68 $Y2=0.905
r111 31 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=0.68 $Y2=0.4
r112 27 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.16
r113 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.985
r114 23 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=1.16
r115 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=0.56
r116 19 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.16
r117 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.985
r118 15 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=1.16
r119 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=0.56
r120 11 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.16
r121 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.985
r122 7 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.16
r123 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r124 2 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.63
r125 2 37 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.31
r126 1 33 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_8%A_215_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 79 83 87 88 89 90 93 97 102 104 110 114 117 119 130
c245 130 0 1.44067e-19 $X=5.61 $Y=1.16
r246 127 128 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.16
+ $X2=5.19 $Y2=1.16
r247 126 127 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.35 $Y=1.16
+ $X2=4.77 $Y2=1.16
r248 125 126 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.35 $Y2=1.16
r249 124 125 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.51 $Y=1.16
+ $X2=3.93 $Y2=1.16
r250 123 124 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.09 $Y=1.16
+ $X2=3.51 $Y2=1.16
r251 111 130 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.52 $Y=1.16
+ $X2=5.61 $Y2=1.16
r252 111 128 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=5.52 $Y=1.16
+ $X2=5.19 $Y2=1.16
r253 110 111 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=5.52
+ $Y=1.16 $X2=5.52 $Y2=1.16
r254 108 123 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=2.8 $Y=1.16
+ $X2=3.09 $Y2=1.16
r255 108 120 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=2.8 $Y=1.16
+ $X2=2.67 $Y2=1.16
r256 107 110 150.836 $w=1.98e-07 $l=2.72e-06 $layer=LI1_cond $X=2.8 $Y=1.175
+ $X2=5.52 $Y2=1.175
r257 107 108 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=2.8
+ $Y=1.16 $X2=2.8 $Y2=1.16
r258 105 119 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=1.175
+ $X2=2.46 $Y2=1.175
r259 105 107 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.545 $Y=1.175
+ $X2=2.8 $Y2=1.175
r260 104 117 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.445
+ $X2=2.46 $Y2=1.53
r261 103 119 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.46 $Y=1.275
+ $X2=2.46 $Y2=1.175
r262 103 104 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.46 $Y=1.275
+ $X2=2.46 $Y2=1.445
r263 102 119 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.46 $Y=1.075
+ $X2=2.46 $Y2=1.175
r264 101 114 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.905
+ $X2=2.46 $Y2=0.82
r265 101 102 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.46 $Y=0.905
+ $X2=2.46 $Y2=1.075
r266 97 99 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.04 $Y=1.63
+ $X2=2.04 $Y2=2.31
r267 95 117 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.04 $Y=1.53
+ $X2=2.46 $Y2=1.53
r268 95 97 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.04 $Y=1.615
+ $X2=2.04 $Y2=1.63
r269 91 114 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.04 $Y=0.82
+ $X2=2.46 $Y2=0.82
r270 91 93 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=0.735
+ $X2=2.04 $Y2=0.4
r271 89 95 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.53
+ $X2=2.04 $Y2=1.53
r272 89 90 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.875 $Y=1.53
+ $X2=1.365 $Y2=1.53
r273 87 91 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.82
+ $X2=2.04 $Y2=0.82
r274 87 88 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.875 $Y=0.82
+ $X2=1.365 $Y2=0.82
r275 83 85 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.63 $X2=1.2
+ $Y2=2.31
r276 81 90 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.365 $Y2=1.53
r277 81 83 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.2 $Y2=1.63
r278 77 88 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.365 $Y2=0.82
r279 77 79 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.2 $Y2=0.4
r280 73 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.16
r281 73 75 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.985
r282 69 130 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=1.16
r283 69 71 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=0.56
r284 65 128 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.16
r285 65 67 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.985
r286 61 128 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=1.16
r287 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=0.56
r288 57 127 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.16
r289 57 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.985
r290 53 127 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=1.16
r291 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=0.56
r292 49 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.16
r293 49 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.985
r294 45 126 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=1.16
r295 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
r296 41 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.16
r297 41 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.985
r298 37 125 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=1.16
r299 37 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=0.56
r300 33 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.16
r301 33 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.985
r302 29 124 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=1.16
r303 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=0.56
r304 25 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.16
r305 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.985
r306 21 123 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=1.16
r307 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=0.56
r308 17 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.16
r309 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.985
r310 13 120 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=1.16
r311 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=0.56
r312 4 99 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2.31
r313 4 97 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=1.63
r314 3 85 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.31
r315 3 83 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.63
r316 2 93 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.4
r317 1 79 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_8%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 46 48
+ 52 55 56 58 59 61 62 63 64 65 67 87 88 94 97
r95 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r96 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r97 88 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r98 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r99 85 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=5.82 $Y2=2.72
r100 85 87 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=2.72
+ $X2=6.21 $Y2=2.72
r101 84 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r102 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r103 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r104 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r105 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r107 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r108 75 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 72 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=1.62 $Y2=2.72
r111 72 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=2.72
+ $X2=2.07 $Y2=2.72
r112 71 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r113 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 68 91 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r115 68 70 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r116 67 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=1.62 $Y2=2.72
r117 67 70 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 65 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 65 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r120 63 83 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.83 $Y2=2.72
r121 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=2.72
+ $X2=4.98 $Y2=2.72
r122 61 80 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.055 $Y=2.72
+ $X2=3.91 $Y2=2.72
r123 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=2.72
+ $X2=4.14 $Y2=2.72
r124 60 83 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.83 $Y2=2.72
r125 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.14 $Y2=2.72
r126 58 77 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=2.99 $Y2=2.72
r127 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.3 $Y2=2.72
r128 57 80 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.91 $Y2=2.72
r129 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.3 $Y2=2.72
r130 55 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.07 $Y2=2.72
r131 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.72
+ $X2=2.46 $Y2=2.72
r132 54 77 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.99 $Y2=2.72
r133 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=2.72
+ $X2=2.46 $Y2=2.72
r134 50 97 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.72
r135 50 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2
r136 49 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=4.98 $Y2=2.72
r137 48 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.82 $Y2=2.72
r138 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.065 $Y2=2.72
r139 44 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r140 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2
r141 40 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.72
r142 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2
r143 36 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.635 $X2=3.3
+ $Y2=2.72
r144 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.3 $Y=2.635
+ $X2=3.3 $Y2=2
r145 32 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.72
r146 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2
r147 28 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r148 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2
r149 24 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r150 22 91 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r151 22 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r152 7 52 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2
r153 6 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2
r154 5 42 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2
r155 4 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=2
r156 3 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2
r157 2 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=2
r158 1 27 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r159 1 24 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_8%Y 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 73 77 79 81 82 83 84 85 86 88 89
c168 38 0 1.25206e-19 $X=3.045 $Y=1.53
c169 36 0 1.25206e-19 $X=3.045 $Y=0.82
r170 88 89 6.62929 $w=5.53e-07 $l=2.55e-07 $layer=LI1_cond $X=6.162 $Y=1.19
+ $X2=6.162 $Y2=1.445
r171 87 88 8.53107 $w=3.83e-07 $l=2.85e-07 $layer=LI1_cond $X=6.162 $Y=0.905
+ $X2=6.162 $Y2=1.19
r172 80 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=1.53
+ $X2=5.4 $Y2=1.53
r173 79 89 5.71163 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=5.97 $Y=1.53
+ $X2=6.162 $Y2=1.53
r174 79 80 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.97 $Y=1.53
+ $X2=5.565 $Y2=1.53
r175 78 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=0.82
+ $X2=5.4 $Y2=0.82
r176 77 87 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=5.97 $Y=0.82
+ $X2=6.162 $Y2=0.905
r177 77 78 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.97 $Y=0.82
+ $X2=5.565 $Y2=0.82
r178 73 75 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.4 $Y=1.63 $X2=5.4
+ $Y2=2.31
r179 71 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=1.615 $X2=5.4
+ $Y2=1.53
r180 71 73 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.4 $Y=1.615
+ $X2=5.4 $Y2=1.63
r181 67 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=0.735 $X2=5.4
+ $Y2=0.82
r182 67 69 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.4 $Y=0.735
+ $X2=5.4 $Y2=0.4
r183 66 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=1.53
+ $X2=4.56 $Y2=1.53
r184 65 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=1.53
+ $X2=5.4 $Y2=1.53
r185 65 66 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.235 $Y=1.53
+ $X2=4.725 $Y2=1.53
r186 64 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=0.82
+ $X2=4.56 $Y2=0.82
r187 63 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=0.82
+ $X2=5.4 $Y2=0.82
r188 63 64 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.235 $Y=0.82
+ $X2=4.725 $Y2=0.82
r189 59 61 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.56 $Y=1.63
+ $X2=4.56 $Y2=2.31
r190 57 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.56 $Y2=1.53
r191 57 59 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.56 $Y2=1.63
r192 53 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.735
+ $X2=4.56 $Y2=0.82
r193 53 55 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=0.735
+ $X2=4.56 $Y2=0.4
r194 52 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=1.53
+ $X2=3.72 $Y2=1.53
r195 51 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.53
+ $X2=4.56 $Y2=1.53
r196 51 52 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.395 $Y=1.53
+ $X2=3.885 $Y2=1.53
r197 50 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0.82
+ $X2=3.72 $Y2=0.82
r198 49 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0.82
+ $X2=4.56 $Y2=0.82
r199 49 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.395 $Y=0.82
+ $X2=3.885 $Y2=0.82
r200 45 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.72 $Y=1.63
+ $X2=3.72 $Y2=2.31
r201 43 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.615
+ $X2=3.72 $Y2=1.53
r202 43 45 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.72 $Y=1.615
+ $X2=3.72 $Y2=1.63
r203 39 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.735
+ $X2=3.72 $Y2=0.82
r204 39 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.72 $Y=0.735
+ $X2=3.72 $Y2=0.4
r205 37 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=1.53
+ $X2=3.72 $Y2=1.53
r206 37 38 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.555 $Y=1.53
+ $X2=3.045 $Y2=1.53
r207 35 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0.82
+ $X2=3.72 $Y2=0.82
r208 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.555 $Y=0.82
+ $X2=3.045 $Y2=0.82
r209 31 33 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.88 $Y=1.63
+ $X2=2.88 $Y2=2.31
r210 29 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.88 $Y=1.615
+ $X2=3.045 $Y2=1.53
r211 29 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.88 $Y=1.615
+ $X2=2.88 $Y2=1.63
r212 25 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.88 $Y=0.735
+ $X2=3.045 $Y2=0.82
r213 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.88 $Y=0.735
+ $X2=2.88 $Y2=0.4
r214 8 75 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=2.31
r215 8 73 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.63
r216 7 61 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=2.31
r217 7 59 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.63
r218 6 47 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2.31
r219 6 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=1.63
r220 5 33 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2.31
r221 5 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.63
r222 4 69 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.4
r223 3 55 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.4
r224 2 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.4
r225 1 27 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__BUFINV_8%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46
+ 50 53 54 56 57 59 60 61 62 63 65 85 86 92 95
r110 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r111 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r112 86 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r113 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r114 83 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0 $X2=5.82
+ $Y2=0
r115 83 85 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.21 $Y2=0
r116 82 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r117 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r118 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r119 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r120 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r121 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r122 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r123 73 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r124 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r125 70 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.62
+ $Y2=0
r126 70 72 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r127 69 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r128 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r129 66 89 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r130 66 68 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r131 65 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.62
+ $Y2=0
r132 65 68 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=0.69 $Y2=0
r133 63 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r134 63 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r135 61 81 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.83
+ $Y2=0
r136 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.98
+ $Y2=0
r137 59 78 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.055 $Y=0
+ $X2=3.91 $Y2=0
r138 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0 $X2=4.14
+ $Y2=0
r139 58 81 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.83 $Y2=0
r140 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.14
+ $Y2=0
r141 56 75 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=0
+ $X2=2.99 $Y2=0
r142 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.3
+ $Y2=0
r143 55 78 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.385 $Y=0
+ $X2=3.91 $Y2=0
r144 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.3
+ $Y2=0
r145 53 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.07 $Y2=0
r146 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.46
+ $Y2=0
r147 52 75 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=0
+ $X2=2.99 $Y2=0
r148 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.46
+ $Y2=0
r149 48 95 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r150 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.4
r151 47 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r152 46 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.82
+ $Y2=0
r153 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.065 $Y2=0
r154 42 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r155 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.4
r156 38 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r157 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.4
r158 34 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.085 $X2=3.3
+ $Y2=0
r159 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0.4
r160 30 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0
r161 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.4
r162 26 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r163 26 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.4
r164 22 89 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r165 22 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r166 7 50 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.4
r167 6 44 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.4
r168 5 40 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.4
r169 4 36 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.4
r170 3 32 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.4
r171 2 28 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.4
r172 1 24 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends


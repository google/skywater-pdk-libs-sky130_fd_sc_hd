* File: sky130_fd_sc_hd__a22oi_4.pex.spice
* Created: Tue Sep  1 18:53:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A22OI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 35 41
r81 39 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.64 $Y=1.16 $X2=1.73
+ $Y2=1.16
r82 37 39 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.64 $Y2=1.16
r83 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r84 35 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.64
+ $Y=1.16 $X2=1.64 $Y2=1.16
r85 34 36 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.62 $Y=1.16
+ $X2=0.89 $Y2=1.16
r86 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r87 31 34 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.62 $Y2=1.16
r88 29 35 0.20277 $w=1.803e-06 $l=3e-08 $layer=LI1_cond $X=0.992 $Y=1.19
+ $X2=0.992 $Y2=1.16
r89 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r90 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r91 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r93 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r94 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r95 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r96 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r97 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r98 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r99 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r100 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r101 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r102 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r103 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
c68 1 0 1.56657e-19 $X=2.15 $Y=0.995
r69 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.495
+ $Y=1.16 $X2=3.495 $Y2=1.16
r70 38 40 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=3.41 $Y=1.16
+ $X2=3.495 $Y2=1.16
r71 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.41 $Y2=1.16
r72 35 37 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.815 $Y=1.16
+ $X2=2.99 $Y2=1.16
r73 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.815
+ $Y=1.16 $X2=2.815 $Y2=1.16
r74 33 35 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.815 $Y2=1.16
r75 31 33 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r76 29 41 27.7273 $w=1.98e-07 $l=5e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=3.495 $Y2=1.175
r77 29 36 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=2.995 $Y=1.175
+ $X2=2.815 $Y2=1.175
r78 25 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r79 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r80 22 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r81 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r82 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r83 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r84 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r85 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r86 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r87 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r88 8 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r89 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r90 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r91 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325 $X2=2.15
+ $Y2=1.985
r92 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r93 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995 $X2=2.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r63 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.46 $Y=1.16
+ $X2=5.61 $Y2=1.16
r64 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.46
+ $Y=1.16 $X2=5.46 $Y2=1.16
r65 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.19 $Y=1.16
+ $X2=5.46 $Y2=1.16
r66 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.16
+ $X2=5.19 $Y2=1.16
r67 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.44 $Y=1.16
+ $X2=4.77 $Y2=1.16
r68 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.44
+ $Y=1.16 $X2=4.44 $Y2=1.16
r69 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.35 $Y=1.16 $X2=4.44
+ $Y2=1.16
r70 29 40 31.9524 $w=2.08e-07 $l=6.05e-07 $layer=LI1_cond $X=4.855 $Y=1.18
+ $X2=5.46 $Y2=1.18
r71 29 35 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=4.855 $Y=1.18
+ $X2=4.44 $Y2=1.18
r72 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.16
r73 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.985
r74 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.16
r75 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r76 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.16
r77 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.985
r78 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.16
r79 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r80 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.16
r81 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.985
r82 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.16
r83 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r84 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.16
r85 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.35 $Y=1.325 $X2=4.35
+ $Y2=1.985
r86 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.16
r87 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995 $X2=4.35
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r75 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.14 $Y=1.16
+ $X2=7.29 $Y2=1.16
r76 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.14
+ $Y=1.16 $X2=7.14 $Y2=1.16
r77 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.87 $Y=1.16
+ $X2=7.14 $Y2=1.16
r78 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.45 $Y=1.16
+ $X2=6.87 $Y2=1.16
r79 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=6.12 $Y=1.16
+ $X2=6.45 $Y2=1.16
r80 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.12
+ $Y=1.16 $X2=6.12 $Y2=1.16
r81 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.03 $Y=1.16 $X2=6.12
+ $Y2=1.16
r82 29 40 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=6.695 $Y=1.18
+ $X2=7.14 $Y2=1.18
r83 29 35 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=6.695 $Y=1.18
+ $X2=6.12 $Y2=1.18
r84 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.16
r85 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.985
r86 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=1.16
r87 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=0.56
r88 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.16
r89 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.985
r90 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=1.16
r91 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=0.56
r92 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r93 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r94 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r95 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r96 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r97 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325 $X2=6.03
+ $Y2=1.985
r98 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r99 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995 $X2=6.03
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%A_27_297# 1 2 3 4 5 6 7 8 9 28 30 32 36 38
+ 42 44 48 50 52 53 54 58 60 64 66 70 72 74 76 80 81 82 88 90 92
r115 74 94 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=1.625 $X2=7.5
+ $Y2=1.54
r116 74 76 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.5 $Y=1.625
+ $X2=7.5 $Y2=2.3
r117 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=1.54
+ $X2=6.66 $Y2=1.54
r118 72 94 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.375 $Y=1.54
+ $X2=7.5 $Y2=1.54
r119 72 73 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.375 $Y=1.54
+ $X2=6.785 $Y2=1.54
r120 68 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=1.625
+ $X2=6.66 $Y2=1.54
r121 68 70 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.66 $Y=1.625
+ $X2=6.66 $Y2=2.3
r122 67 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=1.54
+ $X2=5.82 $Y2=1.54
r123 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=1.54
+ $X2=6.66 $Y2=1.54
r124 66 67 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.535 $Y=1.54
+ $X2=5.945 $Y2=1.54
r125 62 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=1.625
+ $X2=5.82 $Y2=1.54
r126 62 64 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.82 $Y=1.625
+ $X2=5.82 $Y2=2.3
r127 61 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=1.54
+ $X2=4.98 $Y2=1.54
r128 60 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.695 $Y=1.54
+ $X2=5.82 $Y2=1.54
r129 60 61 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.695 $Y=1.54
+ $X2=5.105 $Y2=1.54
r130 56 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.625
+ $X2=4.98 $Y2=1.54
r131 56 58 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.98 $Y=1.625
+ $X2=4.98 $Y2=2.3
r132 55 84 9.25644 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=4.265 $Y=1.54
+ $X2=3.88 $Y2=1.54
r133 54 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=1.54
+ $X2=4.98 $Y2=1.54
r134 54 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.855 $Y=1.54
+ $X2=4.265 $Y2=1.54
r135 53 86 2.04363 $w=7.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=2.295
+ $X2=3.88 $Y2=2.38
r136 52 84 2.04363 $w=7.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=1.625
+ $X2=3.88 $Y2=1.54
r137 52 53 10.4074 $w=7.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.88 $Y=1.625
+ $X2=3.88 $Y2=2.295
r138 51 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.905 $Y=2.38
+ $X2=2.78 $Y2=2.38
r139 50 86 9.25644 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=3.495 $Y=2.38
+ $X2=3.88 $Y2=2.38
r140 50 51 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.495 $Y=2.38
+ $X2=2.905 $Y2=2.38
r141 46 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.295
+ $X2=2.78 $Y2=2.38
r142 46 48 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.78 $Y=2.295
+ $X2=2.78 $Y2=1.96
r143 45 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.065 $Y=2.38
+ $X2=1.94 $Y2=2.38
r144 44 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=2.38
+ $X2=2.78 $Y2=2.38
r145 44 45 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.655 $Y=2.38
+ $X2=2.065 $Y2=2.38
r146 40 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=1.94 $Y2=2.38
r147 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=1.94 $Y2=1.96
r148 39 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=2.38
+ $X2=1.1 $Y2=2.38
r149 38 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.38
+ $X2=1.94 $Y2=2.38
r150 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.815 $Y=2.38
+ $X2=1.225 $Y2=2.38
r151 34 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.295
+ $X2=1.1 $Y2=2.38
r152 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=2.295
+ $X2=1.1 $Y2=1.96
r153 33 79 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.257 $Y2=2.38
r154 32 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=2.38
+ $X2=1.1 $Y2=2.38
r155 32 33 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.975 $Y=2.38
+ $X2=0.425 $Y2=2.38
r156 28 79 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=2.295
+ $X2=0.257 $Y2=2.38
r157 28 30 22.5328 $w=3.33e-07 $l=6.55e-07 $layer=LI1_cond $X=0.257 $Y=2.295
+ $X2=0.257 $Y2=1.64
r158 9 94 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=1.62
r159 9 76 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=2.3
r160 8 92 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=1.62
r161 8 70 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=2.3
r162 7 90 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=1.62
r163 7 64 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2.3
r164 6 88 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=1.62
r165 6 58 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=2.3
r166 5 86 200 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=3 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2.3
r167 5 84 200 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=3 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.62
r168 4 48 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.96
r169 3 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r170 2 36 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r171 1 79 400 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.32
r172 1 30 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%Y 1 2 3 4 5 6 7 8 29 31 32 41 43 47 49 53 55
+ 56 57
r97 57 60 21.5657 $w=1.78e-07 $l=3.5e-07 $layer=LI1_cond $X=1.155 $Y=1.535
+ $X2=0.805 $Y2=1.535
r98 56 60 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.7 $Y=1.535
+ $X2=0.805 $Y2=1.535
r99 47 57 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=1.395 $Y=1.535
+ $X2=1.155 $Y2=1.535
r100 47 49 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.395 $Y=1.535
+ $X2=1.52 $Y2=1.535
r101 44 53 4.10651 $w=1.8e-07 $l=1.45e-07 $layer=LI1_cond $X=2.485 $Y=1.535
+ $X2=2.34 $Y2=1.535
r102 43 55 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.075 $Y=1.535
+ $X2=3.2 $Y2=1.535
r103 43 44 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=3.075 $Y=1.535
+ $X2=2.485 $Y2=1.535
r104 39 41 40.3355 $w=2.38e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=0.765
+ $X2=5.4 $Y2=0.765
r105 37 39 65.3051 $w=2.38e-07 $l=1.36e-06 $layer=LI1_cond $X=3.2 $Y=0.765
+ $X2=4.56 $Y2=0.765
r106 35 51 3.47969 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=2.445 $Y=0.765
+ $X2=2.32 $Y2=0.765
r107 35 37 36.2539 $w=2.38e-07 $l=7.55e-07 $layer=LI1_cond $X=2.445 $Y=0.765
+ $X2=3.2 $Y2=0.765
r108 32 53 2.1123 $w=2.5e-07 $l=9.94987e-08 $layer=LI1_cond $X=2.32 $Y=1.445
+ $X2=2.34 $Y2=1.535
r109 31 51 3.3405 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=2.32 $Y=0.885
+ $X2=2.32 $Y2=0.765
r110 31 32 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=2.32 $Y=0.885
+ $X2=2.32 $Y2=1.445
r111 30 49 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.645 $Y=1.535
+ $X2=1.52 $Y2=1.535
r112 29 53 4.10651 $w=1.8e-07 $l=1.45e-07 $layer=LI1_cond $X=2.195 $Y=1.535
+ $X2=2.34 $Y2=1.535
r113 29 30 33.8889 $w=1.78e-07 $l=5.5e-07 $layer=LI1_cond $X=2.195 $Y=1.535
+ $X2=1.645 $Y2=1.535
r114 8 55 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.62
r115 7 53 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.62
r116 6 49 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.62
r117 5 56 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.62
r118 4 41 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.73
r119 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.73
r120 2 37 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.73
r121 1 51 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%VPWR 1 2 3 4 15 17 21 25 29 31 32 34 35 36
+ 45 55 56 59 62
r102 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r103 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r104 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r105 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r106 53 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r107 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r108 50 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.365 $Y=2.72
+ $X2=6.24 $Y2=2.72
r109 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.365 $Y=2.72
+ $X2=6.67 $Y2=2.72
r110 49 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 49 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r112 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r113 46 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.525 $Y=2.72
+ $X2=5.4 $Y2=2.72
r114 46 48 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.525 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 45 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.115 $Y=2.72
+ $X2=6.24 $Y2=2.72
r116 45 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.115 $Y=2.72
+ $X2=5.75 $Y2=2.72
r117 44 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 43 44 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r119 39 43 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=4.37 $Y2=2.72
r120 36 44 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=4.37 $Y2=2.72
r121 36 39 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r122 34 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.955 $Y=2.72
+ $X2=6.67 $Y2=2.72
r123 34 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=2.72
+ $X2=7.08 $Y2=2.72
r124 33 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.205 $Y=2.72
+ $X2=7.59 $Y2=2.72
r125 33 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.205 $Y=2.72
+ $X2=7.08 $Y2=2.72
r126 31 43 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.37 $Y2=2.72
r127 31 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.56 $Y2=2.72
r128 27 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=2.635
+ $X2=7.08 $Y2=2.72
r129 27 29 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.08 $Y=2.635
+ $X2=7.08 $Y2=1.96
r130 23 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=2.635
+ $X2=6.24 $Y2=2.72
r131 23 25 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.24 $Y=2.635
+ $X2=6.24 $Y2=1.96
r132 19 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=2.635
+ $X2=5.4 $Y2=2.72
r133 19 21 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.4 $Y=2.635
+ $X2=5.4 $Y2=1.96
r134 18 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.685 $Y=2.72
+ $X2=4.56 $Y2=2.72
r135 17 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.275 $Y=2.72
+ $X2=5.4 $Y2=2.72
r136 17 18 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.275 $Y=2.72
+ $X2=4.685 $Y2=2.72
r137 13 32 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2.72
r138 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=1.96
r139 4 29 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=1.96
r140 3 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.96
r141 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.96
r142 1 15 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 28 29 34
+ 36
c68 29 0 1.56657e-19 $X=1.9 $Y=0.725
r69 32 34 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=0.365
+ $X2=3.62 $Y2=0.365
r70 30 38 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.025 $Y=0.365
+ $X2=1.9 $Y2=0.365
r71 30 32 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.365
+ $X2=2.78 $Y2=0.365
r72 29 40 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.9 $Y=0.725 $X2=1.9
+ $Y2=0.815
r73 28 38 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.9 $Y=0.475 $X2=1.9
+ $Y2=0.365
r74 28 29 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.9 $Y=0.475 $X2=1.9
+ $Y2=0.725
r75 27 36 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0.815
+ $X2=1.1 $Y2=0.815
r76 26 40 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.775 $Y=0.815
+ $X2=1.9 $Y2=0.815
r77 26 27 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=0.815
+ $X2=1.265 $Y2=0.815
r78 22 36 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.1 $Y=0.725 $X2=1.1
+ $Y2=0.815
r79 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.1 $Y=0.725 $X2=1.1
+ $Y2=0.39
r80 20 36 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0.815
+ $X2=1.1 $Y2=0.815
r81 20 21 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=0.815
+ $X2=0.425 $Y2=0.815
r82 16 21 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.425 $Y2=0.815
r83 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.26 $Y2=0.39
r84 5 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.39
r85 4 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.39
r86 3 40 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.73
r87 3 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.39
r88 2 24 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r89 1 18 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 47 56 57 60
r106 60 61 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r107 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r108 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r109 54 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r110 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r111 51 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=0 $X2=6.24
+ $Y2=0
r112 51 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.325 $Y=0 $X2=6.67
+ $Y2=0
r113 50 61 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=6.21
+ $Y2=0
r114 49 50 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r115 47 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=0 $X2=6.24
+ $Y2=0
r116 47 49 296.519 $w=1.68e-07 $l=4.545e-06 $layer=LI1_cond $X=6.155 $Y=0
+ $X2=1.61 $Y2=0
r117 46 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r118 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r119 38 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r120 38 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r121 36 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.995 $Y=0
+ $X2=6.67 $Y2=0
r122 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=0 $X2=7.08
+ $Y2=0
r123 35 56 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.165 $Y=0
+ $X2=7.59 $Y2=0
r124 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.165 $Y=0 $X2=7.08
+ $Y2=0
r125 33 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=0
+ $X2=1.15 $Y2=0
r126 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.52
+ $Y2=0
r127 32 49 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.61
+ $Y2=0
r128 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.52
+ $Y2=0
r129 30 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r130 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r131 29 45 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0
+ $X2=1.15 $Y2=0
r132 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r133 25 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0
r134 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0.39
r135 21 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=0.085
+ $X2=6.24 $Y2=0
r136 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.24 $Y=0.085
+ $X2=6.24 $Y2=0.39
r137 17 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r138 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.39
r139 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r140 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.39
r141 4 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.39
r142 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.39
r143 2 19 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r144 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A22OI_4%A_803_47# 1 2 3 4 5 16 22 23 24 28 30 34 40
r64 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.5 $Y=0.725 $X2=7.5
+ $Y2=0.39
r65 31 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=0.815
+ $X2=6.66 $Y2=0.815
r66 30 32 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=7.335 $Y=0.815
+ $X2=7.5 $Y2=0.725
r67 30 31 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.335 $Y=0.815
+ $X2=6.825 $Y2=0.815
r68 26 40 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.66 $Y=0.725 $X2=6.66
+ $Y2=0.815
r69 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.66 $Y=0.725
+ $X2=6.66 $Y2=0.39
r70 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=5.985 $Y=0.815
+ $X2=5.86 $Y2=0.815
r71 24 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=0.815
+ $X2=6.66 $Y2=0.815
r72 24 25 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.495 $Y=0.815
+ $X2=5.985 $Y2=0.815
r73 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.86 $Y=0.725 $X2=5.86
+ $Y2=0.815
r74 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=5.86 $Y=0.475
+ $X2=5.86 $Y2=0.365
r75 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.86 $Y=0.475
+ $X2=5.86 $Y2=0.725
r76 18 21 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.365
+ $X2=4.98 $Y2=0.365
r77 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.735 $Y=0.365
+ $X2=5.86 $Y2=0.365
r78 16 21 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=5.735 $Y=0.365
+ $X2=4.98 $Y2=0.365
r79 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.365
+ $Y=0.235 $X2=7.5 $Y2=0.39
r80 4 28 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.39
r81 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.73
r82 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.39
r83 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.39
r84 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.39
.ends


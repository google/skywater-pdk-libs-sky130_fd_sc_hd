* File: sky130_fd_sc_hd__a21o_1.spice
* Created: Thu Aug 27 14:00:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21o_1.spice.pex"
.subckt sky130_fd_sc_hd__a21o_1  VNB VPB B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_81_21#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.25675 AS=0.169 PD=1.44 PS=1.82 NRD=15.684 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1005 N_A_81_21#_M1005_d N_B1_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.089375 AS=0.25675 PD=0.925 PS=1.44 NRD=0 NRS=15.684 M=1 R=4.33333
+ SA=75001.1 SB=75001 A=0.0975 P=1.6 MULT=1
MM1002 A_384_47# N_A1_M1002_g N_A_81_21#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.089375 PD=0.93 PS=0.925 NRD=15.684 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g A_384_47# VNB NSHORT L=0.15 W=0.65 AD=0.17225
+ AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75002 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_81_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_A_299_297#_M1007_d N_B1_M1007_g N_A_81_21#_M1007_s VPB PHIGHVT L=0.15
+ W=1 AD=0.1375 AS=0.26 PD=1.275 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_299_297#_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.1375 PD=1.28 PS=1.275 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_A_299_297#_M1001_d N_A2_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__a21o_1.spice.SKY130_FD_SC_HD__A21O_1.pxi"
*
.ends
*
*

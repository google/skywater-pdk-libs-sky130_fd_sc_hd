* File: sky130_fd_sc_hd__nor4b_1.pxi.spice
* Created: Thu Aug 27 14:33:02 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4B_1%A_91_199# N_A_91_199#_M1007_d N_A_91_199#_M1009_d
+ N_A_91_199#_M1006_g N_A_91_199#_M1005_g N_A_91_199#_c_56_n N_A_91_199#_c_57_n
+ N_A_91_199#_c_64_n N_A_91_199#_c_92_p N_A_91_199#_c_58_n N_A_91_199#_c_59_n
+ N_A_91_199#_c_60_n PM_SKY130_FD_SC_HD__NOR4B_1%A_91_199#
x_PM_SKY130_FD_SC_HD__NOR4B_1%C N_C_c_119_n N_C_M1001_g N_C_M1003_g C
+ N_C_c_121_n PM_SKY130_FD_SC_HD__NOR4B_1%C
x_PM_SKY130_FD_SC_HD__NOR4B_1%B N_B_c_155_n N_B_M1002_g N_B_M1008_g B
+ N_B_c_157_n PM_SKY130_FD_SC_HD__NOR4B_1%B
x_PM_SKY130_FD_SC_HD__NOR4B_1%A N_A_M1000_g N_A_M1004_g A N_A_c_192_n
+ N_A_c_193_n PM_SKY130_FD_SC_HD__NOR4B_1%A
x_PM_SKY130_FD_SC_HD__NOR4B_1%D_N N_D_N_M1007_g N_D_N_M1009_g D_N N_D_N_c_225_n
+ N_D_N_c_226_n PM_SKY130_FD_SC_HD__NOR4B_1%D_N
x_PM_SKY130_FD_SC_HD__NOR4B_1%Y N_Y_M1006_d N_Y_M1002_d N_Y_M1005_s N_Y_c_254_n
+ N_Y_c_255_n N_Y_c_285_p N_Y_c_268_n N_Y_c_288_p N_Y_c_271_n Y
+ PM_SKY130_FD_SC_HD__NOR4B_1%Y
x_PM_SKY130_FD_SC_HD__NOR4B_1%VPWR N_VPWR_M1004_d N_VPWR_c_307_n N_VPWR_c_308_n
+ N_VPWR_c_309_n VPWR N_VPWR_c_310_n N_VPWR_c_306_n
+ PM_SKY130_FD_SC_HD__NOR4B_1%VPWR
x_PM_SKY130_FD_SC_HD__NOR4B_1%VGND N_VGND_M1006_s N_VGND_M1001_d N_VGND_M1000_d
+ N_VGND_c_339_n N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n
+ N_VGND_c_344_n N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n VGND
+ N_VGND_c_348_n N_VGND_c_349_n PM_SKY130_FD_SC_HD__NOR4B_1%VGND
cc_1 VNB N_A_91_199#_c_56_n 0.00121137f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_2 VNB N_A_91_199#_c_57_n 0.0293852f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_3 VNB N_A_91_199#_c_58_n 0.0232461f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=1.795
cc_4 VNB N_A_91_199#_c_59_n 0.0195245f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=0.66
cc_5 VNB N_A_91_199#_c_60_n 0.018872f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.995
cc_6 VNB N_C_c_119_n 0.017021f $X=-0.19 $Y=-0.24 $X2=2.61 $Y2=0.465
cc_7 VNB C 0.00348804f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_8 VNB N_C_c_121_n 0.020506f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_9 VNB N_B_c_155_n 0.017021f $X=-0.19 $Y=-0.24 $X2=2.61 $Y2=0.465
cc_10 VNB B 0.0054343f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_11 VNB N_B_c_157_n 0.0185871f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_12 VNB A 0.00485483f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_13 VNB N_A_c_192_n 0.0180732f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_14 VNB N_A_c_193_n 0.0185094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB D_N 0.00582678f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_16 VNB N_D_N_c_225_n 0.0252438f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_17 VNB N_D_N_c_226_n 0.020276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_254_n 0.00144477f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.325
cc_19 VNB N_Y_c_255_n 0.0120961f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_20 VNB Y 0.0256889f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=1.795
cc_21 VNB N_VPWR_c_306_n 0.136896f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=1.9
cc_22 VNB N_VGND_c_339_n 0.0120907f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_23 VNB N_VGND_c_340_n 0.00423911f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_24 VNB N_VGND_c_341_n 0.00773408f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.9
cc_25 VNB N_VGND_c_342_n 0.0122893f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=0.825
cc_26 VNB N_VGND_c_343_n 0.00507259f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=1.795
cc_27 VNB N_VGND_c_344_n 0.0128988f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=0.66
cc_28 VNB N_VGND_c_345_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=0.655
cc_29 VNB N_VGND_c_346_n 0.0136663f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.995
cc_30 VNB N_VGND_c_347_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.325
cc_31 VNB N_VGND_c_348_n 0.0249448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_349_n 0.193506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A_91_199#_M1005_g 0.0233057f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_34 VPB N_A_91_199#_c_56_n 0.00150521f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_35 VPB N_A_91_199#_c_57_n 0.00885875f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_36 VPB N_A_91_199#_c_64_n 0.017699f $X=-0.19 $Y=1.305 $X2=2.965 $Y2=1.9
cc_37 VPB N_A_91_199#_c_58_n 0.0238942f $X=-0.19 $Y=1.305 $X2=3.05 $Y2=1.795
cc_38 VPB N_C_M1003_g 0.0179385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB C 0.00224746f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_40 VPB N_C_c_121_n 0.00450845f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_41 VPB N_B_M1008_g 0.0179385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB B 0.0022251f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_43 VPB N_B_c_157_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_44 VPB N_A_M1004_g 0.01942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB A 0.0022218f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_46 VPB N_A_c_192_n 0.00441099f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_47 VPB N_D_N_M1009_g 0.0369743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB D_N 0.00682299f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_49 VPB N_D_N_c_225_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_50 VPB Y 0.0464574f $X=-0.19 $Y=1.305 $X2=3.05 $Y2=1.795
cc_51 VPB N_VPWR_c_307_n 0.013447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_308_n 0.0594614f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.56
cc_53 VPB N_VPWR_c_309_n 0.00507571f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.325
cc_54 VPB N_VPWR_c_310_n 0.0247367f $X=-0.19 $Y=1.305 $X2=2.745 $Y2=1.9
cc_55 VPB N_VPWR_c_306_n 0.052187f $X=-0.19 $Y=1.305 $X2=2.745 $Y2=1.9
cc_56 N_A_91_199#_c_60_n N_C_c_119_n 0.0248545f $X=0.63 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_57 N_A_91_199#_M1005_g N_C_M1003_g 0.0626524f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_58 N_A_91_199#_c_56_n N_C_M1003_g 0.00130099f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_91_199#_c_64_n N_C_M1003_g 0.0139524f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_60 N_A_91_199#_c_56_n C 0.0363495f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_91_199#_c_57_n C 0.00400813f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_91_199#_c_64_n C 0.0135001f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_63 N_A_91_199#_c_56_n N_C_c_121_n 3.62522e-19 $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_91_199#_c_57_n N_C_c_121_n 0.0207278f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_91_199#_c_64_n N_B_M1008_g 0.0139524f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_66 N_A_91_199#_c_64_n B 0.0160118f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_67 N_A_91_199#_c_64_n N_B_c_157_n 2.96745e-19 $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_68 N_A_91_199#_c_64_n N_A_M1004_g 0.0136464f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_69 N_A_91_199#_c_64_n A 0.0182043f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_70 N_A_91_199#_c_64_n N_A_c_192_n 3.76101e-19 $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_71 N_A_91_199#_c_64_n N_D_N_M1009_g 0.0109277f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_72 N_A_91_199#_c_58_n N_D_N_M1009_g 0.0051527f $X=3.05 $Y=1.795 $X2=0 $Y2=0
cc_73 N_A_91_199#_c_64_n D_N 0.024299f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_74 N_A_91_199#_c_58_n D_N 0.0494524f $X=3.05 $Y=1.795 $X2=0 $Y2=0
cc_75 N_A_91_199#_c_59_n D_N 0.0112662f $X=2.745 $Y=0.66 $X2=0 $Y2=0
cc_76 N_A_91_199#_c_64_n N_D_N_c_225_n 3.57126e-19 $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_77 N_A_91_199#_c_58_n N_D_N_c_225_n 0.00192894f $X=3.05 $Y=1.795 $X2=0 $Y2=0
cc_78 N_A_91_199#_c_59_n N_D_N_c_225_n 0.00147244f $X=2.745 $Y=0.66 $X2=0 $Y2=0
cc_79 N_A_91_199#_c_58_n N_D_N_c_226_n 0.00433654f $X=3.05 $Y=1.795 $X2=0 $Y2=0
cc_80 N_A_91_199#_c_59_n N_D_N_c_226_n 0.00137912f $X=2.745 $Y=0.66 $X2=0 $Y2=0
cc_81 N_A_91_199#_c_56_n N_Y_M1005_s 0.00339944f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_91_199#_c_92_p N_Y_M1005_s 0.00382305f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_83 N_A_91_199#_c_56_n N_Y_c_254_n 0.0148398f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_91_199#_c_57_n N_Y_c_254_n 0.00345222f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_91_199#_c_60_n N_Y_c_254_n 0.0148631f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_91_199#_M1005_g Y 0.0174337f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_91_199#_c_56_n Y 0.0587007f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_91_199#_c_57_n Y 0.00817048f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_91_199#_c_92_p Y 0.0168523f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_90 N_A_91_199#_c_60_n Y 0.00524227f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_91_199#_c_64_n A_161_297# 0.00815962f $X=2.965 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_91_199#_c_64_n A_245_297# 0.011259f $X=2.965 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_91_199#_c_64_n A_341_297# 0.00844147f $X=2.965 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_91_199#_c_64_n N_VPWR_M1004_d 0.00830647f $X=2.965 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_91_199#_c_64_n N_VPWR_c_307_n 0.0196046f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_96 N_A_91_199#_M1005_g N_VPWR_c_308_n 0.00436404f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_97 N_A_91_199#_c_64_n N_VPWR_c_308_n 0.0172676f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_98 N_A_91_199#_c_92_p N_VPWR_c_308_n 0.00299109f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_99 N_A_91_199#_c_64_n N_VPWR_c_310_n 0.0102641f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_100 N_A_91_199#_M1005_g N_VPWR_c_306_n 0.00727084f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_101 N_A_91_199#_c_64_n N_VPWR_c_306_n 0.0543541f $X=2.965 $Y=1.9 $X2=0 $Y2=0
cc_102 N_A_91_199#_c_92_p N_VPWR_c_306_n 0.00576409f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_103 N_A_91_199#_c_60_n N_VGND_c_339_n 0.00831615f $X=0.63 $Y=0.995 $X2=0
+ $Y2=0
cc_104 N_A_91_199#_c_59_n N_VGND_c_341_n 0.00374012f $X=2.745 $Y=0.66 $X2=0
+ $Y2=0
cc_105 N_A_91_199#_c_60_n N_VGND_c_344_n 0.00341689f $X=0.63 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_A_91_199#_c_59_n N_VGND_c_348_n 0.0116646f $X=2.745 $Y=0.66 $X2=0 $Y2=0
cc_107 N_A_91_199#_c_59_n N_VGND_c_349_n 0.0147176f $X=2.745 $Y=0.66 $X2=0 $Y2=0
cc_108 N_A_91_199#_c_60_n N_VGND_c_349_n 0.00405445f $X=0.63 $Y=0.995 $X2=0
+ $Y2=0
cc_109 N_C_c_119_n N_B_c_155_n 0.0214284f $X=1.15 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_110 N_C_M1003_g N_B_M1008_g 0.0524945f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_111 C N_B_M1008_g 8.23281e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_112 N_C_M1003_g B 9.18301e-19 $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_113 C B 0.0495147f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_114 N_C_c_121_n B 0.00181407f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_115 C N_B_c_157_n 3.82144e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_116 N_C_c_121_n N_B_c_157_n 0.0203108f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_117 N_C_c_119_n N_Y_c_268_n 0.0116657f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_118 C N_Y_c_268_n 0.0146924f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_119 N_C_c_121_n N_Y_c_268_n 2.91548e-19 $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_120 C N_Y_c_271_n 0.00439754f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_121 N_C_c_121_n N_Y_c_271_n 2.03831e-19 $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_122 C A_161_297# 0.00163656f $X=1.065 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_123 C A_245_297# 0.00114086f $X=1.065 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_124 N_C_M1003_g N_VPWR_c_308_n 0.00436487f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_125 N_C_M1003_g N_VPWR_c_306_n 0.00627599f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C_c_119_n N_VGND_c_339_n 6.85849e-19 $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_127 N_C_c_119_n N_VGND_c_340_n 0.0016712f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_128 N_C_c_119_n N_VGND_c_344_n 0.00427293f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_129 N_C_c_119_n N_VGND_c_349_n 0.00582284f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B_M1008_g N_A_M1004_g 0.0634554f $X=1.63 $Y=1.985 $X2=0 $Y2=0
cc_131 N_B_M1008_g A 5.46577e-19 $X=1.63 $Y=1.985 $X2=0 $Y2=0
cc_132 B A 0.0459536f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B_c_157_n A 0.00102705f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_134 B N_A_c_192_n 0.00198677f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_135 N_B_c_157_n N_A_c_192_n 0.021372f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B_c_155_n N_A_c_193_n 0.0241532f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B_c_155_n N_Y_c_268_n 0.0113209f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_138 B N_Y_c_268_n 0.0214863f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_139 N_B_c_157_n N_Y_c_268_n 5.02391e-19 $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_140 B A_245_297# 0.00161095f $X=1.525 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_141 B A_341_297# 0.00135642f $X=1.525 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_142 N_B_M1008_g N_VPWR_c_307_n 0.00252342f $X=1.63 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B_M1008_g N_VPWR_c_308_n 0.00436487f $X=1.63 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B_M1008_g N_VPWR_c_306_n 0.00627599f $X=1.63 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B_c_155_n N_VGND_c_340_n 0.0016712f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B_c_155_n N_VGND_c_341_n 8.53588e-19 $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B_c_155_n N_VGND_c_346_n 0.00427293f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_148 N_B_c_155_n N_VGND_c_349_n 0.00582284f $X=1.63 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_M1004_g N_D_N_M1009_g 0.0315743f $X=2.05 $Y=1.985 $X2=0 $Y2=0
cc_150 A N_D_N_M1009_g 0.00101886f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A_M1004_g D_N 7.52786e-19 $X=2.05 $Y=1.985 $X2=0 $Y2=0
cc_152 A D_N 0.0518413f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A_c_192_n D_N 0.0010144f $X=2.11 $Y=1.16 $X2=0 $Y2=0
cc_154 A N_D_N_c_225_n 0.00104813f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_c_192_n N_D_N_c_225_n 0.0213757f $X=2.11 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_193_n N_D_N_c_226_n 0.0125721f $X=2.11 $Y=0.995 $X2=0 $Y2=0
cc_157 A N_VPWR_M1004_d 0.00215779f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_158 N_A_M1004_g N_VPWR_c_307_n 0.0123797f $X=2.05 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_M1004_g N_VPWR_c_308_n 0.00348405f $X=2.05 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_M1004_g N_VPWR_c_306_n 0.00417382f $X=2.05 $Y=1.985 $X2=0 $Y2=0
cc_161 A N_VGND_c_341_n 0.0129188f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A_c_192_n N_VGND_c_341_n 0.00262179f $X=2.11 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_c_193_n N_VGND_c_341_n 0.0119667f $X=2.11 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_193_n N_VGND_c_346_n 0.0046653f $X=2.11 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_193_n N_VGND_c_349_n 0.00799591f $X=2.11 $Y=0.995 $X2=0 $Y2=0
cc_166 N_D_N_M1009_g N_VPWR_c_307_n 0.00128404f $X=2.535 $Y=1.89 $X2=0 $Y2=0
cc_167 N_D_N_M1009_g N_VPWR_c_310_n 0.0032767f $X=2.535 $Y=1.89 $X2=0 $Y2=0
cc_168 N_D_N_M1009_g N_VPWR_c_306_n 0.0046803f $X=2.535 $Y=1.89 $X2=0 $Y2=0
cc_169 N_D_N_c_226_n N_VGND_c_341_n 0.00441624f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_170 N_D_N_c_226_n N_VGND_c_348_n 0.00510437f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_171 N_D_N_c_226_n N_VGND_c_349_n 0.00512902f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_172 Y N_VPWR_c_308_n 0.0166143f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_173 N_Y_M1005_s N_VPWR_c_306_n 0.0111456f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_174 Y N_VPWR_c_306_n 0.00986501f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_175 N_Y_c_254_n N_VGND_M1006_s 0.00767279f $X=0.855 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_176 N_Y_c_268_n N_VGND_M1001_d 0.00919431f $X=1.725 $Y=0.74 $X2=0 $Y2=0
cc_177 N_Y_c_254_n N_VGND_c_339_n 0.0201523f $X=0.855 $Y=0.74 $X2=0 $Y2=0
cc_178 N_Y_c_268_n N_VGND_c_340_n 0.0165818f $X=1.725 $Y=0.74 $X2=0 $Y2=0
cc_179 N_Y_c_255_n N_VGND_c_342_n 0.00506771f $X=0.345 $Y=0.74 $X2=0 $Y2=0
cc_180 N_Y_c_254_n N_VGND_c_344_n 0.00232396f $X=0.855 $Y=0.74 $X2=0 $Y2=0
cc_181 N_Y_c_285_p N_VGND_c_344_n 0.00952714f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_182 N_Y_c_268_n N_VGND_c_344_n 0.00251419f $X=1.725 $Y=0.74 $X2=0 $Y2=0
cc_183 N_Y_c_268_n N_VGND_c_346_n 0.00251419f $X=1.725 $Y=0.74 $X2=0 $Y2=0
cc_184 N_Y_c_288_p N_VGND_c_346_n 0.00906533f $X=1.84 $Y=0.495 $X2=0 $Y2=0
cc_185 N_Y_M1006_d N_VGND_c_349_n 0.00244833f $X=0.805 $Y=0.235 $X2=0 $Y2=0
cc_186 N_Y_M1002_d N_VGND_c_349_n 0.00403782f $X=1.705 $Y=0.235 $X2=0 $Y2=0
cc_187 N_Y_c_254_n N_VGND_c_349_n 0.00588597f $X=0.855 $Y=0.74 $X2=0 $Y2=0
cc_188 N_Y_c_255_n N_VGND_c_349_n 0.00770874f $X=0.345 $Y=0.74 $X2=0 $Y2=0
cc_189 N_Y_c_285_p N_VGND_c_349_n 0.00739742f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_190 N_Y_c_268_n N_VGND_c_349_n 0.00936051f $X=1.725 $Y=0.74 $X2=0 $Y2=0
cc_191 N_Y_c_288_p N_VGND_c_349_n 0.00735151f $X=1.84 $Y=0.495 $X2=0 $Y2=0
cc_192 A_161_297# N_VPWR_c_306_n 0.00347015f $X=0.805 $Y=1.485 $X2=2.745 $Y2=1.9
cc_193 A_245_297# N_VPWR_c_306_n 0.0042413f $X=1.225 $Y=1.485 $X2=2.745 $Y2=1.9
cc_194 A_341_297# N_VPWR_c_306_n 0.00347015f $X=1.705 $Y=1.485 $X2=2.745 $Y2=1.9

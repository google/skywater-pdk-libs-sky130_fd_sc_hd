* File: sky130_fd_sc_hd__lpflow_isobufsrc_16.pxi.spice
* Created: Tue Sep  1 19:12:33 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A N_A_M1025_g N_A_c_248_n N_A_M1038_g
+ N_A_M1036_g N_A_c_249_n N_A_M1043_g N_A_M1047_g N_A_c_250_n N_A_M1049_g
+ N_A_M1059_g N_A_c_251_n N_A_M1064_g A N_A_c_253_n N_A_c_254_n N_A_c_255_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A_143_297# N_A_143_297#_M1038_s
+ N_A_143_297#_M1049_s N_A_143_297#_M1025_d N_A_143_297#_M1047_d
+ N_A_143_297#_c_327_n N_A_143_297#_M1002_g N_A_143_297#_M1000_g
+ N_A_143_297#_c_328_n N_A_143_297#_M1003_g N_A_143_297#_M1001_g
+ N_A_143_297#_c_329_n N_A_143_297#_M1007_g N_A_143_297#_M1004_g
+ N_A_143_297#_c_330_n N_A_143_297#_M1008_g N_A_143_297#_M1005_g
+ N_A_143_297#_c_331_n N_A_143_297#_M1010_g N_A_143_297#_M1009_g
+ N_A_143_297#_c_332_n N_A_143_297#_M1015_g N_A_143_297#_M1011_g
+ N_A_143_297#_c_333_n N_A_143_297#_M1016_g N_A_143_297#_M1019_g
+ N_A_143_297#_c_334_n N_A_143_297#_M1021_g N_A_143_297#_M1020_g
+ N_A_143_297#_c_335_n N_A_143_297#_M1022_g N_A_143_297#_M1023_g
+ N_A_143_297#_c_336_n N_A_143_297#_M1027_g N_A_143_297#_M1031_g
+ N_A_143_297#_c_337_n N_A_143_297#_M1028_g N_A_143_297#_M1032_g
+ N_A_143_297#_c_338_n N_A_143_297#_M1055_g N_A_143_297#_M1039_g
+ N_A_143_297#_c_339_n N_A_143_297#_M1062_g N_A_143_297#_M1048_g
+ N_A_143_297#_c_340_n N_A_143_297#_M1065_g N_A_143_297#_M1053_g
+ N_A_143_297#_c_341_n N_A_143_297#_M1067_g N_A_143_297#_M1057_g
+ N_A_143_297#_c_342_n N_A_143_297#_M1068_g N_A_143_297#_M1060_g
+ N_A_143_297#_c_366_n N_A_143_297#_c_343_n N_A_143_297#_c_373_n
+ N_A_143_297#_c_374_n N_A_143_297#_c_376_n N_A_143_297#_c_344_n
+ N_A_143_297#_c_345_n N_A_143_297#_c_384_n N_A_143_297#_c_363_n
+ N_A_143_297#_c_392_n N_A_143_297#_c_346_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A_143_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%SLEEP N_SLEEP_c_663_n N_SLEEP_M1018_g
+ N_SLEEP_M1006_g N_SLEEP_c_664_n N_SLEEP_M1029_g N_SLEEP_M1012_g
+ N_SLEEP_c_665_n N_SLEEP_M1030_g N_SLEEP_M1013_g N_SLEEP_c_666_n
+ N_SLEEP_M1033_g N_SLEEP_M1014_g N_SLEEP_c_667_n N_SLEEP_M1035_g
+ N_SLEEP_M1017_g N_SLEEP_c_668_n N_SLEEP_M1041_g N_SLEEP_M1024_g
+ N_SLEEP_c_669_n N_SLEEP_M1042_g N_SLEEP_M1026_g N_SLEEP_c_670_n
+ N_SLEEP_M1044_g N_SLEEP_M1034_g N_SLEEP_c_671_n N_SLEEP_M1045_g
+ N_SLEEP_M1037_g N_SLEEP_c_672_n N_SLEEP_M1046_g N_SLEEP_M1040_g
+ N_SLEEP_c_673_n N_SLEEP_M1051_g N_SLEEP_M1050_g N_SLEEP_c_674_n
+ N_SLEEP_M1052_g N_SLEEP_M1054_g N_SLEEP_c_675_n N_SLEEP_M1056_g
+ N_SLEEP_M1061_g N_SLEEP_c_676_n N_SLEEP_M1058_g N_SLEEP_M1069_g
+ N_SLEEP_c_677_n N_SLEEP_M1063_g N_SLEEP_M1070_g N_SLEEP_c_678_n
+ N_SLEEP_M1066_g N_SLEEP_M1071_g SLEEP N_SLEEP_c_679_n N_SLEEP_c_680_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%SLEEP
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%VPWR N_VPWR_M1025_s N_VPWR_M1036_s
+ N_VPWR_M1059_s N_VPWR_M1000_d N_VPWR_M1004_d N_VPWR_M1009_d N_VPWR_M1019_d
+ N_VPWR_M1023_d N_VPWR_M1032_d N_VPWR_M1048_d N_VPWR_M1057_d N_VPWR_c_945_n
+ N_VPWR_c_946_n N_VPWR_c_947_n N_VPWR_c_948_n N_VPWR_c_949_n N_VPWR_c_950_n
+ N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_953_n N_VPWR_c_954_n N_VPWR_c_955_n
+ N_VPWR_c_956_n N_VPWR_c_957_n N_VPWR_c_958_n N_VPWR_c_959_n N_VPWR_c_960_n
+ N_VPWR_c_961_n N_VPWR_c_962_n N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n
+ N_VPWR_c_966_n N_VPWR_c_967_n N_VPWR_c_968_n N_VPWR_c_969_n N_VPWR_c_970_n
+ VPWR N_VPWR_c_971_n N_VPWR_c_972_n N_VPWR_c_973_n N_VPWR_c_944_n
+ N_VPWR_c_975_n N_VPWR_c_976_n N_VPWR_c_977_n N_VPWR_c_978_n N_VPWR_c_979_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A_505_297# N_A_505_297#_M1000_s
+ N_A_505_297#_M1001_s N_A_505_297#_M1005_s N_A_505_297#_M1011_s
+ N_A_505_297#_M1020_s N_A_505_297#_M1031_s N_A_505_297#_M1039_s
+ N_A_505_297#_M1053_s N_A_505_297#_M1060_s N_A_505_297#_M1012_d
+ N_A_505_297#_M1014_d N_A_505_297#_M1024_d N_A_505_297#_M1034_d
+ N_A_505_297#_M1040_d N_A_505_297#_M1054_d N_A_505_297#_M1069_d
+ N_A_505_297#_M1071_d N_A_505_297#_c_1180_n N_A_505_297#_c_1181_n
+ N_A_505_297#_c_1182_n N_A_505_297#_c_1287_n N_A_505_297#_c_1183_n
+ N_A_505_297#_c_1291_n N_A_505_297#_c_1184_n N_A_505_297#_c_1295_n
+ N_A_505_297#_c_1185_n N_A_505_297#_c_1299_n N_A_505_297#_c_1186_n
+ N_A_505_297#_c_1303_n N_A_505_297#_c_1187_n N_A_505_297#_c_1307_n
+ N_A_505_297#_c_1188_n N_A_505_297#_c_1311_n N_A_505_297#_c_1189_n
+ N_A_505_297#_c_1190_n N_A_505_297#_c_1315_n N_A_505_297#_c_1248_n
+ N_A_505_297#_c_1358_p N_A_505_297#_c_1250_n N_A_505_297#_c_1362_p
+ N_A_505_297#_c_1252_n N_A_505_297#_c_1366_p N_A_505_297#_c_1254_n
+ N_A_505_297#_c_1370_p N_A_505_297#_c_1256_n N_A_505_297#_c_1374_p
+ N_A_505_297#_c_1258_n N_A_505_297#_c_1378_p N_A_505_297#_c_1260_n
+ N_A_505_297#_c_1382_p N_A_505_297#_c_1262_n N_A_505_297#_c_1394_p
+ N_A_505_297#_c_1191_n N_A_505_297#_c_1192_n N_A_505_297#_c_1193_n
+ N_A_505_297#_c_1194_n N_A_505_297#_c_1195_n N_A_505_297#_c_1196_n
+ N_A_505_297#_c_1197_n N_A_505_297#_c_1333_n N_A_505_297#_c_1335_n
+ N_A_505_297#_c_1337_n N_A_505_297#_c_1339_n N_A_505_297#_c_1341_n
+ N_A_505_297#_c_1343_n N_A_505_297#_c_1345_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%A_505_297#
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%X N_X_M1002_d N_X_M1007_d N_X_M1010_d
+ N_X_M1016_d N_X_M1022_d N_X_M1028_d N_X_M1062_d N_X_M1067_d N_X_M1018_d
+ N_X_M1030_d N_X_M1035_d N_X_M1042_d N_X_M1045_d N_X_M1051_d N_X_M1056_d
+ N_X_M1063_d N_X_M1006_s N_X_M1013_s N_X_M1017_s N_X_M1026_s N_X_M1037_s
+ N_X_M1050_s N_X_M1061_s N_X_M1070_s N_X_c_1442_n N_X_c_1395_n N_X_c_1396_n
+ N_X_c_1453_n N_X_c_1397_n N_X_c_1461_n N_X_c_1398_n N_X_c_1469_n N_X_c_1399_n
+ N_X_c_1477_n N_X_c_1400_n N_X_c_1485_n N_X_c_1401_n N_X_c_1493_n N_X_c_1402_n
+ N_X_c_1501_n N_X_c_1403_n N_X_c_1506_n N_X_c_1427_n N_X_c_1404_n N_X_c_1549_n
+ N_X_c_1428_n N_X_c_1405_n N_X_c_1561_n N_X_c_1429_n N_X_c_1406_n N_X_c_1573_n
+ N_X_c_1430_n N_X_c_1407_n N_X_c_1585_n N_X_c_1431_n N_X_c_1408_n N_X_c_1597_n
+ N_X_c_1432_n N_X_c_1409_n N_X_c_1609_n N_X_c_1433_n N_X_c_1410_n N_X_c_1621_n
+ N_X_c_1411_n N_X_c_1412_n N_X_c_1413_n N_X_c_1414_n N_X_c_1415_n N_X_c_1416_n
+ N_X_c_1417_n N_X_c_1418_n N_X_c_1434_n N_X_c_1419_n N_X_c_1435_n N_X_c_1420_n
+ N_X_c_1436_n N_X_c_1421_n N_X_c_1437_n N_X_c_1422_n N_X_c_1438_n N_X_c_1423_n
+ N_X_c_1439_n N_X_c_1424_n N_X_c_1440_n N_X_c_1425_n X
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%X
x_PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%VGND N_VGND_M1038_d N_VGND_M1043_d
+ N_VGND_M1064_d N_VGND_M1003_s N_VGND_M1008_s N_VGND_M1015_s N_VGND_M1021_s
+ N_VGND_M1027_s N_VGND_M1055_s N_VGND_M1065_s N_VGND_M1068_s N_VGND_M1029_s
+ N_VGND_M1033_s N_VGND_M1041_s N_VGND_M1044_s N_VGND_M1046_s N_VGND_M1052_s
+ N_VGND_M1058_s N_VGND_M1066_s N_VGND_c_1862_n N_VGND_c_1863_n N_VGND_c_1864_n
+ N_VGND_c_1865_n N_VGND_c_1866_n N_VGND_c_1867_n N_VGND_c_1868_n
+ N_VGND_c_1869_n N_VGND_c_1870_n N_VGND_c_1871_n N_VGND_c_1872_n
+ N_VGND_c_1873_n N_VGND_c_1874_n N_VGND_c_1875_n N_VGND_c_1876_n
+ N_VGND_c_1877_n N_VGND_c_1878_n N_VGND_c_1879_n N_VGND_c_1880_n
+ N_VGND_c_1881_n N_VGND_c_1882_n N_VGND_c_1883_n N_VGND_c_1884_n
+ N_VGND_c_1885_n N_VGND_c_1886_n N_VGND_c_1887_n N_VGND_c_1888_n
+ N_VGND_c_1889_n N_VGND_c_1890_n N_VGND_c_1891_n N_VGND_c_1892_n
+ N_VGND_c_1893_n N_VGND_c_1894_n N_VGND_c_1895_n N_VGND_c_1896_n
+ N_VGND_c_1897_n N_VGND_c_1898_n N_VGND_c_1899_n N_VGND_c_1900_n
+ N_VGND_c_1901_n N_VGND_c_1902_n N_VGND_c_1903_n N_VGND_c_1904_n
+ N_VGND_c_1905_n N_VGND_c_1906_n N_VGND_c_1907_n N_VGND_c_1908_n
+ N_VGND_c_1909_n N_VGND_c_1910_n VGND N_VGND_c_1911_n N_VGND_c_1912_n
+ N_VGND_c_1913_n N_VGND_c_1914_n N_VGND_c_1915_n N_VGND_c_1916_n
+ N_VGND_c_1917_n N_VGND_c_1918_n N_VGND_c_1919_n
+ PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_16%VGND
cc_1 VNB N_A_c_248_n 0.018935f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=0.995
cc_2 VNB N_A_c_249_n 0.0159635f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=0.995
cc_3 VNB N_A_c_250_n 0.0159635f $X=-0.19 $Y=-0.24 $X2=1.7 $Y2=0.995
cc_4 VNB N_A_c_251_n 0.0186566f $X=-0.19 $Y=-0.24 $X2=2.12 $Y2=0.995
cc_5 VNB A 0.0389074f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.105
cc_6 VNB N_A_c_253_n 0.0405569f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_7 VNB N_A_c_254_n 0.0123977f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_8 VNB N_A_c_255_n 0.0745978f $X=-0.19 $Y=-0.24 $X2=2.12 $Y2=1.16
cc_9 VNB N_A_143_297#_c_327_n 0.0185904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_143_297#_c_328_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_143_297#_c_329_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_143_297#_c_330_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_143_297#_c_331_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=1.16
cc_14 VNB N_A_143_297#_c_332_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_143_297#_c_333_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_143_297#_c_334_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_143_297#_c_335_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_143_297#_c_336_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_143_297#_c_337_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_143_297#_c_338_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_143_297#_c_339_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_143_297#_c_340_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_143_297#_c_341_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_143_297#_c_342_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_143_297#_c_343_n 0.00189436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_143_297#_c_344_n 0.00181573f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_143_297#_c_345_n 0.0219196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_143_297#_c_346_n 0.256123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_SLEEP_c_663_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_SLEEP_c_664_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=0.56
cc_31 VNB N_SLEEP_c_665_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.28 $Y2=0.56
cc_32 VNB N_SLEEP_c_666_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.7 $Y2=0.56
cc_33 VNB N_SLEEP_c_667_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.12 $Y2=0.56
cc_34 VNB N_SLEEP_c_668_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_35 VNB N_SLEEP_c_669_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.7 $Y2=1.16
cc_36 VNB N_SLEEP_c_670_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_SLEEP_c_671_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_SLEEP_c_672_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_SLEEP_c_673_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_SLEEP_c_674_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_SLEEP_c_675_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_SLEEP_c_676_n 0.0157999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_SLEEP_c_677_n 0.0157944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_SLEEP_c_678_n 0.019415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_SLEEP_c_679_n 0.00291463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_SLEEP_c_680_n 0.257129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VPWR_c_944_n 0.687231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_1395_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_X_c_1396_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_X_c_1397_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_X_c_1398_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_X_c_1399_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_X_c_1400_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_X_c_1401_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_X_c_1402_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_X_c_1403_n 0.00350899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_X_c_1404_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_X_c_1405_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_X_c_1406_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_X_c_1407_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_X_c_1408_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_X_c_1409_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_X_c_1410_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_X_c_1411_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_X_c_1412_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_X_c_1413_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_X_c_1414_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_X_c_1415_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_X_c_1416_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_X_c_1417_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_X_c_1418_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_X_c_1419_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_X_c_1420_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_X_c_1421_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_X_c_1422_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_X_c_1423_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_X_c_1424_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_X_c_1425_n 0.014806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB X 0.0213757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1862_n 0.00972945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1863_n 0.00600292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1864_n 0.0113004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1865_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1866_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1867_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1868_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1869_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1870_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1871_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1872_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1873_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1874_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1875_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1876_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1877_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1878_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1879_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1880_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1881_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1882_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1883_n 0.0151454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1884_n 0.0174928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1885_n 0.0144349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1886_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1887_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1888_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1889_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1890_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1891_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1892_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1893_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1894_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1895_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1896_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1897_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1898_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1899_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1900_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1901_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1902_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1903_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1904_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1905_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1906_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1907_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1908_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1909_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1910_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1911_n 0.015432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1912_n 0.0163782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1913_n 0.0166671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1914_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1915_n 0.0105758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1916_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1917_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1918_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1919_n 0.742627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VPB N_A_M1025_g 0.0259429f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.985
cc_139 VPB N_A_M1036_g 0.0178058f $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.985
cc_140 VPB N_A_M1047_g 0.0178058f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.985
cc_141 VPB N_A_M1059_g 0.0245269f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.985
cc_142 VPB N_A_c_253_n 0.0192162f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_143 VPB N_A_c_254_n 0.00150435f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_144 VPB N_A_c_255_n 0.0185697f $X=-0.19 $Y=1.305 $X2=2.12 $Y2=1.16
cc_145 VPB N_A_143_297#_M1000_g 0.0252703f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.985
cc_146 VPB N_A_143_297#_M1001_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.985
cc_147 VPB N_A_143_297#_M1004_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_143_297#_M1005_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=1.16
cc_149 VPB N_A_143_297#_M1009_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_143_297#_M1011_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_143_297#_M1019_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_143_297#_M1020_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_143_297#_M1023_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_143_297#_M1031_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_143_297#_M1032_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_143_297#_M1039_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_143_297#_M1048_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_143_297#_M1053_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_143_297#_M1057_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_143_297#_M1060_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_143_297#_c_363_n 0.00150087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_143_297#_c_346_n 0.0466477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_SLEEP_M1006_g 0.018818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_SLEEP_M1012_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_SLEEP_M1013_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_SLEEP_M1014_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_SLEEP_M1017_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_SLEEP_M1024_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.28 $Y2=1.16
cc_169 VPB N_SLEEP_M1026_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_SLEEP_M1034_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_SLEEP_M1037_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_SLEEP_M1040_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_SLEEP_M1050_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_SLEEP_M1054_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_SLEEP_M1061_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_SLEEP_M1069_g 0.0182211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_SLEEP_M1070_g 0.01821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_SLEEP_M1071_g 0.022286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_SLEEP_c_680_n 0.0465992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_945_n 0.0394562f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_181 VPB N_VPWR_c_946_n 0.00531853f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.16
cc_182 VPB N_VPWR_c_947_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_948_n 0.0152805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_949_n 0.019061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_950_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_951_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_952_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_953_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_954_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_955_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_956_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_957_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_958_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_959_n 0.0116899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_960_n 0.00410625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_961_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_962_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_963_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_964_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_965_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_966_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_967_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_968_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_969_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_970_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_971_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_972_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_973_n 0.172195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_944_n 0.0717783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_975_n 0.00468329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_976_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_977_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_978_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_979_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_A_505_297#_c_1180_n 0.00513784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_505_297#_c_1181_n 0.00795082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_505_297#_c_1182_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_505_297#_c_1183_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_505_297#_c_1184_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_505_297#_c_1185_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_505_297#_c_1186_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_505_297#_c_1187_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_505_297#_c_1188_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_505_297#_c_1189_n 0.00235943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_505_297#_c_1190_n 0.00364086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_505_297#_c_1191_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_505_297#_c_1192_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_505_297#_c_1193_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_505_297#_c_1194_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_A_505_297#_c_1195_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_505_297#_c_1196_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_505_297#_c_1197_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_X_c_1427_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_X_c_1428_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_X_c_1429_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_X_c_1430_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_X_c_1431_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_X_c_1432_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_X_c_1433_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_X_c_1434_n 0.00224497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_X_c_1435_n 0.0020229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_X_c_1436_n 0.0020229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_X_c_1437_n 0.0020229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_X_c_1438_n 0.0020229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_X_c_1439_n 0.0020229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_X_c_1440_n 0.0020229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB X 0.0291233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 N_A_c_251_n N_A_143_297#_c_327_n 0.0057288f $X=2.12 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_M1025_g N_A_143_297#_c_366_n 0.00907982f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_M1036_g N_A_143_297#_c_366_n 0.00862502f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A_c_248_n N_A_143_297#_c_343_n 0.00146787f $X=0.86 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_c_249_n N_A_143_297#_c_343_n 0.00143714f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_253 A N_A_143_297#_c_343_n 0.00415255f $X=0.295 $Y=1.105 $X2=0 $Y2=0
cc_254 N_A_c_254_n N_A_143_297#_c_343_n 0.0031658f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_c_255_n N_A_143_297#_c_343_n 0.0074827f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_c_255_n N_A_143_297#_c_373_n 0.0253502f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_c_254_n N_A_143_297#_c_374_n 0.0182332f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_c_255_n N_A_143_297#_c_374_n 0.026587f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_M1036_g N_A_143_297#_c_376_n 6.76316e-19 $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_M1047_g N_A_143_297#_c_376_n 0.0148618f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A_M1059_g N_A_143_297#_c_376_n 0.0188314f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A_c_255_n N_A_143_297#_c_376_n 0.00611296f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_c_250_n N_A_143_297#_c_344_n 0.00147598f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_c_251_n N_A_143_297#_c_344_n 0.00258381f $X=2.12 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_c_255_n N_A_143_297#_c_344_n 0.00847892f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_c_255_n N_A_143_297#_c_345_n 0.0154386f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A_M1025_g N_A_143_297#_c_384_n 0.00253838f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A_M1036_g N_A_143_297#_c_384_n 0.00172083f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A_c_255_n N_A_143_297#_c_384_n 0.00132308f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_M1025_g N_A_143_297#_c_363_n 0.00370237f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_M1036_g N_A_143_297#_c_363_n 0.00379809f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_M1047_g N_A_143_297#_c_363_n 6.77474e-19 $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_c_254_n N_A_143_297#_c_363_n 0.00294328f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A_c_255_n N_A_143_297#_c_363_n 0.00421806f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_275 N_A_c_255_n N_A_143_297#_c_392_n 0.0296064f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_c_255_n N_A_143_297#_c_346_n 0.0057288f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_M1025_g N_VPWR_c_945_n 0.00319321f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A_c_253_n N_VPWR_c_945_n 0.00494369f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A_c_254_n N_VPWR_c_945_n 0.0173274f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_M1036_g N_VPWR_c_946_n 0.00166947f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_M1047_g N_VPWR_c_946_n 0.00166947f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A_c_255_n N_VPWR_c_946_n 0.00257112f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A_M1047_g N_VPWR_c_947_n 0.00541359f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A_M1059_g N_VPWR_c_947_n 0.00541359f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A_M1059_g N_VPWR_c_948_n 0.00387648f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A_c_255_n N_VPWR_c_948_n 0.00482783f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A_M1025_g N_VPWR_c_961_n 0.00541359f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A_M1036_g N_VPWR_c_961_n 0.00541359f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A_M1025_g N_VPWR_c_944_n 0.0105836f $X=0.64 $Y=1.985 $X2=0 $Y2=0
cc_290 N_A_M1036_g N_VPWR_c_944_n 0.00950154f $X=1.06 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_M1047_g N_VPWR_c_944_n 0.00950154f $X=1.48 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A_M1059_g N_VPWR_c_944_n 0.0108276f $X=1.9 $Y=1.985 $X2=0 $Y2=0
cc_293 N_A_c_248_n N_VGND_c_1862_n 0.0120101f $X=0.86 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_c_249_n N_VGND_c_1862_n 6.31592e-19 $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_295 A N_VGND_c_1862_n 0.0462006f $X=0.295 $Y=1.105 $X2=0 $Y2=0
cc_296 N_A_c_253_n N_VGND_c_1862_n 0.00837176f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A_c_254_n N_VGND_c_1862_n 0.0148126f $X=0.58 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A_c_249_n N_VGND_c_1863_n 0.00159847f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A_c_250_n N_VGND_c_1863_n 0.00165327f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A_c_255_n N_VGND_c_1863_n 0.00266542f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A_c_251_n N_VGND_c_1864_n 0.00242763f $X=2.12 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A_c_248_n N_VGND_c_1885_n 0.0046653f $X=0.86 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A_c_249_n N_VGND_c_1885_n 0.00585385f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_304 A N_VGND_c_1911_n 0.0163465f $X=0.295 $Y=1.105 $X2=0 $Y2=0
cc_305 N_A_c_250_n N_VGND_c_1912_n 0.00585385f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_c_251_n N_VGND_c_1912_n 0.00585385f $X=2.12 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_c_248_n N_VGND_c_1919_n 0.00789179f $X=0.86 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_c_249_n N_VGND_c_1919_n 0.0104367f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_c_250_n N_VGND_c_1919_n 0.0104367f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A_c_251_n N_VGND_c_1919_n 0.0110911f $X=2.12 $Y=0.995 $X2=0 $Y2=0
cc_311 A N_VGND_c_1919_n 0.00878068f $X=0.295 $Y=1.105 $X2=0 $Y2=0
cc_312 N_A_143_297#_c_342_n N_SLEEP_c_663_n 0.0195911f $X=9.18 $Y=0.995
+ $X2=-0.19 $Y2=-0.24
cc_313 N_A_143_297#_M1060_g N_SLEEP_M1006_g 0.0195911f $X=9.18 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_143_297#_c_345_n N_SLEEP_c_679_n 0.0194016f $X=9.09 $Y=1.16 $X2=0
+ $Y2=0
cc_315 N_A_143_297#_c_346_n N_SLEEP_c_679_n 7.73302e-19 $X=9.18 $Y=1.16 $X2=0
+ $Y2=0
cc_316 N_A_143_297#_c_345_n N_SLEEP_c_680_n 6.90123e-19 $X=9.09 $Y=1.16 $X2=0
+ $Y2=0
cc_317 N_A_143_297#_c_346_n N_SLEEP_c_680_n 0.0195911f $X=9.18 $Y=1.16 $X2=0
+ $Y2=0
cc_318 N_A_143_297#_c_374_n N_VPWR_c_946_n 0.0137165f $X=1.195 $Y=1.175 $X2=0
+ $Y2=0
cc_319 N_A_143_297#_c_376_n N_VPWR_c_946_n 0.0389887f $X=1.69 $Y=1.62 $X2=0
+ $Y2=0
cc_320 N_A_143_297#_c_363_n N_VPWR_c_946_n 0.0387837f $X=0.85 $Y=1.495 $X2=0
+ $Y2=0
cc_321 N_A_143_297#_c_376_n N_VPWR_c_947_n 0.0189039f $X=1.69 $Y=1.62 $X2=0
+ $Y2=0
cc_322 N_A_143_297#_M1000_g N_VPWR_c_948_n 0.00365775f $X=2.88 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_143_297#_c_376_n N_VPWR_c_948_n 0.0390509f $X=1.69 $Y=1.62 $X2=0
+ $Y2=0
cc_324 N_A_143_297#_c_345_n N_VPWR_c_948_n 0.0193948f $X=9.09 $Y=1.16 $X2=0
+ $Y2=0
cc_325 N_A_143_297#_c_392_n N_VPWR_c_948_n 7.60021e-19 $X=1.78 $Y=1.175 $X2=0
+ $Y2=0
cc_326 N_A_143_297#_M1000_g N_VPWR_c_949_n 0.00585385f $X=2.88 $Y=1.985 $X2=0
+ $Y2=0
cc_327 N_A_143_297#_M1000_g N_VPWR_c_950_n 0.00302074f $X=2.88 $Y=1.985 $X2=0
+ $Y2=0
cc_328 N_A_143_297#_M1001_g N_VPWR_c_950_n 0.00157837f $X=3.3 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A_143_297#_M1004_g N_VPWR_c_951_n 0.00157837f $X=3.72 $Y=1.985 $X2=0
+ $Y2=0
cc_330 N_A_143_297#_M1005_g N_VPWR_c_951_n 0.00157837f $X=4.14 $Y=1.985 $X2=0
+ $Y2=0
cc_331 N_A_143_297#_M1009_g N_VPWR_c_952_n 0.00157837f $X=4.56 $Y=1.985 $X2=0
+ $Y2=0
cc_332 N_A_143_297#_M1011_g N_VPWR_c_952_n 0.00157837f $X=4.98 $Y=1.985 $X2=0
+ $Y2=0
cc_333 N_A_143_297#_M1019_g N_VPWR_c_953_n 0.00157837f $X=5.4 $Y=1.985 $X2=0
+ $Y2=0
cc_334 N_A_143_297#_M1020_g N_VPWR_c_953_n 0.00157837f $X=5.82 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_143_297#_M1023_g N_VPWR_c_954_n 0.00157837f $X=6.24 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A_143_297#_M1031_g N_VPWR_c_954_n 0.00157837f $X=6.66 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A_143_297#_M1032_g N_VPWR_c_955_n 0.00157837f $X=7.08 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A_143_297#_M1039_g N_VPWR_c_955_n 0.00157837f $X=7.5 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A_143_297#_M1039_g N_VPWR_c_956_n 0.00585385f $X=7.5 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_143_297#_M1048_g N_VPWR_c_956_n 0.00585385f $X=7.92 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_143_297#_M1048_g N_VPWR_c_957_n 0.00157837f $X=7.92 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_143_297#_M1053_g N_VPWR_c_957_n 0.00157837f $X=8.34 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_143_297#_M1057_g N_VPWR_c_958_n 0.00157837f $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_143_297#_M1060_g N_VPWR_c_958_n 0.00302074f $X=9.18 $Y=1.985 $X2=0
+ $Y2=0
cc_345 N_A_143_297#_c_366_n N_VPWR_c_961_n 0.0189039f $X=0.85 $Y=2.3 $X2=0 $Y2=0
cc_346 N_A_143_297#_M1005_g N_VPWR_c_963_n 0.00585385f $X=4.14 $Y=1.985 $X2=0
+ $Y2=0
cc_347 N_A_143_297#_M1009_g N_VPWR_c_963_n 0.00585385f $X=4.56 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_A_143_297#_M1011_g N_VPWR_c_965_n 0.00585385f $X=4.98 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_143_297#_M1019_g N_VPWR_c_965_n 0.00585385f $X=5.4 $Y=1.985 $X2=0
+ $Y2=0
cc_350 N_A_143_297#_M1020_g N_VPWR_c_967_n 0.00585385f $X=5.82 $Y=1.985 $X2=0
+ $Y2=0
cc_351 N_A_143_297#_M1023_g N_VPWR_c_967_n 0.00585385f $X=6.24 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A_143_297#_M1031_g N_VPWR_c_969_n 0.00585385f $X=6.66 $Y=1.985 $X2=0
+ $Y2=0
cc_353 N_A_143_297#_M1032_g N_VPWR_c_969_n 0.00585385f $X=7.08 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_143_297#_M1001_g N_VPWR_c_971_n 0.00585385f $X=3.3 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A_143_297#_M1004_g N_VPWR_c_971_n 0.00585385f $X=3.72 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A_143_297#_M1053_g N_VPWR_c_972_n 0.00585385f $X=8.34 $Y=1.985 $X2=0
+ $Y2=0
cc_357 N_A_143_297#_M1057_g N_VPWR_c_972_n 0.00585385f $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_358 N_A_143_297#_M1060_g N_VPWR_c_973_n 0.00585385f $X=9.18 $Y=1.985 $X2=0
+ $Y2=0
cc_359 N_A_143_297#_M1025_d N_VPWR_c_944_n 0.00215201f $X=0.715 $Y=1.485 $X2=0
+ $Y2=0
cc_360 N_A_143_297#_M1047_d N_VPWR_c_944_n 0.00215201f $X=1.555 $Y=1.485 $X2=0
+ $Y2=0
cc_361 N_A_143_297#_M1000_g N_VPWR_c_944_n 0.0117628f $X=2.88 $Y=1.985 $X2=0
+ $Y2=0
cc_362 N_A_143_297#_M1001_g N_VPWR_c_944_n 0.0104367f $X=3.3 $Y=1.985 $X2=0
+ $Y2=0
cc_363 N_A_143_297#_M1004_g N_VPWR_c_944_n 0.0104367f $X=3.72 $Y=1.985 $X2=0
+ $Y2=0
cc_364 N_A_143_297#_M1005_g N_VPWR_c_944_n 0.0104367f $X=4.14 $Y=1.985 $X2=0
+ $Y2=0
cc_365 N_A_143_297#_M1009_g N_VPWR_c_944_n 0.0104367f $X=4.56 $Y=1.985 $X2=0
+ $Y2=0
cc_366 N_A_143_297#_M1011_g N_VPWR_c_944_n 0.0104367f $X=4.98 $Y=1.985 $X2=0
+ $Y2=0
cc_367 N_A_143_297#_M1019_g N_VPWR_c_944_n 0.0104367f $X=5.4 $Y=1.985 $X2=0
+ $Y2=0
cc_368 N_A_143_297#_M1020_g N_VPWR_c_944_n 0.0104367f $X=5.82 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_A_143_297#_M1023_g N_VPWR_c_944_n 0.0104367f $X=6.24 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A_143_297#_M1031_g N_VPWR_c_944_n 0.0104367f $X=6.66 $Y=1.985 $X2=0
+ $Y2=0
cc_371 N_A_143_297#_M1032_g N_VPWR_c_944_n 0.0104367f $X=7.08 $Y=1.985 $X2=0
+ $Y2=0
cc_372 N_A_143_297#_M1039_g N_VPWR_c_944_n 0.0104367f $X=7.5 $Y=1.985 $X2=0
+ $Y2=0
cc_373 N_A_143_297#_M1048_g N_VPWR_c_944_n 0.0104367f $X=7.92 $Y=1.985 $X2=0
+ $Y2=0
cc_374 N_A_143_297#_M1053_g N_VPWR_c_944_n 0.0104367f $X=8.34 $Y=1.985 $X2=0
+ $Y2=0
cc_375 N_A_143_297#_M1057_g N_VPWR_c_944_n 0.0104367f $X=8.76 $Y=1.985 $X2=0
+ $Y2=0
cc_376 N_A_143_297#_M1060_g N_VPWR_c_944_n 0.010464f $X=9.18 $Y=1.985 $X2=0
+ $Y2=0
cc_377 N_A_143_297#_c_366_n N_VPWR_c_944_n 0.0122217f $X=0.85 $Y=2.3 $X2=0 $Y2=0
cc_378 N_A_143_297#_c_376_n N_VPWR_c_944_n 0.0122217f $X=1.69 $Y=1.62 $X2=0
+ $Y2=0
cc_379 N_A_143_297#_c_345_n N_A_505_297#_c_1180_n 0.0274221f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_380 N_A_143_297#_M1000_g N_A_505_297#_c_1182_n 0.0147299f $X=2.88 $Y=1.985
+ $X2=0 $Y2=0
cc_381 N_A_143_297#_M1001_g N_A_505_297#_c_1182_n 0.0144778f $X=3.3 $Y=1.985
+ $X2=0 $Y2=0
cc_382 N_A_143_297#_c_345_n N_A_505_297#_c_1182_n 0.0423927f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_383 N_A_143_297#_c_346_n N_A_505_297#_c_1182_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_384 N_A_143_297#_M1004_g N_A_505_297#_c_1183_n 0.0144778f $X=3.72 $Y=1.985
+ $X2=0 $Y2=0
cc_385 N_A_143_297#_M1005_g N_A_505_297#_c_1183_n 0.0144778f $X=4.14 $Y=1.985
+ $X2=0 $Y2=0
cc_386 N_A_143_297#_c_345_n N_A_505_297#_c_1183_n 0.042354f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_387 N_A_143_297#_c_346_n N_A_505_297#_c_1183_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_388 N_A_143_297#_M1009_g N_A_505_297#_c_1184_n 0.0144778f $X=4.56 $Y=1.985
+ $X2=0 $Y2=0
cc_389 N_A_143_297#_M1011_g N_A_505_297#_c_1184_n 0.0144778f $X=4.98 $Y=1.985
+ $X2=0 $Y2=0
cc_390 N_A_143_297#_c_345_n N_A_505_297#_c_1184_n 0.042354f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_391 N_A_143_297#_c_346_n N_A_505_297#_c_1184_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_392 N_A_143_297#_M1019_g N_A_505_297#_c_1185_n 0.0144778f $X=5.4 $Y=1.985
+ $X2=0 $Y2=0
cc_393 N_A_143_297#_M1020_g N_A_505_297#_c_1185_n 0.0144778f $X=5.82 $Y=1.985
+ $X2=0 $Y2=0
cc_394 N_A_143_297#_c_345_n N_A_505_297#_c_1185_n 0.042354f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_395 N_A_143_297#_c_346_n N_A_505_297#_c_1185_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_396 N_A_143_297#_M1023_g N_A_505_297#_c_1186_n 0.0144778f $X=6.24 $Y=1.985
+ $X2=0 $Y2=0
cc_397 N_A_143_297#_M1031_g N_A_505_297#_c_1186_n 0.0144778f $X=6.66 $Y=1.985
+ $X2=0 $Y2=0
cc_398 N_A_143_297#_c_345_n N_A_505_297#_c_1186_n 0.042354f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_399 N_A_143_297#_c_346_n N_A_505_297#_c_1186_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_400 N_A_143_297#_M1032_g N_A_505_297#_c_1187_n 0.0144778f $X=7.08 $Y=1.985
+ $X2=0 $Y2=0
cc_401 N_A_143_297#_M1039_g N_A_505_297#_c_1187_n 0.0144778f $X=7.5 $Y=1.985
+ $X2=0 $Y2=0
cc_402 N_A_143_297#_c_345_n N_A_505_297#_c_1187_n 0.042354f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_403 N_A_143_297#_c_346_n N_A_505_297#_c_1187_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_404 N_A_143_297#_M1048_g N_A_505_297#_c_1188_n 0.0144778f $X=7.92 $Y=1.985
+ $X2=0 $Y2=0
cc_405 N_A_143_297#_M1053_g N_A_505_297#_c_1188_n 0.0144778f $X=8.34 $Y=1.985
+ $X2=0 $Y2=0
cc_406 N_A_143_297#_c_345_n N_A_505_297#_c_1188_n 0.042354f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_407 N_A_143_297#_c_346_n N_A_505_297#_c_1188_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_408 N_A_143_297#_M1057_g N_A_505_297#_c_1189_n 0.0144232f $X=8.76 $Y=1.985
+ $X2=0 $Y2=0
cc_409 N_A_143_297#_M1060_g N_A_505_297#_c_1189_n 0.0144195f $X=9.18 $Y=1.985
+ $X2=0 $Y2=0
cc_410 N_A_143_297#_c_345_n N_A_505_297#_c_1189_n 0.0423927f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_411 N_A_143_297#_c_346_n N_A_505_297#_c_1189_n 0.00212577f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_412 N_A_143_297#_c_345_n N_A_505_297#_c_1190_n 0.00128541f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_413 N_A_143_297#_c_345_n N_A_505_297#_c_1191_n 0.0204549f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_414 N_A_143_297#_c_346_n N_A_505_297#_c_1191_n 0.00220041f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_415 N_A_143_297#_c_345_n N_A_505_297#_c_1192_n 0.0204549f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_416 N_A_143_297#_c_346_n N_A_505_297#_c_1192_n 0.00220041f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_417 N_A_143_297#_c_345_n N_A_505_297#_c_1193_n 0.0204549f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_418 N_A_143_297#_c_346_n N_A_505_297#_c_1193_n 0.00220041f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_419 N_A_143_297#_c_345_n N_A_505_297#_c_1194_n 0.0204549f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_420 N_A_143_297#_c_346_n N_A_505_297#_c_1194_n 0.00220041f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_421 N_A_143_297#_c_345_n N_A_505_297#_c_1195_n 0.0204549f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_422 N_A_143_297#_c_346_n N_A_505_297#_c_1195_n 0.00220041f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_423 N_A_143_297#_c_345_n N_A_505_297#_c_1196_n 0.0204549f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_424 N_A_143_297#_c_346_n N_A_505_297#_c_1196_n 0.00220041f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_425 N_A_143_297#_c_345_n N_A_505_297#_c_1197_n 0.0204549f $X=9.09 $Y=1.16
+ $X2=0 $Y2=0
cc_426 N_A_143_297#_c_346_n N_A_505_297#_c_1197_n 0.00220041f $X=9.18 $Y=1.16
+ $X2=0 $Y2=0
cc_427 N_A_143_297#_c_327_n N_X_c_1442_n 0.00539651f $X=2.88 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A_143_297#_c_328_n N_X_c_1442_n 0.00630972f $X=3.3 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A_143_297#_c_329_n N_X_c_1442_n 5.22228e-19 $X=3.72 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A_143_297#_c_328_n N_X_c_1395_n 0.00870364f $X=3.3 $Y=0.995 $X2=0 $Y2=0
cc_431 N_A_143_297#_c_329_n N_X_c_1395_n 0.00870364f $X=3.72 $Y=0.995 $X2=0
+ $Y2=0
cc_432 N_A_143_297#_c_345_n N_X_c_1395_n 0.0362443f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_433 N_A_143_297#_c_346_n N_X_c_1395_n 0.00222133f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_434 N_A_143_297#_c_327_n N_X_c_1396_n 0.00262807f $X=2.88 $Y=0.995 $X2=0
+ $Y2=0
cc_435 N_A_143_297#_c_328_n N_X_c_1396_n 0.00113286f $X=3.3 $Y=0.995 $X2=0 $Y2=0
cc_436 N_A_143_297#_c_345_n N_X_c_1396_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_143_297#_c_346_n N_X_c_1396_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_438 N_A_143_297#_c_328_n N_X_c_1453_n 5.22228e-19 $X=3.3 $Y=0.995 $X2=0 $Y2=0
cc_439 N_A_143_297#_c_329_n N_X_c_1453_n 0.00630972f $X=3.72 $Y=0.995 $X2=0
+ $Y2=0
cc_440 N_A_143_297#_c_330_n N_X_c_1453_n 0.00630972f $X=4.14 $Y=0.995 $X2=0
+ $Y2=0
cc_441 N_A_143_297#_c_331_n N_X_c_1453_n 5.22228e-19 $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_442 N_A_143_297#_c_330_n N_X_c_1397_n 0.00870364f $X=4.14 $Y=0.995 $X2=0
+ $Y2=0
cc_443 N_A_143_297#_c_331_n N_X_c_1397_n 0.00870364f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_444 N_A_143_297#_c_345_n N_X_c_1397_n 0.0362443f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_445 N_A_143_297#_c_346_n N_X_c_1397_n 0.00222133f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_446 N_A_143_297#_c_330_n N_X_c_1461_n 5.22228e-19 $X=4.14 $Y=0.995 $X2=0
+ $Y2=0
cc_447 N_A_143_297#_c_331_n N_X_c_1461_n 0.00630972f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_448 N_A_143_297#_c_332_n N_X_c_1461_n 0.00630972f $X=4.98 $Y=0.995 $X2=0
+ $Y2=0
cc_449 N_A_143_297#_c_333_n N_X_c_1461_n 5.22228e-19 $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_450 N_A_143_297#_c_332_n N_X_c_1398_n 0.00870364f $X=4.98 $Y=0.995 $X2=0
+ $Y2=0
cc_451 N_A_143_297#_c_333_n N_X_c_1398_n 0.00870364f $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_452 N_A_143_297#_c_345_n N_X_c_1398_n 0.0362443f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_453 N_A_143_297#_c_346_n N_X_c_1398_n 0.00222133f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_454 N_A_143_297#_c_332_n N_X_c_1469_n 5.22228e-19 $X=4.98 $Y=0.995 $X2=0
+ $Y2=0
cc_455 N_A_143_297#_c_333_n N_X_c_1469_n 0.00630972f $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_456 N_A_143_297#_c_334_n N_X_c_1469_n 0.00630972f $X=5.82 $Y=0.995 $X2=0
+ $Y2=0
cc_457 N_A_143_297#_c_335_n N_X_c_1469_n 5.22228e-19 $X=6.24 $Y=0.995 $X2=0
+ $Y2=0
cc_458 N_A_143_297#_c_334_n N_X_c_1399_n 0.00870364f $X=5.82 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_A_143_297#_c_335_n N_X_c_1399_n 0.00870364f $X=6.24 $Y=0.995 $X2=0
+ $Y2=0
cc_460 N_A_143_297#_c_345_n N_X_c_1399_n 0.0362443f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_461 N_A_143_297#_c_346_n N_X_c_1399_n 0.00222133f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_143_297#_c_334_n N_X_c_1477_n 5.22228e-19 $X=5.82 $Y=0.995 $X2=0
+ $Y2=0
cc_463 N_A_143_297#_c_335_n N_X_c_1477_n 0.00630972f $X=6.24 $Y=0.995 $X2=0
+ $Y2=0
cc_464 N_A_143_297#_c_336_n N_X_c_1477_n 0.00630972f $X=6.66 $Y=0.995 $X2=0
+ $Y2=0
cc_465 N_A_143_297#_c_337_n N_X_c_1477_n 5.22228e-19 $X=7.08 $Y=0.995 $X2=0
+ $Y2=0
cc_466 N_A_143_297#_c_336_n N_X_c_1400_n 0.00870364f $X=6.66 $Y=0.995 $X2=0
+ $Y2=0
cc_467 N_A_143_297#_c_337_n N_X_c_1400_n 0.00870364f $X=7.08 $Y=0.995 $X2=0
+ $Y2=0
cc_468 N_A_143_297#_c_345_n N_X_c_1400_n 0.0362443f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_143_297#_c_346_n N_X_c_1400_n 0.00222133f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_470 N_A_143_297#_c_336_n N_X_c_1485_n 5.22228e-19 $X=6.66 $Y=0.995 $X2=0
+ $Y2=0
cc_471 N_A_143_297#_c_337_n N_X_c_1485_n 0.00630972f $X=7.08 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_143_297#_c_338_n N_X_c_1485_n 0.00630972f $X=7.5 $Y=0.995 $X2=0 $Y2=0
cc_473 N_A_143_297#_c_339_n N_X_c_1485_n 5.22228e-19 $X=7.92 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_143_297#_c_338_n N_X_c_1401_n 0.00870364f $X=7.5 $Y=0.995 $X2=0 $Y2=0
cc_475 N_A_143_297#_c_339_n N_X_c_1401_n 0.00870364f $X=7.92 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_A_143_297#_c_345_n N_X_c_1401_n 0.0362443f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_477 N_A_143_297#_c_346_n N_X_c_1401_n 0.00222133f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_478 N_A_143_297#_c_338_n N_X_c_1493_n 5.22228e-19 $X=7.5 $Y=0.995 $X2=0 $Y2=0
cc_479 N_A_143_297#_c_339_n N_X_c_1493_n 0.00630972f $X=7.92 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_A_143_297#_c_340_n N_X_c_1493_n 0.00630972f $X=8.34 $Y=0.995 $X2=0
+ $Y2=0
cc_481 N_A_143_297#_c_341_n N_X_c_1493_n 5.22228e-19 $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_482 N_A_143_297#_c_340_n N_X_c_1402_n 0.00870364f $X=8.34 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_143_297#_c_341_n N_X_c_1402_n 0.00870364f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_484 N_A_143_297#_c_345_n N_X_c_1402_n 0.0362443f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_485 N_A_143_297#_c_346_n N_X_c_1402_n 0.00222133f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_486 N_A_143_297#_c_340_n N_X_c_1501_n 5.22228e-19 $X=8.34 $Y=0.995 $X2=0
+ $Y2=0
cc_487 N_A_143_297#_c_341_n N_X_c_1501_n 0.00630972f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_A_143_297#_c_342_n N_X_c_1501_n 0.00630972f $X=9.18 $Y=0.995 $X2=0
+ $Y2=0
cc_489 N_A_143_297#_c_342_n N_X_c_1403_n 0.00865686f $X=9.18 $Y=0.995 $X2=0
+ $Y2=0
cc_490 N_A_143_297#_c_345_n N_X_c_1403_n 0.0101912f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_491 N_A_143_297#_c_342_n N_X_c_1506_n 5.22228e-19 $X=9.18 $Y=0.995 $X2=0
+ $Y2=0
cc_492 N_A_143_297#_c_329_n N_X_c_1411_n 0.00113286f $X=3.72 $Y=0.995 $X2=0
+ $Y2=0
cc_493 N_A_143_297#_c_330_n N_X_c_1411_n 0.00113286f $X=4.14 $Y=0.995 $X2=0
+ $Y2=0
cc_494 N_A_143_297#_c_345_n N_X_c_1411_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_495 N_A_143_297#_c_346_n N_X_c_1411_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_496 N_A_143_297#_c_331_n N_X_c_1412_n 0.00113286f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_497 N_A_143_297#_c_332_n N_X_c_1412_n 0.00113286f $X=4.98 $Y=0.995 $X2=0
+ $Y2=0
cc_498 N_A_143_297#_c_345_n N_X_c_1412_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_499 N_A_143_297#_c_346_n N_X_c_1412_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_500 N_A_143_297#_c_333_n N_X_c_1413_n 0.00113286f $X=5.4 $Y=0.995 $X2=0 $Y2=0
cc_501 N_A_143_297#_c_334_n N_X_c_1413_n 0.00113286f $X=5.82 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_A_143_297#_c_345_n N_X_c_1413_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_503 N_A_143_297#_c_346_n N_X_c_1413_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_504 N_A_143_297#_c_335_n N_X_c_1414_n 0.00113286f $X=6.24 $Y=0.995 $X2=0
+ $Y2=0
cc_505 N_A_143_297#_c_336_n N_X_c_1414_n 0.00113286f $X=6.66 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_143_297#_c_345_n N_X_c_1414_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_507 N_A_143_297#_c_346_n N_X_c_1414_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_508 N_A_143_297#_c_337_n N_X_c_1415_n 0.00113286f $X=7.08 $Y=0.995 $X2=0
+ $Y2=0
cc_509 N_A_143_297#_c_338_n N_X_c_1415_n 0.00113286f $X=7.5 $Y=0.995 $X2=0 $Y2=0
cc_510 N_A_143_297#_c_345_n N_X_c_1415_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_511 N_A_143_297#_c_346_n N_X_c_1415_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_512 N_A_143_297#_c_339_n N_X_c_1416_n 0.00113286f $X=7.92 $Y=0.995 $X2=0
+ $Y2=0
cc_513 N_A_143_297#_c_340_n N_X_c_1416_n 0.00113286f $X=8.34 $Y=0.995 $X2=0
+ $Y2=0
cc_514 N_A_143_297#_c_345_n N_X_c_1416_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_515 N_A_143_297#_c_346_n N_X_c_1416_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_516 N_A_143_297#_c_341_n N_X_c_1417_n 0.00113286f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_517 N_A_143_297#_c_342_n N_X_c_1417_n 0.00113286f $X=9.18 $Y=0.995 $X2=0
+ $Y2=0
cc_518 N_A_143_297#_c_345_n N_X_c_1417_n 0.0266272f $X=9.09 $Y=1.16 $X2=0 $Y2=0
cc_519 N_A_143_297#_c_346_n N_X_c_1417_n 0.00230339f $X=9.18 $Y=1.16 $X2=0 $Y2=0
cc_520 N_A_143_297#_c_384_n N_VGND_c_1862_n 0.00207986f $X=0.85 $Y=1.62 $X2=0
+ $Y2=0
cc_521 N_A_143_297#_c_343_n N_VGND_c_1863_n 7.08675e-19 $X=1.07 $Y=0.42 $X2=0
+ $Y2=0
cc_522 N_A_143_297#_c_373_n N_VGND_c_1863_n 0.0130132f $X=1.525 $Y=1.175 $X2=0
+ $Y2=0
cc_523 N_A_143_297#_c_344_n N_VGND_c_1863_n 7.18045e-19 $X=1.91 $Y=0.42 $X2=0
+ $Y2=0
cc_524 N_A_143_297#_c_392_n N_VGND_c_1863_n 0.00793623f $X=1.78 $Y=1.175 $X2=0
+ $Y2=0
cc_525 N_A_143_297#_c_327_n N_VGND_c_1864_n 0.00229632f $X=2.88 $Y=0.995 $X2=0
+ $Y2=0
cc_526 N_A_143_297#_c_344_n N_VGND_c_1864_n 0.00161183f $X=1.91 $Y=0.42 $X2=0
+ $Y2=0
cc_527 N_A_143_297#_c_345_n N_VGND_c_1864_n 0.0469604f $X=9.09 $Y=1.16 $X2=0
+ $Y2=0
cc_528 N_A_143_297#_c_327_n N_VGND_c_1865_n 0.00541359f $X=2.88 $Y=0.995 $X2=0
+ $Y2=0
cc_529 N_A_143_297#_c_328_n N_VGND_c_1865_n 0.00423334f $X=3.3 $Y=0.995 $X2=0
+ $Y2=0
cc_530 N_A_143_297#_c_328_n N_VGND_c_1866_n 0.00146448f $X=3.3 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_143_297#_c_329_n N_VGND_c_1866_n 0.00146448f $X=3.72 $Y=0.995 $X2=0
+ $Y2=0
cc_532 N_A_143_297#_c_330_n N_VGND_c_1867_n 0.00146448f $X=4.14 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_A_143_297#_c_331_n N_VGND_c_1867_n 0.00146448f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_534 N_A_143_297#_c_332_n N_VGND_c_1868_n 0.00146448f $X=4.98 $Y=0.995 $X2=0
+ $Y2=0
cc_535 N_A_143_297#_c_333_n N_VGND_c_1868_n 0.00146448f $X=5.4 $Y=0.995 $X2=0
+ $Y2=0
cc_536 N_A_143_297#_c_334_n N_VGND_c_1869_n 0.00146448f $X=5.82 $Y=0.995 $X2=0
+ $Y2=0
cc_537 N_A_143_297#_c_335_n N_VGND_c_1869_n 0.00146448f $X=6.24 $Y=0.995 $X2=0
+ $Y2=0
cc_538 N_A_143_297#_c_336_n N_VGND_c_1870_n 0.00146448f $X=6.66 $Y=0.995 $X2=0
+ $Y2=0
cc_539 N_A_143_297#_c_337_n N_VGND_c_1870_n 0.00146448f $X=7.08 $Y=0.995 $X2=0
+ $Y2=0
cc_540 N_A_143_297#_c_338_n N_VGND_c_1871_n 0.00146448f $X=7.5 $Y=0.995 $X2=0
+ $Y2=0
cc_541 N_A_143_297#_c_339_n N_VGND_c_1871_n 0.00146448f $X=7.92 $Y=0.995 $X2=0
+ $Y2=0
cc_542 N_A_143_297#_c_339_n N_VGND_c_1872_n 0.00423334f $X=7.92 $Y=0.995 $X2=0
+ $Y2=0
cc_543 N_A_143_297#_c_340_n N_VGND_c_1872_n 0.00423334f $X=8.34 $Y=0.995 $X2=0
+ $Y2=0
cc_544 N_A_143_297#_c_340_n N_VGND_c_1873_n 0.00146448f $X=8.34 $Y=0.995 $X2=0
+ $Y2=0
cc_545 N_A_143_297#_c_341_n N_VGND_c_1873_n 0.00146448f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_546 N_A_143_297#_c_342_n N_VGND_c_1874_n 0.00146448f $X=9.18 $Y=0.995 $X2=0
+ $Y2=0
cc_547 N_A_143_297#_c_343_n N_VGND_c_1885_n 0.012815f $X=1.07 $Y=0.42 $X2=0
+ $Y2=0
cc_548 N_A_143_297#_c_329_n N_VGND_c_1887_n 0.00423334f $X=3.72 $Y=0.995 $X2=0
+ $Y2=0
cc_549 N_A_143_297#_c_330_n N_VGND_c_1887_n 0.00423334f $X=4.14 $Y=0.995 $X2=0
+ $Y2=0
cc_550 N_A_143_297#_c_331_n N_VGND_c_1889_n 0.00423334f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_551 N_A_143_297#_c_332_n N_VGND_c_1889_n 0.00423334f $X=4.98 $Y=0.995 $X2=0
+ $Y2=0
cc_552 N_A_143_297#_c_333_n N_VGND_c_1891_n 0.00423334f $X=5.4 $Y=0.995 $X2=0
+ $Y2=0
cc_553 N_A_143_297#_c_334_n N_VGND_c_1891_n 0.00423334f $X=5.82 $Y=0.995 $X2=0
+ $Y2=0
cc_554 N_A_143_297#_c_335_n N_VGND_c_1893_n 0.00423334f $X=6.24 $Y=0.995 $X2=0
+ $Y2=0
cc_555 N_A_143_297#_c_336_n N_VGND_c_1893_n 0.00423334f $X=6.66 $Y=0.995 $X2=0
+ $Y2=0
cc_556 N_A_143_297#_c_337_n N_VGND_c_1895_n 0.00423334f $X=7.08 $Y=0.995 $X2=0
+ $Y2=0
cc_557 N_A_143_297#_c_338_n N_VGND_c_1895_n 0.00423334f $X=7.5 $Y=0.995 $X2=0
+ $Y2=0
cc_558 N_A_143_297#_c_341_n N_VGND_c_1897_n 0.00423334f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_559 N_A_143_297#_c_342_n N_VGND_c_1897_n 0.00423334f $X=9.18 $Y=0.995 $X2=0
+ $Y2=0
cc_560 N_A_143_297#_c_344_n N_VGND_c_1912_n 0.0142343f $X=1.91 $Y=0.42 $X2=0
+ $Y2=0
cc_561 N_A_143_297#_M1038_s N_VGND_c_1919_n 0.00423495f $X=0.935 $Y=0.235 $X2=0
+ $Y2=0
cc_562 N_A_143_297#_M1049_s N_VGND_c_1919_n 0.00284632f $X=1.775 $Y=0.235 $X2=0
+ $Y2=0
cc_563 N_A_143_297#_c_327_n N_VGND_c_1919_n 0.0101559f $X=2.88 $Y=0.995 $X2=0
+ $Y2=0
cc_564 N_A_143_297#_c_328_n N_VGND_c_1919_n 0.0057163f $X=3.3 $Y=0.995 $X2=0
+ $Y2=0
cc_565 N_A_143_297#_c_329_n N_VGND_c_1919_n 0.0057163f $X=3.72 $Y=0.995 $X2=0
+ $Y2=0
cc_566 N_A_143_297#_c_330_n N_VGND_c_1919_n 0.0057163f $X=4.14 $Y=0.995 $X2=0
+ $Y2=0
cc_567 N_A_143_297#_c_331_n N_VGND_c_1919_n 0.0057163f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_568 N_A_143_297#_c_332_n N_VGND_c_1919_n 0.0057163f $X=4.98 $Y=0.995 $X2=0
+ $Y2=0
cc_569 N_A_143_297#_c_333_n N_VGND_c_1919_n 0.0057163f $X=5.4 $Y=0.995 $X2=0
+ $Y2=0
cc_570 N_A_143_297#_c_334_n N_VGND_c_1919_n 0.0057163f $X=5.82 $Y=0.995 $X2=0
+ $Y2=0
cc_571 N_A_143_297#_c_335_n N_VGND_c_1919_n 0.0057163f $X=6.24 $Y=0.995 $X2=0
+ $Y2=0
cc_572 N_A_143_297#_c_336_n N_VGND_c_1919_n 0.0057163f $X=6.66 $Y=0.995 $X2=0
+ $Y2=0
cc_573 N_A_143_297#_c_337_n N_VGND_c_1919_n 0.0057163f $X=7.08 $Y=0.995 $X2=0
+ $Y2=0
cc_574 N_A_143_297#_c_338_n N_VGND_c_1919_n 0.0057163f $X=7.5 $Y=0.995 $X2=0
+ $Y2=0
cc_575 N_A_143_297#_c_339_n N_VGND_c_1919_n 0.0057163f $X=7.92 $Y=0.995 $X2=0
+ $Y2=0
cc_576 N_A_143_297#_c_340_n N_VGND_c_1919_n 0.0057163f $X=8.34 $Y=0.995 $X2=0
+ $Y2=0
cc_577 N_A_143_297#_c_341_n N_VGND_c_1919_n 0.0057163f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_578 N_A_143_297#_c_342_n N_VGND_c_1919_n 0.0057435f $X=9.18 $Y=0.995 $X2=0
+ $Y2=0
cc_579 N_A_143_297#_c_343_n N_VGND_c_1919_n 0.00801045f $X=1.07 $Y=0.42 $X2=0
+ $Y2=0
cc_580 N_A_143_297#_c_344_n N_VGND_c_1919_n 0.00955092f $X=1.91 $Y=0.42 $X2=0
+ $Y2=0
cc_581 N_SLEEP_M1006_g N_VPWR_c_973_n 0.00357877f $X=9.6 $Y=1.985 $X2=0 $Y2=0
cc_582 N_SLEEP_M1012_g N_VPWR_c_973_n 0.00357877f $X=10.02 $Y=1.985 $X2=0 $Y2=0
cc_583 N_SLEEP_M1013_g N_VPWR_c_973_n 0.00357877f $X=10.44 $Y=1.985 $X2=0 $Y2=0
cc_584 N_SLEEP_M1014_g N_VPWR_c_973_n 0.00357877f $X=10.86 $Y=1.985 $X2=0 $Y2=0
cc_585 N_SLEEP_M1017_g N_VPWR_c_973_n 0.00357877f $X=11.28 $Y=1.985 $X2=0 $Y2=0
cc_586 N_SLEEP_M1024_g N_VPWR_c_973_n 0.00357877f $X=11.7 $Y=1.985 $X2=0 $Y2=0
cc_587 N_SLEEP_M1026_g N_VPWR_c_973_n 0.00357877f $X=12.12 $Y=1.985 $X2=0 $Y2=0
cc_588 N_SLEEP_M1034_g N_VPWR_c_973_n 0.00357877f $X=12.54 $Y=1.985 $X2=0 $Y2=0
cc_589 N_SLEEP_M1037_g N_VPWR_c_973_n 0.00357877f $X=12.96 $Y=1.985 $X2=0 $Y2=0
cc_590 N_SLEEP_M1040_g N_VPWR_c_973_n 0.00357877f $X=13.38 $Y=1.985 $X2=0 $Y2=0
cc_591 N_SLEEP_M1050_g N_VPWR_c_973_n 0.00357877f $X=13.8 $Y=1.985 $X2=0 $Y2=0
cc_592 N_SLEEP_M1054_g N_VPWR_c_973_n 0.00357877f $X=14.22 $Y=1.985 $X2=0 $Y2=0
cc_593 N_SLEEP_M1061_g N_VPWR_c_973_n 0.00357877f $X=14.64 $Y=1.985 $X2=0 $Y2=0
cc_594 N_SLEEP_M1069_g N_VPWR_c_973_n 0.00357877f $X=15.06 $Y=1.985 $X2=0 $Y2=0
cc_595 N_SLEEP_M1070_g N_VPWR_c_973_n 0.00357877f $X=15.48 $Y=1.985 $X2=0 $Y2=0
cc_596 N_SLEEP_M1071_g N_VPWR_c_973_n 0.00357877f $X=15.9 $Y=1.985 $X2=0 $Y2=0
cc_597 N_SLEEP_M1006_g N_VPWR_c_944_n 0.00525237f $X=9.6 $Y=1.985 $X2=0 $Y2=0
cc_598 N_SLEEP_M1012_g N_VPWR_c_944_n 0.00522516f $X=10.02 $Y=1.985 $X2=0 $Y2=0
cc_599 N_SLEEP_M1013_g N_VPWR_c_944_n 0.00522516f $X=10.44 $Y=1.985 $X2=0 $Y2=0
cc_600 N_SLEEP_M1014_g N_VPWR_c_944_n 0.00522516f $X=10.86 $Y=1.985 $X2=0 $Y2=0
cc_601 N_SLEEP_M1017_g N_VPWR_c_944_n 0.00522516f $X=11.28 $Y=1.985 $X2=0 $Y2=0
cc_602 N_SLEEP_M1024_g N_VPWR_c_944_n 0.00522516f $X=11.7 $Y=1.985 $X2=0 $Y2=0
cc_603 N_SLEEP_M1026_g N_VPWR_c_944_n 0.00522516f $X=12.12 $Y=1.985 $X2=0 $Y2=0
cc_604 N_SLEEP_M1034_g N_VPWR_c_944_n 0.00522516f $X=12.54 $Y=1.985 $X2=0 $Y2=0
cc_605 N_SLEEP_M1037_g N_VPWR_c_944_n 0.00522516f $X=12.96 $Y=1.985 $X2=0 $Y2=0
cc_606 N_SLEEP_M1040_g N_VPWR_c_944_n 0.00522516f $X=13.38 $Y=1.985 $X2=0 $Y2=0
cc_607 N_SLEEP_M1050_g N_VPWR_c_944_n 0.00522516f $X=13.8 $Y=1.985 $X2=0 $Y2=0
cc_608 N_SLEEP_M1054_g N_VPWR_c_944_n 0.00522516f $X=14.22 $Y=1.985 $X2=0 $Y2=0
cc_609 N_SLEEP_M1061_g N_VPWR_c_944_n 0.00522516f $X=14.64 $Y=1.985 $X2=0 $Y2=0
cc_610 N_SLEEP_M1069_g N_VPWR_c_944_n 0.00522516f $X=15.06 $Y=1.985 $X2=0 $Y2=0
cc_611 N_SLEEP_M1070_g N_VPWR_c_944_n 0.00522516f $X=15.48 $Y=1.985 $X2=0 $Y2=0
cc_612 N_SLEEP_M1071_g N_VPWR_c_944_n 0.00631837f $X=15.9 $Y=1.985 $X2=0 $Y2=0
cc_613 N_SLEEP_M1006_g N_A_505_297#_c_1190_n 2.57315e-19 $X=9.6 $Y=1.985 $X2=0
+ $Y2=0
cc_614 N_SLEEP_c_679_n N_A_505_297#_c_1190_n 0.0055111f $X=9.69 $Y=1.16 $X2=0
+ $Y2=0
cc_615 N_SLEEP_M1006_g N_A_505_297#_c_1248_n 0.0121747f $X=9.6 $Y=1.985 $X2=0
+ $Y2=0
cc_616 N_SLEEP_M1012_g N_A_505_297#_c_1248_n 0.00984328f $X=10.02 $Y=1.985 $X2=0
+ $Y2=0
cc_617 N_SLEEP_M1013_g N_A_505_297#_c_1250_n 0.00988743f $X=10.44 $Y=1.985 $X2=0
+ $Y2=0
cc_618 N_SLEEP_M1014_g N_A_505_297#_c_1250_n 0.00988743f $X=10.86 $Y=1.985 $X2=0
+ $Y2=0
cc_619 N_SLEEP_M1017_g N_A_505_297#_c_1252_n 0.00988743f $X=11.28 $Y=1.985 $X2=0
+ $Y2=0
cc_620 N_SLEEP_M1024_g N_A_505_297#_c_1252_n 0.00988743f $X=11.7 $Y=1.985 $X2=0
+ $Y2=0
cc_621 N_SLEEP_M1026_g N_A_505_297#_c_1254_n 0.00988743f $X=12.12 $Y=1.985 $X2=0
+ $Y2=0
cc_622 N_SLEEP_M1034_g N_A_505_297#_c_1254_n 0.00988743f $X=12.54 $Y=1.985 $X2=0
+ $Y2=0
cc_623 N_SLEEP_M1037_g N_A_505_297#_c_1256_n 0.00988743f $X=12.96 $Y=1.985 $X2=0
+ $Y2=0
cc_624 N_SLEEP_M1040_g N_A_505_297#_c_1256_n 0.00988743f $X=13.38 $Y=1.985 $X2=0
+ $Y2=0
cc_625 N_SLEEP_M1050_g N_A_505_297#_c_1258_n 0.00988743f $X=13.8 $Y=1.985 $X2=0
+ $Y2=0
cc_626 N_SLEEP_M1054_g N_A_505_297#_c_1258_n 0.00988743f $X=14.22 $Y=1.985 $X2=0
+ $Y2=0
cc_627 N_SLEEP_M1061_g N_A_505_297#_c_1260_n 0.00988743f $X=14.64 $Y=1.985 $X2=0
+ $Y2=0
cc_628 N_SLEEP_M1069_g N_A_505_297#_c_1260_n 0.00988743f $X=15.06 $Y=1.985 $X2=0
+ $Y2=0
cc_629 N_SLEEP_M1070_g N_A_505_297#_c_1262_n 0.00984328f $X=15.48 $Y=1.985 $X2=0
+ $Y2=0
cc_630 N_SLEEP_M1071_g N_A_505_297#_c_1262_n 0.00988421f $X=15.9 $Y=1.985 $X2=0
+ $Y2=0
cc_631 N_SLEEP_c_663_n N_X_c_1501_n 5.22228e-19 $X=9.6 $Y=0.995 $X2=0 $Y2=0
cc_632 N_SLEEP_c_663_n N_X_c_1403_n 0.00865195f $X=9.6 $Y=0.995 $X2=0 $Y2=0
cc_633 N_SLEEP_c_679_n N_X_c_1403_n 0.0140306f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_634 N_SLEEP_c_663_n N_X_c_1506_n 0.00630972f $X=9.6 $Y=0.995 $X2=0 $Y2=0
cc_635 N_SLEEP_c_664_n N_X_c_1506_n 0.00630972f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_636 N_SLEEP_c_665_n N_X_c_1506_n 5.22228e-19 $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_637 N_SLEEP_M1012_g N_X_c_1427_n 0.0109196f $X=10.02 $Y=1.985 $X2=0 $Y2=0
cc_638 N_SLEEP_M1013_g N_X_c_1427_n 0.0109338f $X=10.44 $Y=1.985 $X2=0 $Y2=0
cc_639 N_SLEEP_c_679_n N_X_c_1427_n 0.0418862f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_640 N_SLEEP_c_680_n N_X_c_1427_n 0.00211393f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_641 N_SLEEP_c_664_n N_X_c_1404_n 0.00869873f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_642 N_SLEEP_c_665_n N_X_c_1404_n 0.00869873f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_643 N_SLEEP_c_679_n N_X_c_1404_n 0.0364367f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_644 N_SLEEP_c_680_n N_X_c_1404_n 0.00222006f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_645 N_SLEEP_c_664_n N_X_c_1549_n 5.22228e-19 $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_646 N_SLEEP_c_665_n N_X_c_1549_n 0.00630972f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_647 N_SLEEP_c_666_n N_X_c_1549_n 0.00630972f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_648 N_SLEEP_c_667_n N_X_c_1549_n 5.22228e-19 $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_649 N_SLEEP_M1014_g N_X_c_1428_n 0.010978f $X=10.86 $Y=1.985 $X2=0 $Y2=0
cc_650 N_SLEEP_M1017_g N_X_c_1428_n 0.010978f $X=11.28 $Y=1.985 $X2=0 $Y2=0
cc_651 N_SLEEP_c_679_n N_X_c_1428_n 0.0418862f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_652 N_SLEEP_c_680_n N_X_c_1428_n 0.00211393f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_653 N_SLEEP_c_666_n N_X_c_1405_n 0.00869873f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_654 N_SLEEP_c_667_n N_X_c_1405_n 0.00869873f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_655 N_SLEEP_c_679_n N_X_c_1405_n 0.0364367f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_656 N_SLEEP_c_680_n N_X_c_1405_n 0.00222006f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_657 N_SLEEP_c_666_n N_X_c_1561_n 5.22228e-19 $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_658 N_SLEEP_c_667_n N_X_c_1561_n 0.00630972f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_659 N_SLEEP_c_668_n N_X_c_1561_n 0.00630972f $X=11.7 $Y=0.995 $X2=0 $Y2=0
cc_660 N_SLEEP_c_669_n N_X_c_1561_n 5.22228e-19 $X=12.12 $Y=0.995 $X2=0 $Y2=0
cc_661 N_SLEEP_M1024_g N_X_c_1429_n 0.010978f $X=11.7 $Y=1.985 $X2=0 $Y2=0
cc_662 N_SLEEP_M1026_g N_X_c_1429_n 0.010978f $X=12.12 $Y=1.985 $X2=0 $Y2=0
cc_663 N_SLEEP_c_679_n N_X_c_1429_n 0.0418862f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_664 N_SLEEP_c_680_n N_X_c_1429_n 0.00211393f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_665 N_SLEEP_c_668_n N_X_c_1406_n 0.00869873f $X=11.7 $Y=0.995 $X2=0 $Y2=0
cc_666 N_SLEEP_c_669_n N_X_c_1406_n 0.00869873f $X=12.12 $Y=0.995 $X2=0 $Y2=0
cc_667 N_SLEEP_c_679_n N_X_c_1406_n 0.0364367f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_668 N_SLEEP_c_680_n N_X_c_1406_n 0.00222006f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_669 N_SLEEP_c_668_n N_X_c_1573_n 5.22228e-19 $X=11.7 $Y=0.995 $X2=0 $Y2=0
cc_670 N_SLEEP_c_669_n N_X_c_1573_n 0.00630972f $X=12.12 $Y=0.995 $X2=0 $Y2=0
cc_671 N_SLEEP_c_670_n N_X_c_1573_n 0.00630972f $X=12.54 $Y=0.995 $X2=0 $Y2=0
cc_672 N_SLEEP_c_671_n N_X_c_1573_n 5.22228e-19 $X=12.96 $Y=0.995 $X2=0 $Y2=0
cc_673 N_SLEEP_M1034_g N_X_c_1430_n 0.010978f $X=12.54 $Y=1.985 $X2=0 $Y2=0
cc_674 N_SLEEP_M1037_g N_X_c_1430_n 0.010978f $X=12.96 $Y=1.985 $X2=0 $Y2=0
cc_675 N_SLEEP_c_679_n N_X_c_1430_n 0.0418862f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_676 N_SLEEP_c_680_n N_X_c_1430_n 0.00211393f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_677 N_SLEEP_c_670_n N_X_c_1407_n 0.00869873f $X=12.54 $Y=0.995 $X2=0 $Y2=0
cc_678 N_SLEEP_c_671_n N_X_c_1407_n 0.00869873f $X=12.96 $Y=0.995 $X2=0 $Y2=0
cc_679 N_SLEEP_c_679_n N_X_c_1407_n 0.0364367f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_680 N_SLEEP_c_680_n N_X_c_1407_n 0.00222006f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_681 N_SLEEP_c_670_n N_X_c_1585_n 5.22228e-19 $X=12.54 $Y=0.995 $X2=0 $Y2=0
cc_682 N_SLEEP_c_671_n N_X_c_1585_n 0.00630972f $X=12.96 $Y=0.995 $X2=0 $Y2=0
cc_683 N_SLEEP_c_672_n N_X_c_1585_n 0.00630972f $X=13.38 $Y=0.995 $X2=0 $Y2=0
cc_684 N_SLEEP_c_673_n N_X_c_1585_n 5.22228e-19 $X=13.8 $Y=0.995 $X2=0 $Y2=0
cc_685 N_SLEEP_M1040_g N_X_c_1431_n 0.010978f $X=13.38 $Y=1.985 $X2=0 $Y2=0
cc_686 N_SLEEP_M1050_g N_X_c_1431_n 0.010978f $X=13.8 $Y=1.985 $X2=0 $Y2=0
cc_687 N_SLEEP_c_679_n N_X_c_1431_n 0.0418862f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_688 N_SLEEP_c_680_n N_X_c_1431_n 0.00211393f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_689 N_SLEEP_c_672_n N_X_c_1408_n 0.00869873f $X=13.38 $Y=0.995 $X2=0 $Y2=0
cc_690 N_SLEEP_c_673_n N_X_c_1408_n 0.00869873f $X=13.8 $Y=0.995 $X2=0 $Y2=0
cc_691 N_SLEEP_c_679_n N_X_c_1408_n 0.0364367f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_692 N_SLEEP_c_680_n N_X_c_1408_n 0.00222006f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_693 N_SLEEP_c_672_n N_X_c_1597_n 5.22228e-19 $X=13.38 $Y=0.995 $X2=0 $Y2=0
cc_694 N_SLEEP_c_673_n N_X_c_1597_n 0.00630972f $X=13.8 $Y=0.995 $X2=0 $Y2=0
cc_695 N_SLEEP_c_674_n N_X_c_1597_n 0.00630972f $X=14.22 $Y=0.995 $X2=0 $Y2=0
cc_696 N_SLEEP_c_675_n N_X_c_1597_n 5.22228e-19 $X=14.64 $Y=0.995 $X2=0 $Y2=0
cc_697 N_SLEEP_M1054_g N_X_c_1432_n 0.010978f $X=14.22 $Y=1.985 $X2=0 $Y2=0
cc_698 N_SLEEP_M1061_g N_X_c_1432_n 0.010978f $X=14.64 $Y=1.985 $X2=0 $Y2=0
cc_699 N_SLEEP_c_679_n N_X_c_1432_n 0.0418862f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_700 N_SLEEP_c_680_n N_X_c_1432_n 0.00211393f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_701 N_SLEEP_c_674_n N_X_c_1409_n 0.00869873f $X=14.22 $Y=0.995 $X2=0 $Y2=0
cc_702 N_SLEEP_c_675_n N_X_c_1409_n 0.00869873f $X=14.64 $Y=0.995 $X2=0 $Y2=0
cc_703 N_SLEEP_c_679_n N_X_c_1409_n 0.0364367f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_704 N_SLEEP_c_680_n N_X_c_1409_n 0.00222006f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_705 N_SLEEP_c_674_n N_X_c_1609_n 5.22228e-19 $X=14.22 $Y=0.995 $X2=0 $Y2=0
cc_706 N_SLEEP_c_675_n N_X_c_1609_n 0.00630972f $X=14.64 $Y=0.995 $X2=0 $Y2=0
cc_707 N_SLEEP_c_676_n N_X_c_1609_n 0.00630972f $X=15.06 $Y=0.995 $X2=0 $Y2=0
cc_708 N_SLEEP_c_677_n N_X_c_1609_n 5.22228e-19 $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_709 N_SLEEP_M1069_g N_X_c_1433_n 0.010978f $X=15.06 $Y=1.985 $X2=0 $Y2=0
cc_710 N_SLEEP_M1070_g N_X_c_1433_n 0.010978f $X=15.48 $Y=1.985 $X2=0 $Y2=0
cc_711 N_SLEEP_c_679_n N_X_c_1433_n 0.0418862f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_712 N_SLEEP_c_680_n N_X_c_1433_n 0.00211393f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_713 N_SLEEP_c_676_n N_X_c_1410_n 0.00869873f $X=15.06 $Y=0.995 $X2=0 $Y2=0
cc_714 N_SLEEP_c_677_n N_X_c_1410_n 0.00869873f $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_715 N_SLEEP_c_679_n N_X_c_1410_n 0.0364367f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_716 N_SLEEP_c_680_n N_X_c_1410_n 0.00222006f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_717 N_SLEEP_c_676_n N_X_c_1621_n 5.22228e-19 $X=15.06 $Y=0.995 $X2=0 $Y2=0
cc_718 N_SLEEP_c_677_n N_X_c_1621_n 0.00630972f $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_719 N_SLEEP_c_678_n N_X_c_1621_n 0.0109314f $X=15.9 $Y=0.995 $X2=0 $Y2=0
cc_720 N_SLEEP_c_663_n N_X_c_1418_n 0.00113159f $X=9.6 $Y=0.995 $X2=0 $Y2=0
cc_721 N_SLEEP_c_664_n N_X_c_1418_n 0.00113159f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_722 N_SLEEP_c_679_n N_X_c_1418_n 0.0267643f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_723 N_SLEEP_c_680_n N_X_c_1418_n 0.00230167f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_724 N_SLEEP_M1006_g N_X_c_1434_n 2.57315e-19 $X=9.6 $Y=1.985 $X2=0 $Y2=0
cc_725 N_SLEEP_c_679_n N_X_c_1434_n 0.020533f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_726 N_SLEEP_c_680_n N_X_c_1434_n 0.00219397f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_727 N_SLEEP_c_665_n N_X_c_1419_n 0.00113159f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_728 N_SLEEP_c_666_n N_X_c_1419_n 0.00113159f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_729 N_SLEEP_c_679_n N_X_c_1419_n 0.0267643f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_730 N_SLEEP_c_680_n N_X_c_1419_n 0.00230167f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_731 N_SLEEP_c_679_n N_X_c_1435_n 0.020533f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_732 N_SLEEP_c_680_n N_X_c_1435_n 0.00219397f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_733 N_SLEEP_c_667_n N_X_c_1420_n 0.00113159f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_734 N_SLEEP_c_668_n N_X_c_1420_n 0.00113159f $X=11.7 $Y=0.995 $X2=0 $Y2=0
cc_735 N_SLEEP_c_679_n N_X_c_1420_n 0.0267643f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_736 N_SLEEP_c_680_n N_X_c_1420_n 0.00230167f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_737 N_SLEEP_c_679_n N_X_c_1436_n 0.020533f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_738 N_SLEEP_c_680_n N_X_c_1436_n 0.00219397f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_739 N_SLEEP_c_669_n N_X_c_1421_n 0.00113159f $X=12.12 $Y=0.995 $X2=0 $Y2=0
cc_740 N_SLEEP_c_670_n N_X_c_1421_n 0.00113159f $X=12.54 $Y=0.995 $X2=0 $Y2=0
cc_741 N_SLEEP_c_679_n N_X_c_1421_n 0.0267643f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_742 N_SLEEP_c_680_n N_X_c_1421_n 0.00230167f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_743 N_SLEEP_c_679_n N_X_c_1437_n 0.020533f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_744 N_SLEEP_c_680_n N_X_c_1437_n 0.00219397f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_745 N_SLEEP_c_671_n N_X_c_1422_n 0.00113159f $X=12.96 $Y=0.995 $X2=0 $Y2=0
cc_746 N_SLEEP_c_672_n N_X_c_1422_n 0.00113159f $X=13.38 $Y=0.995 $X2=0 $Y2=0
cc_747 N_SLEEP_c_679_n N_X_c_1422_n 0.0267643f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_748 N_SLEEP_c_680_n N_X_c_1422_n 0.00230167f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_749 N_SLEEP_c_679_n N_X_c_1438_n 0.020533f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_750 N_SLEEP_c_680_n N_X_c_1438_n 0.00219397f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_751 N_SLEEP_c_673_n N_X_c_1423_n 0.00113159f $X=13.8 $Y=0.995 $X2=0 $Y2=0
cc_752 N_SLEEP_c_674_n N_X_c_1423_n 0.00113159f $X=14.22 $Y=0.995 $X2=0 $Y2=0
cc_753 N_SLEEP_c_679_n N_X_c_1423_n 0.0267643f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_754 N_SLEEP_c_680_n N_X_c_1423_n 0.00230167f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_755 N_SLEEP_c_679_n N_X_c_1439_n 0.020533f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_756 N_SLEEP_c_680_n N_X_c_1439_n 0.00219397f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_757 N_SLEEP_c_675_n N_X_c_1424_n 0.00113159f $X=14.64 $Y=0.995 $X2=0 $Y2=0
cc_758 N_SLEEP_c_676_n N_X_c_1424_n 0.00113159f $X=15.06 $Y=0.995 $X2=0 $Y2=0
cc_759 N_SLEEP_c_679_n N_X_c_1424_n 0.0267643f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_760 N_SLEEP_c_680_n N_X_c_1424_n 0.00230167f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_761 N_SLEEP_c_679_n N_X_c_1440_n 0.020533f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_762 N_SLEEP_c_680_n N_X_c_1440_n 0.00219397f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_763 N_SLEEP_c_677_n N_X_c_1425_n 0.00113159f $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_764 N_SLEEP_c_678_n N_X_c_1425_n 0.00983958f $X=15.9 $Y=0.995 $X2=0 $Y2=0
cc_765 N_SLEEP_c_679_n N_X_c_1425_n 0.0100243f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_766 N_SLEEP_c_680_n N_X_c_1425_n 0.00283317f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_767 N_SLEEP_c_677_n X 9.58958e-19 $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_768 N_SLEEP_M1070_g X 0.00192061f $X=15.48 $Y=1.985 $X2=0 $Y2=0
cc_769 N_SLEEP_c_678_n X 0.00389713f $X=15.9 $Y=0.995 $X2=0 $Y2=0
cc_770 N_SLEEP_M1071_g X 0.0166118f $X=15.9 $Y=1.985 $X2=0 $Y2=0
cc_771 N_SLEEP_c_679_n X 0.0244542f $X=9.69 $Y=1.16 $X2=0 $Y2=0
cc_772 N_SLEEP_c_680_n X 0.024155f $X=15.9 $Y=1.16 $X2=0 $Y2=0
cc_773 N_SLEEP_c_663_n N_VGND_c_1874_n 0.00146448f $X=9.6 $Y=0.995 $X2=0 $Y2=0
cc_774 N_SLEEP_c_664_n N_VGND_c_1875_n 0.00146448f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_775 N_SLEEP_c_665_n N_VGND_c_1875_n 0.00146448f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_776 N_SLEEP_c_666_n N_VGND_c_1876_n 0.00146448f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_777 N_SLEEP_c_667_n N_VGND_c_1876_n 0.00146448f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_778 N_SLEEP_c_668_n N_VGND_c_1877_n 0.00146448f $X=11.7 $Y=0.995 $X2=0 $Y2=0
cc_779 N_SLEEP_c_669_n N_VGND_c_1877_n 0.00146448f $X=12.12 $Y=0.995 $X2=0 $Y2=0
cc_780 N_SLEEP_c_670_n N_VGND_c_1878_n 0.00146448f $X=12.54 $Y=0.995 $X2=0 $Y2=0
cc_781 N_SLEEP_c_671_n N_VGND_c_1878_n 0.00146448f $X=12.96 $Y=0.995 $X2=0 $Y2=0
cc_782 N_SLEEP_c_671_n N_VGND_c_1879_n 0.00423334f $X=12.96 $Y=0.995 $X2=0 $Y2=0
cc_783 N_SLEEP_c_672_n N_VGND_c_1879_n 0.00423334f $X=13.38 $Y=0.995 $X2=0 $Y2=0
cc_784 N_SLEEP_c_672_n N_VGND_c_1880_n 0.00146448f $X=13.38 $Y=0.995 $X2=0 $Y2=0
cc_785 N_SLEEP_c_673_n N_VGND_c_1880_n 0.00146448f $X=13.8 $Y=0.995 $X2=0 $Y2=0
cc_786 N_SLEEP_c_674_n N_VGND_c_1881_n 0.00146448f $X=14.22 $Y=0.995 $X2=0 $Y2=0
cc_787 N_SLEEP_c_675_n N_VGND_c_1881_n 0.00146448f $X=14.64 $Y=0.995 $X2=0 $Y2=0
cc_788 N_SLEEP_c_676_n N_VGND_c_1882_n 0.00146448f $X=15.06 $Y=0.995 $X2=0 $Y2=0
cc_789 N_SLEEP_c_677_n N_VGND_c_1882_n 0.00146448f $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_790 N_SLEEP_c_678_n N_VGND_c_1884_n 0.00322276f $X=15.9 $Y=0.995 $X2=0 $Y2=0
cc_791 N_SLEEP_c_663_n N_VGND_c_1899_n 0.00423334f $X=9.6 $Y=0.995 $X2=0 $Y2=0
cc_792 N_SLEEP_c_664_n N_VGND_c_1899_n 0.00423334f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_793 N_SLEEP_c_665_n N_VGND_c_1901_n 0.00423334f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_794 N_SLEEP_c_666_n N_VGND_c_1901_n 0.00423334f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_795 N_SLEEP_c_667_n N_VGND_c_1903_n 0.00423334f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_796 N_SLEEP_c_668_n N_VGND_c_1903_n 0.00423334f $X=11.7 $Y=0.995 $X2=0 $Y2=0
cc_797 N_SLEEP_c_669_n N_VGND_c_1905_n 0.00423334f $X=12.12 $Y=0.995 $X2=0 $Y2=0
cc_798 N_SLEEP_c_670_n N_VGND_c_1905_n 0.00423334f $X=12.54 $Y=0.995 $X2=0 $Y2=0
cc_799 N_SLEEP_c_673_n N_VGND_c_1907_n 0.00423334f $X=13.8 $Y=0.995 $X2=0 $Y2=0
cc_800 N_SLEEP_c_674_n N_VGND_c_1907_n 0.00423334f $X=14.22 $Y=0.995 $X2=0 $Y2=0
cc_801 N_SLEEP_c_675_n N_VGND_c_1909_n 0.00423334f $X=14.64 $Y=0.995 $X2=0 $Y2=0
cc_802 N_SLEEP_c_676_n N_VGND_c_1909_n 0.00423334f $X=15.06 $Y=0.995 $X2=0 $Y2=0
cc_803 N_SLEEP_c_677_n N_VGND_c_1913_n 0.00423334f $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_804 N_SLEEP_c_678_n N_VGND_c_1913_n 0.00423225f $X=15.9 $Y=0.995 $X2=0 $Y2=0
cc_805 N_SLEEP_c_663_n N_VGND_c_1919_n 0.0057435f $X=9.6 $Y=0.995 $X2=0 $Y2=0
cc_806 N_SLEEP_c_664_n N_VGND_c_1919_n 0.0057163f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_807 N_SLEEP_c_665_n N_VGND_c_1919_n 0.0057163f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_808 N_SLEEP_c_666_n N_VGND_c_1919_n 0.0057163f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_809 N_SLEEP_c_667_n N_VGND_c_1919_n 0.0057163f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_810 N_SLEEP_c_668_n N_VGND_c_1919_n 0.0057163f $X=11.7 $Y=0.995 $X2=0 $Y2=0
cc_811 N_SLEEP_c_669_n N_VGND_c_1919_n 0.0057163f $X=12.12 $Y=0.995 $X2=0 $Y2=0
cc_812 N_SLEEP_c_670_n N_VGND_c_1919_n 0.0057163f $X=12.54 $Y=0.995 $X2=0 $Y2=0
cc_813 N_SLEEP_c_671_n N_VGND_c_1919_n 0.0057163f $X=12.96 $Y=0.995 $X2=0 $Y2=0
cc_814 N_SLEEP_c_672_n N_VGND_c_1919_n 0.0057163f $X=13.38 $Y=0.995 $X2=0 $Y2=0
cc_815 N_SLEEP_c_673_n N_VGND_c_1919_n 0.0057163f $X=13.8 $Y=0.995 $X2=0 $Y2=0
cc_816 N_SLEEP_c_674_n N_VGND_c_1919_n 0.0057163f $X=14.22 $Y=0.995 $X2=0 $Y2=0
cc_817 N_SLEEP_c_675_n N_VGND_c_1919_n 0.0057163f $X=14.64 $Y=0.995 $X2=0 $Y2=0
cc_818 N_SLEEP_c_676_n N_VGND_c_1919_n 0.0057163f $X=15.06 $Y=0.995 $X2=0 $Y2=0
cc_819 N_SLEEP_c_677_n N_VGND_c_1919_n 0.0057163f $X=15.48 $Y=0.995 $X2=0 $Y2=0
cc_820 N_SLEEP_c_678_n N_VGND_c_1919_n 0.00680753f $X=15.9 $Y=0.995 $X2=0 $Y2=0
cc_821 N_VPWR_c_944_n N_A_505_297#_M1000_s 0.00260431f $X=16.33 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_822 N_VPWR_c_944_n N_A_505_297#_M1001_s 0.00284632f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_823 N_VPWR_c_944_n N_A_505_297#_M1005_s 0.00284632f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_824 N_VPWR_c_944_n N_A_505_297#_M1011_s 0.00284632f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_825 N_VPWR_c_944_n N_A_505_297#_M1020_s 0.00284632f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_826 N_VPWR_c_944_n N_A_505_297#_M1031_s 0.00284632f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_827 N_VPWR_c_944_n N_A_505_297#_M1039_s 0.00284632f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_828 N_VPWR_c_944_n N_A_505_297#_M1053_s 0.00284632f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_829 N_VPWR_c_944_n N_A_505_297#_M1060_s 0.00246446f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_830 N_VPWR_c_944_n N_A_505_297#_M1012_d 0.00215203f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_831 N_VPWR_c_944_n N_A_505_297#_M1014_d 0.00215203f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_832 N_VPWR_c_944_n N_A_505_297#_M1024_d 0.00215203f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_833 N_VPWR_c_944_n N_A_505_297#_M1034_d 0.00215203f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_834 N_VPWR_c_944_n N_A_505_297#_M1040_d 0.00215203f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_835 N_VPWR_c_944_n N_A_505_297#_M1054_d 0.00215203f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_836 N_VPWR_c_944_n N_A_505_297#_M1069_d 0.00215203f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_837 N_VPWR_c_944_n N_A_505_297#_M1071_d 0.00252233f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_838 N_VPWR_c_948_n N_A_505_297#_c_1180_n 0.0159391f $X=2.11 $Y=1.64 $X2=0
+ $Y2=0
cc_839 N_VPWR_c_948_n N_A_505_297#_c_1181_n 0.0569581f $X=2.11 $Y=1.64 $X2=0
+ $Y2=0
cc_840 N_VPWR_c_949_n N_A_505_297#_c_1181_n 0.0208267f $X=2.965 $Y=2.72 $X2=0
+ $Y2=0
cc_841 N_VPWR_c_944_n N_A_505_297#_c_1181_n 0.0122467f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_842 N_VPWR_M1000_d N_A_505_297#_c_1182_n 0.00166915f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_843 N_VPWR_c_950_n N_A_505_297#_c_1182_n 0.0128751f $X=3.09 $Y=2 $X2=0 $Y2=0
cc_844 N_VPWR_c_971_n N_A_505_297#_c_1287_n 0.0142343f $X=3.805 $Y=2.72 $X2=0
+ $Y2=0
cc_845 N_VPWR_c_944_n N_A_505_297#_c_1287_n 0.00955092f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_846 N_VPWR_M1004_d N_A_505_297#_c_1183_n 0.00166915f $X=3.795 $Y=1.485 $X2=0
+ $Y2=0
cc_847 N_VPWR_c_951_n N_A_505_297#_c_1183_n 0.0128751f $X=3.93 $Y=2 $X2=0 $Y2=0
cc_848 N_VPWR_c_963_n N_A_505_297#_c_1291_n 0.0142343f $X=4.645 $Y=2.72 $X2=0
+ $Y2=0
cc_849 N_VPWR_c_944_n N_A_505_297#_c_1291_n 0.00955092f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_850 N_VPWR_M1009_d N_A_505_297#_c_1184_n 0.00166915f $X=4.635 $Y=1.485 $X2=0
+ $Y2=0
cc_851 N_VPWR_c_952_n N_A_505_297#_c_1184_n 0.0128751f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_852 N_VPWR_c_965_n N_A_505_297#_c_1295_n 0.0142343f $X=5.485 $Y=2.72 $X2=0
+ $Y2=0
cc_853 N_VPWR_c_944_n N_A_505_297#_c_1295_n 0.00955092f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_854 N_VPWR_M1019_d N_A_505_297#_c_1185_n 0.00166915f $X=5.475 $Y=1.485 $X2=0
+ $Y2=0
cc_855 N_VPWR_c_953_n N_A_505_297#_c_1185_n 0.0128751f $X=5.61 $Y=2 $X2=0 $Y2=0
cc_856 N_VPWR_c_967_n N_A_505_297#_c_1299_n 0.0142343f $X=6.325 $Y=2.72 $X2=0
+ $Y2=0
cc_857 N_VPWR_c_944_n N_A_505_297#_c_1299_n 0.00955092f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_858 N_VPWR_M1023_d N_A_505_297#_c_1186_n 0.00166915f $X=6.315 $Y=1.485 $X2=0
+ $Y2=0
cc_859 N_VPWR_c_954_n N_A_505_297#_c_1186_n 0.0128751f $X=6.45 $Y=2 $X2=0 $Y2=0
cc_860 N_VPWR_c_969_n N_A_505_297#_c_1303_n 0.0142343f $X=7.165 $Y=2.72 $X2=0
+ $Y2=0
cc_861 N_VPWR_c_944_n N_A_505_297#_c_1303_n 0.00955092f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_862 N_VPWR_M1032_d N_A_505_297#_c_1187_n 0.00166915f $X=7.155 $Y=1.485 $X2=0
+ $Y2=0
cc_863 N_VPWR_c_955_n N_A_505_297#_c_1187_n 0.0128751f $X=7.29 $Y=2 $X2=0 $Y2=0
cc_864 N_VPWR_c_956_n N_A_505_297#_c_1307_n 0.0142343f $X=8.005 $Y=2.72 $X2=0
+ $Y2=0
cc_865 N_VPWR_c_944_n N_A_505_297#_c_1307_n 0.00955092f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_866 N_VPWR_M1048_d N_A_505_297#_c_1188_n 0.00166915f $X=7.995 $Y=1.485 $X2=0
+ $Y2=0
cc_867 N_VPWR_c_957_n N_A_505_297#_c_1188_n 0.0128751f $X=8.13 $Y=2 $X2=0 $Y2=0
cc_868 N_VPWR_c_972_n N_A_505_297#_c_1311_n 0.0142343f $X=8.845 $Y=2.72 $X2=0
+ $Y2=0
cc_869 N_VPWR_c_944_n N_A_505_297#_c_1311_n 0.00955092f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_870 N_VPWR_M1057_d N_A_505_297#_c_1189_n 0.00166915f $X=8.835 $Y=1.485 $X2=0
+ $Y2=0
cc_871 N_VPWR_c_958_n N_A_505_297#_c_1189_n 0.0128751f $X=8.97 $Y=2 $X2=0 $Y2=0
cc_872 N_VPWR_c_973_n N_A_505_297#_c_1315_n 0.0143053f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_873 N_VPWR_c_944_n N_A_505_297#_c_1315_n 0.00962794f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_874 N_VPWR_c_973_n N_A_505_297#_c_1248_n 0.0330174f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_875 N_VPWR_c_944_n N_A_505_297#_c_1248_n 0.0204627f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_876 N_VPWR_c_973_n N_A_505_297#_c_1250_n 0.0330174f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_877 N_VPWR_c_944_n N_A_505_297#_c_1250_n 0.0204627f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_878 N_VPWR_c_973_n N_A_505_297#_c_1252_n 0.0330174f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_879 N_VPWR_c_944_n N_A_505_297#_c_1252_n 0.0204627f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_880 N_VPWR_c_973_n N_A_505_297#_c_1254_n 0.0330174f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_881 N_VPWR_c_944_n N_A_505_297#_c_1254_n 0.0204627f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_882 N_VPWR_c_973_n N_A_505_297#_c_1256_n 0.0330174f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_883 N_VPWR_c_944_n N_A_505_297#_c_1256_n 0.0204627f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_884 N_VPWR_c_973_n N_A_505_297#_c_1258_n 0.0330174f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_885 N_VPWR_c_944_n N_A_505_297#_c_1258_n 0.0204627f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_886 N_VPWR_c_973_n N_A_505_297#_c_1260_n 0.0330174f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_887 N_VPWR_c_944_n N_A_505_297#_c_1260_n 0.0204627f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_973_n N_A_505_297#_c_1262_n 0.0489446f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_944_n N_A_505_297#_c_1262_n 0.0300869f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_973_n N_A_505_297#_c_1333_n 0.0142933f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_944_n N_A_505_297#_c_1333_n 0.00962421f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_973_n N_A_505_297#_c_1335_n 0.0142933f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_944_n N_A_505_297#_c_1335_n 0.00962421f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_973_n N_A_505_297#_c_1337_n 0.0142933f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_944_n N_A_505_297#_c_1337_n 0.00962421f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_973_n N_A_505_297#_c_1339_n 0.0142933f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_944_n N_A_505_297#_c_1339_n 0.00962421f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_973_n N_A_505_297#_c_1341_n 0.0142933f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_944_n N_A_505_297#_c_1341_n 0.00962421f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_973_n N_A_505_297#_c_1343_n 0.0142933f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_944_n N_A_505_297#_c_1343_n 0.00962421f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_973_n N_A_505_297#_c_1345_n 0.0142933f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_903 N_VPWR_c_944_n N_A_505_297#_c_1345_n 0.00962421f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_944_n N_X_M1006_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_905 N_VPWR_c_944_n N_X_M1013_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_906 N_VPWR_c_944_n N_X_M1017_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_907 N_VPWR_c_944_n N_X_M1026_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_908 N_VPWR_c_944_n N_X_M1037_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_909 N_VPWR_c_944_n N_X_M1050_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_910 N_VPWR_c_944_n N_X_M1061_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_911 N_VPWR_c_944_n N_X_M1070_s 0.00216833f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_912 N_A_505_297#_c_1248_n N_X_M1006_s 0.00312348f $X=10.105 $Y=2.38 $X2=0
+ $Y2=0
cc_913 N_A_505_297#_c_1250_n N_X_M1013_s 0.00312348f $X=10.945 $Y=2.38 $X2=0
+ $Y2=0
cc_914 N_A_505_297#_c_1252_n N_X_M1017_s 0.00312348f $X=11.785 $Y=2.38 $X2=0
+ $Y2=0
cc_915 N_A_505_297#_c_1254_n N_X_M1026_s 0.00312348f $X=12.625 $Y=2.38 $X2=0
+ $Y2=0
cc_916 N_A_505_297#_c_1256_n N_X_M1037_s 0.00312348f $X=13.465 $Y=2.38 $X2=0
+ $Y2=0
cc_917 N_A_505_297#_c_1258_n N_X_M1050_s 0.00312348f $X=14.305 $Y=2.38 $X2=0
+ $Y2=0
cc_918 N_A_505_297#_c_1260_n N_X_M1061_s 0.00312348f $X=15.145 $Y=2.38 $X2=0
+ $Y2=0
cc_919 N_A_505_297#_c_1262_n N_X_M1070_s 0.00312348f $X=15.985 $Y=2.38 $X2=0
+ $Y2=0
cc_920 N_A_505_297#_c_1190_n N_X_c_1403_n 0.00640581f $X=9.39 $Y=1.665 $X2=0
+ $Y2=0
cc_921 N_A_505_297#_M1012_d N_X_c_1427_n 0.00165831f $X=10.095 $Y=1.485 $X2=0
+ $Y2=0
cc_922 N_A_505_297#_c_1248_n N_X_c_1427_n 0.00320918f $X=10.105 $Y=2.38 $X2=0
+ $Y2=0
cc_923 N_A_505_297#_c_1358_p N_X_c_1427_n 0.0126766f $X=10.23 $Y=1.96 $X2=0
+ $Y2=0
cc_924 N_A_505_297#_c_1250_n N_X_c_1427_n 0.00320918f $X=10.945 $Y=2.38 $X2=0
+ $Y2=0
cc_925 N_A_505_297#_M1014_d N_X_c_1428_n 0.00165831f $X=10.935 $Y=1.485 $X2=0
+ $Y2=0
cc_926 N_A_505_297#_c_1250_n N_X_c_1428_n 0.00320918f $X=10.945 $Y=2.38 $X2=0
+ $Y2=0
cc_927 N_A_505_297#_c_1362_p N_X_c_1428_n 0.0126766f $X=11.07 $Y=1.96 $X2=0
+ $Y2=0
cc_928 N_A_505_297#_c_1252_n N_X_c_1428_n 0.00320918f $X=11.785 $Y=2.38 $X2=0
+ $Y2=0
cc_929 N_A_505_297#_M1024_d N_X_c_1429_n 0.00165831f $X=11.775 $Y=1.485 $X2=0
+ $Y2=0
cc_930 N_A_505_297#_c_1252_n N_X_c_1429_n 0.00320918f $X=11.785 $Y=2.38 $X2=0
+ $Y2=0
cc_931 N_A_505_297#_c_1366_p N_X_c_1429_n 0.0126766f $X=11.91 $Y=1.96 $X2=0
+ $Y2=0
cc_932 N_A_505_297#_c_1254_n N_X_c_1429_n 0.00320918f $X=12.625 $Y=2.38 $X2=0
+ $Y2=0
cc_933 N_A_505_297#_M1034_d N_X_c_1430_n 0.00165831f $X=12.615 $Y=1.485 $X2=0
+ $Y2=0
cc_934 N_A_505_297#_c_1254_n N_X_c_1430_n 0.00320918f $X=12.625 $Y=2.38 $X2=0
+ $Y2=0
cc_935 N_A_505_297#_c_1370_p N_X_c_1430_n 0.0126766f $X=12.75 $Y=1.96 $X2=0
+ $Y2=0
cc_936 N_A_505_297#_c_1256_n N_X_c_1430_n 0.00320918f $X=13.465 $Y=2.38 $X2=0
+ $Y2=0
cc_937 N_A_505_297#_M1040_d N_X_c_1431_n 0.00165831f $X=13.455 $Y=1.485 $X2=0
+ $Y2=0
cc_938 N_A_505_297#_c_1256_n N_X_c_1431_n 0.00320918f $X=13.465 $Y=2.38 $X2=0
+ $Y2=0
cc_939 N_A_505_297#_c_1374_p N_X_c_1431_n 0.0126766f $X=13.59 $Y=1.96 $X2=0
+ $Y2=0
cc_940 N_A_505_297#_c_1258_n N_X_c_1431_n 0.00320918f $X=14.305 $Y=2.38 $X2=0
+ $Y2=0
cc_941 N_A_505_297#_M1054_d N_X_c_1432_n 0.00165831f $X=14.295 $Y=1.485 $X2=0
+ $Y2=0
cc_942 N_A_505_297#_c_1258_n N_X_c_1432_n 0.00320918f $X=14.305 $Y=2.38 $X2=0
+ $Y2=0
cc_943 N_A_505_297#_c_1378_p N_X_c_1432_n 0.0126766f $X=14.43 $Y=1.96 $X2=0
+ $Y2=0
cc_944 N_A_505_297#_c_1260_n N_X_c_1432_n 0.00320918f $X=15.145 $Y=2.38 $X2=0
+ $Y2=0
cc_945 N_A_505_297#_M1069_d N_X_c_1433_n 0.00165831f $X=15.135 $Y=1.485 $X2=0
+ $Y2=0
cc_946 N_A_505_297#_c_1260_n N_X_c_1433_n 0.00320918f $X=15.145 $Y=2.38 $X2=0
+ $Y2=0
cc_947 N_A_505_297#_c_1382_p N_X_c_1433_n 0.0126766f $X=15.27 $Y=1.96 $X2=0
+ $Y2=0
cc_948 N_A_505_297#_c_1262_n N_X_c_1433_n 0.00320918f $X=15.985 $Y=2.38 $X2=0
+ $Y2=0
cc_949 N_A_505_297#_c_1190_n N_X_c_1434_n 0.00271526f $X=9.39 $Y=1.665 $X2=0
+ $Y2=0
cc_950 N_A_505_297#_c_1248_n N_X_c_1434_n 0.0118729f $X=10.105 $Y=2.38 $X2=0
+ $Y2=0
cc_951 N_A_505_297#_c_1250_n N_X_c_1435_n 0.0118729f $X=10.945 $Y=2.38 $X2=0
+ $Y2=0
cc_952 N_A_505_297#_c_1252_n N_X_c_1436_n 0.0118729f $X=11.785 $Y=2.38 $X2=0
+ $Y2=0
cc_953 N_A_505_297#_c_1254_n N_X_c_1437_n 0.0118729f $X=12.625 $Y=2.38 $X2=0
+ $Y2=0
cc_954 N_A_505_297#_c_1256_n N_X_c_1438_n 0.0118729f $X=13.465 $Y=2.38 $X2=0
+ $Y2=0
cc_955 N_A_505_297#_c_1258_n N_X_c_1439_n 0.0118729f $X=14.305 $Y=2.38 $X2=0
+ $Y2=0
cc_956 N_A_505_297#_c_1260_n N_X_c_1440_n 0.0118729f $X=15.145 $Y=2.38 $X2=0
+ $Y2=0
cc_957 N_A_505_297#_M1071_d X 0.00342901f $X=15.975 $Y=1.485 $X2=0 $Y2=0
cc_958 N_A_505_297#_c_1262_n X 0.0154676f $X=15.985 $Y=2.38 $X2=0 $Y2=0
cc_959 N_A_505_297#_c_1394_p X 0.0181927f $X=16.11 $Y=1.96 $X2=0 $Y2=0
cc_960 N_X_c_1395_n N_VGND_M1003_s 0.00162089f $X=3.765 $Y=0.815 $X2=0 $Y2=0
cc_961 N_X_c_1397_n N_VGND_M1008_s 0.00162089f $X=4.605 $Y=0.815 $X2=0 $Y2=0
cc_962 N_X_c_1398_n N_VGND_M1015_s 0.00162089f $X=5.445 $Y=0.815 $X2=0 $Y2=0
cc_963 N_X_c_1399_n N_VGND_M1021_s 0.00162089f $X=6.285 $Y=0.815 $X2=0 $Y2=0
cc_964 N_X_c_1400_n N_VGND_M1027_s 0.00162089f $X=7.125 $Y=0.815 $X2=0 $Y2=0
cc_965 N_X_c_1401_n N_VGND_M1055_s 0.00162089f $X=7.965 $Y=0.815 $X2=0 $Y2=0
cc_966 N_X_c_1402_n N_VGND_M1065_s 0.00162089f $X=8.805 $Y=0.815 $X2=0 $Y2=0
cc_967 N_X_c_1403_n N_VGND_M1068_s 0.00162089f $X=9.645 $Y=0.815 $X2=0 $Y2=0
cc_968 N_X_c_1404_n N_VGND_M1029_s 0.00162089f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_969 N_X_c_1405_n N_VGND_M1033_s 0.00162089f $X=11.325 $Y=0.815 $X2=0 $Y2=0
cc_970 N_X_c_1406_n N_VGND_M1041_s 0.00162089f $X=12.165 $Y=0.815 $X2=0 $Y2=0
cc_971 N_X_c_1407_n N_VGND_M1044_s 0.00162089f $X=13.005 $Y=0.815 $X2=0 $Y2=0
cc_972 N_X_c_1408_n N_VGND_M1046_s 0.00162089f $X=13.845 $Y=0.815 $X2=0 $Y2=0
cc_973 N_X_c_1409_n N_VGND_M1052_s 0.00162089f $X=14.685 $Y=0.815 $X2=0 $Y2=0
cc_974 N_X_c_1410_n N_VGND_M1058_s 0.00162089f $X=15.525 $Y=0.815 $X2=0 $Y2=0
cc_975 N_X_c_1425_n N_VGND_M1066_s 0.00290026f $X=16 $Y=0.815 $X2=0 $Y2=0
cc_976 N_X_c_1396_n N_VGND_c_1864_n 0.00843985f $X=3.255 $Y=0.815 $X2=0 $Y2=0
cc_977 N_X_c_1442_n N_VGND_c_1865_n 0.0188551f $X=3.09 $Y=0.39 $X2=0 $Y2=0
cc_978 N_X_c_1395_n N_VGND_c_1865_n 0.00198695f $X=3.765 $Y=0.815 $X2=0 $Y2=0
cc_979 N_X_c_1395_n N_VGND_c_1866_n 0.0122559f $X=3.765 $Y=0.815 $X2=0 $Y2=0
cc_980 N_X_c_1397_n N_VGND_c_1867_n 0.0122559f $X=4.605 $Y=0.815 $X2=0 $Y2=0
cc_981 N_X_c_1398_n N_VGND_c_1868_n 0.0122559f $X=5.445 $Y=0.815 $X2=0 $Y2=0
cc_982 N_X_c_1399_n N_VGND_c_1869_n 0.0122559f $X=6.285 $Y=0.815 $X2=0 $Y2=0
cc_983 N_X_c_1400_n N_VGND_c_1870_n 0.0122559f $X=7.125 $Y=0.815 $X2=0 $Y2=0
cc_984 N_X_c_1401_n N_VGND_c_1871_n 0.0122559f $X=7.965 $Y=0.815 $X2=0 $Y2=0
cc_985 N_X_c_1401_n N_VGND_c_1872_n 0.00198695f $X=7.965 $Y=0.815 $X2=0 $Y2=0
cc_986 N_X_c_1493_n N_VGND_c_1872_n 0.0188551f $X=8.13 $Y=0.39 $X2=0 $Y2=0
cc_987 N_X_c_1402_n N_VGND_c_1872_n 0.00198695f $X=8.805 $Y=0.815 $X2=0 $Y2=0
cc_988 N_X_c_1402_n N_VGND_c_1873_n 0.0122559f $X=8.805 $Y=0.815 $X2=0 $Y2=0
cc_989 N_X_c_1403_n N_VGND_c_1874_n 0.0122559f $X=9.645 $Y=0.815 $X2=0 $Y2=0
cc_990 N_X_c_1404_n N_VGND_c_1875_n 0.0122559f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_991 N_X_c_1405_n N_VGND_c_1876_n 0.0122559f $X=11.325 $Y=0.815 $X2=0 $Y2=0
cc_992 N_X_c_1406_n N_VGND_c_1877_n 0.0122559f $X=12.165 $Y=0.815 $X2=0 $Y2=0
cc_993 N_X_c_1407_n N_VGND_c_1878_n 0.0122559f $X=13.005 $Y=0.815 $X2=0 $Y2=0
cc_994 N_X_c_1407_n N_VGND_c_1879_n 0.00198695f $X=13.005 $Y=0.815 $X2=0 $Y2=0
cc_995 N_X_c_1585_n N_VGND_c_1879_n 0.0188551f $X=13.17 $Y=0.39 $X2=0 $Y2=0
cc_996 N_X_c_1408_n N_VGND_c_1879_n 0.00198695f $X=13.845 $Y=0.815 $X2=0 $Y2=0
cc_997 N_X_c_1408_n N_VGND_c_1880_n 0.0122559f $X=13.845 $Y=0.815 $X2=0 $Y2=0
cc_998 N_X_c_1409_n N_VGND_c_1881_n 0.0122559f $X=14.685 $Y=0.815 $X2=0 $Y2=0
cc_999 N_X_c_1410_n N_VGND_c_1882_n 0.0122559f $X=15.525 $Y=0.815 $X2=0 $Y2=0
cc_1000 N_X_c_1425_n N_VGND_c_1883_n 0.00307208f $X=16 $Y=0.815 $X2=0 $Y2=0
cc_1001 N_X_c_1425_n N_VGND_c_1884_n 0.0228574f $X=16 $Y=0.815 $X2=0 $Y2=0
cc_1002 N_X_c_1395_n N_VGND_c_1887_n 0.00198695f $X=3.765 $Y=0.815 $X2=0 $Y2=0
cc_1003 N_X_c_1453_n N_VGND_c_1887_n 0.0188551f $X=3.93 $Y=0.39 $X2=0 $Y2=0
cc_1004 N_X_c_1397_n N_VGND_c_1887_n 0.00198695f $X=4.605 $Y=0.815 $X2=0 $Y2=0
cc_1005 N_X_c_1397_n N_VGND_c_1889_n 0.00198695f $X=4.605 $Y=0.815 $X2=0 $Y2=0
cc_1006 N_X_c_1461_n N_VGND_c_1889_n 0.0188551f $X=4.77 $Y=0.39 $X2=0 $Y2=0
cc_1007 N_X_c_1398_n N_VGND_c_1889_n 0.00198695f $X=5.445 $Y=0.815 $X2=0 $Y2=0
cc_1008 N_X_c_1398_n N_VGND_c_1891_n 0.00198695f $X=5.445 $Y=0.815 $X2=0 $Y2=0
cc_1009 N_X_c_1469_n N_VGND_c_1891_n 0.0188551f $X=5.61 $Y=0.39 $X2=0 $Y2=0
cc_1010 N_X_c_1399_n N_VGND_c_1891_n 0.00198695f $X=6.285 $Y=0.815 $X2=0 $Y2=0
cc_1011 N_X_c_1399_n N_VGND_c_1893_n 0.00198695f $X=6.285 $Y=0.815 $X2=0 $Y2=0
cc_1012 N_X_c_1477_n N_VGND_c_1893_n 0.0188551f $X=6.45 $Y=0.39 $X2=0 $Y2=0
cc_1013 N_X_c_1400_n N_VGND_c_1893_n 0.00198695f $X=7.125 $Y=0.815 $X2=0 $Y2=0
cc_1014 N_X_c_1400_n N_VGND_c_1895_n 0.00198695f $X=7.125 $Y=0.815 $X2=0 $Y2=0
cc_1015 N_X_c_1485_n N_VGND_c_1895_n 0.0188551f $X=7.29 $Y=0.39 $X2=0 $Y2=0
cc_1016 N_X_c_1401_n N_VGND_c_1895_n 0.00198695f $X=7.965 $Y=0.815 $X2=0 $Y2=0
cc_1017 N_X_c_1402_n N_VGND_c_1897_n 0.00198695f $X=8.805 $Y=0.815 $X2=0 $Y2=0
cc_1018 N_X_c_1501_n N_VGND_c_1897_n 0.0188551f $X=8.97 $Y=0.39 $X2=0 $Y2=0
cc_1019 N_X_c_1403_n N_VGND_c_1897_n 0.00198695f $X=9.645 $Y=0.815 $X2=0 $Y2=0
cc_1020 N_X_c_1403_n N_VGND_c_1899_n 0.00198695f $X=9.645 $Y=0.815 $X2=0 $Y2=0
cc_1021 N_X_c_1506_n N_VGND_c_1899_n 0.0188551f $X=9.81 $Y=0.39 $X2=0 $Y2=0
cc_1022 N_X_c_1404_n N_VGND_c_1899_n 0.00198695f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_1023 N_X_c_1404_n N_VGND_c_1901_n 0.00198695f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_1024 N_X_c_1549_n N_VGND_c_1901_n 0.0188551f $X=10.65 $Y=0.39 $X2=0 $Y2=0
cc_1025 N_X_c_1405_n N_VGND_c_1901_n 0.00198695f $X=11.325 $Y=0.815 $X2=0 $Y2=0
cc_1026 N_X_c_1405_n N_VGND_c_1903_n 0.00198695f $X=11.325 $Y=0.815 $X2=0 $Y2=0
cc_1027 N_X_c_1561_n N_VGND_c_1903_n 0.0188551f $X=11.49 $Y=0.39 $X2=0 $Y2=0
cc_1028 N_X_c_1406_n N_VGND_c_1903_n 0.00198695f $X=12.165 $Y=0.815 $X2=0 $Y2=0
cc_1029 N_X_c_1406_n N_VGND_c_1905_n 0.00198695f $X=12.165 $Y=0.815 $X2=0 $Y2=0
cc_1030 N_X_c_1573_n N_VGND_c_1905_n 0.0188551f $X=12.33 $Y=0.39 $X2=0 $Y2=0
cc_1031 N_X_c_1407_n N_VGND_c_1905_n 0.00198695f $X=13.005 $Y=0.815 $X2=0 $Y2=0
cc_1032 N_X_c_1408_n N_VGND_c_1907_n 0.00198695f $X=13.845 $Y=0.815 $X2=0 $Y2=0
cc_1033 N_X_c_1597_n N_VGND_c_1907_n 0.0188551f $X=14.01 $Y=0.39 $X2=0 $Y2=0
cc_1034 N_X_c_1409_n N_VGND_c_1907_n 0.00198695f $X=14.685 $Y=0.815 $X2=0 $Y2=0
cc_1035 N_X_c_1409_n N_VGND_c_1909_n 0.00198695f $X=14.685 $Y=0.815 $X2=0 $Y2=0
cc_1036 N_X_c_1609_n N_VGND_c_1909_n 0.0188551f $X=14.85 $Y=0.39 $X2=0 $Y2=0
cc_1037 N_X_c_1410_n N_VGND_c_1909_n 0.00198695f $X=15.525 $Y=0.815 $X2=0 $Y2=0
cc_1038 N_X_c_1410_n N_VGND_c_1913_n 0.00198695f $X=15.525 $Y=0.815 $X2=0 $Y2=0
cc_1039 N_X_c_1621_n N_VGND_c_1913_n 0.0188614f $X=15.69 $Y=0.39 $X2=0 $Y2=0
cc_1040 N_X_c_1425_n N_VGND_c_1913_n 0.00215161f $X=16 $Y=0.815 $X2=0 $Y2=0
cc_1041 N_X_M1002_d N_VGND_c_1919_n 0.00215201f $X=2.955 $Y=0.235 $X2=0 $Y2=0
cc_1042 N_X_M1007_d N_VGND_c_1919_n 0.00215201f $X=3.795 $Y=0.235 $X2=0 $Y2=0
cc_1043 N_X_M1010_d N_VGND_c_1919_n 0.00215201f $X=4.635 $Y=0.235 $X2=0 $Y2=0
cc_1044 N_X_M1016_d N_VGND_c_1919_n 0.00215201f $X=5.475 $Y=0.235 $X2=0 $Y2=0
cc_1045 N_X_M1022_d N_VGND_c_1919_n 0.00215201f $X=6.315 $Y=0.235 $X2=0 $Y2=0
cc_1046 N_X_M1028_d N_VGND_c_1919_n 0.00215201f $X=7.155 $Y=0.235 $X2=0 $Y2=0
cc_1047 N_X_M1062_d N_VGND_c_1919_n 0.00215201f $X=7.995 $Y=0.235 $X2=0 $Y2=0
cc_1048 N_X_M1067_d N_VGND_c_1919_n 0.00215201f $X=8.835 $Y=0.235 $X2=0 $Y2=0
cc_1049 N_X_M1018_d N_VGND_c_1919_n 0.00215201f $X=9.675 $Y=0.235 $X2=0 $Y2=0
cc_1050 N_X_M1030_d N_VGND_c_1919_n 0.00215201f $X=10.515 $Y=0.235 $X2=0 $Y2=0
cc_1051 N_X_M1035_d N_VGND_c_1919_n 0.00215201f $X=11.355 $Y=0.235 $X2=0 $Y2=0
cc_1052 N_X_M1042_d N_VGND_c_1919_n 0.00215201f $X=12.195 $Y=0.235 $X2=0 $Y2=0
cc_1053 N_X_M1045_d N_VGND_c_1919_n 0.00215201f $X=13.035 $Y=0.235 $X2=0 $Y2=0
cc_1054 N_X_M1051_d N_VGND_c_1919_n 0.00215201f $X=13.875 $Y=0.235 $X2=0 $Y2=0
cc_1055 N_X_M1056_d N_VGND_c_1919_n 0.00215201f $X=14.715 $Y=0.235 $X2=0 $Y2=0
cc_1056 N_X_M1063_d N_VGND_c_1919_n 0.00215201f $X=15.555 $Y=0.235 $X2=0 $Y2=0
cc_1057 N_X_c_1442_n N_VGND_c_1919_n 0.0122069f $X=3.09 $Y=0.39 $X2=0 $Y2=0
cc_1058 N_X_c_1395_n N_VGND_c_1919_n 0.00835832f $X=3.765 $Y=0.815 $X2=0 $Y2=0
cc_1059 N_X_c_1453_n N_VGND_c_1919_n 0.0122069f $X=3.93 $Y=0.39 $X2=0 $Y2=0
cc_1060 N_X_c_1397_n N_VGND_c_1919_n 0.00835832f $X=4.605 $Y=0.815 $X2=0 $Y2=0
cc_1061 N_X_c_1461_n N_VGND_c_1919_n 0.0122069f $X=4.77 $Y=0.39 $X2=0 $Y2=0
cc_1062 N_X_c_1398_n N_VGND_c_1919_n 0.00835832f $X=5.445 $Y=0.815 $X2=0 $Y2=0
cc_1063 N_X_c_1469_n N_VGND_c_1919_n 0.0122069f $X=5.61 $Y=0.39 $X2=0 $Y2=0
cc_1064 N_X_c_1399_n N_VGND_c_1919_n 0.00835832f $X=6.285 $Y=0.815 $X2=0 $Y2=0
cc_1065 N_X_c_1477_n N_VGND_c_1919_n 0.0122069f $X=6.45 $Y=0.39 $X2=0 $Y2=0
cc_1066 N_X_c_1400_n N_VGND_c_1919_n 0.00835832f $X=7.125 $Y=0.815 $X2=0 $Y2=0
cc_1067 N_X_c_1485_n N_VGND_c_1919_n 0.0122069f $X=7.29 $Y=0.39 $X2=0 $Y2=0
cc_1068 N_X_c_1401_n N_VGND_c_1919_n 0.00835832f $X=7.965 $Y=0.815 $X2=0 $Y2=0
cc_1069 N_X_c_1493_n N_VGND_c_1919_n 0.0122069f $X=8.13 $Y=0.39 $X2=0 $Y2=0
cc_1070 N_X_c_1402_n N_VGND_c_1919_n 0.00835832f $X=8.805 $Y=0.815 $X2=0 $Y2=0
cc_1071 N_X_c_1501_n N_VGND_c_1919_n 0.0122069f $X=8.97 $Y=0.39 $X2=0 $Y2=0
cc_1072 N_X_c_1403_n N_VGND_c_1919_n 0.00835832f $X=9.645 $Y=0.815 $X2=0 $Y2=0
cc_1073 N_X_c_1506_n N_VGND_c_1919_n 0.0122069f $X=9.81 $Y=0.39 $X2=0 $Y2=0
cc_1074 N_X_c_1404_n N_VGND_c_1919_n 0.00835832f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_1075 N_X_c_1549_n N_VGND_c_1919_n 0.0122069f $X=10.65 $Y=0.39 $X2=0 $Y2=0
cc_1076 N_X_c_1405_n N_VGND_c_1919_n 0.00835832f $X=11.325 $Y=0.815 $X2=0 $Y2=0
cc_1077 N_X_c_1561_n N_VGND_c_1919_n 0.0122069f $X=11.49 $Y=0.39 $X2=0 $Y2=0
cc_1078 N_X_c_1406_n N_VGND_c_1919_n 0.00835832f $X=12.165 $Y=0.815 $X2=0 $Y2=0
cc_1079 N_X_c_1573_n N_VGND_c_1919_n 0.0122069f $X=12.33 $Y=0.39 $X2=0 $Y2=0
cc_1080 N_X_c_1407_n N_VGND_c_1919_n 0.00835832f $X=13.005 $Y=0.815 $X2=0 $Y2=0
cc_1081 N_X_c_1585_n N_VGND_c_1919_n 0.0122069f $X=13.17 $Y=0.39 $X2=0 $Y2=0
cc_1082 N_X_c_1408_n N_VGND_c_1919_n 0.00835832f $X=13.845 $Y=0.815 $X2=0 $Y2=0
cc_1083 N_X_c_1597_n N_VGND_c_1919_n 0.0122069f $X=14.01 $Y=0.39 $X2=0 $Y2=0
cc_1084 N_X_c_1409_n N_VGND_c_1919_n 0.00835832f $X=14.685 $Y=0.815 $X2=0 $Y2=0
cc_1085 N_X_c_1609_n N_VGND_c_1919_n 0.0122069f $X=14.85 $Y=0.39 $X2=0 $Y2=0
cc_1086 N_X_c_1410_n N_VGND_c_1919_n 0.00835832f $X=15.525 $Y=0.815 $X2=0 $Y2=0
cc_1087 N_X_c_1621_n N_VGND_c_1919_n 0.0122084f $X=15.69 $Y=0.39 $X2=0 $Y2=0
cc_1088 N_X_c_1425_n N_VGND_c_1919_n 0.0104f $X=16 $Y=0.815 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__dlygate4sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
M1000 VGND a_193_47# a_299_93# VNB nshort w=420000u l=150000u
+  ad=3.139e+11p pd=3.35e+06u as=1.092e+11p ps=1.36e+06u
M1001 X a_299_93# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1002 VPWR A a_27_47# VPB phighvt w=420000u l=150000u
+  ad=3.949e+11p pd=4.03e+06u as=1.092e+11p ps=1.36e+06u
M1003 X a_299_93# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1004 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1005 VPWR a_193_47# a_299_93# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1006 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1007 a_193_47# a_27_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends


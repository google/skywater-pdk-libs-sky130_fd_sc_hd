* File: sky130_fd_sc_hd__dlxtn_4.pxi.spice
* Created: Tue Sep  1 19:06:19 2020
* 
x_PM_SKY130_FD_SC_HD__DLXTN_4%GATE_N N_GATE_N_c_150_n N_GATE_N_c_145_n
+ N_GATE_N_M1021_g N_GATE_N_c_151_n N_GATE_N_M1011_g N_GATE_N_c_146_n
+ N_GATE_N_c_152_n GATE_N GATE_N N_GATE_N_c_148_n N_GATE_N_c_149_n
+ PM_SKY130_FD_SC_HD__DLXTN_4%GATE_N
x_PM_SKY130_FD_SC_HD__DLXTN_4%A_27_47# N_A_27_47#_M1021_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1013_g N_A_27_47#_M1000_g N_A_27_47#_M1017_g N_A_27_47#_M1004_g
+ N_A_27_47#_c_342_p N_A_27_47#_c_189_n N_A_27_47#_c_190_n N_A_27_47#_c_200_n
+ N_A_27_47#_c_201_n N_A_27_47#_c_202_n N_A_27_47#_c_191_n N_A_27_47#_c_192_n
+ N_A_27_47#_c_193_n N_A_27_47#_c_194_n N_A_27_47#_c_204_n N_A_27_47#_c_205_n
+ N_A_27_47#_c_206_n N_A_27_47#_c_207_n N_A_27_47#_c_208_n N_A_27_47#_c_195_n
+ N_A_27_47#_c_196_n N_A_27_47#_c_210_n N_A_27_47#_c_197_n
+ PM_SKY130_FD_SC_HD__DLXTN_4%A_27_47#
x_PM_SKY130_FD_SC_HD__DLXTN_4%D N_D_M1005_g N_D_M1020_g D N_D_c_357_n
+ N_D_c_358_n PM_SKY130_FD_SC_HD__DLXTN_4%D
x_PM_SKY130_FD_SC_HD__DLXTN_4%A_299_47# N_A_299_47#_M1005_s N_A_299_47#_M1020_s
+ N_A_299_47#_M1010_g N_A_299_47#_M1015_g N_A_299_47#_c_403_n
+ N_A_299_47#_c_396_n N_A_299_47#_c_404_n N_A_299_47#_c_405_n
+ N_A_299_47#_c_397_n N_A_299_47#_c_398_n N_A_299_47#_c_399_n
+ N_A_299_47#_c_400_n N_A_299_47#_c_401_n PM_SKY130_FD_SC_HD__DLXTN_4%A_299_47#
x_PM_SKY130_FD_SC_HD__DLXTN_4%A_193_47# N_A_193_47#_M1013_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1001_g N_A_193_47#_c_478_n N_A_193_47#_c_479_n
+ N_A_193_47#_M1008_g N_A_193_47#_c_485_n N_A_193_47#_c_481_n
+ N_A_193_47#_c_487_n N_A_193_47#_c_488_n N_A_193_47#_c_489_n
+ N_A_193_47#_c_490_n N_A_193_47#_c_491_n N_A_193_47#_c_492_n
+ N_A_193_47#_c_493_n PM_SKY130_FD_SC_HD__DLXTN_4%A_193_47#
x_PM_SKY130_FD_SC_HD__DLXTN_4%A_724_21# N_A_724_21#_M1009_s N_A_724_21#_M1006_s
+ N_A_724_21#_M1018_g N_A_724_21#_M1007_g N_A_724_21#_c_591_n
+ N_A_724_21#_M1002_g N_A_724_21#_M1003_g N_A_724_21#_c_592_n
+ N_A_724_21#_M1012_g N_A_724_21#_M1014_g N_A_724_21#_c_593_n
+ N_A_724_21#_M1019_g N_A_724_21#_M1016_g N_A_724_21#_c_594_n
+ N_A_724_21#_M1022_g N_A_724_21#_M1023_g N_A_724_21#_c_604_n
+ N_A_724_21#_c_605_n N_A_724_21#_c_644_p N_A_724_21#_c_595_n
+ N_A_724_21#_c_606_n N_A_724_21#_c_596_n N_A_724_21#_c_624_p
+ N_A_724_21#_c_620_p N_A_724_21#_c_626_p N_A_724_21#_c_597_n
+ PM_SKY130_FD_SC_HD__DLXTN_4%A_724_21#
x_PM_SKY130_FD_SC_HD__DLXTN_4%A_561_413# N_A_561_413#_M1017_d
+ N_A_561_413#_M1001_d N_A_561_413#_c_714_n N_A_561_413#_M1009_g
+ N_A_561_413#_M1006_g N_A_561_413#_c_715_n N_A_561_413#_c_716_n
+ N_A_561_413#_c_725_n N_A_561_413#_c_728_n N_A_561_413#_c_717_n
+ N_A_561_413#_c_718_n N_A_561_413#_c_723_n N_A_561_413#_c_719_n
+ PM_SKY130_FD_SC_HD__DLXTN_4%A_561_413#
x_PM_SKY130_FD_SC_HD__DLXTN_4%VPWR N_VPWR_M1011_d N_VPWR_M1020_d N_VPWR_M1007_d
+ N_VPWR_M1006_d N_VPWR_M1014_s N_VPWR_M1023_s N_VPWR_c_797_n N_VPWR_c_798_n
+ N_VPWR_c_799_n N_VPWR_c_800_n N_VPWR_c_801_n N_VPWR_c_802_n N_VPWR_c_803_n
+ N_VPWR_c_804_n N_VPWR_c_805_n VPWR N_VPWR_c_806_n N_VPWR_c_807_n
+ N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n N_VPWR_c_812_n
+ N_VPWR_c_813_n N_VPWR_c_814_n N_VPWR_c_796_n PM_SKY130_FD_SC_HD__DLXTN_4%VPWR
x_PM_SKY130_FD_SC_HD__DLXTN_4%Q N_Q_M1002_s N_Q_M1019_s N_Q_M1003_d N_Q_M1016_d
+ N_Q_c_913_n N_Q_c_922_n N_Q_c_916_n N_Q_c_928_n Q Q Q Q Q Q Q Q Q Q
+ N_Q_c_937_n N_Q_c_918_n PM_SKY130_FD_SC_HD__DLXTN_4%Q
x_PM_SKY130_FD_SC_HD__DLXTN_4%VGND N_VGND_M1021_d N_VGND_M1005_d N_VGND_M1018_d
+ N_VGND_M1009_d N_VGND_M1012_d N_VGND_M1022_d N_VGND_c_958_n N_VGND_c_959_n
+ N_VGND_c_960_n N_VGND_c_961_n N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n
+ N_VGND_c_965_n N_VGND_c_966_n VGND N_VGND_c_967_n N_VGND_c_968_n
+ N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n
+ N_VGND_c_974_n N_VGND_c_975_n N_VGND_c_976_n PM_SKY130_FD_SC_HD__DLXTN_4%VGND
cc_1 VNB N_GATE_N_c_145_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_N_c_146_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE_N 0.0156215f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_N_c_148_n 0.0212744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_N_c_149_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1013_g 0.0397896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_189_n 0.00225054f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_8 VNB N_A_27_47#_c_190_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_191_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_192_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_193_n 0.0271287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_194_n 0.00378508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_195_n 0.0230671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_196_n 0.0176114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_197_n 0.00469707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1005_g 0.025905f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_17 VNB N_D_M1020_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_357_n 0.00407935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_19 VNB N_D_c_358_n 0.0421785f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_20 VNB N_A_299_47#_M1015_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_299_47#_c_396_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_397_n 0.00496114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_47#_c_398_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_24 VNB N_A_299_47#_c_399_n 0.00265154f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_25 VNB N_A_299_47#_c_400_n 0.0274388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_299_47#_c_401_n 0.01709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_478_n 0.0133385f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_28 VNB N_A_193_47#_c_479_n 0.00520223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_193_47#_M1008_g 0.0464035f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_30 VNB N_A_193_47#_c_481_n 0.0140955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_724_21#_M1018_g 0.0483758f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_32 VNB N_A_724_21#_c_591_n 0.0160878f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_33 VNB N_A_724_21#_c_592_n 0.0158665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_724_21#_c_593_n 0.0162704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_724_21#_c_594_n 0.0217074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_724_21#_c_595_n 0.00258236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_724_21#_c_596_n 0.00316203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_724_21#_c_597_n 0.0730409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_561_413#_c_714_n 0.0195151f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_40 VNB N_A_561_413#_c_715_n 0.0485485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_561_413#_c_716_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_42 VNB N_A_561_413#_c_717_n 0.00738412f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_A_561_413#_c_718_n 0.0118438f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_44 VNB N_A_561_413#_c_719_n 0.00297535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VPWR_c_796_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Q_c_913_n 0.00104267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB Q 8.70049e-19 $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_48 VNB Q 0.0188636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_958_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_959_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_51 VNB N_VGND_c_960_n 0.00728254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_961_n 0.0211773f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_53 VNB N_VGND_c_962_n 0.0024799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_963_n 0.0168323f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_964_n 0.00171738f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_965_n 0.0099134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_966_n 0.0233189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_967_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_968_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_969_n 0.0412073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_970_n 0.0163463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_971_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_972_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_973_n 0.00507544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_974_n 0.00423916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_975_n 0.00356594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_976_n 0.356435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VPB N_GATE_N_c_150_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_69 VPB N_GATE_N_c_151_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_70 VPB N_GATE_N_c_152_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_71 VPB GATE_N 0.0156114f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_72 VPB N_GATE_N_c_148_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_73 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_74 VPB N_A_27_47#_M1004_g 0.0212472f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_75 VPB N_A_27_47#_c_200_n 0.00126271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_201_n 0.00556025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_202_n 0.00361484f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_191_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_204_n 0.0280095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_205_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_206_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_207_n 0.0035222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_208_n 0.0037442f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_195_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_210_n 0.0330434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_47#_c_197_n 2.971e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_D_M1020_g 0.0462846f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_88 VPB N_D_c_357_n 0.00235013f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_89 VPB N_A_299_47#_M1015_g 0.0366887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_299_47#_c_403_n 0.00712099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_299_47#_c_404_n 0.00415091f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_92 VPB N_A_299_47#_c_405_n 0.00290124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_299_47#_c_398_n 0.00361895f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_94 VPB N_A_193_47#_M1001_g 0.0316829f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_95 VPB N_A_193_47#_c_478_n 0.0172364f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_96 VPB N_A_193_47#_c_479_n 0.00687211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_193_47#_c_485_n 0.0117991f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_98 VPB N_A_193_47#_c_481_n 0.00804665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_193_47#_c_487_n 0.00293933f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_100 VPB N_A_193_47#_c_488_n 0.00515533f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_101 VPB N_A_193_47#_c_489_n 0.00238602f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_102 VPB N_A_193_47#_c_490_n 0.00711634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_193_47#_c_491_n 0.00114133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_193_47#_c_492_n 0.0104341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_193_47#_c_493_n 0.0126899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_724_21#_M1018_g 0.0157271f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_107 VPB N_A_724_21#_M1007_g 0.0242212f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_108 VPB N_A_724_21#_M1003_g 0.0186895f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_109 VPB N_A_724_21#_M1014_g 0.0182275f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_110 VPB N_A_724_21#_M1016_g 0.0188626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_724_21#_M1023_g 0.0255427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_724_21#_c_604_n 0.00867028f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_724_21#_c_605_n 0.0416927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_724_21#_c_606_n 0.00377107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_724_21#_c_596_n 0.00281539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_724_21#_c_597_n 0.0142196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_561_413#_M1006_g 0.0223351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_561_413#_c_715_n 0.0169629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_561_413#_c_716_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_120 VPB N_A_561_413#_c_723_n 0.00517422f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_121 VPB N_A_561_413#_c_719_n 0.00167692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_797_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_798_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_124 VPB N_VPWR_c_799_n 0.00996035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_800_n 0.0191511f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_126 VPB N_VPWR_c_801_n 0.00194735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_802_n 0.0161675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_803_n 0.00167329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_804_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_805_n 0.0425709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_806_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_807_n 0.0295132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_808_n 0.0406078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_809_n 0.0158285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_810_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_811_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_812_n 0.00574408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_813_n 0.00421326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_814_n 0.00354005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_796_n 0.058359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_Q_c_916_n 0.00152096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB Q 0.0051586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_Q_c_918_n 0.00127285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 N_GATE_N_c_145_n N_A_27_47#_M1013_g 0.0187834f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_145 N_GATE_N_c_149_n N_A_27_47#_M1013_g 0.0041981f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_146 N_GATE_N_c_152_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_147 N_GATE_N_c_148_n N_A_27_47#_M1000_g 0.00527228f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_148 N_GATE_N_c_145_n N_A_27_47#_c_189_n 0.00663556f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_149 N_GATE_N_c_146_n N_A_27_47#_c_189_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_150 N_GATE_N_c_146_n N_A_27_47#_c_190_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_151 GATE_N N_A_27_47#_c_190_n 0.0125186f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_152 N_GATE_N_c_148_n N_A_27_47#_c_190_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_153 N_GATE_N_c_151_n N_A_27_47#_c_200_n 0.0135489f $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_154 N_GATE_N_c_152_n N_A_27_47#_c_200_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_155 N_GATE_N_c_151_n N_A_27_47#_c_202_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0
+ $Y2=0
cc_156 N_GATE_N_c_152_n N_A_27_47#_c_202_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_157 GATE_N N_A_27_47#_c_202_n 0.0139005f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_158 N_GATE_N_c_148_n N_A_27_47#_c_202_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_159 N_GATE_N_c_148_n N_A_27_47#_c_191_n 0.00319708f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_160 N_GATE_N_c_146_n N_A_27_47#_c_192_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_161 GATE_N N_A_27_47#_c_192_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_162 N_GATE_N_c_149_n N_A_27_47#_c_192_n 0.0015185f $X=0.242 $Y=1.07 $X2=0
+ $Y2=0
cc_163 N_GATE_N_c_150_n N_A_27_47#_c_205_n 0.0033897f $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_164 N_GATE_N_c_152_n N_A_27_47#_c_205_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_165 GATE_N N_A_27_47#_c_205_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_166 N_GATE_N_c_150_n N_A_27_47#_c_206_n 7.60515e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_167 N_GATE_N_c_152_n N_A_27_47#_c_206_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_168 GATE_N N_A_27_47#_c_195_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_169 N_GATE_N_c_148_n N_A_27_47#_c_195_n 0.0165992f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_170 N_GATE_N_c_151_n N_VPWR_c_797_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_171 N_GATE_N_c_151_n N_VPWR_c_806_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_172 N_GATE_N_c_151_n N_VPWR_c_796_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_173 N_GATE_N_c_145_n N_VGND_c_958_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_174 N_GATE_N_c_145_n N_VGND_c_967_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_175 N_GATE_N_c_146_n N_VGND_c_967_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_176 N_GATE_N_c_145_n N_VGND_c_976_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_204_n N_D_M1020_g 0.00583826f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_204_n N_D_c_357_n 0.0087134f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_179 N_A_27_47#_M1013_g N_D_c_358_n 0.00520956f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_204_n N_A_299_47#_M1015_g 0.00493352f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_197_n N_A_299_47#_M1015_g 0.00369716f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_182 N_A_27_47#_c_204_n N_A_299_47#_c_404_n 0.0116478f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_204_n N_A_299_47#_c_405_n 0.0115067f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_193_n N_A_299_47#_c_397_n 9.56555e-19 $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_194_n N_A_299_47#_c_397_n 0.0129081f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_204_n N_A_299_47#_c_397_n 0.00675641f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_197_n N_A_299_47#_c_397_n 0.00178567f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_188 N_A_27_47#_c_204_n N_A_299_47#_c_398_n 0.0108506f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_193_n N_A_299_47#_c_400_n 0.0117556f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_194_n N_A_299_47#_c_400_n 9.50608e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_204_n N_A_299_47#_c_400_n 0.00107604f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_197_n N_A_299_47#_c_400_n 9.9633e-19 $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_193_n N_A_299_47#_c_401_n 0.00200147f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_194_n N_A_299_47#_c_401_n 2.04855e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_196_n N_A_299_47#_c_401_n 0.0197936f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_M1004_g N_A_193_47#_M1001_g 0.014011f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_201_n N_A_193_47#_M1001_g 0.00220245f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_194_n N_A_193_47#_c_478_n 7.03475e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_204_n N_A_193_47#_c_478_n 0.00144279f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_207_n N_A_193_47#_c_478_n 0.00140497f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_208_n N_A_193_47#_c_478_n 0.0049391f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_210_n N_A_193_47#_c_478_n 0.0184089f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_197_n N_A_193_47#_c_478_n 0.01293f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_193_n N_A_193_47#_c_479_n 0.0186665f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_194_n N_A_193_47#_c_479_n 0.00136525f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_193_n N_A_193_47#_M1008_g 0.0192792f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_194_n N_A_193_47#_M1008_g 0.00256371f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_196_n N_A_193_47#_M1008_g 0.0126141f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_197_n N_A_193_47#_M1008_g 0.0049729f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_204_n N_A_193_47#_c_485_n 0.00274258f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_207_n N_A_193_47#_c_485_n 7.88621e-19 $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_208_n N_A_193_47#_c_485_n 0.00220245f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_210_n N_A_193_47#_c_485_n 0.0160512f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1013_g N_A_193_47#_c_481_n 0.00779983f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_189_n N_A_193_47#_c_481_n 0.00991525f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_191_n N_A_193_47#_c_481_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_192_n N_A_193_47#_c_481_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_204_n N_A_193_47#_c_481_n 0.0184539f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_205_n N_A_193_47#_c_481_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_206_n N_A_193_47#_c_481_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_200_n N_A_193_47#_c_487_n 0.00293827f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_204_n N_A_193_47#_c_487_n 0.00195186f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_195_n N_A_193_47#_c_487_n 0.00779983f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_204_n N_A_193_47#_c_488_n 0.0871075f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_M1000_g N_A_193_47#_c_489_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_200_n N_A_193_47#_c_489_n 0.00549495f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_204_n N_A_193_47#_c_489_n 0.0259095f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_c_206_n N_A_193_47#_c_489_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_M1000_g N_A_193_47#_c_490_n 0.00779983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_201_n N_A_193_47#_c_491_n 0.00155445f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_204_n N_A_193_47#_c_491_n 0.0255946f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_204_n N_A_193_47#_c_492_n 0.00169866f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_207_n N_A_193_47#_c_492_n 0.00124306f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_197_n N_A_193_47#_c_492_n 0.00220245f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_235 N_A_27_47#_c_193_n N_A_193_47#_c_493_n 4.0812e-19 $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_194_n N_A_193_47#_c_493_n 0.00161882f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_204_n N_A_193_47#_c_493_n 0.0240266f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_207_n N_A_193_47#_c_493_n 0.00272314f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_210_n N_A_193_47#_c_493_n 2.5966e-19 $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_197_n N_A_193_47#_c_493_n 0.0454941f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_208_n N_A_724_21#_M1018_g 4.9921e-19 $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_197_n N_A_724_21#_M1018_g 2.17095e-19 $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_243 N_A_27_47#_M1004_g N_A_724_21#_M1007_g 0.0313447f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_201_n N_A_724_21#_c_605_n 8.09252e-19 $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_210_n N_A_724_21#_c_605_n 0.0313447f $X=3.335 $Y=1.74 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_193_n N_A_561_413#_c_725_n 0.00144439f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_194_n N_A_561_413#_c_725_n 0.0162478f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_196_n N_A_561_413#_c_725_n 0.00412044f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1004_g N_A_561_413#_c_728_n 0.0116262f $X=3.335 $Y=2.275
+ $X2=0 $Y2=0
cc_250 N_A_27_47#_c_201_n N_A_561_413#_c_728_n 0.016081f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_207_n N_A_561_413#_c_728_n 0.00173361f $X=3.015 $Y=1.53
+ $X2=0 $Y2=0
cc_252 N_A_27_47#_c_210_n N_A_561_413#_c_728_n 0.00111122f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_194_n N_A_561_413#_c_717_n 0.0184898f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_194_n N_A_561_413#_c_718_n 0.0027819f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_210_n N_A_561_413#_c_718_n 0.00291146f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_256 N_A_27_47#_c_197_n N_A_561_413#_c_718_n 0.016104f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_207_n N_A_561_413#_c_723_n 0.00130345f $X=3.015 $Y=1.53
+ $X2=0 $Y2=0
cc_258 N_A_27_47#_c_208_n N_A_561_413#_c_723_n 0.0359174f $X=3.015 $Y=1.53 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_210_n N_A_561_413#_c_723_n 0.00856317f $X=3.335 $Y=1.74
+ $X2=0 $Y2=0
cc_260 N_A_27_47#_c_197_n N_A_561_413#_c_723_n 0.00353544f $X=3.095 $Y=1.415
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_200_n N_VPWR_M1011_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_262 N_A_27_47#_M1000_g N_VPWR_c_797_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_200_n N_VPWR_c_797_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_202_n N_VPWR_c_797_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_205_n N_VPWR_c_797_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_204_n N_VPWR_c_798_n 0.0019389f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_200_n N_VPWR_c_806_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_202_n N_VPWR_c_806_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1000_g N_VPWR_c_807_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1004_g N_VPWR_c_808_n 0.00366111f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1000_g N_VPWR_c_796_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1004_g N_VPWR_c_796_n 0.00549379f $X=3.335 $Y=2.275 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_200_n N_VPWR_c_796_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_202_n N_VPWR_c_796_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_189_n N_VGND_M1021_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_276 N_A_27_47#_M1013_g N_VGND_c_958_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_189_n N_VGND_c_958_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_191_n N_VGND_c_958_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_195_n N_VGND_c_958_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_196_n N_VGND_c_959_n 0.00174223f $X=2.8 $Y=0.705 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_342_p N_VGND_c_967_n 0.00713694f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_189_n N_VGND_c_967_n 0.00243651f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_283 N_A_27_47#_M1013_g N_VGND_c_968_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_193_n N_VGND_c_969_n 9.43262e-19 $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_194_n N_VGND_c_969_n 0.00182549f $X=3.01 $Y=0.87 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_196_n N_VGND_c_969_n 0.00425892f $X=2.8 $Y=0.705 $X2=0 $Y2=0
cc_287 N_A_27_47#_M1021_s N_VGND_c_976_n 0.003754f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_288 N_A_27_47#_M1013_g N_VGND_c_976_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_342_p N_VGND_c_976_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_189_n N_VGND_c_976_n 0.00549708f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_193_n N_VGND_c_976_n 0.00121904f $X=2.8 $Y=0.87 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_194_n N_VGND_c_976_n 0.00328555f $X=3.01 $Y=0.87 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_196_n N_VGND_c_976_n 0.00628992f $X=2.8 $Y=0.705 $X2=0 $Y2=0
cc_294 N_D_c_358_n N_A_299_47#_M1015_g 0.0382098f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_295 N_D_M1020_g N_A_299_47#_c_403_n 0.012851f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_296 N_D_M1005_g N_A_299_47#_c_396_n 0.0144498f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_297 N_D_c_357_n N_A_299_47#_c_396_n 0.00627239f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_298 N_D_c_358_n N_A_299_47#_c_396_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_299 N_D_M1020_g N_A_299_47#_c_404_n 0.00794545f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_300 N_D_M1020_g N_A_299_47#_c_405_n 0.00412429f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_301 N_D_c_357_n N_A_299_47#_c_405_n 0.0229667f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_302 N_D_c_358_n N_A_299_47#_c_405_n 0.00131849f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_303 N_D_M1005_g N_A_299_47#_c_397_n 0.00563568f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_304 N_D_c_357_n N_A_299_47#_c_397_n 0.0107593f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_305 N_D_c_357_n N_A_299_47#_c_398_n 0.0164827f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_306 N_D_c_358_n N_A_299_47#_c_398_n 0.00552652f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_307 N_D_M1005_g N_A_299_47#_c_399_n 0.00120855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_308 N_D_c_357_n N_A_299_47#_c_399_n 0.0138491f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_309 N_D_c_358_n N_A_299_47#_c_399_n 0.0042466f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_310 N_D_M1005_g N_A_299_47#_c_400_n 0.0197208f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_311 N_D_M1005_g N_A_299_47#_c_401_n 0.015283f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_312 N_D_M1005_g N_A_193_47#_c_481_n 0.00203374f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_313 N_D_M1020_g N_A_193_47#_c_481_n 0.00459933f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_314 N_D_c_357_n N_A_193_47#_c_481_n 0.0209974f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_315 N_D_c_358_n N_A_193_47#_c_481_n 0.00256393f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_316 N_D_M1020_g N_A_193_47#_c_487_n 0.00134564f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_317 N_D_M1020_g N_A_193_47#_c_488_n 0.00294239f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_318 N_D_M1020_g N_VPWR_c_798_n 0.00304701f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_319 N_D_M1020_g N_VPWR_c_807_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_320 N_D_M1020_g N_VPWR_c_796_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_321 N_D_M1005_g N_VGND_c_959_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_322 N_D_M1005_g N_VGND_c_968_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_323 N_D_M1005_g N_VGND_c_976_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_324 N_D_c_358_n N_VGND_c_976_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_325 N_A_299_47#_M1015_g N_A_193_47#_M1001_g 0.0342299f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_326 N_A_299_47#_M1015_g N_A_193_47#_c_479_n 0.0248238f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_327 N_A_299_47#_c_403_n N_A_193_47#_c_481_n 0.0010921f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_328 N_A_299_47#_c_405_n N_A_193_47#_c_481_n 0.00859001f $X=1.785 $Y=1.58
+ $X2=0 $Y2=0
cc_329 N_A_299_47#_c_399_n N_A_193_47#_c_481_n 0.0191833f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_330 N_A_299_47#_c_403_n N_A_193_47#_c_487_n 0.0471072f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_331 N_A_299_47#_M1015_g N_A_193_47#_c_488_n 0.00365242f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_332 N_A_299_47#_c_403_n N_A_193_47#_c_488_n 0.022748f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_333 N_A_299_47#_c_404_n N_A_193_47#_c_488_n 0.00551435f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_334 N_A_299_47#_c_403_n N_A_193_47#_c_489_n 0.00273055f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_M1015_g N_A_193_47#_c_491_n 0.00149195f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_336 N_A_299_47#_M1015_g N_A_193_47#_c_493_n 0.00673436f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_337 N_A_299_47#_c_404_n N_A_193_47#_c_493_n 0.00754519f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_398_n N_A_193_47#_c_493_n 0.00645446f $X=2.055 $Y=1.495
+ $X2=0 $Y2=0
cc_339 N_A_299_47#_c_401_n N_A_561_413#_c_725_n 6.54613e-19 $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_340 N_A_299_47#_M1015_g N_VPWR_c_798_n 0.0223997f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_341 N_A_299_47#_c_403_n N_VPWR_c_798_n 0.0232987f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_342 N_A_299_47#_c_404_n N_VPWR_c_798_n 0.013562f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_343 N_A_299_47#_c_403_n N_VPWR_c_807_n 0.0159418f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_344 N_A_299_47#_M1015_g N_VPWR_c_808_n 0.00212864f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_345 N_A_299_47#_M1020_s N_VPWR_c_796_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_M1015_g N_VPWR_c_796_n 0.00262666f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_347 N_A_299_47#_c_403_n N_VPWR_c_796_n 0.00576627f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_348 N_A_299_47#_c_397_n N_VGND_M1005_d 0.00156939f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_349 N_A_299_47#_c_396_n N_VGND_c_959_n 0.00259081f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_350 N_A_299_47#_c_397_n N_VGND_c_959_n 0.0141976f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_351 N_A_299_47#_c_401_n N_VGND_c_959_n 0.00964732f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_352 N_A_299_47#_c_396_n N_VGND_c_968_n 0.00255672f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_353 N_A_299_47#_c_399_n N_VGND_c_968_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_354 N_A_299_47#_c_400_n N_VGND_c_969_n 9.84895e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_355 N_A_299_47#_c_401_n N_VGND_c_969_n 0.0046653f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_356 N_A_299_47#_M1005_s N_VGND_c_976_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_357 N_A_299_47#_c_396_n N_VGND_c_976_n 0.00473142f $X=1.97 $Y=0.7 $X2=0 $Y2=0
cc_358 N_A_299_47#_c_397_n N_VGND_c_976_n 0.00552372f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_359 N_A_299_47#_c_399_n N_VGND_c_976_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_360 N_A_299_47#_c_400_n N_VGND_c_976_n 0.00117722f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_361 N_A_299_47#_c_401_n N_VGND_c_976_n 0.00454932f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_362 N_A_193_47#_M1008_g N_A_724_21#_M1018_g 0.0429816f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_363 N_A_193_47#_M1008_g N_A_561_413#_c_725_n 0.0125275f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_364 N_A_193_47#_M1001_g N_A_561_413#_c_728_n 0.00281839f $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_365 N_A_193_47#_M1008_g N_A_561_413#_c_717_n 0.00562201f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_366 N_A_193_47#_M1008_g N_A_561_413#_c_718_n 0.00348305f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_367 N_A_193_47#_M1001_g N_A_561_413#_c_723_n 8.05921e-19 $X=2.73 $Y=2.275
+ $X2=0 $Y2=0
cc_368 N_A_193_47#_c_478_n N_A_561_413#_c_723_n 6.71539e-19 $X=3.145 $Y=1.32
+ $X2=0 $Y2=0
cc_369 N_A_193_47#_c_488_n N_VPWR_M1020_d 6.81311e-19 $X=2.41 $Y=1.87 $X2=0
+ $Y2=0
cc_370 N_A_193_47#_c_490_n N_VPWR_c_797_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_M1001_g N_VPWR_c_798_n 0.00357414f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_372 N_A_193_47#_c_488_n N_VPWR_c_798_n 0.0171797f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_373 N_A_193_47#_c_491_n N_VPWR_c_798_n 0.0013481f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_493_n N_VPWR_c_798_n 0.00972665f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_375 N_A_193_47#_c_490_n N_VPWR_c_807_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_376 N_A_193_47#_M1001_g N_VPWR_c_808_n 0.00487021f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_377 N_A_193_47#_c_493_n N_VPWR_c_808_n 0.00456724f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_378 N_A_193_47#_M1001_g N_VPWR_c_796_n 0.00815857f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_488_n N_VPWR_c_796_n 0.0516753f $X=2.41 $Y=1.87 $X2=0 $Y2=0
cc_380 N_A_193_47#_c_489_n N_VPWR_c_796_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_381 N_A_193_47#_c_490_n N_VPWR_c_796_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_382 N_A_193_47#_c_491_n N_VPWR_c_796_n 0.0151013f $X=2.555 $Y=1.87 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_c_493_n N_VPWR_c_796_n 0.00403974f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_384 N_A_193_47#_c_488_n A_465_369# 0.00119229f $X=2.41 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_385 N_A_193_47#_c_491_n A_465_369# 0.00120144f $X=2.555 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_386 N_A_193_47#_c_493_n A_465_369# 0.0030615f $X=2.67 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_387 N_A_193_47#_M1008_g N_VGND_c_960_n 0.0017297f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_388 N_A_193_47#_c_481_n N_VGND_c_968_n 0.00732874f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_389 N_A_193_47#_M1008_g N_VGND_c_969_n 0.0037981f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_390 N_A_193_47#_M1013_d N_VGND_c_976_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_391 N_A_193_47#_M1008_g N_VGND_c_976_n 0.00555936f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_392 N_A_193_47#_c_481_n N_VGND_c_976_n 0.00616598f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_393 N_A_724_21#_c_591_n N_A_561_413#_c_714_n 0.0211139f $X=5.115 $Y=0.995
+ $X2=0 $Y2=0
cc_394 N_A_724_21#_c_595_n N_A_561_413#_c_714_n 0.00671379f $X=4.52 $Y=0.995
+ $X2=0 $Y2=0
cc_395 N_A_724_21#_M1003_g N_A_561_413#_M1006_g 0.0230216f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_396 N_A_724_21#_c_605_n N_A_561_413#_M1006_g 0.00295738f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_397 N_A_724_21#_c_606_n N_A_561_413#_M1006_g 0.00755466f $X=4.52 $Y=1.535
+ $X2=0 $Y2=0
cc_398 N_A_724_21#_c_620_p N_A_561_413#_M1006_g 3.19411e-19 $X=4.47 $Y=1.755
+ $X2=0 $Y2=0
cc_399 N_A_724_21#_M1018_g N_A_561_413#_c_715_n 0.0214321f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_400 N_A_724_21#_c_604_n N_A_561_413#_c_715_n 0.0105366f $X=4.385 $Y=1.7 $X2=0
+ $Y2=0
cc_401 N_A_724_21#_c_605_n N_A_561_413#_c_715_n 0.00487525f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_402 N_A_724_21#_c_624_p N_A_561_413#_c_715_n 0.00182108f $X=4.47 $Y=0.58
+ $X2=0 $Y2=0
cc_403 N_A_724_21#_c_620_p N_A_561_413#_c_715_n 0.00212837f $X=4.47 $Y=1.755
+ $X2=0 $Y2=0
cc_404 N_A_724_21#_c_626_p N_A_561_413#_c_715_n 0.018768f $X=4.52 $Y=1.16 $X2=0
+ $Y2=0
cc_405 N_A_724_21#_c_596_n N_A_561_413#_c_716_n 0.0218433f $X=5.1 $Y=1.16 $X2=0
+ $Y2=0
cc_406 N_A_724_21#_c_597_n N_A_561_413#_c_716_n 0.0216214f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_407 N_A_724_21#_M1018_g N_A_561_413#_c_725_n 0.00158904f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_408 N_A_724_21#_M1007_g N_A_561_413#_c_728_n 0.00369776f $X=3.695 $Y=2.275
+ $X2=0 $Y2=0
cc_409 N_A_724_21#_M1018_g N_A_561_413#_c_717_n 0.010318f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_724_21#_M1018_g N_A_561_413#_c_718_n 0.00570022f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_411 N_A_724_21#_M1018_g N_A_561_413#_c_723_n 0.0114233f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_412 N_A_724_21#_M1007_g N_A_561_413#_c_723_n 0.0143765f $X=3.695 $Y=2.275
+ $X2=0 $Y2=0
cc_413 N_A_724_21#_c_604_n N_A_561_413#_c_723_n 0.0228437f $X=4.385 $Y=1.7 $X2=0
+ $Y2=0
cc_414 N_A_724_21#_c_605_n N_A_561_413#_c_723_n 0.00824307f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_415 N_A_724_21#_M1018_g N_A_561_413#_c_719_n 0.0173045f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_416 N_A_724_21#_c_604_n N_A_561_413#_c_719_n 0.02399f $X=4.385 $Y=1.7 $X2=0
+ $Y2=0
cc_417 N_A_724_21#_c_605_n N_A_561_413#_c_719_n 0.006103f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_418 N_A_724_21#_c_626_p N_A_561_413#_c_719_n 0.0214234f $X=4.52 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A_724_21#_M1007_g N_VPWR_c_799_n 0.00454869f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_420 N_A_724_21#_c_604_n N_VPWR_c_799_n 0.0154822f $X=4.385 $Y=1.7 $X2=0 $Y2=0
cc_421 N_A_724_21#_c_605_n N_VPWR_c_799_n 0.00545641f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_422 N_A_724_21#_c_644_p N_VPWR_c_799_n 0.0172074f $X=4.47 $Y=2.27 $X2=0 $Y2=0
cc_423 N_A_724_21#_c_644_p N_VPWR_c_800_n 0.0112378f $X=4.47 $Y=2.27 $X2=0 $Y2=0
cc_424 N_A_724_21#_M1003_g N_VPWR_c_801_n 0.0172087f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_425 N_A_724_21#_M1014_g N_VPWR_c_801_n 8.84439e-19 $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_A_724_21#_c_596_n N_VPWR_c_801_n 0.020301f $X=5.1 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A_724_21#_c_597_n N_VPWR_c_801_n 0.00157349f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_428 N_A_724_21#_M1003_g N_VPWR_c_802_n 0.0046653f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_429 N_A_724_21#_M1014_g N_VPWR_c_802_n 0.00489117f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_430 N_A_724_21#_M1014_g N_VPWR_c_803_n 0.00525059f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_431 N_A_724_21#_M1016_g N_VPWR_c_803_n 0.0166964f $X=5.99 $Y=1.985 $X2=0
+ $Y2=0
cc_432 N_A_724_21#_M1023_g N_VPWR_c_803_n 8.45569e-19 $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_433 N_A_724_21#_c_597_n N_VPWR_c_803_n 0.00291196f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_434 N_A_724_21#_M1023_g N_VPWR_c_805_n 0.0071918f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_435 N_A_724_21#_M1007_g N_VPWR_c_808_n 0.00541489f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_436 N_A_724_21#_M1016_g N_VPWR_c_809_n 0.0046653f $X=5.99 $Y=1.985 $X2=0
+ $Y2=0
cc_437 N_A_724_21#_M1023_g N_VPWR_c_809_n 0.00541763f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_438 N_A_724_21#_M1006_s N_VPWR_c_796_n 0.0023739f $X=4.345 $Y=1.485 $X2=0
+ $Y2=0
cc_439 N_A_724_21#_M1007_g N_VPWR_c_796_n 0.0106979f $X=3.695 $Y=2.275 $X2=0
+ $Y2=0
cc_440 N_A_724_21#_M1003_g N_VPWR_c_796_n 0.00789179f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_441 N_A_724_21#_M1014_g N_VPWR_c_796_n 0.00838592f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_442 N_A_724_21#_M1016_g N_VPWR_c_796_n 0.00794405f $X=5.99 $Y=1.985 $X2=0
+ $Y2=0
cc_443 N_A_724_21#_M1023_g N_VPWR_c_796_n 0.0105084f $X=6.43 $Y=1.985 $X2=0
+ $Y2=0
cc_444 N_A_724_21#_c_604_n N_VPWR_c_796_n 0.0106057f $X=4.385 $Y=1.7 $X2=0 $Y2=0
cc_445 N_A_724_21#_c_605_n N_VPWR_c_796_n 0.00110429f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_446 N_A_724_21#_c_644_p N_VPWR_c_796_n 0.00827281f $X=4.47 $Y=2.27 $X2=0
+ $Y2=0
cc_447 N_A_724_21#_c_591_n N_Q_c_913_n 0.00503846f $X=5.115 $Y=0.995 $X2=0 $Y2=0
cc_448 N_A_724_21#_c_592_n N_Q_c_913_n 0.00592887f $X=5.535 $Y=0.995 $X2=0 $Y2=0
cc_449 N_A_724_21#_c_593_n N_Q_c_913_n 5.58257e-19 $X=5.99 $Y=0.995 $X2=0 $Y2=0
cc_450 N_A_724_21#_M1014_g N_Q_c_922_n 0.00307509f $X=5.535 $Y=1.985 $X2=0 $Y2=0
cc_451 N_A_724_21#_M1016_g N_Q_c_922_n 3.9102e-19 $X=5.99 $Y=1.985 $X2=0 $Y2=0
cc_452 N_A_724_21#_c_597_n N_Q_c_922_n 0.0033331f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_453 N_A_724_21#_M1003_g N_Q_c_916_n 0.00348055f $X=5.115 $Y=1.985 $X2=0 $Y2=0
cc_454 N_A_724_21#_M1014_g N_Q_c_916_n 0.00458323f $X=5.535 $Y=1.985 $X2=0 $Y2=0
cc_455 N_A_724_21#_M1016_g N_Q_c_916_n 5.57351e-19 $X=5.99 $Y=1.985 $X2=0 $Y2=0
cc_456 N_A_724_21#_c_596_n N_Q_c_928_n 0.0277655f $X=5.1 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_724_21#_c_597_n N_Q_c_928_n 0.0105619f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_458 N_A_724_21#_c_592_n Q 0.0052048f $X=5.535 $Y=0.995 $X2=0 $Y2=0
cc_459 N_A_724_21#_c_597_n Q 0.00278736f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_460 N_A_724_21#_M1014_g Q 0.0116355f $X=5.535 $Y=1.985 $X2=0 $Y2=0
cc_461 N_A_724_21#_c_597_n Q 0.0136637f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_724_21#_c_593_n Q 0.00206535f $X=5.99 $Y=0.995 $X2=0 $Y2=0
cc_463 N_A_724_21#_c_594_n Q 0.0183717f $X=6.43 $Y=0.995 $X2=0 $Y2=0
cc_464 N_A_724_21#_c_597_n Q 0.0216925f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_465 N_A_724_21#_c_597_n N_Q_c_937_n 0.0551622f $X=6.43 $Y=1.16 $X2=0 $Y2=0
cc_466 N_A_724_21#_M1016_g N_Q_c_918_n 0.0030861f $X=5.99 $Y=1.985 $X2=0 $Y2=0
cc_467 N_A_724_21#_M1023_g N_Q_c_918_n 0.0217052f $X=6.43 $Y=1.985 $X2=0 $Y2=0
cc_468 N_A_724_21#_M1018_g N_VGND_c_960_n 0.0115145f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_469 N_A_724_21#_c_624_p N_VGND_c_960_n 0.00588176f $X=4.47 $Y=0.58 $X2=0
+ $Y2=0
cc_470 N_A_724_21#_c_624_p N_VGND_c_961_n 0.00650283f $X=4.47 $Y=0.58 $X2=0
+ $Y2=0
cc_471 N_A_724_21#_c_591_n N_VGND_c_962_n 0.0119984f $X=5.115 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_724_21#_c_592_n N_VGND_c_962_n 9.5832e-19 $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_473 N_A_724_21#_c_596_n N_VGND_c_962_n 0.0140068f $X=5.1 $Y=1.16 $X2=0 $Y2=0
cc_474 N_A_724_21#_c_597_n N_VGND_c_962_n 0.00142002f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_A_724_21#_c_591_n N_VGND_c_963_n 0.0046653f $X=5.115 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_A_724_21#_c_592_n N_VGND_c_963_n 0.00501545f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_477 N_A_724_21#_c_592_n N_VGND_c_964_n 0.00493342f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_724_21#_c_593_n N_VGND_c_964_n 0.0134596f $X=5.99 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_A_724_21#_c_594_n N_VGND_c_964_n 0.00100593f $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_A_724_21#_c_597_n N_VGND_c_964_n 0.00291196f $X=6.43 $Y=1.16 $X2=0
+ $Y2=0
cc_481 N_A_724_21#_c_594_n N_VGND_c_966_n 0.00544514f $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_482 N_A_724_21#_M1018_g N_VGND_c_969_n 0.0046653f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_483 N_A_724_21#_c_593_n N_VGND_c_970_n 0.0046653f $X=5.99 $Y=0.995 $X2=0
+ $Y2=0
cc_484 N_A_724_21#_c_594_n N_VGND_c_970_n 0.0054633f $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_485 N_A_724_21#_M1009_s N_VGND_c_976_n 0.00370868f $X=4.345 $Y=0.235 $X2=0
+ $Y2=0
cc_486 N_A_724_21#_M1018_g N_VGND_c_976_n 0.00813035f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_487 N_A_724_21#_c_591_n N_VGND_c_976_n 0.00796766f $X=5.115 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_A_724_21#_c_592_n N_VGND_c_976_n 0.00856637f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_489 N_A_724_21#_c_593_n N_VGND_c_976_n 0.00802193f $X=5.99 $Y=0.995 $X2=0
+ $Y2=0
cc_490 N_A_724_21#_c_594_n N_VGND_c_976_n 0.0106813f $X=6.43 $Y=0.995 $X2=0
+ $Y2=0
cc_491 N_A_724_21#_c_624_p N_VGND_c_976_n 0.00761394f $X=4.47 $Y=0.58 $X2=0
+ $Y2=0
cc_492 N_A_561_413#_c_728_n N_VPWR_c_798_n 0.00489615f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_493 N_A_561_413#_M1006_g N_VPWR_c_799_n 0.0024426f $X=4.68 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_A_561_413#_M1006_g N_VPWR_c_800_n 0.00585385f $X=4.68 $Y=1.985 $X2=0
+ $Y2=0
cc_495 N_A_561_413#_M1006_g N_VPWR_c_801_n 0.00277946f $X=4.68 $Y=1.985 $X2=0
+ $Y2=0
cc_496 N_A_561_413#_c_728_n N_VPWR_c_808_n 0.0343719f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_497 N_A_561_413#_M1001_d N_VPWR_c_796_n 0.00699187f $X=2.805 $Y=2.065 $X2=0
+ $Y2=0
cc_498 N_A_561_413#_M1006_g N_VPWR_c_796_n 0.0120037f $X=4.68 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A_561_413#_c_728_n N_VPWR_c_796_n 0.0265731f $X=3.48 $Y=2.34 $X2=0
+ $Y2=0
cc_500 N_A_561_413#_c_728_n A_682_413# 0.00145479f $X=3.48 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_501 N_A_561_413#_c_723_n A_682_413# 0.00208506f $X=3.565 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_502 N_A_561_413#_c_725_n N_VGND_c_959_n 0.00209539f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_503 N_A_561_413#_c_714_n N_VGND_c_960_n 0.00635953f $X=4.68 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_561_413#_c_715_n N_VGND_c_960_n 0.00169847f $X=4.605 $Y=1.16 $X2=0
+ $Y2=0
cc_505 N_A_561_413#_c_725_n N_VGND_c_960_n 0.010424f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_506 N_A_561_413#_c_719_n N_VGND_c_960_n 0.0119873f $X=4.115 $Y=1.16 $X2=0
+ $Y2=0
cc_507 N_A_561_413#_c_714_n N_VGND_c_961_n 0.00585385f $X=4.68 $Y=0.995 $X2=0
+ $Y2=0
cc_508 N_A_561_413#_c_714_n N_VGND_c_962_n 0.00350707f $X=4.68 $Y=0.995 $X2=0
+ $Y2=0
cc_509 N_A_561_413#_c_725_n N_VGND_c_969_n 0.0221606f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_510 N_A_561_413#_M1017_d N_VGND_c_976_n 0.00237979f $X=2.865 $Y=0.235 $X2=0
+ $Y2=0
cc_511 N_A_561_413#_c_714_n N_VGND_c_976_n 0.0120818f $X=4.68 $Y=0.995 $X2=0
+ $Y2=0
cc_512 N_A_561_413#_c_725_n N_VGND_c_976_n 0.0222941f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_513 N_A_561_413#_c_725_n A_659_47# 0.00365607f $X=3.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_514 N_A_561_413#_c_717_n A_659_47# 0.00149829f $X=3.415 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_515 N_VPWR_c_796_n A_465_369# 0.00373974f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_516 N_VPWR_c_796_n A_682_413# 0.00170472f $X=6.67 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_517 N_VPWR_c_796_n N_Q_M1003_d 0.00389051f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_518 N_VPWR_c_796_n N_Q_M1016_d 0.00405136f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_519 N_VPWR_c_803_n N_Q_c_922_n 0.0721194f $X=5.78 $Y=1.835 $X2=0 $Y2=0
cc_520 N_VPWR_c_802_n Q 0.0164828f $X=5.695 $Y=2.72 $X2=0 $Y2=0
cc_521 N_VPWR_c_796_n Q 0.0104806f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_522 N_VPWR_c_805_n Q 0.0221837f $X=6.64 $Y=1.835 $X2=0 $Y2=0
cc_523 N_VPWR_c_803_n N_Q_c_937_n 0.017842f $X=5.78 $Y=1.835 $X2=0 $Y2=0
cc_524 N_VPWR_c_809_n N_Q_c_918_n 0.0155653f $X=6.555 $Y=2.72 $X2=0 $Y2=0
cc_525 N_VPWR_c_796_n N_Q_c_918_n 0.0100668f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_526 Q N_VGND_c_963_n 0.00840617f $X=5.295 $Y=0.425 $X2=0 $Y2=0
cc_527 Q N_VGND_c_964_n 0.0305589f $X=5.295 $Y=0.425 $X2=0 $Y2=0
cc_528 N_Q_c_937_n N_VGND_c_964_n 0.017842f $X=6.115 $Y=1.16 $X2=0 $Y2=0
cc_529 Q N_VGND_c_966_n 0.0155287f $X=6.62 $Y=1.105 $X2=0 $Y2=0
cc_530 Q N_VGND_c_970_n 0.00900416f $X=6.215 $Y=0.425 $X2=0 $Y2=0
cc_531 N_Q_M1002_s N_VGND_c_976_n 0.0041316f $X=5.19 $Y=0.235 $X2=0 $Y2=0
cc_532 N_Q_M1019_s N_VGND_c_976_n 0.00424646f $X=6.065 $Y=0.235 $X2=0 $Y2=0
cc_533 Q N_VGND_c_976_n 0.00950977f $X=5.295 $Y=0.425 $X2=0 $Y2=0
cc_534 Q N_VGND_c_976_n 0.00944386f $X=6.215 $Y=0.425 $X2=0 $Y2=0
cc_535 N_VGND_c_976_n A_465_47# 0.0139156f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24
cc_536 N_VGND_c_976_n A_659_47# 0.00687059f $X=6.67 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__lpflow_inputiso0n_1.pxi.spice
* Created: Tue Sep  1 19:12:03 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%A N_A_M1004_g N_A_M1000_g A A A
+ N_A_c_49_n N_A_c_50_n PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%A
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%SLEEP_B N_SLEEP_B_M1002_g
+ N_SLEEP_B_M1005_g SLEEP_B N_SLEEP_B_c_83_n
+ PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%SLEEP_B
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%A_59_75# N_A_59_75#_M1004_s
+ N_A_59_75#_M1000_d N_A_59_75#_M1003_g N_A_59_75#_M1001_g N_A_59_75#_c_117_n
+ N_A_59_75#_c_118_n N_A_59_75#_c_119_n N_A_59_75#_c_124_n N_A_59_75#_c_125_n
+ N_A_59_75#_c_126_n N_A_59_75#_c_120_n N_A_59_75#_c_128_n N_A_59_75#_c_121_n
+ N_A_59_75#_c_122_n PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%A_59_75#
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%VPWR N_VPWR_M1000_s N_VPWR_M1005_d
+ N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_196_n N_VPWR_c_197_n N_VPWR_c_198_n
+ N_VPWR_c_199_n VPWR N_VPWR_c_200_n N_VPWR_c_193_n
+ PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%X N_X_M1003_d N_X_M1001_d N_X_c_228_n
+ X X X X X X N_X_c_225_n X PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%X
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%VGND N_VGND_M1002_d N_VGND_c_250_n
+ N_VGND_c_251_n N_VGND_c_252_n VGND N_VGND_c_253_n N_VGND_c_254_n
+ PM_SKY130_FD_SC_HD__LPFLOW_INPUTISO0N_1%VGND
cc_1 VNB N_A_M1004_g 0.0276828f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.585
cc_2 VNB A 0.00202634f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_3 VNB N_A_c_49_n 0.0362409f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_4 VNB N_A_c_50_n 0.0168455f $X=-0.19 $Y=-0.24 $X2=0.232 $Y2=1.325
cc_5 VNB N_SLEEP_B_M1002_g 0.0214739f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.585
cc_6 VNB SLEEP_B 0.00149897f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_7 VNB N_SLEEP_B_c_83_n 0.0246237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_59_75#_c_117_n 0.0160682f $X=-0.19 $Y=-0.24 $X2=0.455 $Y2=1.16
cc_9 VNB N_A_59_75#_c_118_n 0.0075306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_59_75#_c_119_n 0.00986719f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_11 VNB N_A_59_75#_c_120_n 0.00477226f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.2
cc_12 VNB N_A_59_75#_c_121_n 0.0264677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_59_75#_c_122_n 0.0221591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_193_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB X 0.0399604f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_16 VNB N_X_c_225_n 0.0159574f $X=-0.19 $Y=-0.24 $X2=0.455 $Y2=1.2
cc_17 VNB N_VGND_c_250_n 0.00682552f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=2.065
cc_18 VNB N_VGND_c_251_n 0.0365485f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_VGND_c_252_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_20 VNB N_VGND_c_253_n 0.0220624f $X=-0.19 $Y=-0.24 $X2=0.232 $Y2=1.325
cc_21 VNB N_VGND_c_254_n 0.162389f $X=-0.19 $Y=-0.24 $X2=0.232 $Y2=1.53
cc_22 VPB N_A_M1000_g 0.0457983f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=2.065
cc_23 VPB A 0.0266413f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_24 VPB A 9.15659e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_25 VPB N_A_c_49_n 0.0110863f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_26 VPB N_A_c_50_n 7.73127e-19 $X=-0.19 $Y=1.305 $X2=0.232 $Y2=1.325
cc_27 VPB N_SLEEP_B_M1005_g 0.0392126f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=2.065
cc_28 VPB SLEEP_B 0.00213477f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_29 VPB N_SLEEP_B_c_83_n 0.00641101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A_59_75#_M1001_g 0.0241244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_59_75#_c_124_n 0.00405675f $X=-0.19 $Y=1.305 $X2=0.232 $Y2=1.53
cc_32 VPB N_A_59_75#_c_125_n 0.00331457f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.2
cc_33 VPB N_A_59_75#_c_126_n 0.00575937f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.2
cc_34 VPB N_A_59_75#_c_120_n 0.00339207f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.2
cc_35 VPB N_A_59_75#_c_128_n 0.00178053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_59_75#_c_121_n 0.00679043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_194_n 0.0282531f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_38 VPB N_VPWR_c_195_n 0.00485351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_196_n 0.0112126f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.16
cc_40 VPB N_VPWR_c_197_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.16
cc_41 VPB N_VPWR_c_198_n 0.0192479f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_42 VPB N_VPWR_c_199_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_200_n 0.0201769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_193_n 0.062916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB X 0.0257284f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_46 VPB X 0.0228396f $X=-0.19 $Y=1.305 $X2=0.455 $Y2=1.16
cc_47 N_A_M1004_g N_SLEEP_B_M1002_g 0.0281599f $X=0.65 $Y=0.585 $X2=0 $Y2=0
cc_48 N_A_M1000_g N_SLEEP_B_M1005_g 0.0281599f $X=0.65 $Y=2.065 $X2=0 $Y2=0
cc_49 A SLEEP_B 0.0172688f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A_c_49_n SLEEP_B 2.90338e-19 $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_51 A N_SLEEP_B_c_83_n 0.00172917f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_52 N_A_c_49_n N_SLEEP_B_c_83_n 0.0281599f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_M1004_g N_A_59_75#_c_117_n 0.00778418f $X=0.65 $Y=0.585 $X2=0 $Y2=0
cc_54 N_A_M1004_g N_A_59_75#_c_118_n 0.00817062f $X=0.65 $Y=0.585 $X2=0 $Y2=0
cc_55 A N_A_59_75#_c_118_n 0.011624f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_M1004_g N_A_59_75#_c_119_n 0.00507008f $X=0.65 $Y=0.585 $X2=0 $Y2=0
cc_57 A N_A_59_75#_c_119_n 0.0201127f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_49_n N_A_59_75#_c_119_n 0.00725535f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_c_50_n N_A_59_75#_c_119_n 0.00698309f $X=0.232 $Y=1.325 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_A_59_75#_c_124_n 0.0035497f $X=0.65 $Y=2.065 $X2=0 $Y2=0
cc_61 N_A_M1000_g N_A_59_75#_c_126_n 0.00342053f $X=0.65 $Y=2.065 $X2=0 $Y2=0
cc_62 A N_A_59_75#_c_126_n 0.00556272f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_63 A N_A_59_75#_c_126_n 0.00266042f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_VPWR_c_194_n 0.0038689f $X=0.65 $Y=2.065 $X2=0 $Y2=0
cc_65 A N_VPWR_c_194_n 0.00497766f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_66 A N_VPWR_c_194_n 0.00489599f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_c_49_n N_VPWR_c_194_n 0.0034325f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_M1000_g N_VPWR_c_198_n 0.00523993f $X=0.65 $Y=2.065 $X2=0 $Y2=0
cc_69 N_A_M1000_g N_VPWR_c_193_n 0.00519019f $X=0.65 $Y=2.065 $X2=0 $Y2=0
cc_70 N_A_M1004_g N_VGND_c_251_n 0.00438605f $X=0.65 $Y=0.585 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_VGND_c_254_n 0.00541051f $X=0.65 $Y=0.585 $X2=0 $Y2=0
cc_72 N_SLEEP_B_M1005_g N_A_59_75#_M1001_g 0.0208544f $X=1.07 $Y=2.065 $X2=0
+ $Y2=0
cc_73 N_SLEEP_B_M1002_g N_A_59_75#_c_117_n 0.00144969f $X=1.07 $Y=0.585 $X2=0
+ $Y2=0
cc_74 N_SLEEP_B_M1002_g N_A_59_75#_c_118_n 0.0132517f $X=1.07 $Y=0.585 $X2=0
+ $Y2=0
cc_75 SLEEP_B N_A_59_75#_c_118_n 0.024687f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_76 N_SLEEP_B_c_83_n N_A_59_75#_c_118_n 0.004446f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_77 N_SLEEP_B_M1005_g N_A_59_75#_c_124_n 0.0105249f $X=1.07 $Y=2.065 $X2=0
+ $Y2=0
cc_78 N_SLEEP_B_M1005_g N_A_59_75#_c_125_n 0.0107487f $X=1.07 $Y=2.065 $X2=0
+ $Y2=0
cc_79 SLEEP_B N_A_59_75#_c_125_n 0.0159907f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_80 N_SLEEP_B_c_83_n N_A_59_75#_c_125_n 0.00117002f $X=1.16 $Y=1.16 $X2=0
+ $Y2=0
cc_81 N_SLEEP_B_M1005_g N_A_59_75#_c_126_n 0.00293143f $X=1.07 $Y=2.065 $X2=0
+ $Y2=0
cc_82 SLEEP_B N_A_59_75#_c_126_n 0.00225797f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_83 N_SLEEP_B_M1002_g N_A_59_75#_c_120_n 0.00156065f $X=1.07 $Y=0.585 $X2=0
+ $Y2=0
cc_84 SLEEP_B N_A_59_75#_c_120_n 0.0207523f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_85 N_SLEEP_B_c_83_n N_A_59_75#_c_120_n 0.00258311f $X=1.16 $Y=1.16 $X2=0
+ $Y2=0
cc_86 N_SLEEP_B_M1005_g N_A_59_75#_c_128_n 0.00302249f $X=1.07 $Y=2.065 $X2=0
+ $Y2=0
cc_87 SLEEP_B N_A_59_75#_c_121_n 7.6667e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_88 N_SLEEP_B_c_83_n N_A_59_75#_c_121_n 0.0212295f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_89 N_SLEEP_B_M1002_g N_A_59_75#_c_122_n 0.0169123f $X=1.07 $Y=0.585 $X2=0
+ $Y2=0
cc_90 N_SLEEP_B_M1005_g N_VPWR_c_195_n 0.00493973f $X=1.07 $Y=2.065 $X2=0 $Y2=0
cc_91 N_SLEEP_B_M1005_g N_VPWR_c_198_n 0.00486831f $X=1.07 $Y=2.065 $X2=0 $Y2=0
cc_92 N_SLEEP_B_M1005_g N_VPWR_c_193_n 0.00519019f $X=1.07 $Y=2.065 $X2=0 $Y2=0
cc_93 N_SLEEP_B_M1002_g N_VGND_c_250_n 0.00545678f $X=1.07 $Y=0.585 $X2=0 $Y2=0
cc_94 N_SLEEP_B_M1002_g N_VGND_c_251_n 0.0044865f $X=1.07 $Y=0.585 $X2=0 $Y2=0
cc_95 N_SLEEP_B_M1002_g N_VGND_c_254_n 0.00541051f $X=1.07 $Y=0.585 $X2=0 $Y2=0
cc_96 N_A_59_75#_c_125_n N_VPWR_M1005_d 0.00727495f $X=1.505 $Y=1.66 $X2=0 $Y2=0
cc_97 N_A_59_75#_c_124_n N_VPWR_c_194_n 0.00155022f $X=0.86 $Y=2.13 $X2=0 $Y2=0
cc_98 N_A_59_75#_M1001_g N_VPWR_c_195_n 0.0134748f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_59_75#_c_124_n N_VPWR_c_195_n 0.0258781f $X=0.86 $Y=2.13 $X2=0 $Y2=0
cc_100 N_A_59_75#_c_125_n N_VPWR_c_195_n 0.0221013f $X=1.505 $Y=1.66 $X2=0 $Y2=0
cc_101 N_A_59_75#_c_124_n N_VPWR_c_198_n 0.0101586f $X=0.86 $Y=2.13 $X2=0 $Y2=0
cc_102 N_A_59_75#_M1001_g N_VPWR_c_200_n 0.0046653f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_59_75#_M1001_g N_VPWR_c_193_n 0.00911899f $X=1.61 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_A_59_75#_c_124_n N_VPWR_c_193_n 0.0103862f $X=0.86 $Y=2.13 $X2=0 $Y2=0
cc_105 N_A_59_75#_c_120_n N_X_c_228_n 0.00473793f $X=1.59 $Y=1.325 $X2=0 $Y2=0
cc_106 N_A_59_75#_c_121_n N_X_c_228_n 0.00253834f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_59_75#_c_122_n N_X_c_228_n 0.00381469f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_59_75#_M1001_g X 0.0130173f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_59_75#_c_125_n X 0.00909028f $X=1.505 $Y=1.66 $X2=0 $Y2=0
cc_110 N_A_59_75#_c_120_n X 0.0403489f $X=1.59 $Y=1.325 $X2=0 $Y2=0
cc_111 N_A_59_75#_c_128_n X 0.0122276f $X=1.59 $Y=1.575 $X2=0 $Y2=0
cc_112 N_A_59_75#_c_121_n X 0.0081095f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_59_75#_c_122_n X 0.0100211f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_59_75#_M1001_g X 0.0124231f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_59_75#_c_120_n X 0.00119426f $X=1.59 $Y=1.325 $X2=0 $Y2=0
cc_116 N_A_59_75#_c_121_n X 0.00218271f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_59_75#_c_118_n A_145_75# 0.00297727f $X=1.505 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_59_75#_c_118_n N_VGND_M1002_d 0.0034258f $X=1.505 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_59_75#_c_117_n N_VGND_c_250_n 0.00521167f $X=0.44 $Y=0.52 $X2=0 $Y2=0
cc_120 N_A_59_75#_c_118_n N_VGND_c_250_n 0.0190303f $X=1.505 $Y=0.81 $X2=0 $Y2=0
cc_121 N_A_59_75#_c_122_n N_VGND_c_250_n 0.0044954f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_59_75#_c_117_n N_VGND_c_251_n 0.0140337f $X=0.44 $Y=0.52 $X2=0 $Y2=0
cc_123 N_A_59_75#_c_118_n N_VGND_c_251_n 0.00774346f $X=1.505 $Y=0.81 $X2=0
+ $Y2=0
cc_124 N_A_59_75#_c_120_n N_VGND_c_253_n 0.00204758f $X=1.59 $Y=1.325 $X2=0
+ $Y2=0
cc_125 N_A_59_75#_c_122_n N_VGND_c_253_n 0.00420655f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_59_75#_c_117_n N_VGND_c_254_n 0.0118489f $X=0.44 $Y=0.52 $X2=0 $Y2=0
cc_127 N_A_59_75#_c_118_n N_VGND_c_254_n 0.0178214f $X=1.505 $Y=0.81 $X2=0 $Y2=0
cc_128 N_A_59_75#_c_120_n N_VGND_c_254_n 0.00363577f $X=1.59 $Y=1.325 $X2=0
+ $Y2=0
cc_129 N_A_59_75#_c_122_n N_VGND_c_254_n 0.00813845f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_130 N_VPWR_c_193_n N_X_M1001_d 0.0063286f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_131 N_VPWR_c_195_n X 0.0402167f $X=1.4 $Y=2 $X2=0 $Y2=0
cc_132 N_VPWR_c_200_n X 0.0320555f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_133 N_VPWR_c_193_n X 0.0175942f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_134 N_X_c_228_n N_VGND_c_253_n 0.0185228f $X=1.965 $Y=0.4 $X2=0 $Y2=0
cc_135 N_X_c_225_n N_VGND_c_253_n 0.0179238f $X=2.09 $Y=0.545 $X2=0 $Y2=0
cc_136 N_X_M1003_d N_VGND_c_254_n 0.00225742f $X=1.685 $Y=0.235 $X2=0 $Y2=0
cc_137 N_X_c_228_n N_VGND_c_254_n 0.0114709f $X=1.965 $Y=0.4 $X2=0 $Y2=0
cc_138 N_X_c_225_n N_VGND_c_254_n 0.00962794f $X=2.09 $Y=0.545 $X2=0 $Y2=0

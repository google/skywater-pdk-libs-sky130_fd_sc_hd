* File: sky130_fd_sc_hd__einvn_4.spice.SKY130_FD_SC_HD__EINVN_4.pxi
* Created: Thu Aug 27 14:20:21 2020
* 
x_PM_SKY130_FD_SC_HD__EINVN_4%TE_B N_TE_B_c_89_n N_TE_B_M1015_g N_TE_B_M1011_g
+ N_TE_B_c_90_n N_TE_B_c_96_n N_TE_B_M1000_g N_TE_B_c_97_n N_TE_B_c_98_n
+ N_TE_B_M1001_g N_TE_B_c_99_n N_TE_B_c_100_n N_TE_B_M1005_g N_TE_B_c_101_n
+ N_TE_B_c_102_n N_TE_B_M1008_g N_TE_B_c_91_n N_TE_B_c_104_n N_TE_B_c_105_n TE_B
+ N_TE_B_c_93_n PM_SKY130_FD_SC_HD__EINVN_4%TE_B
x_PM_SKY130_FD_SC_HD__EINVN_4%A_27_47# N_A_27_47#_M1015_s N_A_27_47#_M1011_s
+ N_A_27_47#_c_168_n N_A_27_47#_M1002_g N_A_27_47#_c_169_n N_A_27_47#_c_170_n
+ N_A_27_47#_c_171_n N_A_27_47#_M1003_g N_A_27_47#_c_172_n N_A_27_47#_c_173_n
+ N_A_27_47#_M1006_g N_A_27_47#_c_174_n N_A_27_47#_c_175_n N_A_27_47#_M1010_g
+ N_A_27_47#_c_176_n N_A_27_47#_c_177_n N_A_27_47#_c_178_n N_A_27_47#_c_183_n
+ N_A_27_47#_c_179_n N_A_27_47#_c_180_n N_A_27_47#_c_184_n N_A_27_47#_c_181_n
+ N_A_27_47#_c_209_n N_A_27_47#_c_182_n PM_SKY130_FD_SC_HD__EINVN_4%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVN_4%A N_A_c_270_n N_A_M1013_g N_A_M1004_g N_A_c_271_n
+ N_A_M1014_g N_A_M1007_g N_A_c_272_n N_A_M1016_g N_A_M1009_g N_A_c_273_n
+ N_A_M1017_g N_A_M1012_g N_A_c_274_n A A N_A_c_276_n
+ PM_SKY130_FD_SC_HD__EINVN_4%A
x_PM_SKY130_FD_SC_HD__EINVN_4%VPWR N_VPWR_M1011_d N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n VPWR N_VPWR_c_343_n
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_339_n N_VPWR_c_348_n
+ N_VPWR_c_349_n N_VPWR_c_350_n PM_SKY130_FD_SC_HD__EINVN_4%VPWR
x_PM_SKY130_FD_SC_HD__EINVN_4%A_204_309# N_A_204_309#_M1000_s
+ N_A_204_309#_M1005_s N_A_204_309#_M1004_s N_A_204_309#_M1007_s
+ N_A_204_309#_M1012_s N_A_204_309#_c_415_n N_A_204_309#_c_408_n
+ N_A_204_309#_c_409_n N_A_204_309#_c_450_n N_A_204_309#_c_410_n
+ N_A_204_309#_c_423_n N_A_204_309#_c_434_n N_A_204_309#_c_411_n
+ N_A_204_309#_c_436_n N_A_204_309#_c_412_n N_A_204_309#_c_413_n
+ N_A_204_309#_c_414_n N_A_204_309#_c_462_n
+ PM_SKY130_FD_SC_HD__EINVN_4%A_204_309#
x_PM_SKY130_FD_SC_HD__EINVN_4%Z N_Z_M1013_d N_Z_M1016_d N_Z_M1004_d N_Z_M1009_d
+ N_Z_c_469_n N_Z_c_470_n Z Z N_Z_c_471_n PM_SKY130_FD_SC_HD__EINVN_4%Z
x_PM_SKY130_FD_SC_HD__EINVN_4%VGND N_VGND_M1015_d N_VGND_M1002_s N_VGND_M1006_s
+ N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n VGND N_VGND_c_511_n
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n
+ N_VGND_c_517_n N_VGND_c_518_n PM_SKY130_FD_SC_HD__EINVN_4%VGND
x_PM_SKY130_FD_SC_HD__EINVN_4%A_215_47# N_A_215_47#_M1002_d N_A_215_47#_M1003_d
+ N_A_215_47#_M1010_d N_A_215_47#_M1014_s N_A_215_47#_M1017_s
+ N_A_215_47#_c_582_n N_A_215_47#_c_588_n N_A_215_47#_c_583_n
+ N_A_215_47#_c_630_n N_A_215_47#_c_594_n N_A_215_47#_c_613_n
+ N_A_215_47#_c_598_n N_A_215_47#_c_584_n N_A_215_47#_c_600_n
+ PM_SKY130_FD_SC_HD__EINVN_4%A_215_47#
cc_1 VNB N_TE_B_c_89_n 0.0250205f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_TE_B_c_90_n 0.0136319f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.25
cc_3 VNB N_TE_B_c_91_n 0.0100604f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.25
cc_4 VNB TE_B 0.0136135f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_TE_B_c_93_n 0.0362295f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_6 VNB N_A_27_47#_c_168_n 0.0175424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_169_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.47
cc_8 VNB N_A_27_47#_c_170_n 0.00831588f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=2.015
cc_9 VNB N_A_27_47#_c_171_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=2.015
cc_10 VNB N_A_27_47#_c_172_n 0.00891962f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.47
cc_11 VNB N_A_27_47#_c_173_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_12 VNB N_A_27_47#_c_174_n 0.00887388f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.47
cc_13 VNB N_A_27_47#_c_175_n 0.0146322f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=2.015
cc_14 VNB N_A_27_47#_c_176_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=1.47
cc_15 VNB N_A_27_47#_c_177_n 0.00473803f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=2.015
cc_16 VNB N_A_27_47#_c_178_n 0.0156779f $X=-0.19 $Y=-0.24 $X2=2.205 $Y2=2.015
cc_17 VNB N_A_27_47#_c_179_n 0.00951289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_180_n 0.0030044f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_19 VNB N_A_27_47#_c_181_n 0.0144552f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_20 VNB N_A_27_47#_c_182_n 0.0213729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_c_270_n 0.0162767f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_22 VNB N_A_c_271_n 0.0150503f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.25
cc_23 VNB N_A_c_272_n 0.0150503f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=1.47
cc_24 VNB N_A_c_273_n 0.0186926f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=2.015
cc_25 VNB N_A_c_274_n 0.0605328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB A 0.0304598f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_27 VNB N_A_c_276_n 0.0381416f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_28 VNB N_VPWR_c_339_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_508_n 0.00474451f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=2.015
cc_30 VNB N_VGND_c_509_n 3.18775e-19 $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_31 VNB N_VGND_c_510_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.47
cc_32 VNB N_VGND_c_511_n 0.014319f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.395
cc_33 VNB N_VGND_c_512_n 0.0150454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_513_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_514_n 0.0570164f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_515_n 0.265511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_516_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_517_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_518_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_215_47#_c_582_n 0.00496433f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_41 VNB N_A_215_47#_c_583_n 0.00198743f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.47
cc_42 VNB N_A_215_47#_c_584_n 0.012533f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_TE_B_M1011_g 0.0257066f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_44 VPB N_TE_B_c_90_n 0.00483829f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.25
cc_45 VPB N_TE_B_c_96_n 0.0144321f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.47
cc_46 VPB N_TE_B_c_97_n 0.013715f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.395
cc_47 VPB N_TE_B_c_98_n 0.0135568f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.47
cc_48 VPB N_TE_B_c_99_n 0.0088967f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=1.395
cc_49 VPB N_TE_B_c_100_n 0.013575f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.47
cc_50 VPB N_TE_B_c_101_n 0.0207809f $X=-0.19 $Y=1.305 $X2=2.13 $Y2=1.395
cc_51 VPB N_TE_B_c_102_n 0.0171184f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=1.47
cc_52 VPB N_TE_B_c_91_n 0.00578605f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.25
cc_53 VPB N_TE_B_c_104_n 0.00473803f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.395
cc_54 VPB N_TE_B_c_105_n 0.00391059f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.395
cc_55 VPB TE_B 0.00311688f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_56 VPB N_TE_B_c_93_n 0.00941639f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_57 VPB N_A_27_47#_c_183_n 0.0308842f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.395
cc_58 VPB N_A_27_47#_c_184_n 0.00992248f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_59 VPB N_A_27_47#_c_181_n 0.00452491f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_60 VPB N_A_27_47#_c_182_n 0.00828812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_M1004_g 0.0252376f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_62 VPB N_A_M1007_g 0.0171014f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.395
cc_63 VPB N_A_M1009_g 0.0171014f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.47
cc_64 VPB N_A_M1012_g 0.0252376f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=2.015
cc_65 VPB N_A_c_274_n 0.0111069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB A 0.00614372f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_67 VPB N_A_c_276_n 0.0162504f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_68 VPB N_VPWR_c_340_n 0.00210688f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=2.015
cc_69 VPB N_VPWR_c_341_n 3.11529e-19 $X=-0.19 $Y=1.305 $X2=1.365 $Y2=2.015
cc_70 VPB N_VPWR_c_342_n 0.0108326f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.47
cc_71 VPB N_VPWR_c_343_n 0.0150576f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=1.395
cc_72 VPB N_VPWR_c_344_n 0.0146397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_345_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_346_n 0.0582824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_339_n 0.0523552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_348_n 0.0050755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_349_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_350_n 0.00623291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_204_309#_c_408_n 0.00251378f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.47
cc_80 VPB N_A_204_309#_c_409_n 0.0017513f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=2.015
cc_81 VPB N_A_204_309#_c_410_n 0.0122803f $X=-0.19 $Y=1.305 $X2=2.205 $Y2=2.015
cc_82 VPB N_A_204_309#_c_411_n 0.00126293f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_83 VPB N_A_204_309#_c_412_n 0.0101051f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_204_309#_c_413_n 0.0324936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_204_309#_c_414_n 0.00108194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_Z_c_469_n 6.87213e-19 $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.47
cc_87 VPB N_Z_c_470_n 6.87213e-19 $X=-0.19 $Y=1.305 $X2=1.44 $Y2=1.395
cc_88 VPB N_Z_c_471_n 0.00727359f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_89 N_TE_B_c_99_n N_A_27_47#_c_169_n 0.0153404f $X=1.71 $Y=1.395 $X2=0 $Y2=0
cc_90 N_TE_B_c_104_n N_A_27_47#_c_170_n 0.0153404f $X=1.365 $Y=1.395 $X2=0 $Y2=0
cc_91 N_TE_B_c_101_n N_A_27_47#_c_172_n 0.0153404f $X=2.13 $Y=1.395 $X2=0 $Y2=0
cc_92 N_TE_B_c_105_n N_A_27_47#_c_176_n 0.0153404f $X=1.785 $Y=1.395 $X2=0 $Y2=0
cc_93 N_TE_B_c_89_n N_A_27_47#_c_179_n 0.0138591f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_94 N_TE_B_c_90_n N_A_27_47#_c_179_n 9.15163e-19 $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_95 TE_B N_A_27_47#_c_179_n 0.0190911f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_96 N_TE_B_c_93_n N_A_27_47#_c_179_n 0.00163649f $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_97 N_TE_B_c_89_n N_A_27_47#_c_180_n 0.0108991f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_98 N_TE_B_M1011_g N_A_27_47#_c_184_n 0.0254636f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_99 N_TE_B_c_90_n N_A_27_47#_c_184_n 7.21838e-19 $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_100 N_TE_B_c_96_n N_A_27_47#_c_184_n 0.00105498f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_101 N_TE_B_c_91_n N_A_27_47#_c_184_n 0.00517984f $X=0.945 $Y=1.25 $X2=0 $Y2=0
cc_102 TE_B N_A_27_47#_c_184_n 0.0190911f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_103 N_TE_B_c_93_n N_A_27_47#_c_184_n 0.00163649f $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_104 N_TE_B_c_90_n N_A_27_47#_c_181_n 0.00183428f $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_105 N_TE_B_c_97_n N_A_27_47#_c_181_n 0.00881838f $X=1.29 $Y=1.395 $X2=0 $Y2=0
cc_106 N_TE_B_c_99_n N_A_27_47#_c_181_n 0.0058575f $X=1.71 $Y=1.395 $X2=0 $Y2=0
cc_107 N_TE_B_c_101_n N_A_27_47#_c_181_n 0.00936175f $X=2.13 $Y=1.395 $X2=0
+ $Y2=0
cc_108 N_TE_B_c_91_n N_A_27_47#_c_181_n 0.0154391f $X=0.945 $Y=1.25 $X2=0 $Y2=0
cc_109 N_TE_B_c_104_n N_A_27_47#_c_181_n 0.00405558f $X=1.365 $Y=1.395 $X2=0
+ $Y2=0
cc_110 N_TE_B_c_105_n N_A_27_47#_c_181_n 0.00354669f $X=1.785 $Y=1.395 $X2=0
+ $Y2=0
cc_111 N_TE_B_c_90_n N_A_27_47#_c_209_n 0.0130163f $X=0.87 $Y=1.25 $X2=0 $Y2=0
cc_112 TE_B N_A_27_47#_c_209_n 0.0258959f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_113 N_TE_B_c_93_n N_A_27_47#_c_209_n 0.0101792f $X=0.545 $Y=1.16 $X2=0 $Y2=0
cc_114 N_TE_B_c_101_n N_A_27_47#_c_182_n 3.38171e-19 $X=2.13 $Y=1.395 $X2=0
+ $Y2=0
cc_115 N_TE_B_M1011_g N_VPWR_c_340_n 0.0129471f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_116 N_TE_B_c_96_n N_VPWR_c_340_n 0.0016047f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_117 N_TE_B_c_96_n N_VPWR_c_341_n 7.4754e-19 $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_118 N_TE_B_c_98_n N_VPWR_c_341_n 0.0111574f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_119 N_TE_B_c_100_n N_VPWR_c_341_n 0.0110282f $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_120 N_TE_B_c_102_n N_VPWR_c_341_n 6.72101e-19 $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_121 N_TE_B_c_100_n N_VPWR_c_342_n 6.75043e-19 $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_122 N_TE_B_c_102_n N_VPWR_c_342_n 0.0122412f $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_123 N_TE_B_M1011_g N_VPWR_c_343_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_124 N_TE_B_c_96_n N_VPWR_c_344_n 0.00579312f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_125 N_TE_B_c_98_n N_VPWR_c_344_n 0.0046653f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_126 N_TE_B_c_100_n N_VPWR_c_345_n 0.0046653f $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_127 N_TE_B_c_102_n N_VPWR_c_345_n 0.0046653f $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_128 N_TE_B_M1011_g N_VPWR_c_339_n 0.00895857f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_129 N_TE_B_c_96_n N_VPWR_c_339_n 0.010505f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_130 N_TE_B_c_98_n N_VPWR_c_339_n 0.00796766f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_131 N_TE_B_c_100_n N_VPWR_c_339_n 0.00796766f $X=1.785 $Y=1.47 $X2=0 $Y2=0
cc_132 N_TE_B_c_102_n N_VPWR_c_339_n 0.00796766f $X=2.205 $Y=1.47 $X2=0 $Y2=0
cc_133 N_TE_B_M1011_g N_A_204_309#_c_415_n 4.91309e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_TE_B_c_96_n N_A_204_309#_c_415_n 0.00967786f $X=0.945 $Y=1.47 $X2=0
+ $Y2=0
cc_135 N_TE_B_c_98_n N_A_204_309#_c_408_n 0.0134056f $X=1.365 $Y=1.47 $X2=0
+ $Y2=0
cc_136 N_TE_B_c_99_n N_A_204_309#_c_408_n 0.0020486f $X=1.71 $Y=1.395 $X2=0
+ $Y2=0
cc_137 N_TE_B_c_100_n N_A_204_309#_c_408_n 0.0133633f $X=1.785 $Y=1.47 $X2=0
+ $Y2=0
cc_138 N_TE_B_c_96_n N_A_204_309#_c_409_n 0.00301378f $X=0.945 $Y=1.47 $X2=0
+ $Y2=0
cc_139 N_TE_B_c_97_n N_A_204_309#_c_409_n 0.00215435f $X=1.29 $Y=1.395 $X2=0
+ $Y2=0
cc_140 N_TE_B_c_102_n N_A_204_309#_c_410_n 0.0154663f $X=2.205 $Y=1.47 $X2=0
+ $Y2=0
cc_141 N_TE_B_c_102_n N_A_204_309#_c_423_n 0.00373536f $X=2.205 $Y=1.47 $X2=0
+ $Y2=0
cc_142 N_TE_B_c_101_n N_A_204_309#_c_414_n 0.00215435f $X=2.13 $Y=1.395 $X2=0
+ $Y2=0
cc_143 N_TE_B_c_89_n N_VGND_c_508_n 0.00966951f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_144 N_TE_B_c_89_n N_VGND_c_511_n 0.00341689f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_145 N_TE_B_c_89_n N_VGND_c_515_n 0.0050171f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_146 N_TE_B_c_89_n N_A_215_47#_c_582_n 0.00178374f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_TE_B_c_89_n N_A_215_47#_c_583_n 7.04009e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_TE_B_c_97_n N_A_215_47#_c_583_n 0.00101297f $X=1.29 $Y=1.395 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_175_n N_A_c_270_n 0.0189878f $X=2.67 $Y=0.96 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_27_47#_c_181_n N_A_c_274_n 0.00345774f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_182_n N_A_c_274_n 0.012916f $X=2.625 $Y=1.035 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_184_n N_VPWR_M1011_d 0.00404069f $X=0.68 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_27_47#_c_184_n N_VPWR_c_340_n 0.0193336f $X=0.68 $Y=1.495 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_183_n N_VPWR_c_343_n 0.018001f $X=0.26 $Y=1.815 $X2=0 $Y2=0
cc_155 N_A_27_47#_M1011_s N_VPWR_c_339_n 0.00387172f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_183_n N_VPWR_c_339_n 0.00993603f $X=0.26 $Y=1.815 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_170_n N_A_204_309#_c_408_n 4.28192e-19 $X=1.485 $Y=1.035
+ $X2=0 $Y2=0
cc_158 N_A_27_47#_c_181_n N_A_204_309#_c_408_n 0.0490093f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_184_n N_A_204_309#_c_409_n 0.0093578f $X=0.68 $Y=1.495 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_181_n N_A_204_309#_c_409_n 0.0189161f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_177_n N_A_204_309#_c_410_n 8.9107e-19 $X=2.25 $Y=1.035 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_181_n N_A_204_309#_c_410_n 0.0731545f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_182_n N_A_204_309#_c_410_n 0.00700619f $X=2.625 $Y=1.035
+ $X2=0 $Y2=0
cc_164 N_A_27_47#_c_172_n N_A_204_309#_c_414_n 2.23657e-19 $X=2.175 $Y=1.035
+ $X2=0 $Y2=0
cc_165 N_A_27_47#_c_181_n N_A_204_309#_c_414_n 0.0143368f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_175_n N_Z_c_471_n 9.25498e-19 $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_181_n N_Z_c_471_n 0.0292385f $X=2.625 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_182_n N_Z_c_471_n 2.34249e-19 $X=2.625 $Y=1.035 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_179_n N_VGND_M1015_d 0.00334969f $X=0.68 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_27_47#_c_180_n N_VGND_M1015_d 8.61564e-19 $X=0.68 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A_27_47#_c_168_n N_VGND_c_508_n 0.00195572f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_179_n N_VGND_c_508_n 0.0207342f $X=0.68 $Y=0.825 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_168_n N_VGND_c_509_n 0.00725083f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_171_n N_VGND_c_509_n 0.00685342f $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_173_n N_VGND_c_509_n 5.54209e-19 $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_171_n N_VGND_c_510_n 5.54209e-19 $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_173_n N_VGND_c_510_n 0.00685342f $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_175_n N_VGND_c_510_n 0.00823169f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_178_n N_VGND_c_511_n 0.0173297f $X=0.215 $Y=0.655 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_179_n N_VGND_c_511_n 0.00235077f $X=0.68 $Y=0.825 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_168_n N_VGND_c_512_n 0.00341689f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_171_n N_VGND_c_513_n 0.00341689f $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_173_n N_VGND_c_513_n 0.00341689f $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_175_n N_VGND_c_514_n 0.00341689f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1015_s N_VGND_c_515_n 0.00230206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_168_n N_VGND_c_515_n 0.00540327f $X=1.41 $Y=0.96 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_171_n N_VGND_c_515_n 0.0040262f $X=1.83 $Y=0.96 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_173_n N_VGND_c_515_n 0.0040262f $X=2.25 $Y=0.96 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_175_n N_VGND_c_515_n 0.00418888f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_178_n N_VGND_c_515_n 0.00980382f $X=0.215 $Y=0.655 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_179_n N_VGND_c_515_n 0.00561963f $X=0.68 $Y=0.825 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_168_n N_A_215_47#_c_588_n 0.0108561f $X=1.41 $Y=0.96 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_169_n N_A_215_47#_c_588_n 0.00179137f $X=1.755 $Y=1.035
+ $X2=0 $Y2=0
cc_194 N_A_27_47#_c_171_n N_A_215_47#_c_588_n 0.010245f $X=1.83 $Y=0.96 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_181_n N_A_215_47#_c_588_n 0.0410653f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_179_n N_A_215_47#_c_583_n 0.0157409f $X=0.68 $Y=0.825 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_181_n N_A_215_47#_c_583_n 0.0228911f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_173_n N_A_215_47#_c_594_n 0.0102303f $X=2.25 $Y=0.96 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_174_n N_A_215_47#_c_594_n 0.00183302f $X=2.49 $Y=1.035 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_175_n N_A_215_47#_c_594_n 0.0102733f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_181_n N_A_215_47#_c_594_n 0.057592f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_175_n N_A_215_47#_c_598_n 0.00133088f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_181_n N_A_215_47#_c_584_n 7.29254e-19 $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_172_n N_A_215_47#_c_600_n 0.00186022f $X=2.175 $Y=1.035
+ $X2=0 $Y2=0
cc_205 N_A_27_47#_c_181_n N_A_215_47#_c_600_n 0.0132296f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_206 N_A_M1004_g N_VPWR_c_342_n 0.00345994f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_M1004_g N_VPWR_c_346_n 0.00357877f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_M1007_g N_VPWR_c_346_n 0.00357877f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_M1009_g N_VPWR_c_346_n 0.00357877f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_M1012_g N_VPWR_c_346_n 0.00357877f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_M1004_g N_VPWR_c_339_n 0.00664112f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_M1007_g N_VPWR_c_339_n 0.00526405f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A_M1009_g N_VPWR_c_339_n 0.00526405f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_M1012_g N_VPWR_c_339_n 0.00639647f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_M1004_g N_A_204_309#_c_434_n 0.0135411f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_M1007_g N_A_204_309#_c_434_n 0.0126401f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_c_274_n N_A_204_309#_c_436_n 4.9277e-19 $X=4.48 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_M1009_g N_A_204_309#_c_412_n 0.0126843f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_M1012_g N_A_204_309#_c_412_n 0.0138832f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_220 A N_A_204_309#_c_413_n 0.0238853f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_221 N_A_c_276_n N_A_204_309#_c_413_n 0.00306997f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_M1004_g N_Z_c_469_n 0.00757723f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_M1007_g N_Z_c_469_n 0.00793926f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_M1009_g N_Z_c_469_n 5.59859e-19 $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_c_274_n N_Z_c_469_n 4.65424e-19 $X=4.48 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_M1007_g N_Z_c_470_n 5.59859e-19 $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_M1009_g N_Z_c_470_n 0.00793926f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_M1012_g N_Z_c_470_n 0.012658f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A_c_274_n N_Z_c_470_n 4.65424e-19 $X=4.48 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_c_270_n N_Z_c_471_n 0.00745389f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_M1004_g N_Z_c_471_n 0.00914036f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A_c_271_n N_Z_c_471_n 0.012949f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_M1007_g N_Z_c_471_n 0.0120754f $X=3.565 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_c_272_n N_Z_c_471_n 0.012949f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_M1009_g N_Z_c_471_n 0.0120754f $X=3.985 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A_c_273_n N_Z_c_471_n 0.00579339f $X=4.405 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_M1012_g N_Z_c_471_n 0.00914036f $X=4.405 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A_c_274_n N_Z_c_471_n 0.0541223f $X=4.48 $Y=1.16 $X2=0 $Y2=0
cc_239 A N_Z_c_471_n 0.0474012f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_240 N_A_c_270_n N_VGND_c_510_n 0.0011729f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_c_270_n N_VGND_c_514_n 0.00357877f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_271_n N_VGND_c_514_n 0.00357877f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_272_n N_VGND_c_514_n 0.00357877f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_c_273_n N_VGND_c_514_n 0.00357877f $X=4.405 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_c_270_n N_VGND_c_515_n 0.00542674f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_c_271_n N_VGND_c_515_n 0.00522516f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_c_272_n N_VGND_c_515_n 0.00522516f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_c_273_n N_VGND_c_515_n 0.00631565f $X=4.405 $Y=0.995 $X2=0 $Y2=0
cc_249 A N_A_215_47#_M1017_s 0.00469049f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_250 N_A_c_270_n N_A_215_47#_c_594_n 0.00103287f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_270_n N_A_215_47#_c_584_n 0.0131453f $X=3.145 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_c_271_n N_A_215_47#_c_584_n 0.00822564f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_c_272_n N_A_215_47#_c_584_n 0.00827637f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_c_273_n N_A_215_47#_c_584_n 0.0119853f $X=4.405 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_c_274_n N_A_215_47#_c_584_n 8.77588e-19 $X=4.48 $Y=1.16 $X2=0 $Y2=0
cc_256 A N_A_215_47#_c_584_n 0.0345321f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_257 N_A_c_276_n N_A_215_47#_c_584_n 0.00136866f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_258 N_VPWR_c_339_n N_A_204_309#_M1000_s 0.00393857f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_259 N_VPWR_c_339_n N_A_204_309#_M1005_s 0.00570907f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_339_n N_A_204_309#_M1004_s 0.00210127f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_339_n N_A_204_309#_M1007_s 0.00216817f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_339_n N_A_204_309#_M1012_s 0.00210127f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_344_n N_A_204_309#_c_415_n 0.0134781f $X=1.41 $Y=2.72 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_339_n N_A_204_309#_c_415_n 0.00856983f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_265 N_VPWR_M1001_d N_A_204_309#_c_408_n 0.00165831f $X=1.44 $Y=1.545 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_341_n N_A_204_309#_c_408_n 0.0170258f $X=1.575 $Y=2.02 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_345_n N_A_204_309#_c_450_n 0.0113958f $X=2.25 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_339_n N_A_204_309#_c_450_n 0.00646998f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_VPWR_M1008_d N_A_204_309#_c_410_n 0.00268486f $X=2.28 $Y=1.545 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_342_n N_A_204_309#_c_410_n 0.0270443f $X=2.415 $Y=2 $X2=0 $Y2=0
cc_271 N_VPWR_c_342_n N_A_204_309#_c_423_n 0.0368471f $X=2.415 $Y=2 $X2=0 $Y2=0
cc_272 N_VPWR_c_346_n N_A_204_309#_c_434_n 0.0358916f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_339_n N_A_204_309#_c_434_n 0.0235822f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_342_n N_A_204_309#_c_411_n 0.014919f $X=2.415 $Y=2 $X2=0 $Y2=0
cc_275 N_VPWR_c_346_n N_A_204_309#_c_411_n 0.0145235f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_339_n N_A_204_309#_c_411_n 0.00808747f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_346_n N_A_204_309#_c_412_n 0.0672272f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_339_n N_A_204_309#_c_412_n 0.0407095f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_346_n N_A_204_309#_c_462_n 0.0114668f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_339_n N_A_204_309#_c_462_n 0.006547f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_339_n N_Z_M1004_d 0.00216833f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_339_n N_Z_M1009_d 0.00216833f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_283 N_A_204_309#_c_434_n N_Z_M1004_d 0.00332127f $X=3.69 $Y=2.38 $X2=0 $Y2=0
cc_284 N_A_204_309#_c_412_n N_Z_M1009_d 0.00332127f $X=4.53 $Y=2.38 $X2=0 $Y2=0
cc_285 N_A_204_309#_c_434_n N_Z_c_469_n 0.0126022f $X=3.69 $Y=2.38 $X2=0 $Y2=0
cc_286 N_A_204_309#_c_412_n N_Z_c_470_n 0.0126022f $X=4.53 $Y=2.38 $X2=0 $Y2=0
cc_287 N_A_204_309#_c_436_n N_Z_c_471_n 0.0148392f $X=3.775 $Y=1.815 $X2=0 $Y2=0
cc_288 N_Z_M1013_d N_VGND_c_515_n 0.00216833f $X=3.22 $Y=0.235 $X2=0 $Y2=0
cc_289 N_Z_M1016_d N_VGND_c_515_n 0.00216833f $X=4.06 $Y=0.235 $X2=0 $Y2=0
cc_290 N_Z_c_471_n N_A_215_47#_M1014_s 0.00166399f $X=4.195 $Y=0.74 $X2=0 $Y2=0
cc_291 N_Z_c_471_n N_A_215_47#_c_594_n 0.0133517f $X=4.195 $Y=0.74 $X2=0 $Y2=0
cc_292 N_Z_c_471_n N_A_215_47#_c_613_n 0.0023689f $X=4.195 $Y=0.74 $X2=0 $Y2=0
cc_293 N_Z_M1013_d N_A_215_47#_c_584_n 0.00304533f $X=3.22 $Y=0.235 $X2=0 $Y2=0
cc_294 N_Z_M1016_d N_A_215_47#_c_584_n 0.00304533f $X=4.06 $Y=0.235 $X2=0 $Y2=0
cc_295 N_Z_c_471_n N_A_215_47#_c_584_n 0.0617386f $X=4.195 $Y=0.74 $X2=0 $Y2=0
cc_296 N_VGND_c_515_n N_A_215_47#_M1002_d 0.00229009f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_297 N_VGND_c_515_n N_A_215_47#_M1003_d 0.00254582f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_298 N_VGND_c_515_n N_A_215_47#_M1010_d 0.00292483f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_299 N_VGND_c_515_n N_A_215_47#_M1014_s 0.00215227f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_300 N_VGND_c_515_n N_A_215_47#_M1017_s 0.00225742f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_c_508_n N_A_215_47#_c_582_n 0.0188652f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_302 N_VGND_c_512_n N_A_215_47#_c_582_n 0.0184794f $X=1.455 $Y=0 $X2=0 $Y2=0
cc_303 N_VGND_c_515_n N_A_215_47#_c_582_n 0.0102739f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_M1002_s N_A_215_47#_c_588_n 0.00297022f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_305 N_VGND_c_509_n N_A_215_47#_c_588_n 0.0160613f $X=1.62 $Y=0.36 $X2=0 $Y2=0
cc_306 N_VGND_c_512_n N_A_215_47#_c_588_n 0.00232396f $X=1.455 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_513_n N_A_215_47#_c_588_n 0.00232396f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_308 N_VGND_c_515_n N_A_215_47#_c_588_n 0.00970544f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_513_n N_A_215_47#_c_630_n 0.0112554f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_515_n N_A_215_47#_c_630_n 0.00644035f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_M1006_s N_A_215_47#_c_594_n 0.00304947f $X=2.325 $Y=0.235 $X2=0
+ $Y2=0
cc_312 N_VGND_c_510_n N_A_215_47#_c_594_n 0.0160613f $X=2.46 $Y=0.36 $X2=0 $Y2=0
cc_313 N_VGND_c_513_n N_A_215_47#_c_594_n 0.00232396f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_514_n N_A_215_47#_c_594_n 0.00276686f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_515_n N_A_215_47#_c_594_n 0.0105423f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_510_n N_A_215_47#_c_613_n 0.00224761f $X=2.46 $Y=0.36 $X2=0
+ $Y2=0
cc_317 N_VGND_c_510_n N_A_215_47#_c_598_n 0.0142026f $X=2.46 $Y=0.36 $X2=0 $Y2=0
cc_318 N_VGND_c_514_n N_A_215_47#_c_598_n 0.0118015f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_515_n N_A_215_47#_c_598_n 0.00651702f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_514_n N_A_215_47#_c_584_n 0.112563f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_515_n N_A_215_47#_c_584_n 0.0710168f $X=4.83 $Y=0 $X2=0 $Y2=0

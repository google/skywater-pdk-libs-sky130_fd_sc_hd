* File: sky130_fd_sc_hd__or3_2.pex.spice
* Created: Tue Sep  1 19:27:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR3_2%C 3 7 9 15
r26 12 15 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.255 $Y=1.16
+ $X2=0.485 $Y2=1.16
r27 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r28 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.16
r29 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.695
r30 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.16
r31 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_2%B 4 7 8 9 10 11 15 16
r42 15 17 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.905 $Y=2.28
+ $X2=0.905 $Y2=2.145
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=2.28 $X2=0.905 $Y2=2.28
r44 11 16 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=0.69 $Y=2.27
+ $X2=0.905 $Y2=2.27
r45 10 11 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.23 $Y=2.27
+ $X2=0.69 $Y2=2.27
r46 8 9 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=0.875 $Y=0.76
+ $X2=0.875 $Y2=0.91
r47 7 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.905 $Y=0.475
+ $X2=0.905 $Y2=0.76
r48 4 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.845 $Y=1.695
+ $X2=0.845 $Y2=2.145
r49 4 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.845 $Y=1.695
+ $X2=0.845 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_2%A 3 7 9 10 11 16 17 20
c52 20 0 1.18156e-19 $X=0.717 $Y=1.325
r53 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.31 $Y2=1.325
r54 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.31 $Y2=0.995
r55 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.16 $X2=1.31 $Y2=1.16
r56 11 17 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.31
+ $Y2=1.16
r57 11 24 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=0.83 $Y2=1.16
r58 10 20 10.5 $w=2.23e-07 $l=2.05e-07 $layer=LI1_cond $X=0.717 $Y=1.53
+ $X2=0.717 $Y2=1.325
r59 9 20 4.237 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=0.717 $Y=1.16
+ $X2=0.717 $Y2=1.325
r60 9 24 2.9017 $w=3.3e-07 $l=1.13e-07 $layer=LI1_cond $X=0.717 $Y=1.16 $X2=0.83
+ $Y2=1.16
r61 7 19 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.325 $Y=1.695
+ $X2=1.325 $Y2=1.325
r62 3 18 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.325 $Y=0.475
+ $X2=1.325 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_2%A_30_53# 1 2 3 10 12 15 17 19 22 26 28 29 30
+ 34 36 38 43 45 49 50 55 57 62
c110 55 0 1.14153e-19 $X=1.79 $Y=1.16
c111 43 0 1.06604e-19 $X=1.685 $Y=1.495
c112 36 0 2.93657e-20 $X=1.6 $Y=0.74
r113 61 62 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.815 $Y=1.16
+ $X2=2.235 $Y2=1.16
r114 56 61 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.79 $Y=1.16
+ $X2=1.815 $Y2=1.16
r115 55 58 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.737 $Y=1.16
+ $X2=1.737 $Y2=1.325
r116 55 57 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.737 $Y=1.16
+ $X2=1.737 $Y2=0.995
r117 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.16 $X2=1.79 $Y2=1.16
r118 50 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.185 $Y=1.58
+ $X2=1.185 $Y2=1.87
r119 45 47 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.27 $Y=1.685
+ $X2=0.27 $Y2=1.87
r120 43 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.685 $Y=1.495
+ $X2=1.685 $Y2=1.325
r121 40 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.685 $Y=0.825
+ $X2=1.685 $Y2=0.995
r122 39 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=1.58
+ $X2=1.185 $Y2=1.58
r123 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=1.58
+ $X2=1.685 $Y2=1.495
r124 38 39 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.6 $Y=1.58
+ $X2=1.27 $Y2=1.58
r125 37 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.74
+ $X2=1.115 $Y2=0.74
r126 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=0.74
+ $X2=1.685 $Y2=0.825
r127 36 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.6 $Y=0.74 $X2=1.2
+ $Y2=0.74
r128 32 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.655
+ $X2=1.115 $Y2=0.74
r129 32 34 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.115 $Y=0.655
+ $X2=1.115 $Y2=0.47
r130 31 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=1.87
+ $X2=0.27 $Y2=1.87
r131 30 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.87
+ $X2=1.185 $Y2=1.87
r132 30 31 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.1 $Y=1.87
+ $X2=0.435 $Y2=1.87
r133 28 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=0.74
+ $X2=1.115 $Y2=0.74
r134 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.03 $Y=0.74
+ $X2=0.36 $Y2=0.74
r135 24 29 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.232 $Y=0.655
+ $X2=0.36 $Y2=0.74
r136 24 26 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=0.232 $Y=0.655
+ $X2=0.232 $Y2=0.47
r137 20 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.325
+ $X2=2.235 $Y2=1.16
r138 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.235 $Y=1.325
+ $X2=2.235 $Y2=1.985
r139 17 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=0.995
+ $X2=2.235 $Y2=1.16
r140 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.235 $Y=0.995
+ $X2=2.235 $Y2=0.56
r141 13 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.16
r142 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.985
r143 10 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=1.16
r144 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=0.56
r145 3 45 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.485 $X2=0.275 $Y2=1.685
r146 2 34 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.265 $X2=1.115 $Y2=0.47
r147 1 26 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.265 $X2=0.275 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_2%VPWR 1 2 9 11 13 17 19 27 33 37
c33 1 0 1.06604e-19 $X=1.4 $Y=1.485
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r36 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r37 31 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r38 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 28 33 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.73 $Y=2.72 $X2=1.59
+ $Y2=2.72
r40 28 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.73 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 27 36 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.572 $Y2=2.72
r42 27 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r44 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r45 21 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 19 33 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.45 $Y=2.72 $X2=1.59
+ $Y2=2.72
r47 19 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.45 $Y=2.72 $X2=1.15
+ $Y2=2.72
r48 17 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 17 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r50 13 16 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=2.53 $Y=1.62
+ $X2=2.53 $Y2=2.3
r51 11 36 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.53 $Y=2.635
+ $X2=2.572 $Y2=2.72
r52 11 16 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.53 $Y=2.635
+ $X2=2.53 $Y2=2.3
r53 7 33 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.635
+ $X2=1.59 $Y2=2.72
r54 7 9 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.59 $Y=2.635
+ $X2=1.59 $Y2=2
r55 2 16 400 $w=1.7e-07 $l=8.91417e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=1.485 $X2=2.47 $Y2=2.3
r56 2 13 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=1.485 $X2=2.47 $Y2=1.62
r57 1 9 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=1.4
+ $Y=1.485 $X2=1.6 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_2%X 1 2 12 14 15 16
r25 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=2.077 $Y=1.632
+ $X2=2.077 $Y2=1.845
r26 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.077 $Y=1.632
+ $X2=2.077 $Y2=1.495
r27 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=2.025 $Y=0.587
+ $X2=2.13 $Y2=0.587
r28 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.13 $Y=0.76 $X2=2.13
+ $Y2=0.587
r29 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.13 $Y=0.76
+ $X2=2.13 $Y2=1.495
r30 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=1.485 $X2=2.025 $Y2=1.845
r31 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.235 $X2=2.025 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR3_2%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
c51 20 0 2.93657e-20 $X=2.47 $Y=0.4
r52 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r53 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r54 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r55 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r56 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r57 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r58 35 43 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.75 $Y=0 $X2=1.56
+ $Y2=0
r59 35 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.75 $Y=0 $X2=2.07
+ $Y2=0
r60 34 46 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.572
+ $Y2=0
r61 34 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.07
+ $Y2=0
r62 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r63 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r64 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r65 30 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.695
+ $Y2=0
r66 30 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.15
+ $Y2=0
r67 29 43 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.56
+ $Y2=0
r68 29 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.15
+ $Y2=0
r69 24 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.695
+ $Y2=0
r70 24 26 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.23
+ $Y2=0
r71 22 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r72 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 18 46 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.572 $Y2=0
r74 18 20 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0.4
r75 14 43 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=0.085
+ $X2=1.56 $Y2=0
r76 14 16 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.56 $Y=0.085
+ $X2=1.56 $Y2=0.4
r77 10 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r78 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.4
r79 3 20 91 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=2 $X=2.31
+ $Y=0.235 $X2=2.47 $Y2=0.4
r80 2 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.265 $X2=1.585 $Y2=0.4
r81 1 12 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.265 $X2=0.695 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__sdfstp_2.spice.pex
* Created: Thu Aug 27 14:46:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%SCD 1 2 3 5 6 8 11 13 14
r33 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r34 14 19 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.53
+ $X2=0.212 $Y2=1.16
r35 13 19 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.212 $Y=0.85
+ $X2=0.212 $Y2=1.16
r36 9 11 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.315 $Y=1.695
+ $X2=0.47 $Y2=1.695
r37 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=1.695
r38 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=2.165
r39 3 18 87.63 $w=2.63e-07 $l=4.97242e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.325 $Y2=1.16
r40 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r41 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.315 $Y=1.62
+ $X2=0.315 $Y2=1.695
r42 1 18 39.0634 $w=2.63e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.325 $Y2=1.16
r43 1 2 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.315 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%SCE 3 5 7 11 15 17 19 20 26 33 34
c108 26 0 1.07953e-19 $X=2.53 $Y=1.19
c109 7 0 1.86564e-19 $X=0.89 $Y=2.165
r110 33 36 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.557 $Y=1.16
+ $X2=2.557 $Y2=1.325
r111 33 35 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.557 $Y=1.16
+ $X2=2.557 $Y2=0.995
r112 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=1.16 $X2=2.535 $Y2=1.16
r113 26 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r114 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.19
+ $X2=0.69 $Y2=1.19
r115 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r116 19 20 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.835 $Y2=1.19
r117 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.735
+ $Y=1.25 $X2=0.735 $Y2=1.25
r118 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.19
+ $X2=0.69 $Y2=1.19
r119 15 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.64 $Y=0.445
+ $X2=2.64 $Y2=0.995
r120 11 36 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.61 $Y=2.165
+ $X2=2.61 $Y2=1.325
r121 5 30 38.6139 $w=3.32e-07 $l=2.12238e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.782 $Y2=1.25
r122 5 7 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.89 $Y2=2.165
r123 1 30 38.6139 $w=3.32e-07 $l=1.8747e-07 $layer=POLY_cond $X=0.83 $Y=1.085
+ $X2=0.782 $Y2=1.25
r124 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.83 $Y=1.085 $X2=0.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%D 1 3 6 8 9 13
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=0.93 $X2=1.25 $Y2=0.93
r42 9 14 24.262 $w=2.83e-07 $l=6e-07 $layer=LI1_cond $X=1.192 $Y=1.53 $X2=1.192
+ $Y2=0.93
r43 8 14 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=1.192 $Y=0.85 $X2=1.192
+ $Y2=0.93
r44 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.095
+ $X2=1.25 $Y2=0.93
r45 4 6 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.25 $Y=1.095 $X2=1.25
+ $Y2=2.165
r46 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=0.765
+ $X2=1.25 $Y2=0.93
r47 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.25 $Y=0.765 $X2=1.25
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_319_21# 1 2 9 13 16 20 21 22 24 34 36
c76 21 0 1.4475e-19 $X=1.95 $Y=1.16
r77 34 36 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=2.395 $Y=1.927
+ $X2=2.4 $Y2=1.927
r78 22 24 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=2.39 $Y=0.715
+ $X2=2.39 $Y2=0.44
r79 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.16 $X2=1.95 $Y2=1.16
r80 18 34 13.2805 $w=3.13e-07 $l=3.63e-07 $layer=LI1_cond $X=2.032 $Y=1.927
+ $X2=2.395 $Y2=1.927
r81 18 20 20.9848 $w=3.33e-07 $l=6.1e-07 $layer=LI1_cond $X=2.032 $Y=1.77
+ $X2=2.032 $Y2=1.16
r82 17 22 20.8976 $w=1.88e-07 $l=3.58e-07 $layer=LI1_cond $X=2.032 $Y=0.81
+ $X2=2.39 $Y2=0.81
r83 17 20 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.032 $Y=0.905
+ $X2=2.032 $Y2=1.16
r84 15 21 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.745 $Y=1.16
+ $X2=1.95 $Y2=1.16
r85 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.745 $Y=1.16
+ $X2=1.67 $Y2=1.16
r86 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.325
+ $X2=1.67 $Y2=1.16
r87 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.67 $Y=1.325
+ $X2=1.67 $Y2=2.165
r88 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=0.995
+ $X2=1.67 $Y2=1.16
r89 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.67 $Y=0.995 $X2=1.67
+ $Y2=0.445
r90 2 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.845 $X2=2.4 $Y2=1.99
r91 1 24 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.235 $X2=2.43 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%CLK 7 8 10 13 15 16 17 18 19 20 26 28
c73 20 0 1.05862e-19 $X=3.45 $Y=1.19
c74 15 0 7.67918e-20 $X=3.52 $Y=1.62
c75 13 0 1.07242e-19 $X=3.58 $Y=0.805
r76 41 42 0.14951 $w=5.58e-07 $l=7e-09 $layer=LI1_cond $X=2.995 $Y=1.335
+ $X2=3.002 $Y2=1.335
r77 34 41 7.51078 $w=1.8e-07 $l=2.8e-07 $layer=LI1_cond $X=2.995 $Y=1.615
+ $X2=2.995 $Y2=1.335
r78 30 42 7.01796 $w=1.95e-07 $l=2.8e-07 $layer=LI1_cond $X=3.002 $Y=1.055
+ $X2=3.002 $Y2=1.335
r79 26 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.42
r80 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.09
r81 20 42 9.14146 $w=5.58e-07 $l=4.28e-07 $layer=LI1_cond $X=3.43 $Y=1.335
+ $X2=3.002 $Y2=1.335
r82 20 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.255 $X2=3.43 $Y2=1.255
r83 19 34 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.995 $Y=1.87
+ $X2=2.995 $Y2=1.615
r84 18 41 0.106793 $w=5.58e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=1.335
+ $X2=2.995 $Y2=1.335
r85 17 30 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.002 $Y=0.85
+ $X2=3.002 $Y2=1.055
r86 15 16 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.52 $Y=1.62
+ $X2=3.52 $Y2=1.77
r87 15 29 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.49 $Y=1.62 $X2=3.49
+ $Y2=1.42
r88 11 13 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.49 $Y=0.805 $X2=3.58
+ $Y2=0.805
r89 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.58 $Y=0.73 $X2=3.58
+ $Y2=0.805
r90 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.58 $Y=0.73 $X2=3.58
+ $Y2=0.445
r91 7 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.55 $Y=2.165
+ $X2=3.55 $Y2=1.77
r92 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.88 $X2=3.49
+ $Y2=0.805
r93 1 28 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.49 $Y=0.88 $X2=3.49
+ $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_643_369# 1 2 9 13 15 16 18 20 23 27 31 33
+ 36 40 42 43 44 45 47 49 50 54 55 56 57 60 61 63 64 65 66 67 76 80 83 84
c285 84 0 1.78722e-19 $X=5.33 $Y=1.74
c286 80 0 3.22574e-20 $X=3.917 $Y=1.09
c287 76 0 1.95341e-19 $X=7.645 $Y=1.87
c288 66 0 1.36329e-19 $X=7.5 $Y=1.87
c289 64 0 1.42859e-19 $X=5.145 $Y=1.87
c290 61 0 6.7173e-20 $X=8.94 $Y=1.09
c291 60 0 3.87856e-19 $X=8.94 $Y=1.09
c292 49 0 7.67918e-20 $X=3.91 $Y=1.255
r293 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=1.74 $X2=5.33 $Y2=1.74
r294 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.645 $Y=1.87
+ $X2=7.645 $Y2=1.87
r295 73 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r296 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=1.87
+ $X2=3.91 $Y2=1.87
r297 67 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r298 66 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.5 $Y=1.87
+ $X2=7.645 $Y2=1.87
r299 66 67 2.55569 $w=1.4e-07 $l=2.065e-06 $layer=MET1_cond $X=7.5 $Y=1.87
+ $X2=5.435 $Y2=1.87
r300 65 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=1.87
+ $X2=3.91 $Y2=1.87
r301 64 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r302 64 65 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=4.055 $Y2=1.87
r303 63 77 9.70478 $w=2.83e-07 $l=2.4e-07 $layer=LI1_cond $X=7.885 $Y=1.812
+ $X2=7.645 $Y2=1.812
r304 61 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.94 $Y=1.09
+ $X2=8.94 $Y2=0.925
r305 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.94
+ $Y=1.09 $X2=8.94 $Y2=1.09
r306 58 60 7.48077 $w=2.83e-07 $l=1.85e-07 $layer=LI1_cond $X=8.962 $Y=0.905
+ $X2=8.962 $Y2=1.09
r307 56 58 7.22568 $w=1.85e-07 $l=1.82675e-07 $layer=LI1_cond $X=8.82 $Y=0.812
+ $X2=8.962 $Y2=0.905
r308 56 57 41.0663 $w=1.83e-07 $l=6.85e-07 $layer=LI1_cond $X=8.82 $Y=0.812
+ $X2=8.135 $Y2=0.812
r309 55 88 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.97 $Y=1.16
+ $X2=7.97 $Y2=1.325
r310 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.16 $X2=7.97 $Y2=1.16
r311 52 63 6.85451 $w=2.85e-07 $l=1.94715e-07 $layer=LI1_cond $X=8.01 $Y=1.67
+ $X2=7.885 $Y2=1.812
r312 52 54 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=8.01 $Y=1.67
+ $X2=8.01 $Y2=1.16
r313 51 57 7.01633 $w=1.85e-07 $l=1.65076e-07 $layer=LI1_cond $X=8.01 $Y=0.905
+ $X2=8.135 $Y2=0.812
r314 51 54 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.01 $Y=0.905
+ $X2=8.01 $Y2=1.16
r315 50 81 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.917 $Y=1.255
+ $X2=3.917 $Y2=1.42
r316 50 80 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.917 $Y=1.255
+ $X2=3.917 $Y2=1.09
r317 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.91
+ $Y=1.255 $X2=3.91 $Y2=1.255
r318 47 70 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=1.83
+ $X2=3.865 $Y2=1.915
r319 47 49 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.865 $Y=1.83
+ $X2=3.865 $Y2=1.255
r320 46 49 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.865 $Y=0.885
+ $X2=3.865 $Y2=1.255
r321 44 46 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.865 $Y2=0.885
r322 44 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.455 $Y2=0.8
r323 42 70 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.735 $Y=1.915
+ $X2=3.865 $Y2=1.915
r324 42 43 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.735 $Y=1.915
+ $X2=3.425 $Y2=1.915
r325 38 45 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.362 $Y=0.715
+ $X2=3.455 $Y2=0.8
r326 38 40 16.4865 $w=1.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.362 $Y=0.715
+ $X2=3.362 $Y2=0.44
r327 34 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.34 $Y=2
+ $X2=3.425 $Y2=1.915
r328 34 36 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.34 $Y=2 $X2=3.34
+ $Y2=2.16
r329 31 90 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9 $Y=0.445 $X2=9
+ $Y2=0.925
r330 27 88 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.91 $Y=2.065
+ $X2=7.91 $Y2=1.325
r331 21 83 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.33 $Y=1.905
+ $X2=5.33 $Y2=1.74
r332 21 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.33 $Y=1.905
+ $X2=5.33 $Y2=2.275
r333 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.94 $Y=0.73
+ $X2=4.94 $Y2=0.445
r334 17 33 5.30422 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=4.075 $Y=0.805
+ $X2=3.992 $Y2=0.805
r335 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.94 $Y2=0.73
r336 16 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.075 $Y2=0.805
r337 13 33 20.4101 $w=1.5e-07 $l=7.88987e-08 $layer=POLY_cond $X=4 $Y=0.73
+ $X2=3.992 $Y2=0.805
r338 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4 $Y=0.73 $X2=4
+ $Y2=0.445
r339 11 33 20.4101 $w=1.5e-07 $l=7.84219e-08 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=3.992 $Y2=0.805
r340 11 80 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=3.985 $Y2=1.09
r341 9 81 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.97 $Y=2.165
+ $X2=3.97 $Y2=1.42
r342 2 36 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.845 $X2=3.34 $Y2=2.16
r343 1 40 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.37 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_809_369# 1 2 8 9 11 13 16 20 22 24 28 35
+ 36 39 42 43 46 49 50 57 66
c179 66 0 8.01298e-20 $X=4.327 $Y=1.09
c180 46 0 3.47594e-20 $X=4.37 $Y=1.19
c181 22 0 5.6211e-20 $X=8.54 $Y=1.905
c182 16 0 9.48056e-20 $X=5.36 $Y=0.445
c183 9 0 1.42859e-19 $X=5.285 $Y=1.165
c184 8 0 1.78722e-19 $X=4.615 $Y=1.84
r185 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.56
+ $Y=1.74 $X2=8.56 $Y2=1.74
r186 56 57 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.615 $Y=1.255
+ $X2=4.69 $Y2=1.255
r187 53 56 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.405 $Y=1.255
+ $X2=4.615 $Y2=1.255
r188 50 60 28.1708 $w=2.23e-07 $l=5.5e-07 $layer=LI1_cond $X=8.537 $Y=1.19
+ $X2=8.537 $Y2=1.74
r189 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.565 $Y=1.19
+ $X2=8.565 $Y2=1.19
r190 46 67 8.46186 $w=3.23e-07 $l=2.3e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.42
r191 46 66 6.15528 $w=3.23e-07 $l=1e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.09
r192 46 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.255 $X2=4.405 $Y2=1.255
r193 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=1.19
+ $X2=4.37 $Y2=1.19
r194 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=1.19
+ $X2=4.37 $Y2=1.19
r195 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.42 $Y=1.19
+ $X2=8.565 $Y2=1.19
r196 42 43 4.83291 $w=1.4e-07 $l=3.905e-06 $layer=MET1_cond $X=8.42 $Y=1.19
+ $X2=4.515 $Y2=1.19
r197 41 66 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.25 $Y=0.585
+ $X2=4.25 $Y2=1.09
r198 39 41 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0.42
+ $X2=4.23 $Y2=0.585
r199 36 67 29.9635 $w=2.73e-07 $l=7.15e-07 $layer=LI1_cond $X=4.302 $Y=2.135
+ $X2=4.302 $Y2=1.42
r200 35 36 6.01906 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.267 $Y=2.3
+ $X2=4.267 $Y2=2.135
r201 26 28 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=4.615 $Y=1.915
+ $X2=4.91 $Y2=1.915
r202 22 59 38.5495 $w=3.2e-07 $l=1.81659e-07 $layer=POLY_cond $X=8.54 $Y=1.905
+ $X2=8.505 $Y2=1.74
r203 22 24 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.54 $Y=1.905
+ $X2=8.54 $Y2=2.275
r204 18 59 38.5495 $w=3.2e-07 $l=2.14942e-07 $layer=POLY_cond $X=8.39 $Y=1.575
+ $X2=8.505 $Y2=1.74
r205 18 20 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=8.39 $Y=1.575
+ $X2=8.39 $Y2=0.555
r206 14 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.36 $Y=1.09
+ $X2=5.36 $Y2=0.445
r207 11 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.91 $Y=1.99
+ $X2=4.91 $Y2=1.915
r208 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.91 $Y=1.99
+ $X2=4.91 $Y2=2.275
r209 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.285 $Y=1.165
+ $X2=5.36 $Y2=1.09
r210 9 57 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.285 $Y=1.165
+ $X2=4.69 $Y2=1.165
r211 8 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.615 $Y=1.84
+ $X2=4.615 $Y2=1.915
r212 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.615 $Y=1.42
+ $X2=4.615 $Y2=1.255
r213 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.615 $Y=1.42
+ $X2=4.615 $Y2=1.84
r214 2 35 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.845 $X2=4.18 $Y2=2.3
r215 1 39 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.235 $X2=4.21 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_1129_21# 1 2 9 15 19 20 22 24 25 28 32 34
+ 38 44
c96 34 0 4.32543e-20 $X=5.81 $Y=0.72
c97 22 0 4.56917e-20 $X=6.285 $Y=0.72
c98 20 0 5.68782e-20 $X=6.01 $Y=1.74
r99 42 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.84 $Y=1.065
+ $X2=5.84 $Y2=1.575
r100 38 42 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=1.065
r101 38 41 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=0.795
r102 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.81
+ $Y=0.93 $X2=5.81 $Y2=0.93
r103 34 37 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.81 $Y=0.72
+ $X2=5.81 $Y2=0.93
r104 30 32 9.64836 $w=2.13e-07 $l=1.8e-07 $layer=LI1_cond $X=6.712 $Y=2.105
+ $X2=6.712 $Y2=2.285
r105 26 28 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=0.635
+ $X2=6.41 $Y2=0.51
r106 24 30 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.712 $Y2=2.105
r107 24 25 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.095 $Y2=2.02
r108 23 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=0.72
+ $X2=5.81 $Y2=0.72
r109 22 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.285 $Y=0.72
+ $X2=6.41 $Y2=0.635
r110 22 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.285 $Y=0.72
+ $X2=5.975 $Y2=0.72
r111 20 45 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.74
+ $X2=5.955 $Y2=1.905
r112 20 44 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.74
+ $X2=5.955 $Y2=1.575
r113 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.01
+ $Y=1.74 $X2=6.01 $Y2=1.74
r114 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.01 $Y=1.935
+ $X2=6.095 $Y2=2.02
r115 17 19 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.01 $Y=1.935
+ $X2=6.01 $Y2=1.74
r116 15 45 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.84 $Y=2.275
+ $X2=5.84 $Y2=1.905
r117 9 41 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.72 $Y=0.445
+ $X2=5.72 $Y2=0.795
r118 2 32 600 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_PDIFF $count=1 $X=6.555
+ $Y=2.065 $X2=6.715 $Y2=2.285
r119 1 28 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.325
+ $Y=0.235 $X2=6.45 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_997_413# 1 2 11 13 15 18 21 25 29 31 36
+ 38 39 45 46 47 50 52 55
c145 52 0 4.32543e-20 $X=6.39 $Y=1.095
r146 50 56 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.465 $Y=1.16
+ $X2=7.465 $Y2=1.325
r147 50 55 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.465 $Y=1.16
+ $X2=7.465 $Y2=0.995
r148 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.44
+ $Y=1.16 $X2=7.44 $Y2=1.16
r149 45 53 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.39 $Y=1.23
+ $X2=6.39 $Y2=1.365
r150 45 52 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.39 $Y=1.23
+ $X2=6.39 $Y2=1.095
r151 44 47 3.29018 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.475 $Y2=1.185
r152 44 46 6.54147 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.305 $Y2=1.185
r153 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.39
+ $Y=1.23 $X2=6.39 $Y2=1.23
r154 39 49 3.24611 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.355 $Y=1.125
+ $X2=7.44 $Y2=1.125
r155 39 47 33.805 $w=2.98e-07 $l=8.8e-07 $layer=LI1_cond $X=7.355 $Y=1.125
+ $X2=6.475 $Y2=1.125
r156 38 42 6.20468 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=1.31
+ $X2=5.67 $Y2=1.31
r157 38 46 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.755 $Y=1.31
+ $X2=6.305 $Y2=1.31
r158 35 42 0.18542 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=1.395
+ $X2=5.67 $Y2=1.31
r159 35 36 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.67 $Y=1.395
+ $X2=5.67 $Y2=2.135
r160 31 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.585 $Y=2.3
+ $X2=5.67 $Y2=2.135
r161 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.585 $Y=2.3
+ $X2=5.12 $Y2=2.3
r162 27 42 35.1923 $w=1.56e-07 $l=4.5e-07 $layer=LI1_cond $X=5.22 $Y=1.31
+ $X2=5.67 $Y2=1.31
r163 27 29 21.0845 $w=4.38e-07 $l=8.05e-07 $layer=LI1_cond $X=5.22 $Y=1.225
+ $X2=5.22 $Y2=0.42
r164 23 25 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.48 $Y=0.805
+ $X2=6.66 $Y2=0.805
r165 21 56 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.55 $Y=2.065
+ $X2=7.55 $Y2=1.325
r166 18 55 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.495 $Y=0.555
+ $X2=7.495 $Y2=0.995
r167 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.66 $Y=0.73
+ $X2=6.66 $Y2=0.805
r168 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.66 $Y=0.73
+ $X2=6.66 $Y2=0.445
r169 11 53 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=6.48 $Y=2.275
+ $X2=6.48 $Y2=1.365
r170 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.48 $Y=0.88
+ $X2=6.48 $Y2=0.805
r171 7 52 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.48 $Y=0.88
+ $X2=6.48 $Y2=1.095
r172 2 33 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=2.065 $X2=5.12 $Y2=2.3
r173 1 29 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%SET_B 5 9 13 16 19 22 23 27 28 30 32 33 39
+ 40 44 45 46
c136 45 0 4.11784e-20 $X=6.9 $Y=1.68
c137 22 0 2.22391e-19 $X=9.715 $Y=1.985
c138 9 0 4.56917e-20 $X=7.02 $Y=0.445
c139 5 0 1.54163e-19 $X=6.97 $Y=2.275
r140 44 47 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=1.845
r141 44 46 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=1.515
r142 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.9
+ $Y=1.68 $X2=6.9 $Y2=1.68
r143 40 55 4.74535 $w=2.53e-07 $l=1.05e-07 $layer=LI1_cond $X=9.007 $Y=1.53
+ $X2=9.007 $Y2=1.635
r144 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.025 $Y=1.53
+ $X2=9.025 $Y2=1.53
r145 33 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.87 $Y=1.53
+ $X2=6.725 $Y2=1.53
r146 32 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.88 $Y=1.53
+ $X2=9.025 $Y2=1.53
r147 32 33 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=8.88 $Y=1.53
+ $X2=6.87 $Y2=1.53
r148 30 45 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=6.725 $Y=1.605
+ $X2=6.9 $Y2=1.605
r149 30 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.725 $Y=1.53
+ $X2=6.725 $Y2=1.53
r150 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.63 $X2=9.78 $Y2=1.63
r151 25 55 2.77751 $w=1.8e-07 $l=1.28e-07 $layer=LI1_cond $X=9.135 $Y=1.635
+ $X2=9.007 $Y2=1.635
r152 25 27 39.7424 $w=1.78e-07 $l=6.45e-07 $layer=LI1_cond $X=9.135 $Y=1.635
+ $X2=9.78 $Y2=1.635
r153 23 28 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=9.78 $Y=1.6 $X2=9.78
+ $Y2=1.63
r154 23 24 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=9.78 $Y=1.6
+ $X2=9.78 $Y2=1.465
r155 21 28 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=9.78 $Y=1.835
+ $X2=9.78 $Y2=1.63
r156 21 22 45.0833 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=9.715 $Y=1.835
+ $X2=9.715 $Y2=1.985
r157 19 46 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.97 $Y=1.365
+ $X2=6.97 $Y2=1.515
r158 18 19 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.995 $Y=1.215
+ $X2=6.995 $Y2=1.365
r159 16 24 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=9.84 $Y=0.445
+ $X2=9.84 $Y2=1.465
r160 13 22 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.59 $Y=2.275
+ $X2=9.59 $Y2=1.985
r161 9 18 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.02 $Y=0.445
+ $X2=7.02 $Y2=1.215
r162 5 47 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.97 $Y=2.275
+ $X2=6.97 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_1781_295# 1 2 9 11 12 15 18 21 22 24 25
+ 28 31 33 36
c106 25 0 6.7173e-20 $X=9.53 $Y=1.28
c107 12 0 1.89883e-19 $X=9.055 $Y=1.55
c108 11 0 1.97973e-19 $X=9.285 $Y=1.55
r109 33 35 6.80499 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=0.42
+ $X2=10.745 $Y2=0.585
r110 31 36 3.77418 $w=2.45e-07 $l=9.21954e-08 $layer=LI1_cond $X=10.8 $Y=1.195
+ $X2=10.785 $Y2=1.28
r111 31 35 30.5648 $w=2.28e-07 $l=6.1e-07 $layer=LI1_cond $X=10.8 $Y=1.195
+ $X2=10.8 $Y2=0.585
r112 26 36 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.785 $Y=1.365
+ $X2=10.785 $Y2=1.28
r113 26 28 40.7788 $w=2.58e-07 $l=9.2e-07 $layer=LI1_cond $X=10.785 $Y=1.365
+ $X2=10.785 $Y2=2.285
r114 24 36 2.68609 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.655 $Y=1.28
+ $X2=10.785 $Y2=1.28
r115 24 25 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=10.655 $Y=1.28
+ $X2=9.53 $Y2=1.28
r116 22 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.42 $Y=1.02
+ $X2=9.42 $Y2=1.185
r117 22 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.42 $Y=1.02
+ $X2=9.42 $Y2=0.855
r118 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.42
+ $Y=1.02 $X2=9.42 $Y2=1.02
r119 19 25 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.425 $Y=1.195
+ $X2=9.53 $Y2=1.28
r120 19 21 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=9.425 $Y=1.195
+ $X2=9.425 $Y2=1.02
r121 18 39 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.36 $Y=1.475
+ $X2=9.36 $Y2=1.185
r122 15 38 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.36 $Y=0.445
+ $X2=9.36 $Y2=0.855
r123 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.285 $Y=1.55
+ $X2=9.36 $Y2=1.475
r124 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=9.285 $Y=1.55
+ $X2=9.055 $Y2=1.55
r125 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.98 $Y=1.625
+ $X2=9.055 $Y2=1.55
r126 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=8.98 $Y=1.625
+ $X2=8.98 $Y2=2.275
r127 2 28 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=2.065 $X2=10.74 $Y2=2.285
r128 1 33 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=10.485
+ $Y=0.235 $X2=10.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_1597_329# 1 2 3 12 15 17 21 23 25 26 27
+ 28 29 33 37 41 44 45 47 48 50 52 56 58 69
c148 58 0 1.3574e-19 $X=10.32 $Y=1.69
c149 52 0 1.42862e-19 $X=8.905 $Y=1.98
c150 21 0 1.28536e-19 $X=11.47 $Y=0.445
r151 68 69 28.4203 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=10.53 $Y=1.69
+ $X2=10.605 $Y2=1.69
r152 67 68 39.9913 $w=2.7e-07 $l=1.8e-07 $layer=POLY_cond $X=10.35 $Y=1.69
+ $X2=10.53 $Y2=1.69
r153 63 67 2.83073 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=10.35 $Y=1.555
+ $X2=10.35 $Y2=1.69
r154 59 67 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=10.32 $Y=1.69
+ $X2=10.35 $Y2=1.69
r155 58 61 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=10.32 $Y=1.69
+ $X2=10.32 $Y2=1.98
r156 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.32
+ $Y=1.69 $X2=10.32 $Y2=1.69
r157 51 56 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=9.965 $Y=1.98
+ $X2=9.812 $Y2=1.98
r158 50 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.155 $Y=1.98
+ $X2=10.32 $Y2=1.98
r159 50 51 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.155 $Y=1.98
+ $X2=9.965 $Y2=1.98
r160 48 63 138.859 $w=2.7e-07 $l=6.25e-07 $layer=POLY_cond $X=10.35 $Y=0.93
+ $X2=10.35 $Y2=1.555
r161 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.35
+ $Y=0.93 $X2=10.35 $Y2=0.93
r162 45 47 22.0467 $w=2.28e-07 $l=4.4e-07 $layer=LI1_cond $X=9.91 $Y=0.9
+ $X2=10.35 $Y2=0.9
r163 44 45 6.85974 $w=2.3e-07 $l=1.57242e-07 $layer=LI1_cond $X=9.81 $Y=0.785
+ $X2=9.91 $Y2=0.9
r164 43 44 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=9.81 $Y=0.545
+ $X2=9.81 $Y2=0.785
r165 39 56 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.812 $Y=2.065
+ $X2=9.812 $Y2=1.98
r166 39 41 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=9.812 $Y=2.065
+ $X2=9.812 $Y2=2.285
r167 38 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=1.98
+ $X2=8.905 $Y2=1.98
r168 37 56 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.66 $Y=1.98
+ $X2=9.812 $Y2=1.98
r169 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.66 $Y=1.98
+ $X2=8.99 $Y2=1.98
r170 33 43 7.01501 $w=2.7e-07 $l=1.78115e-07 $layer=LI1_cond $X=9.71 $Y=0.41
+ $X2=9.81 $Y2=0.545
r171 33 35 46.0977 $w=2.68e-07 $l=1.08e-06 $layer=LI1_cond $X=9.71 $Y=0.41
+ $X2=8.63 $Y2=0.41
r172 29 52 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=8.905 $Y=2.292
+ $X2=8.905 $Y2=1.98
r173 29 31 18.9207 $w=3.33e-07 $l=5.5e-07 $layer=LI1_cond $X=8.82 $Y=2.292
+ $X2=8.27 $Y2=2.292
r174 26 48 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=10.35 $Y=0.9
+ $X2=10.35 $Y2=0.93
r175 26 27 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=10.35 $Y=0.9
+ $X2=10.35 $Y2=0.765
r176 23 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.47 $Y=1.705
+ $X2=11.47 $Y2=1.63
r177 23 25 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=11.47 $Y=1.705
+ $X2=11.47 $Y2=2.12
r178 19 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.47 $Y=1.555
+ $X2=11.47 $Y2=1.63
r179 19 21 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=11.47 $Y=1.555
+ $X2=11.47 $Y2=0.445
r180 17 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.395 $Y=1.63
+ $X2=11.47 $Y2=1.63
r181 17 69 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.395 $Y=1.63
+ $X2=10.605 $Y2=1.63
r182 13 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.53 $Y=1.825
+ $X2=10.53 $Y2=1.69
r183 13 15 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=10.53 $Y=1.825
+ $X2=10.53 $Y2=2.275
r184 12 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.41 $Y=0.445
+ $X2=10.41 $Y2=0.765
r185 3 41 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=2.065 $X2=9.8 $Y2=2.285
r186 2 31 600 $w=1.7e-07 $l=7.745e-07 $layer=licon1_PDIFF $count=1 $X=7.985
+ $Y=1.645 $X2=8.27 $Y2=2.29
r187 1 35 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=0.235 $X2=8.63 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_2227_47# 1 2 7 9 12 14 16 19 23 27 31 34
+ 38
r62 37 38 81.3105 $w=3.3e-07 $l=4.65e-07 $layer=POLY_cond $X=11.945 $Y=1.16
+ $X2=12.41 $Y2=1.16
r63 32 37 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=11.89 $Y=1.16
+ $X2=11.945 $Y2=1.16
r64 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.89
+ $Y=1.16 $X2=11.89 $Y2=1.16
r65 29 34 0.499868 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=11.345 $Y=1.16
+ $X2=11.215 $Y2=1.16
r66 29 31 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=11.345 $Y=1.16
+ $X2=11.89 $Y2=1.16
r67 25 34 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=11.215 $Y=1.325
+ $X2=11.215 $Y2=1.16
r68 25 27 27.9246 $w=2.58e-07 $l=6.3e-07 $layer=LI1_cond $X=11.215 $Y=1.325
+ $X2=11.215 $Y2=1.955
r69 21 34 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=11.215 $Y=0.995
+ $X2=11.215 $Y2=1.16
r70 21 23 25.2651 $w=2.58e-07 $l=5.7e-07 $layer=LI1_cond $X=11.215 $Y=0.995
+ $X2=11.215 $Y2=0.425
r71 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.41 $Y=1.325
+ $X2=12.41 $Y2=1.16
r72 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.41 $Y=1.325
+ $X2=12.41 $Y2=1.985
r73 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.41 $Y2=1.16
r74 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.41 $Y2=0.56
r75 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.945 $Y=1.325
+ $X2=11.945 $Y2=1.16
r76 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.945 $Y=1.325
+ $X2=11.945 $Y2=1.985
r77 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.945 $Y=0.995
+ $X2=11.945 $Y2=1.16
r78 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.945 $Y=0.995
+ $X2=11.945 $Y2=0.56
r79 2 27 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=11.135
+ $Y=1.8 $X2=11.26 $Y2=1.955
r80 1 23 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=11.135
+ $Y=0.235 $X2=11.26 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_27_369# 1 2 7 10 11 13 14 16
r41 14 16 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=1.125 $Y=2.36
+ $X2=1.88 $Y2=2.36
r42 13 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.04 $Y=2.255
+ $X2=1.125 $Y2=2.36
r43 12 13 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.04 $Y=2.025
+ $X2=1.04 $Y2=2.255
r44 10 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.955 $Y=1.935
+ $X2=1.04 $Y2=2.025
r45 10 11 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=0.955 $Y=1.935
+ $X2=0.345 $Y2=1.935
r46 7 11 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.345 $Y2=1.935
r47 7 9 2.11154 $w=2.6e-07 $l=4.5e-08 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.215 $Y2=2.07
r48 2 16 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=1.845 $X2=1.88 $Y2=2.34
r49 1 9 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 44 48 52 54
+ 56 61 62 64 65 66 68 80 84 96 100 105 111 114 117 126 132 134 137 141
c192 141 0 5.68782e-20 $X=12.65 $Y=2.72
c193 34 0 3.22446e-20 $X=2.82 $Y=2.34
c194 5 0 1.36329e-19 $X=7.045 $Y=2.065
r195 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r196 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r197 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r198 130 132 15.2496 $w=6.78e-07 $l=4.25e-07 $layer=LI1_cond $X=7.59 $Y=2.465
+ $X2=8.015 $Y2=2.465
r199 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r200 128 130 6.42013 $w=6.78e-07 $l=3.65e-07 $layer=LI1_cond $X=7.225 $Y=2.465
+ $X2=7.59 $Y2=2.465
r201 125 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r202 124 128 1.67099 $w=6.78e-07 $l=9.5e-08 $layer=LI1_cond $X=7.13 $Y=2.465
+ $X2=7.225 $Y2=2.465
r203 124 126 9.00537 $w=6.78e-07 $l=7e-08 $layer=LI1_cond $X=7.13 $Y=2.465
+ $X2=7.06 $Y2=2.465
r204 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r205 121 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r206 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r207 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r208 109 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=12.65 $Y2=2.72
r209 109 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r210 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r211 106 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.82 $Y=2.72
+ $X2=11.695 $Y2=2.72
r212 106 108 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.82 $Y=2.72
+ $X2=12.19 $Y2=2.72
r213 105 140 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=12.535 $Y=2.72
+ $X2=12.707 $Y2=2.72
r214 105 108 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.535 $Y=2.72
+ $X2=12.19 $Y2=2.72
r215 104 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r216 104 135 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=10.35 $Y2=2.72
r217 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r218 101 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=2.72
+ $X2=10.32 $Y2=2.72
r219 101 103 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=10.485 $Y=2.72
+ $X2=11.27 $Y2=2.72
r220 100 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.57 $Y=2.72
+ $X2=11.695 $Y2=2.72
r221 100 103 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=11.57 $Y=2.72
+ $X2=11.27 $Y2=2.72
r222 99 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r223 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r224 96 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.155 $Y=2.72
+ $X2=10.32 $Y2=2.72
r225 96 98 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.155 $Y=2.72
+ $X2=9.89 $Y2=2.72
r226 95 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r227 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r228 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r229 92 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r230 91 94 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r231 91 132 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.015 $Y2=2.72
r232 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r233 88 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r234 88 115 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r235 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r236 85 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=3.76 $Y2=2.72
r237 85 87 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r238 84 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r239 84 117 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=6.137 $Y=2.72
+ $X2=6.137 $Y2=2.36
r240 84 87 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=5.75 $Y2=2.72
r241 83 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r242 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r243 80 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.76 $Y2=2.72
r244 80 82 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.45 $Y2=2.72
r245 79 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r246 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r247 76 79 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r248 76 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r249 75 78 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r250 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r251 73 111 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.785 $Y=2.72
+ $X2=0.65 $Y2=2.72
r252 73 75 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=2.72
+ $X2=1.15 $Y2=2.72
r253 68 111 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.65 $Y2=2.72
r254 68 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r255 66 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r256 66 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r257 64 94 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.16 $Y=2.72
+ $X2=8.97 $Y2=2.72
r258 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.16 $Y=2.72
+ $X2=9.325 $Y2=2.72
r259 63 98 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.49 $Y=2.72 $X2=9.89
+ $Y2=2.72
r260 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.49 $Y=2.72
+ $X2=9.325 $Y2=2.72
r261 61 78 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r262 61 62 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.837 $Y2=2.72
r263 60 82 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.985 $Y=2.72
+ $X2=3.45 $Y2=2.72
r264 60 62 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.985 $Y=2.72
+ $X2=2.837 $Y2=2.72
r265 56 59 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=12.665 $Y=1.66
+ $X2=12.665 $Y2=2.34
r266 54 140 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=12.665 $Y=2.635
+ $X2=12.707 $Y2=2.72
r267 54 59 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=12.665 $Y=2.635
+ $X2=12.665 $Y2=2.34
r268 50 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.695 $Y=2.635
+ $X2=11.695 $Y2=2.72
r269 50 52 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=11.695 $Y=2.635
+ $X2=11.695 $Y2=1.955
r270 46 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.32 $Y=2.635
+ $X2=10.32 $Y2=2.72
r271 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.32 $Y=2.635
+ $X2=10.32 $Y2=2.34
r272 42 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=2.635
+ $X2=9.325 $Y2=2.72
r273 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.325 $Y=2.635
+ $X2=9.325 $Y2=2.36
r274 41 84 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=6.137 $Y2=2.72
r275 41 126 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=7.06 $Y2=2.72
r276 36 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=2.635
+ $X2=3.76 $Y2=2.72
r277 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.76 $Y=2.635
+ $X2=3.76 $Y2=2.36
r278 32 62 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.837 $Y=2.635
+ $X2=2.837 $Y2=2.72
r279 32 34 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=2.837 $Y=2.635
+ $X2=2.837 $Y2=2.34
r280 28 111 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=2.635
+ $X2=0.65 $Y2=2.72
r281 28 30 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.65 $Y=2.635
+ $X2=0.65 $Y2=2.36
r282 9 59 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.62 $Y2=2.34
r283 9 56 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.62 $Y2=1.66
r284 8 52 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=11.545
+ $Y=1.8 $X2=11.735 $Y2=1.955
r285 7 48 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=10.195
+ $Y=2.065 $X2=10.32 $Y2=2.34
r286 6 44 600 $w=1.7e-07 $l=4.08258e-07 $layer=licon1_PDIFF $count=1 $X=9.055
+ $Y=2.065 $X2=9.325 $Y2=2.36
r287 5 128 600 $w=1.7e-07 $l=3.74333e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=2.065 $X2=7.225 $Y2=2.36
r288 4 117 600 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_PDIFF $count=1 $X=5.915
+ $Y=2.065 $X2=6.11 $Y2=2.36
r289 3 38 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.845 $X2=3.76 $Y2=2.36
r290 2 34 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.845 $X2=2.82 $Y2=2.34
r291 1 30 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%A_181_47# 1 2 3 4 13 19 21 23 26 30 33 35
+ 36 37 40 43
c137 43 0 3.47594e-20 $X=4.83 $Y=1.53
c138 37 0 1.4475e-19 $X=1.755 $Y=1.53
c139 30 0 1.86564e-19 $X=1.6 $Y=1.965
c140 19 0 9.48056e-20 $X=4.73 $Y=0.42
r141 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.53
+ $X2=4.83 $Y2=1.53
r142 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.53
+ $X2=1.61 $Y2=1.53
r143 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.53
+ $X2=1.61 $Y2=1.53
r144 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.53
+ $X2=4.83 $Y2=1.53
r145 36 37 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=4.685 $Y=1.53
+ $X2=1.755 $Y2=1.53
r146 33 40 42.3206 $w=1.88e-07 $l=7.25e-07 $layer=LI1_cond $X=1.6 $Y=0.805
+ $X2=1.6 $Y2=1.53
r147 31 40 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=1.6 $Y=1.845
+ $X2=1.6 $Y2=1.53
r148 30 31 2.10789 $w=1.9e-07 $l=1.2e-07 $layer=LI1_cond $X=1.6 $Y=1.965 $X2=1.6
+ $Y2=1.845
r149 28 30 6.72258 $w=2.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.46 $Y=1.965
+ $X2=1.6 $Y2=1.965
r150 26 44 5.45457 $w=2.61e-07 $l=9.44722e-08 $layer=LI1_cond $X=4.745 $Y=1.445
+ $X2=4.765 $Y2=1.53
r151 26 35 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.745 $Y=1.445
+ $X2=4.745 $Y2=0.92
r152 21 44 4.38824 $w=2.61e-07 $l=1.04307e-07 $layer=LI1_cond $X=4.722 $Y=1.615
+ $X2=4.765 $Y2=1.53
r153 21 23 36.7174 $w=2.13e-07 $l=6.85e-07 $layer=LI1_cond $X=4.722 $Y=1.615
+ $X2=4.722 $Y2=2.3
r154 17 35 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=4.667 $Y=0.758
+ $X2=4.667 $Y2=0.92
r155 17 19 11.9854 $w=3.23e-07 $l=3.38e-07 $layer=LI1_cond $X=4.667 $Y=0.758
+ $X2=4.667 $Y2=0.42
r156 13 33 20.7082 $w=2.28e-07 $l=4.10293e-07 $layer=LI1_cond $X=1.537 $Y=0.425
+ $X2=1.6 $Y2=0.805
r157 13 15 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.38 $Y=0.425
+ $X2=1.04 $Y2=0.425
r158 4 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=4.575
+ $Y=2.065 $X2=4.7 $Y2=2.3
r159 3 28 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=1.845 $X2=1.46 $Y2=1.97
r160 2 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.605
+ $Y=0.235 $X2=4.73 $Y2=0.42
r161 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.905
+ $Y=0.235 $X2=1.04 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%Q 1 2 7 8 9 10 11 12 23 30 48
c20 30 0 1.28536e-19 $X=12.28 $Y=0.85
r21 48 49 2.50578 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=12.2 $Y=1.53
+ $X2=12.2 $Y2=1.495
r22 30 46 1.30959 $w=2.18e-07 $l=2.5e-08 $layer=LI1_cond $X=12.255 $Y=0.85
+ $X2=12.255 $Y2=0.825
r23 12 43 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=12.2 $Y=2.21
+ $X2=12.2 $Y2=2.34
r24 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=12.2 $Y=1.87
+ $X2=12.2 $Y2=2.21
r25 11 37 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=12.2 $Y=1.87
+ $X2=12.2 $Y2=1.66
r26 10 37 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=12.2 $Y=1.555
+ $X2=12.2 $Y2=1.66
r27 10 48 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=12.2 $Y=1.555
+ $X2=12.2 $Y2=1.53
r28 10 49 1.30959 $w=2.18e-07 $l=2.5e-08 $layer=LI1_cond $X=12.255 $Y=1.47
+ $X2=12.255 $Y2=1.495
r29 9 10 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=12.255 $Y=1.19
+ $X2=12.255 $Y2=1.47
r30 8 46 2.33117 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=12.2 $Y=0.795 $X2=12.2
+ $Y2=0.825
r31 8 21 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=12.2 $Y=0.795
+ $X2=12.2 $Y2=0.66
r32 8 9 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=12.255 $Y=0.88
+ $X2=12.255 $Y2=1.19
r33 8 30 1.57151 $w=2.18e-07 $l=3e-08 $layer=LI1_cond $X=12.255 $Y=0.88
+ $X2=12.255 $Y2=0.85
r34 7 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=12.2 $Y=0.51 $X2=12.2
+ $Y2=0.66
r35 7 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=12.2 $Y=0.51 $X2=12.2
+ $Y2=0.36
r36 2 43 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=12.02
+ $Y=1.485 $X2=12.2 $Y2=2.34
r37 2 37 400 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=12.02
+ $Y=1.485 $X2=12.2 $Y2=1.66
r38 1 23 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=12.02
+ $Y=0.235 $X2=12.2 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 44 47 49
+ 52 53 54 60 64 69 79 87 92 98 105 108 119 123 125 128 132
c176 132 0 2.71124e-20 $X=12.65 $Y=0
c177 34 0 4.13602e-20 $X=2.85 $Y=0.38
r178 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r179 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r180 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r181 121 123 11.6653 $w=8.88e-07 $l=1.25e-07 $layer=LI1_cond $X=7.59 $Y=0.36
+ $X2=7.715 $Y2=0.36
r182 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r183 118 121 4.79775 $w=8.88e-07 $l=3.5e-07 $layer=LI1_cond $X=7.24 $Y=0.36
+ $X2=7.59 $Y2=0.36
r184 118 119 17.2855 $w=8.88e-07 $l=5.35e-07 $layer=LI1_cond $X=7.24 $Y=0.36
+ $X2=6.705 $Y2=0.36
r185 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r186 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r187 98 103 8.24843 $w=6.36e-07 $l=4.3e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.35
+ $Y2=0.43
r188 98 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r189 96 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=12.65 $Y2=0
r190 96 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r191 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r192 93 128 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=11.865 $Y=0
+ $X2=11.717 $Y2=0
r193 93 95 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.865 $Y=0
+ $X2=12.19 $Y2=0
r194 92 131 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=12.535 $Y=0
+ $X2=12.707 $Y2=0
r195 92 95 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.535 $Y=0
+ $X2=12.19 $Y2=0
r196 91 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r197 91 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=10.35 $Y2=0
r198 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r199 88 125 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=10.24 $Y2=0
r200 88 90 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=11.27 $Y2=0
r201 87 128 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=11.57 $Y=0
+ $X2=11.717 $Y2=0
r202 87 90 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=11.57 $Y=0 $X2=11.27
+ $Y2=0
r203 86 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r204 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r205 83 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.89 $Y2=0
r206 83 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r207 82 85 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=8.05 $Y=0 $X2=9.89
+ $Y2=0
r208 82 123 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=7.715 $Y2=0
r209 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r210 79 125 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.24 $Y2=0
r211 79 85 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.89 $Y2=0
r212 78 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r213 78 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=5.75 $Y2=0
r214 77 119 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=6.705 $Y2=0
r215 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r216 75 77 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.67 $Y2=0
r217 73 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r218 73 109 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=3.91 $Y2=0
r219 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r220 70 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=3.79 $Y2=0
r221 70 72 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=5.29 $Y2=0
r222 69 115 9.37134 $w=4.83e-07 $l=3.8e-07 $layer=LI1_cond $X=5.852 $Y=0
+ $X2=5.852 $Y2=0.38
r223 69 75 6.96588 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=5.852 $Y=0
+ $X2=6.095 $Y2=0
r224 69 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r225 69 72 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.29
+ $Y2=0
r226 68 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r227 68 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.99 $Y2=0
r228 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r229 65 105 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.895
+ $Y2=0
r230 65 67 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.45
+ $Y2=0
r231 64 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0
+ $X2=3.79 $Y2=0
r232 64 67 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.625 $Y=0
+ $X2=3.45 $Y2=0
r233 63 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.99 $Y2=0
r234 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r235 60 105 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.69 $Y=0
+ $X2=2.895 $Y2=0
r236 60 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.53
+ $Y2=0
r237 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r238 59 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=0.69 $Y2=0
r239 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r240 56 98 8.69404 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=0.7 $Y=0 $X2=0.35
+ $Y2=0
r241 56 58 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.7 $Y=0 $X2=1.61
+ $Y2=0
r242 54 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r243 54 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r244 52 58 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=1.61 $Y2=0
r245 52 53 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=1.957 $Y2=0
r246 51 62 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.53
+ $Y2=0
r247 51 53 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.957
+ $Y2=0
r248 47 131 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=12.665 $Y=0.085
+ $X2=12.707 $Y2=0
r249 47 49 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=12.665 $Y=0.085
+ $X2=12.665 $Y2=0.38
r250 44 128 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=11.717 $Y=0.085
+ $X2=11.717 $Y2=0
r251 44 46 11.3729 $w=2.95e-07 $l=2.75e-07 $layer=LI1_cond $X=11.717 $Y=0.085
+ $X2=11.717 $Y2=0.36
r252 40 125 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.24 $Y=0.085
+ $X2=10.24 $Y2=0
r253 40 42 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=10.24 $Y=0.085
+ $X2=10.24 $Y2=0.36
r254 36 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0
r255 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0.36
r256 32 105 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0
r257 32 34 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0.38
r258 28 53 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.957 $Y=0.085
+ $X2=1.957 $Y2=0
r259 28 30 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.957 $Y=0.085
+ $X2=1.957 $Y2=0.38
r260 9 49 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.485
+ $Y=0.235 $X2=12.62 $Y2=0.38
r261 8 46 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=11.545
+ $Y=0.235 $X2=11.735 $Y2=0.36
r262 7 42 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=9.915
+ $Y=0.235 $X2=10.2 $Y2=0.36
r263 6 118 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.095
+ $Y=0.235 $X2=7.24 $Y2=0.36
r264 5 115 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.235 $X2=5.93 $Y2=0.38
r265 4 38 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.235 $X2=3.79 $Y2=0.36
r266 3 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.85 $Y2=0.38
r267 2 30 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=1.745
+ $Y=0.235 $X2=1.91 $Y2=0.38
r268 1 103 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends


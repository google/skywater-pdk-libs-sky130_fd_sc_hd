* File: sky130_fd_sc_hd__dlymetal6s6s_1.spice.SKY130_FD_SC_HD__DLYMETAL6S6S_1.pxi
* Created: Thu Aug 27 14:19:12 2020
* 
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A N_A_M1002_g N_A_M1011_g A A N_A_c_92_n
+ N_A_c_93_n PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_63_47# N_A_63_47#_M1002_s
+ N_A_63_47#_M1011_s N_A_63_47#_M1006_g N_A_63_47#_M1009_g N_A_63_47#_c_122_n
+ N_A_63_47#_c_129_n N_A_63_47#_c_130_n N_A_63_47#_c_123_n N_A_63_47#_c_131_n
+ N_A_63_47#_c_124_n N_A_63_47#_c_125_n N_A_63_47#_c_126_n N_A_63_47#_c_127_n
+ PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_63_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_240_47# N_A_240_47#_M1006_d
+ N_A_240_47#_M1009_d N_A_240_47#_M1000_g N_A_240_47#_M1010_g
+ N_A_240_47#_c_183_n N_A_240_47#_c_184_n N_A_240_47#_c_190_n
+ N_A_240_47#_c_185_n N_A_240_47#_c_186_n N_A_240_47#_c_187_n
+ PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_240_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_346_47# N_A_346_47#_M1000_s
+ N_A_346_47#_M1010_s N_A_346_47#_M1005_g N_A_346_47#_M1007_g
+ N_A_346_47#_c_237_n N_A_346_47#_c_244_n N_A_346_47#_c_238_n
+ N_A_346_47#_c_239_n N_A_346_47#_c_245_n N_A_346_47#_c_246_n
+ N_A_346_47#_c_240_n N_A_346_47#_c_247_n N_A_346_47#_c_241_n
+ N_A_346_47#_c_242_n PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_346_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_523_47# N_A_523_47#_M1005_d
+ N_A_523_47#_M1007_d N_A_523_47#_M1003_g N_A_523_47#_M1001_g
+ N_A_523_47#_c_307_n N_A_523_47#_c_308_n N_A_523_47#_c_314_n
+ N_A_523_47#_c_309_n N_A_523_47#_c_310_n N_A_523_47#_c_311_n
+ PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_523_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_629_47# N_A_629_47#_M1003_s
+ N_A_629_47#_M1001_s N_A_629_47#_M1008_g N_A_629_47#_M1004_g
+ N_A_629_47#_c_361_n N_A_629_47#_c_368_n N_A_629_47#_c_362_n
+ N_A_629_47#_c_363_n N_A_629_47#_c_369_n N_A_629_47#_c_370_n
+ N_A_629_47#_c_364_n N_A_629_47#_c_371_n N_A_629_47#_c_365_n
+ N_A_629_47#_c_366_n PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%A_629_47#
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%VPWR N_VPWR_M1011_d N_VPWR_M1010_d
+ N_VPWR_M1001_d N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n
+ N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n
+ VPWR N_VPWR_c_437_n N_VPWR_c_427_n VPWR
+ PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%VPWR
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%X N_X_M1008_d N_X_M1004_d X X X X X X X
+ N_X_c_491_n X PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%X
x_PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%VGND N_VGND_M1002_d N_VGND_M1000_d
+ N_VGND_M1003_d N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n
+ N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n
+ VGND N_VGND_c_515_n N_VGND_c_516_n VGND
+ PM_SKY130_FD_SC_HD__DLYMETAL6S6S_1%VGND
cc_1 VNB N_A_M1002_g 0.0375092f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.445
cc_2 VNB N_A_c_92_n 0.0169688f $X=-0.19 $Y=-0.24 $X2=0.425 $Y2=1.16
cc_3 VNB N_A_c_93_n 0.0364194f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_4 VNB N_A_63_47#_c_122_n 0.00223093f $X=-0.19 $Y=-0.24 $X2=0.425 $Y2=1.16
cc_5 VNB N_A_63_47#_c_123_n 0.0325421f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.53
cc_6 VNB N_A_63_47#_c_124_n 0.00181412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_63_47#_c_125_n 0.0236222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_63_47#_c_126_n 0.00164805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_63_47#_c_127_n 0.0190552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_240_47#_M1000_g 0.0342027f $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.105
cc_11 VNB N_A_240_47#_c_183_n 0.00445733f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_12 VNB N_A_240_47#_c_184_n 0.0136496f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_13 VNB N_A_240_47#_c_185_n 0.00354377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_240_47#_c_186_n 0.00124639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_240_47#_c_187_n 0.0338076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_346_47#_c_237_n 0.00372278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_346_47#_c_238_n 9.94839e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_346_47#_c_239_n 0.0035095f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.53
cc_19 VNB N_A_346_47#_c_240_n 0.00356627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_346_47#_c_241_n 0.0236222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_346_47#_c_242_n 0.0190552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_523_47#_M1003_g 0.0342704f $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.105
cc_23 VNB N_A_523_47#_c_307_n 0.00410383f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_24 VNB N_A_523_47#_c_308_n 0.0138223f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_25 VNB N_A_523_47#_c_309_n 0.00345589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_523_47#_c_310_n 0.00106881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_523_47#_c_311_n 0.0338076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_629_47#_c_361_n 0.00413815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_629_47#_c_362_n 9.94839e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_629_47#_c_363_n 0.0038023f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.53
cc_31 VNB N_A_629_47#_c_364_n 0.00358557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_629_47#_c_365_n 0.0227379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_629_47#_c_366_n 0.0190552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_427_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB X 0.0265377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_491_n 0.028327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_506_n 4.8975e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_507_n 4.8975e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_508_n 4.8975e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_509_n 0.0183578f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.53
cc_41 VNB N_VGND_c_510_n 0.00509417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_511_n 0.0250307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_512_n 0.00509417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_513_n 0.0250307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_514_n 0.00509417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_515_n 0.0189802f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_516_n 0.256851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VPB N_A_M1011_g 0.0605617f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=2.275
cc_49 VPB N_A_c_92_n 0.0258557f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.16
cc_50 VPB N_A_c_93_n 0.00991829f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_51 VPB N_A_63_47#_M1009_g 0.0216941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_63_47#_c_129_n 0.00279153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_63_47#_c_130_n 0.00421703f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.19
cc_54 VPB N_A_63_47#_c_131_n 0.0344591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_63_47#_c_125_n 0.00483834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_240_47#_M1010_g 0.057273f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.16
cc_57 VPB N_A_240_47#_c_184_n 0.0173651f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_58 VPB N_A_240_47#_c_190_n 0.0085186f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.19
cc_59 VPB N_A_240_47#_c_187_n 0.00984422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_346_47#_M1007_g 0.0216941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_346_47#_c_244_n 0.00422847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_346_47#_c_245_n 0.00171281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_346_47#_c_246_n 0.00414163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_346_47#_c_247_n 0.00412498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_346_47#_c_241_n 0.00483834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_523_47#_M1001_g 0.0573411f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.16
cc_67 VPB N_A_523_47#_c_308_n 0.0175457f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_68 VPB N_A_523_47#_c_314_n 0.00787309f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.19
cc_69 VPB N_A_523_47#_c_311_n 0.00984422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_629_47#_M1004_g 0.0216957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_629_47#_c_368_n 0.00466306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_629_47#_c_369_n 0.00171281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_629_47#_c_370_n 0.00445875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_629_47#_c_371_n 0.00414413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_629_47#_c_365_n 0.00478128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_428_n 4.8975e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_429_n 4.8975e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_430_n 4.8975e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_431_n 0.0183929f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.53
cc_80 VPB N_VPWR_c_432_n 0.00509586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_433_n 0.0250658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_434_n 0.00509586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_435_n 0.0250658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_436_n 0.00509586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_437_n 0.0189802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_427_n 0.0630238f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB X 0.036851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB X 0.0107121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB X 0.0101632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 N_A_M1011_g N_A_63_47#_M1009_g 0.0332384f $X=0.65 $Y=2.275 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_A_63_47#_c_122_n 0.0169506f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_c_92_n N_A_63_47#_c_122_n 0.00392725f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_c_93_n N_A_63_47#_c_122_n 3.45424e-19 $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_M1011_g N_A_63_47#_c_129_n 0.017035f $X=0.65 $Y=2.275 $X2=0 $Y2=0
cc_95 N_A_c_92_n N_A_63_47#_c_129_n 0.00415099f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_M1011_g N_A_63_47#_c_130_n 0.00523842f $X=0.65 $Y=2.275 $X2=0 $Y2=0
cc_97 N_A_M1002_g N_A_63_47#_c_123_n 0.00157467f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_c_92_n N_A_63_47#_c_123_n 0.0395459f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_c_93_n N_A_63_47#_c_123_n 0.00181525f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_M1011_g N_A_63_47#_c_131_n 0.00297922f $X=0.65 $Y=2.275 $X2=0 $Y2=0
cc_101 N_A_c_92_n N_A_63_47#_c_131_n 0.0407433f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_c_93_n N_A_63_47#_c_131_n 8.36308e-19 $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_c_92_n N_A_63_47#_c_124_n 0.0594988f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_c_93_n N_A_63_47#_c_124_n 0.00523842f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_c_92_n N_A_63_47#_c_125_n 2.32992e-19 $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_c_93_n N_A_63_47#_c_125_n 0.0207322f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_M1002_g N_A_63_47#_c_126_n 0.00523842f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_M1002_g N_A_63_47#_c_127_n 0.0194524f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_M1011_g N_VPWR_c_428_n 0.00906078f $X=0.65 $Y=2.275 $X2=0 $Y2=0
cc_110 N_A_M1011_g N_VPWR_c_431_n 0.00344532f $X=0.65 $Y=2.275 $X2=0 $Y2=0
cc_111 N_A_M1011_g N_VPWR_c_427_n 0.00520521f $X=0.65 $Y=2.275 $X2=0 $Y2=0
cc_112 N_A_M1002_g N_VGND_c_506_n 0.00878516f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_M1002_g N_VGND_c_509_n 0.00341689f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_M1002_g N_VGND_c_516_n 0.00515575f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_63_47#_M1009_g N_A_240_47#_c_184_n 0.00377535f $X=1.125 $Y=1.985
+ $X2=0 $Y2=0
cc_116 N_A_63_47#_c_130_n N_A_240_47#_c_184_n 0.0108332f $X=0.912 $Y=1.87 $X2=0
+ $Y2=0
cc_117 N_A_63_47#_c_124_n N_A_240_47#_c_184_n 0.0281441f $X=1.07 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_A_63_47#_c_125_n N_A_240_47#_c_184_n 0.00337067f $X=1.07 $Y=1.16 $X2=0
+ $Y2=0
cc_119 N_A_63_47#_c_126_n N_A_240_47#_c_185_n 0.00963224f $X=0.95 $Y=0.995 $X2=0
+ $Y2=0
cc_120 N_A_63_47#_c_127_n N_A_240_47#_c_185_n 0.00357896f $X=1.07 $Y=0.995 $X2=0
+ $Y2=0
cc_121 N_A_63_47#_c_124_n N_A_240_47#_c_187_n 2.35103e-19 $X=1.07 $Y=1.16 $X2=0
+ $Y2=0
cc_122 N_A_63_47#_c_125_n N_A_240_47#_c_187_n 0.0058474f $X=1.07 $Y=1.16 $X2=0
+ $Y2=0
cc_123 N_A_63_47#_c_129_n N_VPWR_M1011_d 0.00207054f $X=0.745 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_124 N_A_63_47#_c_130_n N_VPWR_M1011_d 7.20661e-19 $X=0.912 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_125 N_A_63_47#_M1009_g N_VPWR_c_428_n 0.00905956f $X=1.125 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_63_47#_c_129_n N_VPWR_c_428_n 0.0245954f $X=0.745 $Y=1.955 $X2=0
+ $Y2=0
cc_127 N_A_63_47#_c_129_n N_VPWR_c_431_n 0.00259647f $X=0.745 $Y=1.955 $X2=0
+ $Y2=0
cc_128 N_A_63_47#_c_131_n N_VPWR_c_431_n 0.0306027f $X=0.305 $Y=1.955 $X2=0
+ $Y2=0
cc_129 N_A_63_47#_M1009_g N_VPWR_c_433_n 0.0046653f $X=1.125 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_63_47#_M1011_s N_VPWR_c_427_n 0.00230841f $X=0.315 $Y=2.065 $X2=0
+ $Y2=0
cc_131 N_A_63_47#_M1009_g N_VPWR_c_427_n 0.00921786f $X=1.125 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_63_47#_c_129_n N_VPWR_c_427_n 0.00581522f $X=0.745 $Y=1.955 $X2=0
+ $Y2=0
cc_133 N_A_63_47#_c_131_n N_VPWR_c_427_n 0.0168095f $X=0.305 $Y=1.955 $X2=0
+ $Y2=0
cc_134 N_A_63_47#_c_122_n N_VGND_M1002_d 0.00264964f $X=0.745 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_63_47#_c_122_n N_VGND_c_506_n 0.024366f $X=0.745 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_63_47#_c_125_n N_VGND_c_506_n 3.47021e-19 $X=1.07 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_63_47#_c_127_n N_VGND_c_506_n 0.00878394f $X=1.07 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_A_63_47#_c_122_n N_VGND_c_509_n 0.00273399f $X=0.745 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_63_47#_c_123_n N_VGND_c_509_n 0.0305064f $X=0.44 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A_63_47#_c_127_n N_VGND_c_511_n 0.0046653f $X=1.07 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_63_47#_M1002_s N_VGND_c_516_n 0.00229009f $X=0.315 $Y=0.235 $X2=0
+ $Y2=0
cc_142 N_A_63_47#_c_122_n N_VGND_c_516_n 0.00598099f $X=0.745 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_63_47#_c_123_n N_VGND_c_516_n 0.0167909f $X=0.44 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_63_47#_c_127_n N_VGND_c_516_n 0.00934473f $X=1.07 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_A_240_47#_M1010_g N_A_346_47#_M1007_g 0.0333474f $X=2.065 $Y=2.275
+ $X2=0 $Y2=0
cc_146 N_A_240_47#_c_183_n N_A_346_47#_c_237_n 0.0320836f $X=1.335 $Y=0.44 $X2=0
+ $Y2=0
cc_147 N_A_240_47#_M1010_g N_A_346_47#_c_244_n 0.00126727f $X=2.065 $Y=2.275
+ $X2=0 $Y2=0
cc_148 N_A_240_47#_c_190_n N_A_346_47#_c_244_n 0.0340913f $X=1.335 $Y=1.96 $X2=0
+ $Y2=0
cc_149 N_A_240_47#_M1000_g N_A_346_47#_c_238_n 0.0178073f $X=2.065 $Y=0.445
+ $X2=0 $Y2=0
cc_150 N_A_240_47#_c_184_n N_A_346_47#_c_238_n 0.00275926f $X=1.385 $Y=1.675
+ $X2=0 $Y2=0
cc_151 N_A_240_47#_c_187_n N_A_346_47#_c_238_n 8.08044e-19 $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_152 N_A_240_47#_c_183_n N_A_346_47#_c_239_n 0.014785f $X=1.335 $Y=0.44 $X2=0
+ $Y2=0
cc_153 N_A_240_47#_c_184_n N_A_346_47#_c_239_n 0.0220527f $X=1.385 $Y=1.675
+ $X2=0 $Y2=0
cc_154 N_A_240_47#_c_187_n N_A_346_47#_c_239_n 0.00182316f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_155 N_A_240_47#_M1010_g N_A_346_47#_c_245_n 0.0191857f $X=2.065 $Y=2.275
+ $X2=0 $Y2=0
cc_156 N_A_240_47#_c_184_n N_A_346_47#_c_245_n 0.00294539f $X=1.385 $Y=1.675
+ $X2=0 $Y2=0
cc_157 N_A_240_47#_c_187_n N_A_346_47#_c_245_n 5.13753e-19 $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_158 N_A_240_47#_c_184_n N_A_346_47#_c_246_n 0.023264f $X=1.385 $Y=1.675 $X2=0
+ $Y2=0
cc_159 N_A_240_47#_c_190_n N_A_346_47#_c_246_n 0.0170057f $X=1.335 $Y=1.96 $X2=0
+ $Y2=0
cc_160 N_A_240_47#_c_187_n N_A_346_47#_c_246_n 8.79705e-19 $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_161 N_A_240_47#_M1000_g N_A_346_47#_c_240_n 0.00553444f $X=2.065 $Y=0.445
+ $X2=0 $Y2=0
cc_162 N_A_240_47#_c_184_n N_A_346_47#_c_240_n 0.0282667f $X=1.385 $Y=1.675
+ $X2=0 $Y2=0
cc_163 N_A_240_47#_c_185_n N_A_346_47#_c_240_n 0.00544075f $X=1.422 $Y=0.995
+ $X2=0 $Y2=0
cc_164 N_A_240_47#_M1010_g N_A_346_47#_c_247_n 0.00587049f $X=2.065 $Y=2.275
+ $X2=0 $Y2=0
cc_165 N_A_240_47#_c_184_n N_A_346_47#_c_247_n 0.0309738f $X=1.385 $Y=1.675
+ $X2=0 $Y2=0
cc_166 N_A_240_47#_c_190_n N_A_346_47#_c_247_n 0.00556293f $X=1.335 $Y=1.96
+ $X2=0 $Y2=0
cc_167 N_A_240_47#_c_184_n N_A_346_47#_c_241_n 2.22114e-19 $X=1.385 $Y=1.675
+ $X2=0 $Y2=0
cc_168 N_A_240_47#_c_187_n N_A_346_47#_c_241_n 0.0207275f $X=2.065 $Y=1.16 $X2=0
+ $Y2=0
cc_169 N_A_240_47#_M1000_g N_A_346_47#_c_242_n 0.0194472f $X=2.065 $Y=0.445
+ $X2=0 $Y2=0
cc_170 N_A_240_47#_M1010_g N_VPWR_c_429_n 0.00906078f $X=2.065 $Y=2.275 $X2=0
+ $Y2=0
cc_171 N_A_240_47#_M1010_g N_VPWR_c_433_n 0.00344532f $X=2.065 $Y=2.275 $X2=0
+ $Y2=0
cc_172 N_A_240_47#_c_190_n N_VPWR_c_433_n 0.018718f $X=1.335 $Y=1.96 $X2=0 $Y2=0
cc_173 N_A_240_47#_M1009_d N_VPWR_c_427_n 0.00382897f $X=1.2 $Y=1.485 $X2=0
+ $Y2=0
cc_174 N_A_240_47#_M1010_g N_VPWR_c_427_n 0.00545273f $X=2.065 $Y=2.275 $X2=0
+ $Y2=0
cc_175 N_A_240_47#_c_190_n N_VPWR_c_427_n 0.0103212f $X=1.335 $Y=1.96 $X2=0
+ $Y2=0
cc_176 N_A_240_47#_M1000_g N_VGND_c_507_n 0.00878516f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_240_47#_M1000_g N_VGND_c_511_n 0.00341689f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A_240_47#_c_183_n N_VGND_c_511_n 0.0186568f $X=1.335 $Y=0.44 $X2=0
+ $Y2=0
cc_179 N_A_240_47#_M1006_d N_VGND_c_516_n 0.00387172f $X=1.2 $Y=0.235 $X2=0
+ $Y2=0
cc_180 N_A_240_47#_M1000_g N_VGND_c_516_n 0.00540327f $X=2.065 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_240_47#_c_183_n N_VGND_c_516_n 0.0103081f $X=1.335 $Y=0.44 $X2=0
+ $Y2=0
cc_182 N_A_346_47#_M1007_g N_A_523_47#_c_308_n 0.00377535f $X=2.54 $Y=1.985
+ $X2=0 $Y2=0
cc_183 N_A_346_47#_c_240_n N_A_523_47#_c_308_n 0.0283504f $X=2.32 $Y=1.325 $X2=0
+ $Y2=0
cc_184 N_A_346_47#_c_247_n N_A_523_47#_c_308_n 0.0108652f $X=2.32 $Y=1.845 $X2=0
+ $Y2=0
cc_185 N_A_346_47#_c_241_n N_A_523_47#_c_308_n 0.00336476f $X=2.485 $Y=1.16
+ $X2=0 $Y2=0
cc_186 N_A_346_47#_c_240_n N_A_523_47#_c_309_n 0.00964625f $X=2.32 $Y=1.325
+ $X2=0 $Y2=0
cc_187 N_A_346_47#_c_242_n N_A_523_47#_c_309_n 0.00356258f $X=2.485 $Y=0.995
+ $X2=0 $Y2=0
cc_188 N_A_346_47#_c_240_n N_A_523_47#_c_311_n 2.35222e-19 $X=2.32 $Y=1.325
+ $X2=0 $Y2=0
cc_189 N_A_346_47#_c_241_n N_A_523_47#_c_311_n 0.0058474f $X=2.485 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_346_47#_c_245_n N_VPWR_M1010_d 0.00207054f $X=2.145 $Y=1.942 $X2=0
+ $Y2=0
cc_191 N_A_346_47#_c_247_n N_VPWR_M1010_d 6.23798e-19 $X=2.32 $Y=1.845 $X2=0
+ $Y2=0
cc_192 N_A_346_47#_M1007_g N_VPWR_c_429_n 0.00905956f $X=2.54 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_346_47#_c_245_n N_VPWR_c_429_n 0.024785f $X=2.145 $Y=1.942 $X2=0
+ $Y2=0
cc_194 N_A_346_47#_c_244_n N_VPWR_c_433_n 0.0171684f $X=1.855 $Y=2.275 $X2=0
+ $Y2=0
cc_195 N_A_346_47#_c_245_n N_VPWR_c_433_n 0.00261227f $X=2.145 $Y=1.942 $X2=0
+ $Y2=0
cc_196 N_A_346_47#_M1007_g N_VPWR_c_435_n 0.0046653f $X=2.54 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A_346_47#_M1010_s N_VPWR_c_427_n 0.00230841f $X=1.73 $Y=2.065 $X2=0
+ $Y2=0
cc_198 N_A_346_47#_M1007_g N_VPWR_c_427_n 0.00921786f $X=2.54 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_346_47#_c_244_n N_VPWR_c_427_n 0.00952784f $X=1.855 $Y=2.275 $X2=0
+ $Y2=0
cc_200 N_A_346_47#_c_245_n N_VPWR_c_427_n 0.005846f $X=2.145 $Y=1.942 $X2=0
+ $Y2=0
cc_201 N_A_346_47#_c_240_n N_VGND_M1000_d 0.0028099f $X=2.32 $Y=1.325 $X2=0
+ $Y2=0
cc_202 N_A_346_47#_c_238_n N_VGND_c_507_n 0.00217981f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_203 N_A_346_47#_c_240_n N_VGND_c_507_n 0.0222857f $X=2.32 $Y=1.325 $X2=0
+ $Y2=0
cc_204 N_A_346_47#_c_241_n N_VGND_c_507_n 3.47021e-19 $X=2.485 $Y=1.16 $X2=0
+ $Y2=0
cc_205 N_A_346_47#_c_242_n N_VGND_c_507_n 0.00878394f $X=2.485 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_346_47#_c_237_n N_VGND_c_511_n 0.0170644f $X=1.855 $Y=0.44 $X2=0
+ $Y2=0
cc_207 N_A_346_47#_c_238_n N_VGND_c_511_n 0.00273399f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A_346_47#_c_242_n N_VGND_c_513_n 0.0046653f $X=2.485 $Y=0.995 $X2=0
+ $Y2=0
cc_209 N_A_346_47#_M1000_s N_VGND_c_516_n 0.00229009f $X=1.73 $Y=0.235 $X2=0
+ $Y2=0
cc_210 N_A_346_47#_c_237_n N_VGND_c_516_n 0.00950719f $X=1.855 $Y=0.44 $X2=0
+ $Y2=0
cc_211 N_A_346_47#_c_238_n N_VGND_c_516_n 0.00430392f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_346_47#_c_240_n N_VGND_c_516_n 0.00168578f $X=2.32 $Y=1.325 $X2=0
+ $Y2=0
cc_213 N_A_346_47#_c_242_n N_VGND_c_516_n 0.00934473f $X=2.485 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_523_47#_M1001_g N_A_629_47#_M1004_g 0.0333474f $X=3.48 $Y=2.275 $X2=0
+ $Y2=0
cc_215 N_A_523_47#_c_307_n N_A_629_47#_c_361_n 0.0320831f $X=2.75 $Y=0.44 $X2=0
+ $Y2=0
cc_216 N_A_523_47#_M1001_g N_A_629_47#_c_368_n 0.00127614f $X=3.48 $Y=2.275
+ $X2=0 $Y2=0
cc_217 N_A_523_47#_c_314_n N_A_629_47#_c_368_n 0.0340908f $X=2.75 $Y=1.96 $X2=0
+ $Y2=0
cc_218 N_A_523_47#_M1003_g N_A_629_47#_c_362_n 0.0178581f $X=3.48 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_A_523_47#_c_308_n N_A_629_47#_c_362_n 0.00275926f $X=2.79 $Y=1.675
+ $X2=0 $Y2=0
cc_220 N_A_523_47#_c_311_n N_A_629_47#_c_362_n 8.08044e-19 $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_221 N_A_523_47#_c_307_n N_A_629_47#_c_363_n 0.0147055f $X=2.75 $Y=0.44 $X2=0
+ $Y2=0
cc_222 N_A_523_47#_c_308_n N_A_629_47#_c_363_n 0.0239021f $X=2.79 $Y=1.675 $X2=0
+ $Y2=0
cc_223 N_A_523_47#_c_311_n N_A_629_47#_c_363_n 0.00182316f $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_224 N_A_523_47#_M1001_g N_A_629_47#_c_369_n 0.019244f $X=3.48 $Y=2.275 $X2=0
+ $Y2=0
cc_225 N_A_523_47#_c_308_n N_A_629_47#_c_369_n 0.00294539f $X=2.79 $Y=1.675
+ $X2=0 $Y2=0
cc_226 N_A_523_47#_c_311_n N_A_629_47#_c_369_n 5.13753e-19 $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_227 N_A_523_47#_c_308_n N_A_629_47#_c_370_n 0.025125f $X=2.79 $Y=1.675 $X2=0
+ $Y2=0
cc_228 N_A_523_47#_c_314_n N_A_629_47#_c_370_n 0.016914f $X=2.75 $Y=1.96 $X2=0
+ $Y2=0
cc_229 N_A_523_47#_c_311_n N_A_629_47#_c_370_n 8.79705e-19 $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_523_47#_M1003_g N_A_629_47#_c_364_n 0.00557763f $X=3.48 $Y=0.445
+ $X2=0 $Y2=0
cc_231 N_A_523_47#_c_308_n N_A_629_47#_c_364_n 0.0282667f $X=2.79 $Y=1.675 $X2=0
+ $Y2=0
cc_232 N_A_523_47#_c_309_n N_A_629_47#_c_364_n 0.00527024f $X=2.827 $Y=0.995
+ $X2=0 $Y2=0
cc_233 N_A_523_47#_M1001_g N_A_629_47#_c_371_n 0.00591327f $X=3.48 $Y=2.275
+ $X2=0 $Y2=0
cc_234 N_A_523_47#_c_308_n N_A_629_47#_c_371_n 0.0309738f $X=2.79 $Y=1.675 $X2=0
+ $Y2=0
cc_235 N_A_523_47#_c_314_n N_A_629_47#_c_371_n 0.00540018f $X=2.75 $Y=1.96 $X2=0
+ $Y2=0
cc_236 N_A_523_47#_c_308_n N_A_629_47#_c_365_n 2.22114e-19 $X=2.79 $Y=1.675
+ $X2=0 $Y2=0
cc_237 N_A_523_47#_c_311_n N_A_629_47#_c_365_n 0.0207275f $X=3.48 $Y=1.16 $X2=0
+ $Y2=0
cc_238 N_A_523_47#_M1003_g N_A_629_47#_c_366_n 0.0194472f $X=3.48 $Y=0.445 $X2=0
+ $Y2=0
cc_239 N_A_523_47#_M1001_g N_VPWR_c_430_n 0.00906078f $X=3.48 $Y=2.275 $X2=0
+ $Y2=0
cc_240 N_A_523_47#_M1001_g N_VPWR_c_435_n 0.00344532f $X=3.48 $Y=2.275 $X2=0
+ $Y2=0
cc_241 N_A_523_47#_c_314_n N_VPWR_c_435_n 0.0172841f $X=2.75 $Y=1.96 $X2=0 $Y2=0
cc_242 N_A_523_47#_M1007_d N_VPWR_c_427_n 0.00382897f $X=2.615 $Y=1.485 $X2=0
+ $Y2=0
cc_243 N_A_523_47#_M1001_g N_VPWR_c_427_n 0.00545273f $X=3.48 $Y=2.275 $X2=0
+ $Y2=0
cc_244 N_A_523_47#_c_314_n N_VPWR_c_427_n 0.00955092f $X=2.75 $Y=1.96 $X2=0
+ $Y2=0
cc_245 N_A_523_47#_M1003_g N_VGND_c_508_n 0.00878516f $X=3.48 $Y=0.445 $X2=0
+ $Y2=0
cc_246 N_A_523_47#_M1003_g N_VGND_c_513_n 0.00341689f $X=3.48 $Y=0.445 $X2=0
+ $Y2=0
cc_247 N_A_523_47#_c_307_n N_VGND_c_513_n 0.0172229f $X=2.75 $Y=0.44 $X2=0 $Y2=0
cc_248 N_A_523_47#_M1005_d N_VGND_c_516_n 0.00387172f $X=2.615 $Y=0.235 $X2=0
+ $Y2=0
cc_249 N_A_523_47#_M1003_g N_VGND_c_516_n 0.00540327f $X=3.48 $Y=0.445 $X2=0
+ $Y2=0
cc_250 N_A_523_47#_c_307_n N_VGND_c_516_n 0.00953787f $X=2.75 $Y=0.44 $X2=0
+ $Y2=0
cc_251 N_A_629_47#_c_369_n N_VPWR_M1001_d 0.00207054f $X=3.56 $Y=1.942 $X2=0
+ $Y2=0
cc_252 N_A_629_47#_c_371_n N_VPWR_M1001_d 6.23798e-19 $X=3.735 $Y=1.845 $X2=0
+ $Y2=0
cc_253 N_A_629_47#_M1004_g N_VPWR_c_430_n 0.00905956f $X=3.955 $Y=1.985 $X2=0
+ $Y2=0
cc_254 N_A_629_47#_c_369_n N_VPWR_c_430_n 0.024785f $X=3.56 $Y=1.942 $X2=0 $Y2=0
cc_255 N_A_629_47#_c_368_n N_VPWR_c_435_n 0.0185923f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_256 N_A_629_47#_c_369_n N_VPWR_c_435_n 0.00261227f $X=3.56 $Y=1.942 $X2=0
+ $Y2=0
cc_257 N_A_629_47#_M1004_g N_VPWR_c_437_n 0.0046653f $X=3.955 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_A_629_47#_M1001_s N_VPWR_c_427_n 0.00230841f $X=3.145 $Y=2.065 $X2=0
+ $Y2=0
cc_259 N_A_629_47#_M1004_g N_VPWR_c_427_n 0.00897671f $X=3.955 $Y=1.985 $X2=0
+ $Y2=0
cc_260 N_A_629_47#_c_368_n N_VPWR_c_427_n 0.0102962f $X=3.27 $Y=2.275 $X2=0
+ $Y2=0
cc_261 N_A_629_47#_c_369_n N_VPWR_c_427_n 0.005846f $X=3.56 $Y=1.942 $X2=0 $Y2=0
cc_262 N_A_629_47#_M1004_g X 0.00367081f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_629_47#_c_364_n X 0.0371498f $X=3.735 $Y=1.325 $X2=0 $Y2=0
cc_264 N_A_629_47#_c_371_n X 0.0102825f $X=3.735 $Y=1.845 $X2=0 $Y2=0
cc_265 N_A_629_47#_c_365_n X 0.00767819f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_629_47#_c_366_n X 0.00366835f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_629_47#_c_364_n N_VGND_M1003_d 0.0028099f $X=3.735 $Y=1.325 $X2=0
+ $Y2=0
cc_268 N_A_629_47#_c_362_n N_VGND_c_508_n 0.00217981f $X=3.56 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_629_47#_c_364_n N_VGND_c_508_n 0.0222857f $X=3.735 $Y=1.325 $X2=0
+ $Y2=0
cc_270 N_A_629_47#_c_365_n N_VGND_c_508_n 3.47021e-19 $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_629_47#_c_366_n N_VGND_c_508_n 0.00878394f $X=3.9 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A_629_47#_c_361_n N_VGND_c_513_n 0.0184794f $X=3.27 $Y=0.44 $X2=0 $Y2=0
cc_273 N_A_629_47#_c_362_n N_VGND_c_513_n 0.00273399f $X=3.56 $Y=0.74 $X2=0
+ $Y2=0
cc_274 N_A_629_47#_c_366_n N_VGND_c_515_n 0.0046653f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A_629_47#_M1003_s N_VGND_c_516_n 0.00229009f $X=3.145 $Y=0.235 $X2=0
+ $Y2=0
cc_276 N_A_629_47#_c_361_n N_VGND_c_516_n 0.0102739f $X=3.27 $Y=0.44 $X2=0 $Y2=0
cc_277 N_A_629_47#_c_362_n N_VGND_c_516_n 0.00430392f $X=3.56 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A_629_47#_c_364_n N_VGND_c_516_n 0.00168578f $X=3.735 $Y=1.325 $X2=0
+ $Y2=0
cc_279 N_A_629_47#_c_366_n N_VGND_c_516_n 0.0090943f $X=3.9 $Y=0.995 $X2=0 $Y2=0
cc_280 N_VPWR_c_427_n N_X_M1004_d 0.00382897f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_437_n X 0.0305477f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_427_n X 0.0166756f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_283 N_X_c_491_n N_VGND_c_515_n 0.0304865f $X=4.165 $Y=0.44 $X2=0 $Y2=0
cc_284 N_X_M1008_d N_VGND_c_516_n 0.00387172f $X=4.03 $Y=0.235 $X2=0 $Y2=0
cc_285 N_X_c_491_n N_VGND_c_516_n 0.0166625f $X=4.165 $Y=0.44 $X2=0 $Y2=0

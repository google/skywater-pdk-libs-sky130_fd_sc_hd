* NGSPICE file created from sky130_fd_sc_hd__o41a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_697_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.28e+12p pd=8.56e+06u as=3.5e+11p ps=2.7e+06u
M1001 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1002 a_393_47# B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=7.3125e+11p pd=6.15e+06u as=2.08e+11p ps=1.94e+06u
M1003 VGND A4 a_393_47# VNB nshort w=650000u l=150000u
+  ad=7.9625e+11p pd=7.65e+06u as=0p ps=0u
M1004 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1005 a_79_21# B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6.05e+11p pd=3.21e+06u as=0p ps=0u
M1006 a_496_297# A4 a_79_21# VPB phighvt w=1e+06u l=150000u
+  ad=3.55e+11p pd=2.71e+06u as=0p ps=0u
M1007 a_597_297# A3 a_496_297# VPB phighvt w=1e+06u l=150000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
M1008 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_393_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_393_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_697_297# A2 a_597_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_393_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


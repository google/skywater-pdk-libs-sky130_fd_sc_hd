* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_79_21# C1 a_585_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1001 a_348_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=2.665e+11p pd=2.12e+06u as=7.8325e+11p ps=6.31e+06u
M1002 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=9.1e+11p pd=7.82e+06u as=2.7e+11p ps=2.54e+06u
M1003 a_299_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1004 VGND B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.9975e+11p ps=3.83e+06u
M1005 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_79_21# C1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A2 a_299_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_79_21# A1 a_348_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_585_297# B1 a_299_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1011 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__decap_12.spice
* Created: Thu Aug 27 14:13:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__decap_12.spice.pex"
.subckt sky130_fd_sc_hd__decap_12  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_VPWR_M1001_g N_VGND_M1001_s VNB NSHORT L=4.73 W=0.55
+ AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 M=1 R=0.116279 SA=2.365e+06
+ SB=2.365e+06 A=2.6015 P=10.56 MULT=1
MM1000 N_VPWR_M1000_s N_VGND_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=4.73 W=0.87
+ AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 M=1 R=0.183932 SA=2.365e+06
+ SB=2.365e+06 A=4.1151 P=11.2 MULT=1
DX2_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__decap_12.spice.SKY130_FD_SC_HD__DECAP_12.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_isobufsrc_4.pex.spice
* Created: Thu Aug 27 14:25:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4%SLEEP 1 3 6 8 10 13 15 17 20 22
+ 24 27 29 40 41
r79 39 41 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.62 $Y=1.16 $X2=1.75
+ $Y2=1.16
r80 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.62
+ $Y=1.16 $X2=1.62 $Y2=1.16
r81 37 39 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.62 $Y2=1.16
r82 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r83 34 36 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.6 $Y=1.16 $X2=0.91
+ $Y2=1.16
r84 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6 $Y=1.16
+ $X2=0.6 $Y2=1.16
r85 31 34 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.49 $Y=1.16 $X2=0.6
+ $Y2=1.16
r86 29 40 51.2955 $w=1.98e-07 $l=9.25e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.62 $Y2=1.175
r87 29 35 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.6 $Y2=1.175
r88 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r89 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r90 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r92 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r93 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r94 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r95 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r96 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r97 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r98 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r99 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r100 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r101 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.985
r102 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4%A_419_21# 1 2 7 9 12 14 16 19 21
+ 23 26 28 30 33 35 42 45 48 53 55 56 58 59 60
c115 59 0 1.68547e-19 $X=4.19 $Y=1.575
c116 42 0 1.86625e-19 $X=3.98 $Y=1.16
c117 19 0 7.39456e-20 $X=2.59 $Y=1.985
r118 67 68 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=3.43 $Y2=1.16
r119 63 65 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.17 $Y=1.16
+ $X2=2.59 $Y2=1.16
r120 60 68 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=1.16
+ $X2=3.43 $Y2=1.16
r121 58 59 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=1.66
+ $X2=4.19 $Y2=1.575
r122 51 58 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.19 $Y=1.74 $X2=4.19
+ $Y2=1.66
r123 51 53 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=4.19 $Y=1.74 $X2=4.19
+ $Y2=2.34
r124 49 56 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=4.15 $Y=1.275 $X2=4.15
+ $Y2=1.175
r125 49 59 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=4.15 $Y=1.275
+ $X2=4.15 $Y2=1.575
r126 48 56 4.27425 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=4.15 $Y=1.075 $X2=4.15
+ $Y2=1.175
r127 48 55 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=4.15 $Y=1.075
+ $X2=4.15 $Y2=0.815
r128 43 55 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=0.65
+ $X2=4.19 $Y2=0.815
r129 43 45 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=4.19 $Y=0.65
+ $X2=4.19 $Y2=0.39
r130 42 60 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=3.98 $Y=1.16
+ $X2=3.505 $Y2=1.16
r131 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.98
+ $Y=1.16 $X2=3.98 $Y2=1.16
r132 38 67 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.96 $Y=1.16 $X2=3.01
+ $Y2=1.16
r133 38 65 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.96 $Y=1.16
+ $X2=2.59 $Y2=1.16
r134 37 41 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=2.96 $Y=1.175
+ $X2=3.98 $Y2=1.175
r135 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.96
+ $Y=1.16 $X2=2.96 $Y2=1.16
r136 35 56 2.15711 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.025 $Y=1.175
+ $X2=4.15 $Y2=1.175
r137 35 41 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=4.025 $Y=1.175
+ $X2=3.98 $Y2=1.175
r138 31 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.16
r139 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.985
r140 28 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.16
r141 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
r142 24 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.16
r143 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.985
r144 21 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=1.16
r145 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r146 17 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.16
r147 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.985
r148 14 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.16
r149 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r150 10 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.16
r151 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.985
r152 7 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r153 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=0.56
r154 2 58 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.485 $X2=4.19 $Y2=1.66
r155 2 53 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.485 $X2=4.19 $Y2=2.34
r156 1 45 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=4.045
+ $Y=0.235 $X2=4.19 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4%A 1 3 6 8 13 19
c27 8 0 1.86625e-19 $X=4.75 $Y=1.105
r28 14 19 10.3485 $w=2.43e-07 $l=2.2e-07 $layer=LI1_cond $X=4.61 $Y=1.197
+ $X2=4.83 $Y2=1.197
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.61
+ $Y=1.16 $X2=4.61 $Y2=1.16
r30 10 13 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.4 $Y=1.16 $X2=4.61
+ $Y2=1.16
r31 8 19 0.235192 $w=2.43e-07 $l=5e-09 $layer=LI1_cond $X=4.835 $Y=1.197
+ $X2=4.83 $Y2=1.197
r32 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.4 $Y=1.325 $X2=4.4
+ $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.4 $Y=1.325 $X2=4.4
+ $Y2=1.985
r34 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.4 $Y=0.995 $X2=4.4
+ $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.4 $Y=0.995 $X2=4.4
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4%A_27_297# 1 2 3 4 5 16 18 20 24
+ 26 28 29 30 34 36 38 40 45 50
c78 28 0 7.39456e-20 $X=1.96 $Y=1.665
r79 38 52 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=2.295
+ $X2=3.665 $Y2=2.38
r80 38 40 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.665 $Y=2.295
+ $X2=3.665 $Y2=1.66
r81 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=2.38
+ $X2=2.8 $Y2=2.38
r82 36 52 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.475 $Y=2.38
+ $X2=3.665 $Y2=2.38
r83 36 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.475 $Y=2.38
+ $X2=2.965 $Y2=2.38
r84 32 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=2.295 $X2=2.8
+ $Y2=2.38
r85 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.8 $Y=2.295
+ $X2=2.8 $Y2=2.02
r86 31 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=2.38
+ $X2=1.96 $Y2=2.38
r87 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=2.38
+ $X2=2.8 $Y2=2.38
r88 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.635 $Y=2.38
+ $X2=2.125 $Y2=2.38
r89 29 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=2.295 $X2=1.96
+ $Y2=2.38
r90 28 47 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=1.56
r91 28 29 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=2.295
r92 27 45 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.56 $X2=1.12
+ $Y2=1.56
r93 26 47 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=1.56
+ $X2=1.96 $Y2=1.56
r94 26 27 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=1.795 $Y=1.56
+ $X2=1.205 $Y2=1.56
r95 22 45 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.56
r96 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=2.3
r97 21 43 3.99943 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.56
+ $X2=0.225 $Y2=1.56
r98 20 45 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=1.56 $X2=1.12
+ $Y2=1.56
r99 20 21 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.035 $Y=1.56
+ $X2=0.365 $Y2=1.56
r100 16 43 2.99957 $w=2.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=1.56
r101 16 18 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=2.3
r102 5 52 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=2.34
r103 5 40 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=1.66
r104 4 34 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=2.02
r105 3 49 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.34
r106 3 47 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r107 2 45 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r108 2 24 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r109 1 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r110 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4%VPWR 1 2 3 12 16 18 20 24 26 31
+ 36 42 45 49
r66 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r67 45 46 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 40 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r70 40 46 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=1.61 $Y2=2.72
r71 39 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r72 37 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=1.5 $Y2=2.72
r73 37 39 179.086 $w=1.68e-07 $l=2.745e-06 $layer=LI1_cond $X=1.625 $Y=2.72
+ $X2=4.37 $Y2=2.72
r74 36 48 5.38769 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.525 $Y=2.72
+ $X2=4.792 $Y2=2.72
r75 36 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.525 $Y=2.72
+ $X2=4.37 $Y2=2.72
r76 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 35 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.7 $Y2=2.72
r80 32 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=1.15 $Y2=2.72
r81 31 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.5 $Y2=2.72
r82 31 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 26 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.7 $Y2=2.72
r84 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 24 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r87 20 23 19.3497 $w=4.03e-07 $l=6.8e-07 $layer=LI1_cond $X=4.727 $Y=1.66
+ $X2=4.727 $Y2=2.34
r88 18 48 3.02679 $w=4.05e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.727 $Y=2.635
+ $X2=4.792 $Y2=2.72
r89 18 23 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=4.727 $Y=2.635
+ $X2=4.727 $Y2=2.34
r90 14 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=2.635
+ $X2=1.5 $Y2=2.72
r91 14 16 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.5 $Y=2.635
+ $X2=1.5 $Y2=2
r92 10 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2.72
r93 10 12 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2
r94 3 23 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.485 $X2=4.61 $Y2=2.34
r95 3 20 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.485 $X2=4.61 $Y2=1.66
r96 2 16 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=2
r97 1 12 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4%X 1 2 3 4 5 6 21 23 24 27 29 33
+ 36 39 41 45 47 49 51 52 55 56 59
r110 56 59 5.37807 $w=2.98e-07 $l=1.4e-07 $layer=LI1_cond $X=3.135 $Y=1.595
+ $X2=2.995 $Y2=1.595
r111 56 58 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=1.595
+ $X2=3.22 $Y2=1.595
r112 53 59 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=1.595
+ $X2=2.995 $Y2=1.595
r113 53 55 0.695019 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=1.595
+ $X2=2.46 $Y2=1.595
r114 47 58 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.22 $Y=1.745
+ $X2=3.22 $Y2=1.595
r115 47 49 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.22 $Y=1.745
+ $X2=3.22 $Y2=1.96
r116 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.39
r117 42 52 5.06882 $w=1.8e-07 $l=2.05e-07 $layer=LI1_cond $X=2.625 $Y=0.815
+ $X2=2.42 $Y2=0.815
r118 41 43 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=3.22 $Y2=0.725
r119 41 42 26.4949 $w=1.78e-07 $l=4.3e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=2.625 $Y2=0.815
r120 37 55 5.99569 $w=2.5e-07 $l=1.85742e-07 $layer=LI1_cond $X=2.38 $Y=1.745
+ $X2=2.46 $Y2=1.595
r121 37 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.38 $Y=1.745
+ $X2=2.38 $Y2=1.96
r122 36 55 5.99569 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=2.46 $Y=1.445
+ $X2=2.46 $Y2=1.595
r123 35 52 1.4294 $w=3.3e-07 $l=1.08167e-07 $layer=LI1_cond $X=2.46 $Y=0.905
+ $X2=2.42 $Y2=0.815
r124 35 36 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.46 $Y=0.905
+ $X2=2.46 $Y2=1.445
r125 31 52 1.4294 $w=3.3e-07 $l=1.08167e-07 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.42 $Y2=0.815
r126 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.39
r127 30 51 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r128 29 52 5.06882 $w=1.8e-07 $l=2.05e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=2.42 $Y2=0.815
r129 29 30 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=1.705 $Y2=0.815
r130 25 51 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.815
r131 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r132 23 51 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r133 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r134 19 24 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r135 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.7 $Y2=0.39
r136 6 58 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.62
r137 6 49 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=1.96
r138 5 55 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.62
r139 5 39 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=1.96
r140 4 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.39
r141 3 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.39
r142 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r143 1 21 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_4%VGND 1 2 3 4 5 6 19 21 25 29 33
+ 37 39 41 44 45 47 48 50 51 53 54 55 70 79
r87 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r88 73 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r89 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r90 70 78 4.18967 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.525 $Y=0 $X2=4.792
+ $Y2=0
r91 70 72 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.525 $Y=0 $X2=4.37
+ $Y2=0
r92 69 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r93 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r94 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r95 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r96 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r97 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r98 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r99 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r100 57 75 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r101 57 59 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.69 $Y2=0
r102 55 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r103 55 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r104 53 68 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.45 $Y2=0
r105 53 54 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.7
+ $Y2=0
r106 52 72 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.845 $Y=0
+ $X2=4.37 $Y2=0
r107 52 54 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.845 $Y=0 $X2=3.7
+ $Y2=0
r108 50 65 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0
+ $X2=2.53 $Y2=0
r109 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.8
+ $Y2=0
r110 49 68 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.45
+ $Y2=0
r111 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.8
+ $Y2=0
r112 47 62 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r113 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r114 46 65 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.53 $Y2=0
r115 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r116 44 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r117 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r118 43 62 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.61 $Y2=0
r119 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r120 39 78 3.24817 $w=2.9e-07 $l=1.58915e-07 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.792 $Y2=0
r121 39 41 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0.39
r122 35 54 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r123 35 37 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.39
r124 31 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r125 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.39
r126 27 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r127 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r128 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r129 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r130 19 75 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.182 $Y2=0
r131 19 21 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.39
r132 6 41 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.475
+ $Y=0.235 $X2=4.61 $Y2=0.39
r133 5 37 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.39
r134 4 33 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.39
r135 3 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r136 2 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r137 1 21 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__inv_2.pxi.spice
* Created: Thu Aug 27 14:22:39 2020
* 
x_PM_SKY130_FD_SC_HD__INV_2%A N_A_c_24_n N_A_M1001_g N_A_M1000_g N_A_c_25_n
+ N_A_M1003_g N_A_M1002_g A N_A_c_27_n PM_SKY130_FD_SC_HD__INV_2%A
x_PM_SKY130_FD_SC_HD__INV_2%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_c_61_n
+ N_VPWR_c_62_n N_VPWR_c_63_n N_VPWR_c_64_n VPWR N_VPWR_c_65_n N_VPWR_c_60_n
+ PM_SKY130_FD_SC_HD__INV_2%VPWR
x_PM_SKY130_FD_SC_HD__INV_2%Y N_Y_M1001_d N_Y_M1000_s N_Y_c_81_n N_Y_c_83_n Y Y
+ Y Y Y PM_SKY130_FD_SC_HD__INV_2%Y
x_PM_SKY130_FD_SC_HD__INV_2%VGND N_VGND_M1001_s N_VGND_M1003_s N_VGND_c_101_n
+ N_VGND_c_102_n N_VGND_c_103_n N_VGND_c_104_n VGND N_VGND_c_105_n
+ N_VGND_c_106_n PM_SKY130_FD_SC_HD__INV_2%VGND
cc_1 VNB N_A_c_24_n 0.0214124f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_2 VNB N_A_c_25_n 0.0209918f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.995
cc_3 VNB A 0.00854082f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_c_27_n 0.0683249f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.16
cc_5 VNB N_VPWR_c_60_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB Y 9.8125e-19 $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_7 VNB N_VGND_c_101_n 0.010609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_VGND_c_102_n 0.030306f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=0.56
cc_9 VNB N_VGND_c_103_n 0.0108622f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.325
cc_10 VNB N_VGND_c_104_n 0.00872689f $X=-0.19 $Y=-0.24 $X2=0.9 $Y2=1.985
cc_11 VNB N_VGND_c_105_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_12 VNB N_VGND_c_106_n 0.106998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VPB N_A_M1000_g 0.0259172f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_14 VPB N_A_M1002_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_15 VPB A 7.08627e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_16 VPB N_A_c_27_n 0.0152489f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.16
cc_17 VPB N_VPWR_c_61_n 0.0105831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_62_n 0.0404906f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=0.56
cc_19 VPB N_VPWR_c_63_n 0.0108363f $X=-0.19 $Y=1.305 $X2=0.9 $Y2=1.985
cc_20 VPB N_VPWR_c_64_n 0.00438892f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_21 VPB N_VPWR_c_65_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_22 VPB N_VPWR_c_60_n 0.0460103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB Y 0.00151227f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_24 N_A_M1000_g N_VPWR_c_62_n 0.00320188f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_25 A N_VPWR_c_62_n 0.0182344f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_26 N_A_c_27_n N_VPWR_c_62_n 0.00529313f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_27 N_A_M1002_g N_VPWR_c_64_n 0.0031902f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_28 N_A_M1000_g N_VPWR_c_65_n 0.00541359f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_29 N_A_M1002_g N_VPWR_c_65_n 0.00541359f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_30 N_A_M1000_g N_VPWR_c_60_n 0.0104652f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_31 N_A_M1002_g N_VPWR_c_60_n 0.0104652f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_32 N_A_c_24_n N_Y_c_81_n 0.00534153f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_33 N_A_c_25_n N_Y_c_81_n 0.00534153f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_34 N_A_M1000_g N_Y_c_83_n 0.00918977f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_35 N_A_M1002_g N_Y_c_83_n 0.00918977f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_36 N_A_c_24_n Y 0.00503194f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_37 N_A_M1000_g Y 0.00408533f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_38 N_A_c_25_n Y 0.00675111f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_39 N_A_M1002_g Y 0.00809641f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_40 A Y 0.0183187f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_41 N_A_c_27_n Y 0.0322431f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_42 N_A_M1000_g Y 0.002888f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_43 N_A_M1002_g Y 0.00214168f $X=0.9 $Y=1.985 $X2=0 $Y2=0
cc_44 N_A_c_24_n N_VGND_c_102_n 0.00366806f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_45 A N_VGND_c_102_n 0.0188678f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_46 N_A_c_27_n N_VGND_c_102_n 0.00585411f $X=0.9 $Y=1.16 $X2=0 $Y2=0
cc_47 N_A_c_25_n N_VGND_c_104_n 0.00363144f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_48 N_A_c_24_n N_VGND_c_105_n 0.00541359f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_49 N_A_c_25_n N_VGND_c_105_n 0.00541359f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_50 N_A_c_24_n N_VGND_c_106_n 0.0104652f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_51 N_A_c_25_n N_VGND_c_106_n 0.0104652f $X=0.9 $Y=0.995 $X2=0 $Y2=0
cc_52 N_VPWR_c_60_n N_Y_M1000_s 0.00215201f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_53 N_VPWR_c_65_n N_Y_c_83_n 0.0189039f $X=1.025 $Y=2.72 $X2=0 $Y2=0
cc_54 N_VPWR_c_60_n N_Y_c_83_n 0.0122217f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_55 N_VPWR_c_64_n N_VGND_c_104_n 0.00765463f $X=1.11 $Y=1.66 $X2=0 $Y2=0
cc_56 Y N_VGND_c_102_n 0.00115029f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_57 N_Y_c_81_n N_VGND_c_104_n 0.025023f $X=0.69 $Y=0.38 $X2=0 $Y2=0
cc_58 N_Y_c_81_n N_VGND_c_105_n 0.0188933f $X=0.69 $Y=0.38 $X2=0 $Y2=0
cc_59 N_Y_M1001_d N_VGND_c_106_n 0.00215201f $X=0.555 $Y=0.235 $X2=0 $Y2=0
cc_60 N_Y_c_81_n N_VGND_c_106_n 0.0122158f $X=0.69 $Y=0.38 $X2=0 $Y2=0

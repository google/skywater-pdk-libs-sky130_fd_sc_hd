* File: sky130_fd_sc_hd__a2bb2o_1.pxi.spice
* Created: Thu Aug 27 14:03:10 2020
* 
x_PM_SKY130_FD_SC_HD__A2BB2O_1%A_76_199# N_A_76_199#_M1001_d N_A_76_199#_M1002_s
+ N_A_76_199#_M1011_g N_A_76_199#_M1005_g N_A_76_199#_c_87_n N_A_76_199#_c_88_n
+ N_A_76_199#_c_145_p N_A_76_199#_c_89_n N_A_76_199#_c_90_n N_A_76_199#_c_91_n
+ N_A_76_199#_c_80_n N_A_76_199#_c_81_n N_A_76_199#_c_82_n N_A_76_199#_c_83_n
+ N_A_76_199#_c_94_n N_A_76_199#_c_84_n N_A_76_199#_c_85_n
+ PM_SKY130_FD_SC_HD__A2BB2O_1%A_76_199#
x_PM_SKY130_FD_SC_HD__A2BB2O_1%A1_N N_A1_N_M1009_g N_A1_N_M1010_g A1_N A1_N
+ N_A1_N_c_178_n N_A1_N_c_179_n PM_SKY130_FD_SC_HD__A2BB2O_1%A1_N
x_PM_SKY130_FD_SC_HD__A2BB2O_1%A2_N N_A2_N_c_213_n N_A2_N_M1000_g N_A2_N_M1007_g
+ A2_N PM_SKY130_FD_SC_HD__A2BB2O_1%A2_N
x_PM_SKY130_FD_SC_HD__A2BB2O_1%A_226_47# N_A_226_47#_M1009_d N_A_226_47#_M1000_d
+ N_A_226_47#_M1001_g N_A_226_47#_c_248_n N_A_226_47#_M1002_g
+ N_A_226_47#_c_250_n N_A_226_47#_c_303_p N_A_226_47#_c_244_n
+ N_A_226_47#_c_245_n N_A_226_47#_c_251_n N_A_226_47#_c_252_n
+ N_A_226_47#_c_246_n N_A_226_47#_c_254_n N_A_226_47#_c_247_n
+ PM_SKY130_FD_SC_HD__A2BB2O_1%A_226_47#
x_PM_SKY130_FD_SC_HD__A2BB2O_1%B2 N_B2_M1004_g N_B2_M1008_g B2 N_B2_c_313_n
+ N_B2_c_314_n PM_SKY130_FD_SC_HD__A2BB2O_1%B2
x_PM_SKY130_FD_SC_HD__A2BB2O_1%B1 N_B1_M1003_g N_B1_M1006_g B1 B1 B1
+ N_B1_c_360_n PM_SKY130_FD_SC_HD__A2BB2O_1%B1
x_PM_SKY130_FD_SC_HD__A2BB2O_1%X N_X_M1011_s N_X_M1005_s N_X_c_388_n N_X_c_391_n
+ N_X_c_389_n X X X N_X_c_393_n PM_SKY130_FD_SC_HD__A2BB2O_1%X
x_PM_SKY130_FD_SC_HD__A2BB2O_1%VPWR N_VPWR_M1005_d N_VPWR_M1008_d N_VPWR_c_406_n
+ N_VPWR_c_407_n VPWR VPWR N_VPWR_c_408_n VPWR N_VPWR_c_409_n N_VPWR_c_410_n
+ N_VPWR_c_405_n N_VPWR_c_412_n N_VPWR_c_413_n PM_SKY130_FD_SC_HD__A2BB2O_1%VPWR
x_PM_SKY130_FD_SC_HD__A2BB2O_1%A_489_413# N_A_489_413#_M1002_d
+ N_A_489_413#_M1006_d N_A_489_413#_c_459_n N_A_489_413#_c_460_n
+ N_A_489_413#_c_461_n N_A_489_413#_c_462_n N_A_489_413#_c_468_n
+ PM_SKY130_FD_SC_HD__A2BB2O_1%A_489_413#
x_PM_SKY130_FD_SC_HD__A2BB2O_1%VGND N_VGND_M1011_d N_VGND_M1007_d N_VGND_M1003_d
+ N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n VGND VGND N_VGND_c_495_n VGND
+ N_VGND_c_496_n N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n
+ PM_SKY130_FD_SC_HD__A2BB2O_1%VGND
cc_1 VNB N_A_76_199#_c_80_n 0.0038174f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=1.895
cc_2 VNB N_A_76_199#_c_81_n 0.00126861f $X=-0.19 $Y=-0.24 $X2=2.495 $Y2=0.445
cc_3 VNB N_A_76_199#_c_82_n 0.00405192f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_4 VNB N_A_76_199#_c_83_n 0.0229624f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_5 VNB N_A_76_199#_c_84_n 0.0090512f $X=-0.19 $Y=-0.24 $X2=2.495 $Y2=0.785
cc_6 VNB N_A_76_199#_c_85_n 0.0205627f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=0.995
cc_7 VNB N_A1_N_M1009_g 0.0314275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_N_c_178_n 0.0208395f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.325
cc_9 VNB N_A1_N_c_179_n 0.00632248f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.805
cc_10 VNB N_A2_N_c_213_n 0.0210975f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=0.235
cc_11 VNB N_A2_N_M1007_g 0.0291169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A2_N 0.00256217f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_A_226_47#_c_244_n 0.0106281f $X=-0.19 $Y=-0.24 $X2=2.495 $Y2=0.7
cc_14 VNB N_A_226_47#_c_245_n 0.00674176f $X=-0.19 $Y=-0.24 $X2=2.495 $Y2=0.445
cc_15 VNB N_A_226_47#_c_246_n 0.0566535f $X=-0.19 $Y=-0.24 $X2=0.557 $Y2=1.325
cc_16 VNB N_A_226_47#_c_247_n 0.0182811f $X=-0.19 $Y=-0.24 $X2=2.495 $Y2=0.785
cc_17 VNB N_B2_M1004_g 0.0454671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B2_c_313_n 0.00452246f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.325
cc_19 VNB N_B2_c_314_n 0.0100925f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=2.285
cc_20 VNB N_B1_M1003_g 0.0328058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB B1 0.0236663f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_22 VNB N_B1_c_360_n 0.0392237f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=1.89
cc_23 VNB N_X_c_388_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_24 VNB N_X_c_389_n 0.0225917f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_25 VNB X 0.016472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_405_n 0.155873f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=2.275
cc_27 VNB N_VGND_c_492_n 0.00271435f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_28 VNB N_VGND_c_493_n 0.0125248f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.325
cc_29 VNB N_VGND_c_494_n 0.0192404f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=1.89
cc_30 VNB N_VGND_c_495_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=2.315 $Y2=0.87
cc_31 VNB N_VGND_c_496_n 0.0246972f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=2.275
cc_32 VNB N_VGND_c_497_n 0.00699789f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_33 VNB N_VGND_c_498_n 0.0148665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_499_n 0.0134177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_500_n 0.20045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A_76_199#_M1005_g 0.0240088f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A_76_199#_c_87_n 0.00111481f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.805
cc_38 VPB N_A_76_199#_c_88_n 0.00311328f $X=-0.19 $Y=1.305 $X2=1.105 $Y2=1.89
cc_39 VPB N_A_76_199#_c_89_n 0.00838989f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=2.2
cc_40 VPB N_A_76_199#_c_90_n 0.0216647f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=2.285
cc_41 VPB N_A_76_199#_c_91_n 0.00416782f $X=-0.19 $Y=1.305 $X2=1.275 $Y2=2.285
cc_42 VPB N_A_76_199#_c_80_n 0.00345937f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.895
cc_43 VPB N_A_76_199#_c_83_n 0.00500576f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_44 VPB N_A_76_199#_c_94_n 0.0152984f $X=-0.19 $Y=1.305 $X2=2.16 $Y2=2.275
cc_45 VPB N_A1_N_M1010_g 0.01833f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_46 VPB N_A1_N_c_178_n 0.0046179f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.325
cc_47 VPB N_A1_N_c_179_n 0.00266137f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.805
cc_48 VPB N_A2_N_c_213_n 0.0271735f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=0.235
cc_49 VPB A2_N 0.00182103f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_50 VPB N_A_226_47#_c_248_n 0.0191389f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_51 VPB N_A_226_47#_M1002_g 0.0233374f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.325
cc_52 VPB N_A_226_47#_c_250_n 0.0173549f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=1.975
cc_53 VPB N_A_226_47#_c_251_n 0.00952294f $X=-0.19 $Y=1.305 $X2=2.495 $Y2=0.445
cc_54 VPB N_A_226_47#_c_252_n 0.00187459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_226_47#_c_246_n 0.022381f $X=-0.19 $Y=1.305 $X2=0.557 $Y2=1.325
cc_56 VPB N_A_226_47#_c_254_n 0.00173986f $X=-0.19 $Y=1.305 $X2=2.195 $Y2=2.285
cc_57 VPB N_B2_M1008_g 0.0313625f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_58 VPB B2 0.00852446f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_59 VPB N_B2_c_313_n 0.025717f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.325
cc_60 VPB N_B2_c_314_n 8.17517e-19 $X=-0.19 $Y=1.305 $X2=1.99 $Y2=2.285
cc_61 VPB N_B1_M1006_g 0.0611811f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_62 VPB B1 0.0162554f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_63 VPB N_B1_c_360_n 0.00784466f $X=-0.19 $Y=1.305 $X2=1.105 $Y2=1.89
cc_64 VPB N_X_c_391_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_65 VPB N_X_c_389_n 0.00991797f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_66 VPB N_X_c_393_n 0.0311049f $X=-0.19 $Y=1.305 $X2=2.495 $Y2=0.7
cc_67 VPB N_VPWR_c_406_n 0.00923837f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_68 VPB N_VPWR_c_407_n 0.00232023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_408_n 0.0150576f $X=-0.19 $Y=1.305 $X2=1.19 $Y2=2.2
cc_70 VPB N_VPWR_c_409_n 0.051396f $X=-0.19 $Y=1.305 $X2=2.495 $Y2=0.445
cc_71 VPB N_VPWR_c_410_n 0.0151573f $X=-0.19 $Y=1.305 $X2=2.195 $Y2=2.275
cc_72 VPB N_VPWR_c_405_n 0.056706f $X=-0.19 $Y=1.305 $X2=2.16 $Y2=2.275
cc_73 VPB N_VPWR_c_412_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_413_n 0.0035381f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_75 VPB N_A_489_413#_c_459_n 3.5109e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_76 VPB N_A_489_413#_c_460_n 0.0148879f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_77 VPB N_A_489_413#_c_461_n 0.00277544f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_78 VPB N_A_489_413#_c_462_n 0.00261535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 N_A_76_199#_c_85_n N_A1_N_M1009_g 0.0182272f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_76_199#_M1005_g N_A1_N_M1010_g 0.0168573f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_76_199#_c_87_n N_A1_N_M1010_g 0.00451623f $X=0.6 $Y=1.805 $X2=0 $Y2=0
cc_82 N_A_76_199#_c_88_n N_A1_N_M1010_g 0.0103819f $X=1.105 $Y=1.89 $X2=0 $Y2=0
cc_83 N_A_76_199#_c_89_n N_A1_N_M1010_g 0.00195951f $X=1.19 $Y=2.2 $X2=0 $Y2=0
cc_84 N_A_76_199#_c_88_n N_A1_N_c_178_n 0.00156259f $X=1.105 $Y=1.89 $X2=0 $Y2=0
cc_85 N_A_76_199#_c_82_n N_A1_N_c_178_n 0.00197826f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_76_199#_c_83_n N_A1_N_c_178_n 0.0203259f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_76_199#_M1005_g N_A1_N_c_179_n 8.79726e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_88 N_A_76_199#_c_88_n N_A1_N_c_179_n 0.0156175f $X=1.105 $Y=1.89 $X2=0 $Y2=0
cc_89 N_A_76_199#_c_82_n N_A1_N_c_179_n 0.0392215f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_76_199#_c_83_n N_A1_N_c_179_n 3.61509e-19 $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_76_199#_c_88_n N_A2_N_c_213_n 0.003006f $X=1.105 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_76_199#_c_89_n N_A2_N_c_213_n 0.00133815f $X=1.19 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_76_199#_c_90_n N_A2_N_c_213_n 0.00625967f $X=1.99 $Y=2.285 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_76_199#_c_94_n N_A2_N_c_213_n 0.00353563f $X=2.16 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_76_199#_c_80_n N_A_226_47#_c_248_n 0.00741354f $X=2.315 $Y=1.895 $X2=0
+ $Y2=0
cc_96 N_A_76_199#_c_94_n N_A_226_47#_M1002_g 0.00815975f $X=2.16 $Y=2.275 $X2=0
+ $Y2=0
cc_97 N_A_76_199#_c_80_n N_A_226_47#_c_250_n 0.00656604f $X=2.315 $Y=1.895 $X2=0
+ $Y2=0
cc_98 N_A_76_199#_c_94_n N_A_226_47#_c_250_n 0.00309485f $X=2.16 $Y=2.275 $X2=0
+ $Y2=0
cc_99 N_A_76_199#_c_81_n N_A_226_47#_c_244_n 0.00227074f $X=2.495 $Y=0.445 $X2=0
+ $Y2=0
cc_100 N_A_76_199#_c_84_n N_A_226_47#_c_244_n 0.010242f $X=2.495 $Y=0.785 $X2=0
+ $Y2=0
cc_101 N_A_76_199#_c_90_n N_A_226_47#_c_251_n 0.0105401f $X=1.99 $Y=2.285 $X2=0
+ $Y2=0
cc_102 N_A_76_199#_c_80_n N_A_226_47#_c_251_n 0.0129713f $X=2.315 $Y=1.895 $X2=0
+ $Y2=0
cc_103 N_A_76_199#_c_94_n N_A_226_47#_c_251_n 0.00621416f $X=2.16 $Y=2.275 $X2=0
+ $Y2=0
cc_104 N_A_76_199#_c_80_n N_A_226_47#_c_252_n 0.0460919f $X=2.315 $Y=1.895 $X2=0
+ $Y2=0
cc_105 N_A_76_199#_c_84_n N_A_226_47#_c_252_n 0.00313949f $X=2.495 $Y=0.785
+ $X2=0 $Y2=0
cc_106 N_A_76_199#_c_80_n N_A_226_47#_c_246_n 0.0170253f $X=2.315 $Y=1.895 $X2=0
+ $Y2=0
cc_107 N_A_76_199#_c_94_n N_A_226_47#_c_246_n 0.00547327f $X=2.16 $Y=2.275 $X2=0
+ $Y2=0
cc_108 N_A_76_199#_c_84_n N_A_226_47#_c_246_n 0.0040021f $X=2.495 $Y=0.785 $X2=0
+ $Y2=0
cc_109 N_A_76_199#_c_90_n N_A_226_47#_c_254_n 0.00792284f $X=1.99 $Y=2.285 $X2=0
+ $Y2=0
cc_110 N_A_76_199#_c_80_n N_A_226_47#_c_254_n 0.00530118f $X=2.315 $Y=1.895
+ $X2=0 $Y2=0
cc_111 N_A_76_199#_c_94_n N_A_226_47#_c_254_n 5.57416e-19 $X=2.16 $Y=2.275 $X2=0
+ $Y2=0
cc_112 N_A_76_199#_c_81_n N_A_226_47#_c_247_n 4.8064e-19 $X=2.495 $Y=0.445 $X2=0
+ $Y2=0
cc_113 N_A_76_199#_c_84_n N_A_226_47#_c_247_n 0.00476789f $X=2.495 $Y=0.785
+ $X2=0 $Y2=0
cc_114 N_A_76_199#_c_80_n N_B2_M1004_g 0.00355563f $X=2.315 $Y=1.895 $X2=0 $Y2=0
cc_115 N_A_76_199#_c_81_n N_B2_M1004_g 0.00111676f $X=2.495 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_76_199#_c_84_n N_B2_M1004_g 0.00266107f $X=2.495 $Y=0.785 $X2=0 $Y2=0
cc_117 N_A_76_199#_c_80_n N_B2_M1008_g 0.00238676f $X=2.315 $Y=1.895 $X2=0 $Y2=0
cc_118 N_A_76_199#_c_80_n B2 0.0217994f $X=2.315 $Y=1.895 $X2=0 $Y2=0
cc_119 N_A_76_199#_c_80_n N_B2_c_313_n 8.3553e-19 $X=2.315 $Y=1.895 $X2=0 $Y2=0
cc_120 N_A_76_199#_c_80_n N_B2_c_314_n 0.0199037f $X=2.315 $Y=1.895 $X2=0 $Y2=0
cc_121 N_A_76_199#_c_84_n N_B2_c_314_n 0.00673007f $X=2.495 $Y=0.785 $X2=0 $Y2=0
cc_122 N_A_76_199#_M1005_g N_X_c_389_n 0.00417382f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_76_199#_c_87_n N_X_c_389_n 0.010489f $X=0.6 $Y=1.805 $X2=0 $Y2=0
cc_124 N_A_76_199#_c_82_n N_X_c_389_n 0.0243753f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_76_199#_c_83_n N_X_c_389_n 0.00753785f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_76_199#_c_85_n N_X_c_389_n 0.00656531f $X=0.515 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_76_199#_c_87_n N_VPWR_M1005_d 0.00369532f $X=0.6 $Y=1.805 $X2=-0.19
+ $Y2=-0.24
cc_128 N_A_76_199#_c_88_n N_VPWR_M1005_d 0.00971438f $X=1.105 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A_76_199#_c_145_p N_VPWR_M1005_d 0.00106957f $X=0.685 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_76_199#_M1005_g N_VPWR_c_406_n 0.00977218f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_76_199#_c_88_n N_VPWR_c_406_n 0.00867614f $X=1.105 $Y=1.89 $X2=0
+ $Y2=0
cc_132 N_A_76_199#_c_145_p N_VPWR_c_406_n 0.00642951f $X=0.685 $Y=1.89 $X2=0
+ $Y2=0
cc_133 N_A_76_199#_c_91_n N_VPWR_c_406_n 0.00887201f $X=1.275 $Y=2.285 $X2=0
+ $Y2=0
cc_134 N_A_76_199#_M1005_g N_VPWR_c_408_n 0.0046653f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_76_199#_c_88_n N_VPWR_c_409_n 0.00357178f $X=1.105 $Y=1.89 $X2=0
+ $Y2=0
cc_136 N_A_76_199#_c_90_n N_VPWR_c_409_n 0.028843f $X=1.99 $Y=2.285 $X2=0 $Y2=0
cc_137 N_A_76_199#_c_91_n N_VPWR_c_409_n 0.00749299f $X=1.275 $Y=2.285 $X2=0
+ $Y2=0
cc_138 N_A_76_199#_c_94_n N_VPWR_c_409_n 0.0202509f $X=2.16 $Y=2.275 $X2=0 $Y2=0
cc_139 N_A_76_199#_M1002_s N_VPWR_c_405_n 0.0022974f $X=2.035 $Y=2.065 $X2=0
+ $Y2=0
cc_140 N_A_76_199#_M1005_g N_VPWR_c_405_n 0.00895857f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_76_199#_c_88_n N_VPWR_c_405_n 0.00736589f $X=1.105 $Y=1.89 $X2=0
+ $Y2=0
cc_142 N_A_76_199#_c_145_p N_VPWR_c_405_n 8.6225e-19 $X=0.685 $Y=1.89 $X2=0
+ $Y2=0
cc_143 N_A_76_199#_c_90_n N_VPWR_c_405_n 0.0250414f $X=1.99 $Y=2.285 $X2=0 $Y2=0
cc_144 N_A_76_199#_c_91_n N_VPWR_c_405_n 0.00618211f $X=1.275 $Y=2.285 $X2=0
+ $Y2=0
cc_145 N_A_76_199#_c_94_n N_VPWR_c_405_n 0.0138272f $X=2.16 $Y=2.275 $X2=0 $Y2=0
cc_146 N_A_76_199#_c_88_n A_226_297# 0.00320261f $X=1.105 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_76_199#_c_94_n N_A_489_413#_c_459_n 0.00447001f $X=2.16 $Y=2.275
+ $X2=0 $Y2=0
cc_148 N_A_76_199#_c_80_n N_A_489_413#_c_461_n 0.00470312f $X=2.315 $Y=1.895
+ $X2=0 $Y2=0
cc_149 N_A_76_199#_c_94_n N_A_489_413#_c_461_n 0.0092171f $X=2.16 $Y=2.275 $X2=0
+ $Y2=0
cc_150 N_A_76_199#_c_82_n N_VGND_c_492_n 0.00551674f $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_76_199#_c_83_n N_VGND_c_492_n 4.58244e-19 $X=0.515 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_76_199#_c_85_n N_VGND_c_492_n 0.0100539f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_76_199#_c_85_n N_VGND_c_495_n 0.0046653f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_A_76_199#_c_81_n N_VGND_c_496_n 0.0110645f $X=2.495 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_A_76_199#_c_84_n N_VGND_c_496_n 0.00251982f $X=2.495 $Y=0.785 $X2=0
+ $Y2=0
cc_156 N_A_76_199#_c_84_n N_VGND_c_499_n 5.80399e-19 $X=2.495 $Y=0.785 $X2=0
+ $Y2=0
cc_157 N_A_76_199#_M1001_d N_VGND_c_500_n 0.00413042f $X=2.36 $Y=0.235 $X2=0
+ $Y2=0
cc_158 N_A_76_199#_c_81_n N_VGND_c_500_n 0.00640047f $X=2.495 $Y=0.445 $X2=0
+ $Y2=0
cc_159 N_A_76_199#_c_84_n N_VGND_c_500_n 0.00407678f $X=2.495 $Y=0.785 $X2=0
+ $Y2=0
cc_160 N_A_76_199#_c_85_n N_VGND_c_500_n 0.00895857f $X=0.515 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A1_N_c_178_n N_A2_N_c_213_n 0.0604884f $X=0.995 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A1_N_c_179_n N_A2_N_c_213_n 0.00503544f $X=0.995 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_163 N_A1_N_M1009_g N_A2_N_M1007_g 0.0240597f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A1_N_c_178_n A2_N 3.51879e-19 $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A1_N_c_179_n A2_N 0.0297809f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_N_M1009_g N_A_226_47#_c_245_n 0.00536216f $X=1.055 $Y=0.445 $X2=0
+ $Y2=0
cc_167 N_A1_N_c_179_n N_A_226_47#_c_245_n 0.00541889f $X=0.995 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A1_N_c_179_n N_A_226_47#_c_252_n 0.00495338f $X=0.995 $Y=1.16 $X2=0
+ $Y2=0
cc_169 N_A1_N_c_179_n N_VPWR_M1005_d 0.00147965f $X=0.995 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A1_N_M1010_g N_VPWR_c_409_n 0.00226132f $X=1.055 $Y=1.695 $X2=0 $Y2=0
cc_171 N_A1_N_M1010_g N_VPWR_c_405_n 0.00349386f $X=1.055 $Y=1.695 $X2=0 $Y2=0
cc_172 N_A1_N_c_179_n A_226_297# 0.0022049f $X=0.995 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_173 N_A1_N_M1009_g N_VGND_c_492_n 0.00364237f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_174 N_A1_N_c_178_n N_VGND_c_492_n 0.00176065f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A1_N_c_179_n N_VGND_c_492_n 8.57019e-19 $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A1_N_M1009_g N_VGND_c_498_n 0.00585385f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A1_N_M1009_g N_VGND_c_499_n 5.89496e-19 $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A1_N_M1009_g N_VGND_c_500_n 0.0110737f $X=1.055 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A2_N_c_213_n N_A_226_47#_c_248_n 0.0025391f $X=1.415 $Y=1.375 $X2=0
+ $Y2=0
cc_180 N_A2_N_c_213_n N_A_226_47#_c_244_n 0.00377055f $X=1.415 $Y=1.375 $X2=0
+ $Y2=0
cc_181 N_A2_N_M1007_g N_A_226_47#_c_244_n 0.0121989f $X=1.475 $Y=0.445 $X2=0
+ $Y2=0
cc_182 A2_N N_A_226_47#_c_244_n 0.0218033f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_183 N_A2_N_c_213_n N_A_226_47#_c_245_n 3.76221e-19 $X=1.415 $Y=1.375 $X2=0
+ $Y2=0
cc_184 N_A2_N_c_213_n N_A_226_47#_c_252_n 0.00149507f $X=1.415 $Y=1.375 $X2=0
+ $Y2=0
cc_185 N_A2_N_M1007_g N_A_226_47#_c_252_n 9.56524e-19 $X=1.475 $Y=0.445 $X2=0
+ $Y2=0
cc_186 A2_N N_A_226_47#_c_252_n 0.0260982f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A2_N_c_213_n N_A_226_47#_c_246_n 0.0254182f $X=1.415 $Y=1.375 $X2=0
+ $Y2=0
cc_188 N_A2_N_M1007_g N_A_226_47#_c_246_n 0.0108133f $X=1.475 $Y=0.445 $X2=0
+ $Y2=0
cc_189 A2_N N_A_226_47#_c_246_n 0.00253557f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_190 N_A2_N_c_213_n N_A_226_47#_c_254_n 7.48305e-19 $X=1.415 $Y=1.375 $X2=0
+ $Y2=0
cc_191 A2_N N_A_226_47#_c_254_n 0.013002f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_192 N_A2_N_M1007_g N_A_226_47#_c_247_n 0.00393414f $X=1.475 $Y=0.445 $X2=0
+ $Y2=0
cc_193 N_A2_N_M1007_g N_VGND_c_498_n 0.00341689f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A2_N_M1007_g N_VGND_c_499_n 0.00815507f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A2_N_M1007_g N_VGND_c_500_n 0.0040385f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_196 N_A_226_47#_c_247_n N_B2_M1004_g 0.0256273f $X=2.1 $Y=0.765 $X2=0 $Y2=0
cc_197 N_A_226_47#_c_248_n N_B2_M1008_g 0.00365421f $X=2.285 $Y=1.755 $X2=0
+ $Y2=0
cc_198 N_A_226_47#_c_250_n N_B2_M1008_g 0.0238667f $X=2.37 $Y=1.83 $X2=0 $Y2=0
cc_199 N_A_226_47#_c_246_n B2 0.00105716f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_200 N_A_226_47#_c_246_n N_B2_c_313_n 0.0256273f $X=1.975 $Y=1.07 $X2=0 $Y2=0
cc_201 N_A_226_47#_M1002_g N_VPWR_c_409_n 0.00431274f $X=2.37 $Y=2.275 $X2=0
+ $Y2=0
cc_202 N_A_226_47#_M1002_g N_VPWR_c_405_n 0.00764842f $X=2.37 $Y=2.275 $X2=0
+ $Y2=0
cc_203 N_A_226_47#_M1002_g N_A_489_413#_c_459_n 0.00144965f $X=2.37 $Y=2.275
+ $X2=0 $Y2=0
cc_204 N_A_226_47#_c_250_n N_A_489_413#_c_461_n 0.00119371f $X=2.37 $Y=1.83
+ $X2=0 $Y2=0
cc_205 N_A_226_47#_M1002_g N_A_489_413#_c_468_n 0.00336318f $X=2.37 $Y=2.275
+ $X2=0 $Y2=0
cc_206 N_A_226_47#_c_244_n N_VGND_M1007_d 0.00182057f $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_226_47#_c_247_n N_VGND_c_496_n 0.0034676f $X=2.1 $Y=0.765 $X2=0 $Y2=0
cc_208 N_A_226_47#_c_303_p N_VGND_c_498_n 0.0112554f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_226_47#_c_244_n N_VGND_c_498_n 0.00273399f $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A_226_47#_c_244_n N_VGND_c_499_n 0.0403001f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_226_47#_c_246_n N_VGND_c_499_n 0.00636187f $X=1.975 $Y=1.07 $X2=0
+ $Y2=0
cc_212 N_A_226_47#_c_247_n N_VGND_c_499_n 0.00993236f $X=2.1 $Y=0.765 $X2=0
+ $Y2=0
cc_213 N_A_226_47#_M1009_d N_VGND_c_500_n 0.00412745f $X=1.13 $Y=0.235 $X2=0
+ $Y2=0
cc_214 N_A_226_47#_c_303_p N_VGND_c_500_n 0.00644035f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_226_47#_c_244_n N_VGND_c_500_n 0.00654297f $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_216 N_A_226_47#_c_247_n N_VGND_c_500_n 0.00412709f $X=2.1 $Y=0.765 $X2=0
+ $Y2=0
cc_217 N_B2_M1004_g N_B1_M1003_g 0.0464258f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_218 N_B2_c_314_n N_B1_M1003_g 0.00547864f $X=2.95 $Y=1.505 $X2=0 $Y2=0
cc_219 N_B2_M1008_g N_B1_M1006_g 0.0307672f $X=2.79 $Y=2.275 $X2=0 $Y2=0
cc_220 B2 N_B1_M1006_g 0.00230104f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_221 B2 B1 0.0212546f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_222 N_B2_c_313_n B1 2.49998e-19 $X=2.765 $Y=1.47 $X2=0 $Y2=0
cc_223 N_B2_c_314_n B1 0.039191f $X=2.95 $Y=1.505 $X2=0 $Y2=0
cc_224 N_B2_M1004_g N_B1_c_360_n 0.00420826f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B2_c_313_n N_B1_c_360_n 0.0167199f $X=2.765 $Y=1.47 $X2=0 $Y2=0
cc_226 N_B2_c_314_n N_B1_c_360_n 0.00651406f $X=2.95 $Y=1.505 $X2=0 $Y2=0
cc_227 N_B2_M1008_g N_VPWR_c_407_n 0.00279634f $X=2.79 $Y=2.275 $X2=0 $Y2=0
cc_228 N_B2_M1008_g N_VPWR_c_409_n 0.00422411f $X=2.79 $Y=2.275 $X2=0 $Y2=0
cc_229 N_B2_M1008_g N_VPWR_c_405_n 0.0057538f $X=2.79 $Y=2.275 $X2=0 $Y2=0
cc_230 N_B2_M1008_g N_A_489_413#_c_459_n 0.00512513f $X=2.79 $Y=2.275 $X2=0
+ $Y2=0
cc_231 N_B2_M1008_g N_A_489_413#_c_460_n 0.00844573f $X=2.79 $Y=2.275 $X2=0
+ $Y2=0
cc_232 B2 N_A_489_413#_c_460_n 0.0243011f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_233 N_B2_c_313_n N_A_489_413#_c_460_n 2.30917e-19 $X=2.765 $Y=1.47 $X2=0
+ $Y2=0
cc_234 N_B2_M1008_g N_A_489_413#_c_461_n 0.00208357f $X=2.79 $Y=2.275 $X2=0
+ $Y2=0
cc_235 B2 N_A_489_413#_c_461_n 0.0115301f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_236 N_B2_c_313_n N_A_489_413#_c_461_n 5.97005e-19 $X=2.765 $Y=1.47 $X2=0
+ $Y2=0
cc_237 N_B2_M1008_g N_A_489_413#_c_468_n 0.00214984f $X=2.79 $Y=2.275 $X2=0
+ $Y2=0
cc_238 N_B2_M1004_g N_VGND_c_494_n 0.00224511f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_239 N_B2_M1004_g N_VGND_c_496_n 0.00585385f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_240 N_B2_M1004_g N_VGND_c_499_n 0.00126121f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_241 N_B2_M1004_g N_VGND_c_500_n 0.0108681f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_242 N_B2_c_314_n N_VGND_c_500_n 0.0104262f $X=2.95 $Y=1.505 $X2=0 $Y2=0
cc_243 N_B1_M1006_g N_VPWR_c_407_n 0.00884045f $X=3.21 $Y=2.275 $X2=0 $Y2=0
cc_244 N_B1_M1006_g N_VPWR_c_410_n 0.00348405f $X=3.21 $Y=2.275 $X2=0 $Y2=0
cc_245 N_B1_M1006_g N_VPWR_c_405_n 0.00513647f $X=3.21 $Y=2.275 $X2=0 $Y2=0
cc_246 N_B1_M1006_g N_A_489_413#_c_459_n 4.53479e-19 $X=3.21 $Y=2.275 $X2=0
+ $Y2=0
cc_247 N_B1_M1006_g N_A_489_413#_c_460_n 0.0172172f $X=3.21 $Y=2.275 $X2=0 $Y2=0
cc_248 B1 N_A_489_413#_c_460_n 0.0204099f $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_249 N_B1_c_360_n N_A_489_413#_c_460_n 0.00216853f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B1_M1006_g N_A_489_413#_c_462_n 0.00192069f $X=3.21 $Y=2.275 $X2=0
+ $Y2=0
cc_251 N_B1_M1003_g N_VGND_c_494_n 0.0157597f $X=3.125 $Y=0.445 $X2=0 $Y2=0
cc_252 B1 N_VGND_c_494_n 0.0230984f $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_253 N_B1_c_360_n N_VGND_c_494_n 0.00301098f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_M1003_g N_VGND_c_496_n 0.00407992f $X=3.125 $Y=0.445 $X2=0 $Y2=0
cc_255 N_B1_M1003_g N_VGND_c_500_n 0.00618209f $X=3.125 $Y=0.445 $X2=0 $Y2=0
cc_256 B1 N_VGND_c_500_n 0.00104546f $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_257 N_X_c_393_n N_VPWR_c_408_n 0.018001f $X=0.26 $Y=1.76 $X2=0 $Y2=0
cc_258 N_X_M1005_s N_VPWR_c_405_n 0.00387172f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_259 N_X_c_393_n N_VPWR_c_405_n 0.00993603f $X=0.26 $Y=1.76 $X2=0 $Y2=0
cc_260 X N_VGND_c_495_n 0.0179204f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_261 N_X_M1011_s N_VGND_c_500_n 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_262 X N_VGND_c_500_n 0.00991903f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_263 N_VPWR_c_405_n N_A_489_413#_M1002_d 0.00217615f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_264 N_VPWR_c_405_n N_A_489_413#_M1006_d 0.0034105f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_407_n N_A_489_413#_c_460_n 0.0166491f $X=3 $Y=2.34 $X2=0 $Y2=0
cc_266 N_VPWR_c_409_n N_A_489_413#_c_460_n 0.00240484f $X=2.915 $Y=2.72 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_410_n N_A_489_413#_c_460_n 0.00240298f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_405_n N_A_489_413#_c_460_n 0.00878585f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_410_n N_A_489_413#_c_462_n 0.0122405f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_405_n N_A_489_413#_c_462_n 0.00684138f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_409_n N_A_489_413#_c_468_n 0.0140432f $X=2.915 $Y=2.72 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_405_n N_A_489_413#_c_468_n 0.011577f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_273 N_VGND_c_500_n A_556_47# 0.00486328f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

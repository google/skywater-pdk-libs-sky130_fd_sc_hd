* File: sky130_fd_sc_hd__o311ai_4.pex.spice
* Created: Thu Aug 27 14:39:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O311AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 54
c74 36 0 1.92558e-19 $X=1.59 $Y=1.19
r75 52 54 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=1.595 $Y=1.16
+ $X2=1.81 $Y2=1.16
r76 50 52 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=1.39 $Y=1.16
+ $X2=1.595 $Y2=1.16
r77 48 50 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.255 $Y=1.16
+ $X2=1.39 $Y2=1.16
r78 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.255
+ $Y=1.16 $X2=1.255 $Y2=1.16
r79 46 48 63.3195 $w=2.7e-07 $l=2.85e-07 $layer=POLY_cond $X=0.97 $Y=1.16
+ $X2=1.255 $Y2=1.16
r80 44 46 12.2196 $w=2.7e-07 $l=5.5e-08 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=0.97 $Y2=1.16
r81 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.915
+ $Y=1.16 $X2=0.915 $Y2=1.16
r82 41 44 81.0934 $w=2.7e-07 $l=3.65e-07 $layer=POLY_cond $X=0.55 $Y=1.16
+ $X2=0.915 $Y2=1.16
r83 36 49 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.59 $Y=1.185
+ $X2=1.255 $Y2=1.185
r84 36 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.595
+ $Y=1.16 $X2=1.595 $Y2=1.16
r85 35 49 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=1.13 $Y=1.185
+ $X2=1.255 $Y2=1.185
r86 35 45 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=1.13 $Y=1.185
+ $X2=0.915 $Y2=1.185
r87 34 45 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=0.67 $Y=1.185
+ $X2=0.915 $Y2=1.185
r88 33 34 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=0.21 $Y=1.185
+ $X2=0.67 $Y2=1.185
r89 29 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.81 $Y=1.295
+ $X2=1.81 $Y2=1.16
r90 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.81 $Y=1.295
+ $X2=1.81 $Y2=1.985
r91 25 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.81 $Y=1.025
+ $X2=1.81 $Y2=1.16
r92 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.81 $Y=1.025
+ $X2=1.81 $Y2=0.56
r93 21 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.39 $Y=1.295
+ $X2=1.39 $Y2=1.16
r94 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.39 $Y=1.295
+ $X2=1.39 $Y2=1.985
r95 17 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.39 $Y=1.025
+ $X2=1.39 $Y2=1.16
r96 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.39 $Y=1.025
+ $X2=1.39 $Y2=0.56
r97 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.97 $Y=1.295
+ $X2=0.97 $Y2=1.16
r98 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.97 $Y=1.295
+ $X2=0.97 $Y2=1.985
r99 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.97 $Y=1.025
+ $X2=0.97 $Y2=1.16
r100 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.97 $Y=1.025
+ $X2=0.97 $Y2=0.56
r101 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.55 $Y2=1.16
r102 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.55 $Y=1.295
+ $X2=0.55 $Y2=1.985
r103 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.55 $Y=1.025
+ $X2=0.55 $Y2=1.16
r104 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.55 $Y=1.025
+ $X2=0.55 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%A2 3 7 11 15 19 23 27 31 33 34 35 36 54
c87 54 0 1.92558e-19 $X=3.49 $Y=1.16
r88 52 54 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.34 $Y=1.16
+ $X2=3.49 $Y2=1.16
r89 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.34
+ $Y=1.16 $X2=3.34 $Y2=1.16
r90 50 52 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=3.07 $Y=1.16
+ $X2=3.34 $Y2=1.16
r91 48 50 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=3 $Y=1.16 $X2=3.07
+ $Y2=1.16
r92 46 48 77.7608 $w=2.7e-07 $l=3.5e-07 $layer=POLY_cond $X=2.65 $Y=1.16 $X2=3
+ $Y2=1.16
r93 44 46 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.32 $Y=1.16
+ $X2=2.65 $Y2=1.16
r94 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.16 $X2=2.32 $Y2=1.16
r95 41 44 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.23 $Y=1.16 $X2=2.32
+ $Y2=1.16
r96 36 53 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=3.43 $Y=1.185 $X2=3.34
+ $Y2=1.185
r97 35 53 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.97 $Y=1.185
+ $X2=3.34 $Y2=1.185
r98 35 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3 $Y=1.16
+ $X2=3 $Y2=1.16
r99 34 35 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=2.51 $Y=1.185
+ $X2=2.97 $Y2=1.185
r100 34 45 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=2.51 $Y=1.185
+ $X2=2.32 $Y2=1.185
r101 33 45 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=2.05 $Y=1.185
+ $X2=2.32 $Y2=1.185
r102 29 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.49 $Y=1.295
+ $X2=3.49 $Y2=1.16
r103 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.49 $Y=1.295
+ $X2=3.49 $Y2=1.985
r104 25 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.49 $Y=1.025
+ $X2=3.49 $Y2=1.16
r105 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.49 $Y=1.025
+ $X2=3.49 $Y2=0.56
r106 21 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.07 $Y=1.295
+ $X2=3.07 $Y2=1.16
r107 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.07 $Y=1.295
+ $X2=3.07 $Y2=1.985
r108 17 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.07 $Y=1.025
+ $X2=3.07 $Y2=1.16
r109 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.07 $Y=1.025
+ $X2=3.07 $Y2=0.56
r110 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.65 $Y=1.295
+ $X2=2.65 $Y2=1.16
r111 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.65 $Y=1.295
+ $X2=2.65 $Y2=1.985
r112 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.65 $Y=1.025
+ $X2=2.65 $Y2=1.16
r113 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.65 $Y=1.025
+ $X2=2.65 $Y2=0.56
r114 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.23 $Y=1.295
+ $X2=2.23 $Y2=1.16
r115 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.23 $Y=1.295
+ $X2=2.23 $Y2=1.985
r116 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.23 $Y=1.025
+ $X2=2.23 $Y2=1.16
r117 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.23 $Y=1.025
+ $X2=2.23 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 37 63
c90 63 0 7.33294e-20 $X=5.69 $Y=1.16
r91 61 63 68.8738 $w=2.7e-07 $l=3.1e-07 $layer=POLY_cond $X=5.38 $Y=1.16
+ $X2=5.69 $Y2=1.16
r92 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.38
+ $Y=1.16 $X2=5.38 $Y2=1.16
r93 59 61 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=5.27 $Y=1.16
+ $X2=5.38 $Y2=1.16
r94 58 59 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=5.19 $Y=1.16 $X2=5.27
+ $Y2=1.16
r95 56 58 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=5.04 $Y=1.16
+ $X2=5.19 $Y2=1.16
r96 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=1.16 $X2=5.04 $Y2=1.16
r97 54 56 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=4.85 $Y=1.16 $X2=5.04
+ $Y2=1.16
r98 53 54 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=4.77 $Y=1.16 $X2=4.85
+ $Y2=1.16
r99 51 53 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=4.7 $Y=1.16 $X2=4.77
+ $Y2=1.16
r100 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.7
+ $Y=1.16 $X2=4.7 $Y2=1.16
r101 49 51 59.9869 $w=2.7e-07 $l=2.7e-07 $layer=POLY_cond $X=4.43 $Y=1.16
+ $X2=4.7 $Y2=1.16
r102 47 49 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=4.36 $Y=1.16 $X2=4.43
+ $Y2=1.16
r103 45 47 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=4.35 $Y=1.16 $X2=4.36
+ $Y2=1.16
r104 43 45 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.35 $Y2=1.16
r105 37 62 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=5.75 $Y=1.185
+ $X2=5.38 $Y2=1.185
r106 36 62 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=5.29 $Y=1.185
+ $X2=5.38 $Y2=1.185
r107 36 57 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=5.29 $Y=1.185
+ $X2=5.04 $Y2=1.185
r108 35 57 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=1.185
+ $X2=5.04 $Y2=1.185
r109 35 52 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=4.83 $Y=1.185
+ $X2=4.7 $Y2=1.185
r110 34 52 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=4.36 $Y=1.185
+ $X2=4.7 $Y2=1.185
r111 34 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.36
+ $Y=1.16 $X2=4.36 $Y2=1.16
r112 33 34 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=3.91 $Y=1.185
+ $X2=4.36 $Y2=1.185
r113 29 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.69 $Y=1.295
+ $X2=5.69 $Y2=1.16
r114 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.69 $Y=1.295
+ $X2=5.69 $Y2=1.985
r115 25 59 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.27 $Y=1.295
+ $X2=5.27 $Y2=1.16
r116 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.27 $Y=1.295
+ $X2=5.27 $Y2=1.985
r117 21 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=1.16
r118 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=0.56
r119 17 54 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.85 $Y=1.295
+ $X2=4.85 $Y2=1.16
r120 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.85 $Y=1.295
+ $X2=4.85 $Y2=1.985
r121 13 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=1.16
r122 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=0.56
r123 9 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.43 $Y=1.295
+ $X2=4.43 $Y2=1.16
r124 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.43 $Y=1.295
+ $X2=4.43 $Y2=1.985
r125 5 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=1.16
r126 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
r127 1 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=1.16
r128 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 58
c72 58 0 1.73414e-19 $X=7.43 $Y=1.16
c73 27 0 1.30541e-20 $X=7.39 $Y=1.985
r74 57 58 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=7.39 $Y=1.16 $X2=7.43
+ $Y2=1.16
r75 55 57 21.1065 $w=2.7e-07 $l=9.5e-08 $layer=POLY_cond $X=7.295 $Y=1.16
+ $X2=7.39 $Y2=1.16
r76 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.295
+ $Y=1.16 $X2=7.295 $Y2=1.16
r77 53 55 63.3195 $w=2.7e-07 $l=2.85e-07 $layer=POLY_cond $X=7.01 $Y=1.16
+ $X2=7.295 $Y2=1.16
r78 52 53 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=6.97 $Y=1.16 $X2=7.01
+ $Y2=1.16
r79 50 52 3.33261 $w=2.7e-07 $l=1.5e-08 $layer=POLY_cond $X=6.955 $Y=1.16
+ $X2=6.97 $Y2=1.16
r80 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.955
+ $Y=1.16 $X2=6.955 $Y2=1.16
r81 48 50 81.0934 $w=2.7e-07 $l=3.65e-07 $layer=POLY_cond $X=6.59 $Y=1.16
+ $X2=6.955 $Y2=1.16
r82 47 48 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=6.55 $Y=1.16 $X2=6.59
+ $Y2=1.16
r83 45 47 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=6.275 $Y=1.16
+ $X2=6.55 $Y2=1.16
r84 43 45 23.3282 $w=2.7e-07 $l=1.05e-07 $layer=POLY_cond $X=6.17 $Y=1.16
+ $X2=6.275 $Y2=1.16
r85 41 43 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=6.13 $Y=1.16 $X2=6.17
+ $Y2=1.16
r86 36 56 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=7.61 $Y=1.185
+ $X2=7.295 $Y2=1.185
r87 35 56 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=7.15 $Y=1.185
+ $X2=7.295 $Y2=1.185
r88 35 51 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=7.15 $Y=1.185
+ $X2=6.955 $Y2=1.185
r89 34 51 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=6.69 $Y=1.185
+ $X2=6.955 $Y2=1.185
r90 33 34 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=6.23 $Y=1.185
+ $X2=6.69 $Y2=1.185
r91 33 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.275
+ $Y=1.16 $X2=6.275 $Y2=1.16
r92 29 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.43 $Y=1.025
+ $X2=7.43 $Y2=1.16
r93 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.43 $Y=1.025
+ $X2=7.43 $Y2=0.56
r94 25 57 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.39 $Y=1.295
+ $X2=7.39 $Y2=1.16
r95 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.39 $Y=1.295
+ $X2=7.39 $Y2=1.985
r96 21 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.01 $Y=1.025
+ $X2=7.01 $Y2=1.16
r97 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.01 $Y=1.025
+ $X2=7.01 $Y2=0.56
r98 17 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.97 $Y=1.295
+ $X2=6.97 $Y2=1.16
r99 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.97 $Y=1.295
+ $X2=6.97 $Y2=1.985
r100 13 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.59 $Y=1.025
+ $X2=6.59 $Y2=1.16
r101 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.59 $Y=1.025
+ $X2=6.59 $Y2=0.56
r102 9 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.16
r103 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.985
r104 5 43 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.17 $Y=1.025
+ $X2=6.17 $Y2=1.16
r105 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.17 $Y=1.025
+ $X2=6.17 $Y2=0.56
r106 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.13 $Y=1.295
+ $X2=6.13 $Y2=1.16
r107 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.13 $Y=1.295
+ $X2=6.13 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%C1 3 7 11 15 19 23 27 31 33 34 35 56
c66 35 0 1.86468e-19 $X=8.99 $Y=1.19
r67 55 56 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=9.07 $Y=1.16 $X2=9.11
+ $Y2=1.16
r68 53 55 79.9825 $w=2.7e-07 $l=3.6e-07 $layer=POLY_cond $X=8.71 $Y=1.16
+ $X2=9.07 $Y2=1.16
r69 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.71
+ $Y=1.16 $X2=8.71 $Y2=1.16
r70 51 53 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=8.69 $Y=1.16 $X2=8.71
+ $Y2=1.16
r71 50 51 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=8.65 $Y=1.16 $X2=8.69
+ $Y2=1.16
r72 48 50 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=8.37 $Y=1.16
+ $X2=8.65 $Y2=1.16
r73 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.37
+ $Y=1.16 $X2=8.37 $Y2=1.16
r74 46 48 22.2174 $w=2.7e-07 $l=1e-07 $layer=POLY_cond $X=8.27 $Y=1.16 $X2=8.37
+ $Y2=1.16
r75 45 46 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=8.23 $Y=1.16 $X2=8.27
+ $Y2=1.16
r76 43 45 44.4347 $w=2.7e-07 $l=2e-07 $layer=POLY_cond $X=8.03 $Y=1.16 $X2=8.23
+ $Y2=1.16
r77 41 43 39.9913 $w=2.7e-07 $l=1.8e-07 $layer=POLY_cond $X=7.85 $Y=1.16
+ $X2=8.03 $Y2=1.16
r78 39 41 8.88695 $w=2.7e-07 $l=4e-08 $layer=POLY_cond $X=7.81 $Y=1.16 $X2=7.85
+ $Y2=1.16
r79 35 54 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=8.99 $Y=1.185
+ $X2=8.71 $Y2=1.185
r80 34 54 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=8.53 $Y=1.185
+ $X2=8.71 $Y2=1.185
r81 34 49 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=8.53 $Y=1.185
+ $X2=8.37 $Y2=1.185
r82 33 49 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=8.03 $Y=1.185
+ $X2=8.37 $Y2=1.185
r83 33 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.03
+ $Y=1.16 $X2=8.03 $Y2=1.16
r84 29 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.11 $Y=1.025
+ $X2=9.11 $Y2=1.16
r85 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.11 $Y=1.025
+ $X2=9.11 $Y2=0.56
r86 25 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.07 $Y=1.295
+ $X2=9.07 $Y2=1.16
r87 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.07 $Y=1.295
+ $X2=9.07 $Y2=1.985
r88 21 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.69 $Y=1.025
+ $X2=8.69 $Y2=1.16
r89 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.69 $Y=1.025
+ $X2=8.69 $Y2=0.56
r90 17 50 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.65 $Y=1.295
+ $X2=8.65 $Y2=1.16
r91 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.65 $Y=1.295
+ $X2=8.65 $Y2=1.985
r92 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.27 $Y=1.025
+ $X2=8.27 $Y2=1.16
r93 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.27 $Y=1.025
+ $X2=8.27 $Y2=0.56
r94 9 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.23 $Y=1.295
+ $X2=8.23 $Y2=1.16
r95 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.23 $Y=1.295
+ $X2=8.23 $Y2=1.985
r96 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.85 $Y=1.025
+ $X2=7.85 $Y2=1.16
r97 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.85 $Y=1.025
+ $X2=7.85 $Y2=0.56
r98 1 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.81 $Y=1.295
+ $X2=7.81 $Y2=1.16
r99 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.81 $Y=1.295 $X2=7.81
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%A_39_297# 1 2 3 4 5 18 20 21 24 26 30 32 34
+ 37 39 42 43 44
c63 43 0 9.67656e-20 $X=2.02 $Y=1.605
c64 37 0 7.33294e-20 $X=3.615 $Y=1.605
r65 39 41 4.392 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=3.74 $Y=1.725 $X2=3.74
+ $Y2=1.815
r66 38 44 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=1.605
+ $X2=2.86 $Y2=1.605
r67 37 39 6.82018 $w=2.4e-07 $l=1.75e-07 $layer=LI1_cond $X=3.615 $Y=1.605
+ $X2=3.74 $Y2=1.725
r68 37 38 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=3.615 $Y=1.605
+ $X2=2.945 $Y2=1.605
r69 34 44 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.86 $Y=1.725
+ $X2=2.86 $Y2=1.605
r70 34 36 6.45882 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.86 $Y=1.725 $X2=2.86
+ $Y2=1.815
r71 33 43 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=1.605
+ $X2=2.02 $Y2=1.605
r72 32 44 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=1.605
+ $X2=2.86 $Y2=1.605
r73 32 33 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=2.775 $Y=1.605
+ $X2=2.105 $Y2=1.605
r74 28 43 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.02 $Y=1.725
+ $X2=2.02 $Y2=1.605
r75 28 30 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.02 $Y=1.725 $X2=2.02
+ $Y2=1.815
r76 27 42 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=1.605
+ $X2=1.18 $Y2=1.605
r77 26 43 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=1.605
+ $X2=2.02 $Y2=1.605
r78 26 27 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=1.935 $Y=1.605
+ $X2=1.265 $Y2=1.605
r79 22 42 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.18 $Y=1.725
+ $X2=1.18 $Y2=1.605
r80 22 24 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.18 $Y=1.725 $X2=1.18
+ $Y2=1.815
r81 20 42 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=1.605
+ $X2=1.18 $Y2=1.605
r82 20 21 33.1327 $w=2.38e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.605
+ $X2=0.405 $Y2=1.605
r83 16 21 6.999 $w=2.4e-07 $l=2.1166e-07 $layer=LI1_cond $X=0.245 $Y=1.725
+ $X2=0.405 $Y2=1.605
r84 16 18 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=0.245 $Y=1.725
+ $X2=0.245 $Y2=1.815
r85 5 41 600 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.485 $X2=3.7 $Y2=1.815
r86 4 36 600 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=1 $X=2.725
+ $Y=1.485 $X2=2.86 $Y2=1.815
r87 3 30 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=1.885
+ $Y=1.485 $X2=2.02 $Y2=1.815
r88 2 24 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.485 $X2=1.18 $Y2=1.815
r89 1 18 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=1.485 $X2=0.32 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 46
+ 48 53 58 63 68 78 79 82 85 88 91 94 99
r140 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r141 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r142 88 89 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r143 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r144 83 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r145 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r147 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r148 76 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r149 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r150 73 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=2.72
+ $X2=8.02 $Y2=2.72
r151 73 75 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.185 $Y=2.72
+ $X2=8.51 $Y2=2.72
r152 72 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r153 72 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r154 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r155 69 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.345 $Y=2.72
+ $X2=7.18 $Y2=2.72
r156 69 71 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.345 $Y=2.72
+ $X2=7.59 $Y2=2.72
r157 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.855 $Y=2.72
+ $X2=8.02 $Y2=2.72
r158 68 71 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.855 $Y=2.72
+ $X2=7.59 $Y2=2.72
r159 67 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r160 67 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r161 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r162 64 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.34 $Y2=2.72
r163 64 66 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.67 $Y2=2.72
r164 63 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=7.18 $Y2=2.72
r165 63 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=6.67 $Y2=2.72
r166 62 89 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=6.21 $Y2=2.72
r167 62 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r168 61 62 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r169 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=2.72
+ $X2=1.6 $Y2=2.72
r170 59 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.765 $Y=2.72
+ $X2=2.07 $Y2=2.72
r171 58 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=2.72
+ $X2=6.34 $Y2=2.72
r172 58 61 267.813 $w=1.68e-07 $l=4.105e-06 $layer=LI1_cond $X=6.175 $Y=2.72
+ $X2=2.07 $Y2=2.72
r173 57 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r174 57 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r175 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r176 54 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.76 $Y2=2.72
r177 54 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.15 $Y2=2.72
r178 53 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.6 $Y2=2.72
r179 53 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.435 $Y=2.72
+ $X2=1.15 $Y2=2.72
r180 50 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r181 48 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.76 $Y2=2.72
r182 48 50 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r183 46 99 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=2.72
+ $X2=0.23 $Y2=2.72
r184 44 75 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.695 $Y=2.72
+ $X2=8.51 $Y2=2.72
r185 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=2.72
+ $X2=8.86 $Y2=2.72
r186 43 78 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=9.025 $Y=2.72
+ $X2=9.43 $Y2=2.72
r187 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=2.72
+ $X2=8.86 $Y2=2.72
r188 39 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=2.635
+ $X2=8.86 $Y2=2.72
r189 39 41 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=8.86 $Y=2.635
+ $X2=8.86 $Y2=2.02
r190 35 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=2.635
+ $X2=8.02 $Y2=2.72
r191 35 37 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=8.02 $Y=2.635
+ $X2=8.02 $Y2=2.02
r192 31 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=2.635
+ $X2=7.18 $Y2=2.72
r193 31 33 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=7.18 $Y=2.635
+ $X2=7.18 $Y2=2.02
r194 27 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.34 $Y=2.635
+ $X2=6.34 $Y2=2.72
r195 27 29 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=6.34 $Y=2.635
+ $X2=6.34 $Y2=2.02
r196 23 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=2.635 $X2=1.6
+ $Y2=2.72
r197 23 25 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.6 $Y=2.635
+ $X2=1.6 $Y2=2.02
r198 19 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=2.72
r199 19 21 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.76 $Y=2.635
+ $X2=0.76 $Y2=2.02
r200 6 41 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=8.725
+ $Y=1.485 $X2=8.86 $Y2=2.02
r201 5 37 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=2.02
r202 4 33 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=7.045
+ $Y=1.485 $X2=7.18 $Y2=2.02
r203 3 29 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=2.02
r204 2 25 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.465
+ $Y=1.485 $X2=1.6 $Y2=2.02
r205 1 21 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=0.625
+ $Y=1.485 $X2=0.76 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%A_461_297# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
r64 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.48 $Y=2.295
+ $X2=5.48 $Y2=2.02
r65 30 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=2.38
+ $X2=4.64 $Y2=2.38
r66 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.315 $Y=2.38
+ $X2=5.48 $Y2=2.295
r67 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.315 $Y=2.38
+ $X2=4.805 $Y2=2.38
r68 25 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=2.295
+ $X2=4.64 $Y2=2.38
r69 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.64 $Y=2.295
+ $X2=4.64 $Y2=2.02
r70 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=2.38
+ $X2=3.28 $Y2=2.38
r71 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=2.38
+ $X2=4.64 $Y2=2.38
r72 23 24 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=4.475 $Y=2.38
+ $X2=3.445 $Y2=2.38
r73 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=2.295
+ $X2=3.28 $Y2=2.38
r74 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.28 $Y=2.295
+ $X2=3.28 $Y2=2.02
r75 17 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=2.38
+ $X2=3.28 $Y2=2.38
r76 17 18 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.115 $Y=2.38
+ $X2=2.605 $Y2=2.38
r77 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.44 $Y=2.295
+ $X2=2.605 $Y2=2.38
r78 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.44 $Y=2.295
+ $X2=2.44 $Y2=2.02
r79 4 33 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=5.345
+ $Y=1.485 $X2=5.48 $Y2=2.02
r80 3 27 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=1.485 $X2=4.64 $Y2=2.02
r81 2 21 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.145
+ $Y=1.485 $X2=3.28 $Y2=2.02
r82 1 15 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.305
+ $Y=1.485 $X2=2.44 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%Y 1 2 3 4 5 6 7 8 9 28 31 32 33 36 40 42 46
+ 48 52 54 56 64 66 68 69 70 71 72 73 74 75 76 77 85 93
r104 91 93 2.72947 $w=3.78e-07 $l=9e-08 $layer=LI1_cond $X=9.385 $Y=1.725
+ $X2=9.385 $Y2=1.815
r105 76 77 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=9.385 $Y=1.87
+ $X2=9.385 $Y2=2.21
r106 76 93 1.66801 $w=3.78e-07 $l=5.5e-08 $layer=LI1_cond $X=9.385 $Y=1.87
+ $X2=9.385 $Y2=1.815
r107 75 86 3.75865 $w=3.47e-07 $l=1.35056e-07 $layer=LI1_cond $X=9.385 $Y=1.605
+ $X2=9.417 $Y2=1.485
r108 75 91 3.75865 $w=3.47e-07 $l=1.2e-07 $layer=LI1_cond $X=9.385 $Y=1.605
+ $X2=9.385 $Y2=1.725
r109 75 86 0.73171 $w=3.13e-07 $l=2e-08 $layer=LI1_cond $X=9.417 $Y=1.465
+ $X2=9.417 $Y2=1.485
r110 74 75 10.061 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=9.417 $Y=1.19
+ $X2=9.417 $Y2=1.465
r111 73 85 2.9741 $w=3.15e-07 $l=1.15e-07 $layer=LI1_cond $X=9.417 $Y=0.77
+ $X2=9.417 $Y2=0.885
r112 73 74 10.2439 $w=3.13e-07 $l=2.8e-07 $layer=LI1_cond $X=9.417 $Y=0.91
+ $X2=9.417 $Y2=1.19
r113 73 85 0.914637 $w=3.13e-07 $l=2.5e-08 $layer=LI1_cond $X=9.417 $Y=0.91
+ $X2=9.417 $Y2=0.885
r114 67 72 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=1.605
+ $X2=8.44 $Y2=1.605
r115 66 75 2.70353 $w=2.4e-07 $l=1.9e-07 $layer=LI1_cond $X=9.195 $Y=1.605
+ $X2=9.385 $Y2=1.605
r116 66 67 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=9.195 $Y=1.605
+ $X2=8.525 $Y2=1.605
r117 62 72 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=8.44 $Y=1.725
+ $X2=8.44 $Y2=1.605
r118 62 64 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.44 $Y=1.725
+ $X2=8.44 $Y2=1.815
r119 58 61 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=8.06 $Y=0.77
+ $X2=8.9 $Y2=0.77
r120 56 73 4.06029 $w=2.3e-07 $l=1.57e-07 $layer=LI1_cond $X=9.26 $Y=0.77
+ $X2=9.417 $Y2=0.77
r121 56 61 18.0382 $w=2.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.26 $Y=0.77
+ $X2=8.9 $Y2=0.77
r122 55 71 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=1.605
+ $X2=7.6 $Y2=1.605
r123 54 72 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=1.605
+ $X2=8.44 $Y2=1.605
r124 54 55 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=8.355 $Y=1.605
+ $X2=7.685 $Y2=1.605
r125 50 71 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.6 $Y=1.725 $X2=7.6
+ $Y2=1.605
r126 50 52 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.6 $Y=1.725 $X2=7.6
+ $Y2=1.815
r127 49 70 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=1.605
+ $X2=6.76 $Y2=1.605
r128 48 71 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=1.605
+ $X2=7.6 $Y2=1.605
r129 48 49 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=7.515 $Y=1.605
+ $X2=6.845 $Y2=1.605
r130 44 70 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.76 $Y=1.725
+ $X2=6.76 $Y2=1.605
r131 44 46 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.76 $Y=1.725
+ $X2=6.76 $Y2=1.815
r132 43 69 4.23567 $w=2.4e-07 $l=9.5e-08 $layer=LI1_cond $X=6.005 $Y=1.605
+ $X2=5.91 $Y2=1.605
r133 42 70 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=1.605
+ $X2=6.76 $Y2=1.605
r134 42 43 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=6.675 $Y=1.605
+ $X2=6.005 $Y2=1.605
r135 38 69 2.19581 $w=1.9e-07 $l=1.2e-07 $layer=LI1_cond $X=5.91 $Y=1.725
+ $X2=5.91 $Y2=1.605
r136 38 40 5.25359 $w=1.88e-07 $l=9e-08 $layer=LI1_cond $X=5.91 $Y=1.725
+ $X2=5.91 $Y2=1.815
r137 37 68 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=1.605
+ $X2=5.06 $Y2=1.605
r138 36 69 4.23567 $w=2.4e-07 $l=9.5e-08 $layer=LI1_cond $X=5.815 $Y=1.605
+ $X2=5.91 $Y2=1.605
r139 36 37 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=5.815 $Y=1.605
+ $X2=5.145 $Y2=1.605
r140 33 68 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.06 $Y=1.725
+ $X2=5.06 $Y2=1.605
r141 33 35 6.45882 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.06 $Y=1.725 $X2=5.06
+ $Y2=1.815
r142 31 68 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=1.605
+ $X2=5.06 $Y2=1.605
r143 31 32 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=1.605
+ $X2=4.305 $Y2=1.605
r144 28 32 6.82018 $w=2.4e-07 $l=1.75e-07 $layer=LI1_cond $X=4.18 $Y=1.725
+ $X2=4.305 $Y2=1.605
r145 28 30 4.392 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=4.18 $Y=1.725 $X2=4.18
+ $Y2=1.815
r146 9 93 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=9.145
+ $Y=1.485 $X2=9.28 $Y2=1.815
r147 8 64 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=1.815
r148 7 52 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=7.465
+ $Y=1.485 $X2=7.6 $Y2=1.815
r149 6 46 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=6.625
+ $Y=1.485 $X2=6.76 $Y2=1.815
r150 5 40 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=5.765
+ $Y=1.485 $X2=5.9 $Y2=1.815
r151 4 35 600 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.485 $X2=5.06 $Y2=1.815
r152 3 30 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=1.485 $X2=4.22 $Y2=1.815
r153 2 61 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=8.765
+ $Y=0.235 $X2=8.9 $Y2=0.76
r154 1 58 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=7.925
+ $Y=0.235 $X2=8.06 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46
+ 50 53 54 56 57 58 59 60 62 67 87 88 94 97 100 105
r153 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r154 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r155 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r156 91 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r157 87 88 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r158 85 88 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r159 85 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r160 84 87 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r161 84 85 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r162 82 100 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.585 $Y=0 $X2=5.41
+ $Y2=0
r163 82 84 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=0
+ $X2=5.75 $Y2=0
r164 81 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r165 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r166 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r167 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r168 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r169 75 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r170 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r171 72 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.02
+ $Y2=0
r172 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.53
+ $Y2=0
r173 71 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r174 71 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r175 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r176 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.18
+ $Y2=0
r177 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.345 $Y=0
+ $X2=1.61 $Y2=0
r178 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.02
+ $Y2=0
r179 67 70 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r180 66 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r181 66 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=0.23 $Y2=0
r182 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r183 63 91 5.67426 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.252 $Y2=0
r184 63 65 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.69 $Y2=0
r185 62 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.18
+ $Y2=0
r186 62 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r187 60 105 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=0
+ $X2=0.23 $Y2=0
r188 58 80 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.37
+ $Y2=0
r189 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.56
+ $Y2=0
r190 56 77 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.45
+ $Y2=0
r191 56 57 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.71
+ $Y2=0
r192 55 80 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=4.37 $Y2=0
r193 55 57 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.71
+ $Y2=0
r194 53 74 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=2.53 $Y2=0
r195 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.86
+ $Y2=0
r196 52 77 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.025 $Y=0
+ $X2=3.45 $Y2=0
r197 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.86
+ $Y2=0
r198 48 100 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=0.085
+ $X2=5.41 $Y2=0
r199 48 50 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.41 $Y=0.085
+ $X2=5.41 $Y2=0.36
r200 47 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=0 $X2=4.56
+ $Y2=0
r201 46 100 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.41
+ $Y2=0
r202 46 47 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.235 $Y=0
+ $X2=4.725 $Y2=0
r203 42 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0
r204 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0.36
r205 38 57 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.71 $Y2=0
r206 38 40 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.71 $Y2=0.36
r207 34 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r208 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.36
r209 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r210 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.36
r211 26 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0
r212 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.36
r213 22 91 2.87077 $w=4.2e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.252 $Y2=0
r214 22 24 7.54576 $w=4.18e-07 $l=2.75e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.36
r215 7 50 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.36
r216 6 44 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.36
r217 5 40 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.235 $X2=3.72 $Y2=0.36
r218 4 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.235 $X2=2.86 $Y2=0.36
r219 3 32 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.885
+ $Y=0.235 $X2=2.02 $Y2=0.36
r220 2 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.235 $X2=1.18 $Y2=0.36
r221 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.195
+ $Y=0.235 $X2=0.34 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%A_125_47# 1 2 3 4 5 6 7 8 25 28 29 30 33 35
+ 38 40 43 45 48 50 57 59 60 61 62 63
c106 33 0 9.67656e-20 $X=2.355 $Y=0.77
r107 55 57 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=6.38 $Y=0.77
+ $X2=7.22 $Y2=0.77
r108 53 63 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0.77
+ $X2=4.98 $Y2=0.77
r109 53 55 65.8897 $w=2.28e-07 $l=1.315e-06 $layer=LI1_cond $X=5.065 $Y=0.77
+ $X2=6.38 $Y2=0.77
r110 50 63 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.98 $Y=0.655
+ $X2=4.98 $Y2=0.77
r111 50 52 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.98 $Y=0.655
+ $X2=4.98 $Y2=0.56
r112 49 62 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0.77
+ $X2=4.14 $Y2=0.77
r113 48 63 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0.77
+ $X2=4.98 $Y2=0.77
r114 48 49 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=4.895 $Y=0.77
+ $X2=4.225 $Y2=0.77
r115 45 62 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.14 $Y=0.655
+ $X2=4.14 $Y2=0.77
r116 45 47 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.14 $Y=0.655
+ $X2=4.14 $Y2=0.56
r117 44 61 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=0.77
+ $X2=3.28 $Y2=0.77
r118 43 62 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0.77
+ $X2=4.14 $Y2=0.77
r119 43 44 34.5733 $w=2.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4.055 $Y=0.77
+ $X2=3.365 $Y2=0.77
r120 40 61 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.28 $Y=0.655
+ $X2=3.28 $Y2=0.77
r121 40 42 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.28 $Y=0.655
+ $X2=3.28 $Y2=0.56
r122 39 60 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.77
+ $X2=2.44 $Y2=0.77
r123 38 61 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=0.77
+ $X2=3.28 $Y2=0.77
r124 38 39 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=3.195 $Y=0.77
+ $X2=2.525 $Y2=0.77
r125 35 60 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.44 $Y=0.655
+ $X2=2.44 $Y2=0.77
r126 35 37 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.44 $Y=0.655
+ $X2=2.44 $Y2=0.56
r127 34 59 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=0.77
+ $X2=1.6 $Y2=0.77
r128 33 60 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=0.77
+ $X2=2.44 $Y2=0.77
r129 33 34 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.355 $Y=0.77
+ $X2=1.685 $Y2=0.77
r130 30 59 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.6 $Y=0.655
+ $X2=1.6 $Y2=0.77
r131 30 32 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.6 $Y=0.655 $X2=1.6
+ $Y2=0.56
r132 28 59 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.515 $Y=0.77
+ $X2=1.6 $Y2=0.77
r133 28 29 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.515 $Y=0.77
+ $X2=0.845 $Y2=0.77
r134 25 29 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.76 $Y=0.655
+ $X2=0.845 $Y2=0.77
r135 25 27 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.76 $Y=0.655
+ $X2=0.76 $Y2=0.56
r136 8 57 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=7.085
+ $Y=0.235 $X2=7.22 $Y2=0.76
r137 7 55 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=6.245
+ $Y=0.235 $X2=6.38 $Y2=0.76
r138 6 52 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.56
r139 5 47 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.56
r140 4 42 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.28 $Y2=0.56
r141 3 37 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.235 $X2=2.44 $Y2=0.56
r142 2 32 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.235 $X2=1.6 $Y2=0.56
r143 1 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.235 $X2=0.76 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311AI_4%A_1163_47# 1 2 3 4 5 16 24 30 33
r38 28 30 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=8.48 $Y=0.37
+ $X2=9.32 $Y2=0.37
r39 26 33 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=0.37
+ $X2=7.64 $Y2=0.37
r40 26 28 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=7.725 $Y=0.37
+ $X2=8.48 $Y2=0.37
r41 22 33 2.45049 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.64 $Y=0.485
+ $X2=7.64 $Y2=0.37
r42 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.64 $Y=0.485
+ $X2=7.64 $Y2=0.7
r43 18 21 42.0892 $w=2.28e-07 $l=8.4e-07 $layer=LI1_cond $X=5.96 $Y=0.37 $X2=6.8
+ $Y2=0.37
r44 16 33 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.37
+ $X2=7.64 $Y2=0.37
r45 16 21 37.8302 $w=2.28e-07 $l=7.55e-07 $layer=LI1_cond $X=7.555 $Y=0.37
+ $X2=6.8 $Y2=0.37
r46 5 30 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=9.185
+ $Y=0.235 $X2=9.32 $Y2=0.36
r47 4 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=8.345
+ $Y=0.235 $X2=8.48 $Y2=0.36
r48 3 33 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.505
+ $Y=0.235 $X2=7.64 $Y2=0.36
r49 3 24 182 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_NDIFF $count=1 $X=7.505
+ $Y=0.235 $X2=7.64 $Y2=0.7
r50 2 21 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.665
+ $Y=0.235 $X2=6.8 $Y2=0.36
r51 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.235 $X2=5.96 $Y2=0.36
.ends


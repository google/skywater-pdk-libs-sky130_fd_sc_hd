* File: sky130_fd_sc_hd__o211a_1.spice.SKY130_FD_SC_HD__O211A_1.pxi
* Created: Thu Aug 27 14:34:27 2020
* 
x_PM_SKY130_FD_SC_HD__O211A_1%A_79_21# N_A_79_21#_M1004_d N_A_79_21#_M1008_d
+ N_A_79_21#_M1003_d N_A_79_21#_M1009_g N_A_79_21#_M1007_g N_A_79_21#_c_68_n
+ N_A_79_21#_c_69_n N_A_79_21#_c_70_n N_A_79_21#_c_80_p N_A_79_21#_c_75_n
+ N_A_79_21#_c_81_p N_A_79_21#_c_97_p N_A_79_21#_c_71_n N_A_79_21#_c_77_n
+ N_A_79_21#_c_92_p N_A_79_21#_c_72_n N_A_79_21#_c_78_n
+ PM_SKY130_FD_SC_HD__O211A_1%A_79_21#
x_PM_SKY130_FD_SC_HD__O211A_1%A1 N_A1_M1002_g N_A1_M1000_g A1 N_A1_c_155_n
+ N_A1_c_156_n PM_SKY130_FD_SC_HD__O211A_1%A1
x_PM_SKY130_FD_SC_HD__O211A_1%A2 N_A2_M1005_g N_A2_M1008_g A2 N_A2_c_191_n
+ N_A2_c_192_n PM_SKY130_FD_SC_HD__O211A_1%A2
x_PM_SKY130_FD_SC_HD__O211A_1%B1 N_B1_M1006_g N_B1_M1001_g B1 N_B1_c_223_n
+ N_B1_c_224_n PM_SKY130_FD_SC_HD__O211A_1%B1
x_PM_SKY130_FD_SC_HD__O211A_1%C1 N_C1_c_252_n N_C1_M1004_g N_C1_M1003_g
+ N_C1_c_253_n C1 N_C1_c_255_n PM_SKY130_FD_SC_HD__O211A_1%C1
x_PM_SKY130_FD_SC_HD__O211A_1%X N_X_M1009_s N_X_M1007_s N_X_c_280_n N_X_c_283_n
+ N_X_c_281_n X X X N_X_c_282_n PM_SKY130_FD_SC_HD__O211A_1%X
x_PM_SKY130_FD_SC_HD__O211A_1%VPWR N_VPWR_M1007_d N_VPWR_M1000_s N_VPWR_M1001_d
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n
+ N_VPWR_c_304_n VPWR N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_298_n
+ N_VPWR_c_308_n N_VPWR_c_309_n PM_SKY130_FD_SC_HD__O211A_1%VPWR
x_PM_SKY130_FD_SC_HD__O211A_1%VGND N_VGND_M1009_d N_VGND_M1002_d N_VGND_c_346_n
+ N_VGND_c_347_n N_VGND_c_348_n VGND N_VGND_c_349_n N_VGND_c_350_n
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n PM_SKY130_FD_SC_HD__O211A_1%VGND
x_PM_SKY130_FD_SC_HD__O211A_1%A_215_47# N_A_215_47#_M1002_s N_A_215_47#_M1005_d
+ N_A_215_47#_c_390_n N_A_215_47#_c_391_n N_A_215_47#_c_392_n
+ N_A_215_47#_c_405_n PM_SKY130_FD_SC_HD__O211A_1%A_215_47#
cc_1 VNB N_A_79_21#_M1009_g 0.0285858f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_79_21#_M1007_g 5.7828e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_3 VNB N_A_79_21#_c_68_n 0.0173624f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=1.16
cc_4 VNB N_A_79_21#_c_69_n 0.036332f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_5 VNB N_A_79_21#_c_70_n 0.00144075f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=1.495
cc_6 VNB N_A_79_21#_c_71_n 0.00625919f $X=-0.19 $Y=-0.24 $X2=2.975 $Y2=1.495
cc_7 VNB N_A_79_21#_c_72_n 0.025334f $X=-0.19 $Y=-0.24 $X2=3.225 $Y2=0.38
cc_8 VNB A1 0.00553426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A1_c_155_n 0.0236488f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_10 VNB N_A1_c_156_n 0.022188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A2 0.00178447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_191_n 0.0269031f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_A2_c_192_n 0.0181251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB B1 0.00414972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_223_n 0.0243798f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_B1_c_224_n 0.0185792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_C1_c_252_n 0.0202414f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=0.235
cc_18 VNB N_C1_c_253_n 0.00806218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB C1 0.00932265f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_20 VNB N_C1_c_255_n 0.0457285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_280_n 0.00778155f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_22 VNB N_X_c_281_n 0.0199656f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.295
cc_23 VNB N_X_c_282_n 0.0183576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_298_n 0.155873f $X=-0.19 $Y=-0.24 $X2=3.14 $Y2=1.58
cc_25 VNB N_VGND_c_346_n 0.0127919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_347_n 0.0180541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_27 VNB N_VGND_c_348_n 0.00493933f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_28 VNB N_VGND_c_349_n 0.0177718f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_29 VNB N_VGND_c_350_n 0.0545477f $X=-0.19 $Y=-0.24 $X2=2.095 $Y2=2.34
cc_30 VNB N_VGND_c_351_n 0.216269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_352_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=2.975 $Y2=0.865
cc_32 VNB N_VGND_c_353_n 0.00429352f $X=-0.19 $Y=-0.24 $X2=3.225 $Y2=2.34
cc_33 VNB N_A_215_47#_c_390_n 0.00455239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_215_47#_c_391_n 0.00571864f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_35 VNB N_A_215_47#_c_392_n 0.00572586f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_36 VPB N_A_79_21#_M1007_g 0.0285309f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_37 VPB N_A_79_21#_c_70_n 0.00516767f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.495
cc_38 VPB N_A_79_21#_c_75_n 0.00555173f $X=-0.19 $Y=1.305 $X2=1.125 $Y2=1.58
cc_39 VPB N_A_79_21#_c_71_n 0.00615736f $X=-0.19 $Y=1.305 $X2=2.975 $Y2=1.495
cc_40 VPB N_A_79_21#_c_77_n 0.0312141f $X=-0.19 $Y=1.305 $X2=3.225 $Y2=2.34
cc_41 VPB N_A_79_21#_c_78_n 0.00740132f $X=-0.19 $Y=1.305 $X2=3.225 $Y2=1.66
cc_42 VPB N_A1_M1000_g 0.023064f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A1_c_155_n 0.00428957f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_44 VPB N_A2_M1008_g 0.0214731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A2_c_191_n 0.00703367f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_46 VPB N_B1_M1001_g 0.021701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_B1_c_223_n 0.0046465f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_48 VPB N_C1_M1003_g 0.0232687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_C1_c_253_n 5.2145e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB C1 0.00143415f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.025
cc_51 VPB N_C1_c_255_n 0.0192956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_283_n 0.00666696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_X_c_281_n 0.00903612f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.295
cc_54 VPB X 0.0316915f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_55 VPB N_VPWR_c_299_n 0.00350665f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_56 VPB N_VPWR_c_300_n 0.0085283f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_57 VPB N_VPWR_c_301_n 0.00953318f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_58 VPB N_VPWR_c_302_n 0.00561441f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.495
cc_59 VPB N_VPWR_c_303_n 0.0372945f $X=-0.19 $Y=1.305 $X2=2.095 $Y2=1.665
cc_60 VPB N_VPWR_c_304_n 0.00632158f $X=-0.19 $Y=1.305 $X2=2.095 $Y2=2.34
cc_61 VPB N_VPWR_c_305_n 0.0177718f $X=-0.19 $Y=1.305 $X2=2.89 $Y2=1.58
cc_62 VPB N_VPWR_c_306_n 0.024197f $X=-0.19 $Y=1.305 $X2=3.14 $Y2=0.865
cc_63 VPB N_VPWR_c_298_n 0.0614792f $X=-0.19 $Y=1.305 $X2=3.14 $Y2=1.58
cc_64 VPB N_VPWR_c_308_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_309_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_70_n N_A1_M1000_g 0.00554206f $X=1.04 $Y=1.495 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_80_p N_A1_M1000_g 0.0171407f $X=1.93 $Y=1.58 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_81_p N_A1_M1000_g 0.00279494f $X=2.095 $Y=2.34 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_68_n A1 0.0149908f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_69_n A1 3.81318e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_70_n A1 0.00226941f $X=1.04 $Y=1.495 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_80_p A1 0.021947f $X=1.93 $Y=1.58 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_68_n N_A1_c_155_n 7.48097e-19 $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_69_n N_A1_c_155_n 0.00478449f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_70_n N_A1_c_155_n 0.00165042f $X=1.04 $Y=1.495 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_80_p N_A1_c_155_n 0.00248719f $X=1.93 $Y=1.58 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_80_p N_A2_M1008_g 0.0121334f $X=1.93 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_81_p N_A2_M1008_g 0.0159806f $X=2.095 $Y=2.34 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_92_p N_A2_M1008_g 9.46316e-19 $X=2.095 $Y=1.66 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_80_p A2 0.00220653f $X=1.93 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_92_p A2 0.0168626f $X=2.095 $Y=1.66 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_92_p N_A2_c_191_n 0.00532551f $X=2.095 $Y=1.66 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_81_p N_B1_M1001_g 0.0105671f $X=2.095 $Y=2.34 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_97_p N_B1_M1001_g 0.016428f $X=2.89 $Y=1.58 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_71_n N_B1_M1001_g 0.00302379f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_97_p B1 0.0169969f $X=2.89 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_71_n B1 0.0158511f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_97_p N_B1_c_223_n 0.00306135f $X=2.89 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_71_n N_B1_c_223_n 0.00309378f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_71_n N_B1_c_224_n 0.00368286f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_71_n N_C1_c_252_n 0.004205f $X=2.975 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_79_21#_c_72_n N_C1_c_252_n 0.0126809f $X=3.225 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_79_21#_c_71_n N_C1_M1003_g 0.00575696f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_78_n N_C1_M1003_g 0.0124876f $X=3.225 $Y=1.66 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_71_n N_C1_c_253_n 0.00511845f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_71_n C1 0.0167085f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_72_n C1 0.00989252f $X=3.225 $Y=0.38 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_78_n C1 0.0118166f $X=3.225 $Y=1.66 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_71_n N_C1_c_255_n 0.00753997f $X=2.975 $Y=1.495 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_72_n N_C1_c_255_n 0.00886679f $X=3.225 $Y=0.38 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_78_n N_C1_c_255_n 0.0084293f $X=3.225 $Y=1.66 $X2=0 $Y2=0
cc_102 N_A_79_21#_M1009_g N_X_c_280_n 0.00262265f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A_79_21#_M1007_g N_X_c_283_n 0.00262265f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_79_21#_M1009_g N_X_c_281_n 0.0165779f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_68_n N_X_c_281_n 0.0134769f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_79_21#_M1007_g X 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_79_21#_M1009_g N_X_c_282_n 0.00528656f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_80_p N_VPWR_M1000_s 0.00488181f $X=1.93 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_75_n N_VPWR_M1000_s 0.00101038f $X=1.125 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_97_p N_VPWR_M1001_d 0.00835181f $X=2.89 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A_79_21#_M1007_g N_VPWR_c_299_n 0.00438629f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A_79_21#_c_68_n N_VPWR_c_299_n 0.00967581f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_69_n N_VPWR_c_299_n 0.00371763f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_75_n N_VPWR_c_299_n 0.0130371f $X=1.125 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_80_p N_VPWR_c_301_n 0.0124114f $X=1.93 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_75_n N_VPWR_c_301_n 0.0080326f $X=1.125 $Y=1.58 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_97_p N_VPWR_c_302_n 0.0192006f $X=2.89 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_81_p N_VPWR_c_303_n 0.0209845f $X=2.095 $Y=2.34 $X2=0 $Y2=0
cc_119 N_A_79_21#_M1007_g N_VPWR_c_305_n 0.00541359f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_79_21#_c_77_n N_VPWR_c_306_n 0.0215162f $X=3.225 $Y=2.34 $X2=0 $Y2=0
cc_121 N_A_79_21#_M1008_d N_VPWR_c_298_n 0.00843348f $X=1.96 $Y=1.485 $X2=0
+ $Y2=0
cc_122 N_A_79_21#_M1003_d N_VPWR_c_298_n 0.00276827f $X=3.05 $Y=1.485 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_M1007_g N_VPWR_c_298_n 0.0117818f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_81_p N_VPWR_c_298_n 0.0124268f $X=2.095 $Y=2.34 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_77_n N_VPWR_c_298_n 0.0126319f $X=3.225 $Y=2.34 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_80_p A_297_297# 0.0106695f $X=1.93 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A_79_21#_M1009_g N_VGND_c_346_n 0.0044954f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_68_n N_VGND_c_346_n 0.0181074f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_69_n N_VGND_c_346_n 0.00384364f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_79_21#_M1009_g N_VGND_c_349_n 0.00541359f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_72_n N_VGND_c_350_n 0.0322619f $X=3.225 $Y=0.38 $X2=0 $Y2=0
cc_132 N_A_79_21#_M1004_d N_VGND_c_351_n 0.00242111f $X=3.05 $Y=0.235 $X2=0
+ $Y2=0
cc_133 N_A_79_21#_M1009_g N_VGND_c_351_n 0.0117818f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_72_n N_VGND_c_351_n 0.0183845f $X=3.225 $Y=0.38 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_80_p N_A_215_47#_c_391_n 0.00384113f $X=1.93 $Y=1.58 $X2=0
+ $Y2=0
cc_136 N_A_79_21#_c_71_n N_A_215_47#_c_391_n 0.00321211f $X=2.975 $Y=1.495 $X2=0
+ $Y2=0
cc_137 N_A_79_21#_c_92_p N_A_215_47#_c_391_n 0.00148729f $X=2.095 $Y=1.66 $X2=0
+ $Y2=0
cc_138 N_A_79_21#_M1009_g N_A_215_47#_c_392_n 8.68203e-19 $X=0.47 $Y=0.56 $X2=0
+ $Y2=0
cc_139 N_A_79_21#_c_68_n N_A_215_47#_c_392_n 0.00831554f $X=0.955 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_79_21#_c_80_p N_A_215_47#_c_392_n 0.00558853f $X=1.93 $Y=1.58 $X2=0
+ $Y2=0
cc_141 N_A1_M1000_g N_A2_M1008_g 0.0479876f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_142 A1 A2 0.0161298f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_143 A1 N_A2_c_191_n 0.00136615f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A1_c_155_n N_A2_c_191_n 0.0220263f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A1_c_156_n N_A2_c_192_n 0.0212272f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A1_M1000_g N_VPWR_c_299_n 0.00524019f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A1_M1000_g N_VPWR_c_301_n 0.0044954f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A1_M1000_g N_VPWR_c_303_n 0.00585385f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A1_M1000_g N_VPWR_c_298_n 0.0121017f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A1_c_156_n N_VGND_c_346_n 0.0022981f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_156_n N_VGND_c_347_n 0.00424416f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A1_c_156_n N_VGND_c_348_n 0.00284731f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_156_n N_VGND_c_351_n 0.0072188f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_c_156_n N_A_215_47#_c_390_n 0.00680383f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_155 A1 N_A_215_47#_c_391_n 0.0256749f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_c_155_n N_A_215_47#_c_391_n 0.00283443f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_c_156_n N_A_215_47#_c_391_n 0.00876939f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_158 A1 N_A_215_47#_c_392_n 0.00526159f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A1_c_156_n N_A_215_47#_c_392_n 0.00126808f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A1_c_156_n N_A_215_47#_c_405_n 5.83925e-19 $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A2_M1008_g N_B1_M1001_g 0.0190229f $X=1.885 $Y=1.985 $X2=0 $Y2=0
cc_162 A2 B1 0.0165577f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A2_c_191_n B1 6.03485e-19 $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_164 A2 N_B1_c_223_n 6.36684e-19 $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_165 N_A2_c_191_n N_B1_c_223_n 0.0226595f $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A2_c_192_n N_B1_c_224_n 0.0132662f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_M1008_g N_VPWR_c_303_n 0.00541359f $X=1.885 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A2_M1008_g N_VPWR_c_298_n 0.0102518f $X=1.885 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A2_c_192_n N_VGND_c_348_n 0.00284731f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A2_c_192_n N_VGND_c_350_n 0.00424416f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A2_c_192_n N_VGND_c_351_n 0.00628166f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_192_n N_A_215_47#_c_390_n 5.83925e-19 $X=2 $Y=0.995 $X2=0 $Y2=0
cc_173 A2 N_A_215_47#_c_391_n 0.026248f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A2_c_191_n N_A_215_47#_c_391_n 0.00588644f $X=2.055 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A2_c_192_n N_A_215_47#_c_391_n 0.0109827f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A2_c_192_n N_A_215_47#_c_405_n 0.00680383f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B1_c_224_n N_C1_c_252_n 0.0289317f $X=2.545 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_178 N_B1_M1001_g N_C1_M1003_g 0.0206405f $X=2.475 $Y=1.985 $X2=0 $Y2=0
cc_179 B1 N_C1_c_253_n 6.40576e-19 $X=2.47 $Y=1.105 $X2=0 $Y2=0
cc_180 N_B1_c_223_n N_C1_c_253_n 0.0211366f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_181 N_B1_M1001_g N_VPWR_c_302_n 0.00323788f $X=2.475 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B1_M1001_g N_VPWR_c_303_n 0.00585385f $X=2.475 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B1_M1001_g N_VPWR_c_298_n 0.0111279f $X=2.475 $Y=1.985 $X2=0 $Y2=0
cc_184 N_B1_c_224_n N_VGND_c_350_n 0.00585385f $X=2.545 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B1_c_224_n N_VGND_c_351_n 0.011435f $X=2.545 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_224_n N_A_215_47#_c_391_n 0.00259343f $X=2.545 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_B1_c_224_n N_A_215_47#_c_405_n 0.00651785f $X=2.545 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_C1_M1003_g N_VPWR_c_302_n 0.00323788f $X=2.975 $Y=1.985 $X2=0 $Y2=0
cc_189 N_C1_M1003_g N_VPWR_c_306_n 0.00585385f $X=2.975 $Y=1.985 $X2=0 $Y2=0
cc_190 N_C1_M1003_g N_VPWR_c_298_n 0.011764f $X=2.975 $Y=1.985 $X2=0 $Y2=0
cc_191 N_C1_c_252_n N_VGND_c_350_n 0.00357668f $X=2.975 $Y=0.995 $X2=0 $Y2=0
cc_192 N_C1_c_252_n N_VGND_c_351_n 0.00656041f $X=2.975 $Y=0.995 $X2=0 $Y2=0
cc_193 X N_VPWR_c_305_n 0.0217551f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_194 N_X_M1007_s N_VPWR_c_298_n 0.00209319f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_195 X N_VPWR_c_298_n 0.0128119f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_196 N_X_c_282_n N_VGND_c_349_n 0.0217139f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_197 N_X_M1009_s N_VGND_c_351_n 0.00209319f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_198 N_X_c_282_n N_VGND_c_351_n 0.0127994f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_199 N_VPWR_c_298_n A_297_297# 0.0138923f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_200 N_VGND_c_351_n N_A_215_47#_M1002_s 0.00209319f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_201 N_VGND_c_351_n N_A_215_47#_M1005_d 0.00843348f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_346_n N_A_215_47#_c_390_n 0.0361618f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_203 N_VGND_c_347_n N_A_215_47#_c_390_n 0.0209752f $X=1.535 $Y=0 $X2=0 $Y2=0
cc_204 N_VGND_c_351_n N_A_215_47#_c_390_n 0.0124119f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_205 N_VGND_M1002_d N_A_215_47#_c_391_n 0.0022938f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_206 N_VGND_c_347_n N_A_215_47#_c_391_n 0.00193763f $X=1.535 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_348_n N_A_215_47#_c_391_n 0.0150374f $X=1.65 $Y=0.38 $X2=0 $Y2=0
cc_208 N_VGND_c_350_n N_A_215_47#_c_391_n 0.00193763f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_c_351_n N_A_215_47#_c_391_n 0.00850387f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_346_n N_A_215_47#_c_392_n 0.0120261f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_211 N_VGND_c_350_n N_A_215_47#_c_405_n 0.020922f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_351_n N_A_215_47#_c_405_n 0.0124119f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_351_n A_510_47# 0.0146485f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

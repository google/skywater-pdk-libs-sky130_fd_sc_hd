* File: sky130_fd_sc_hd__o21bai_1.spice
* Created: Thu Aug 27 14:36:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21bai_1.spice.pex"
.subckt sky130_fd_sc_hd__o21bai_1  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1007 N_A_105_352#_M1007_d N_B1_N_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_297_47#_M1002_d N_A_105_352#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10075 AS=0.169 PD=0.96 PS=1.82 NRD=5.532 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_297_47#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10075 PD=0.92 PS=0.96 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_297_47#_M1004_d N_A1_M1004_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_B1_N_M1005_g N_A_105_352#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.105444 AS=0.1092 PD=0.828169 PS=1.36 NRD=28.1316 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_105_352#_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1525 AS=0.251056 PD=1.305 PS=1.97183 NRD=5.91 NRS=11.8003 M=1 R=6.66667
+ SA=75000.5 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1001 A_388_297# N_A2_M1001_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=1 AD=0.1275
+ AS=0.1525 PD=1.255 PS=1.305 NRD=14.2628 NRS=0 M=1 R=6.66667 SA=75000.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_388_297# VPB PHIGHVT L=0.15 W=1 AD=0.28
+ AS=0.1275 PD=2.56 PS=1.255 NRD=0 NRS=14.2628 M=1 R=6.66667 SA=75001.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__o21bai_1.spice.SKY130_FD_SC_HD__O21BAI_1.pxi"
*
.ends
*
*

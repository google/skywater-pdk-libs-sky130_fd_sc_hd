* File: sky130_fd_sc_hd__nand4b_2.spice.SKY130_FD_SC_HD__NAND4B_2.pxi
* Created: Thu Aug 27 14:30:35 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4B_2%A_N N_A_N_M1017_g N_A_N_M1007_g A_N A_N
+ N_A_N_c_86_n PM_SKY130_FD_SC_HD__NAND4B_2%A_N
x_PM_SKY130_FD_SC_HD__NAND4B_2%A_27_47# N_A_27_47#_M1017_s N_A_27_47#_M1007_s
+ N_A_27_47#_c_113_n N_A_27_47#_M1002_g N_A_27_47#_M1000_g N_A_27_47#_c_114_n
+ N_A_27_47#_M1003_g N_A_27_47#_M1015_g N_A_27_47#_c_115_n N_A_27_47#_c_123_n
+ N_A_27_47#_c_116_n N_A_27_47#_c_117_n N_A_27_47#_c_118_n N_A_27_47#_c_119_n
+ N_A_27_47#_c_125_n N_A_27_47#_c_139_n N_A_27_47#_c_120_n
+ PM_SKY130_FD_SC_HD__NAND4B_2%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND4B_2%B N_B_c_201_n N_B_M1006_g N_B_M1011_g N_B_c_202_n
+ N_B_M1009_g N_B_M1013_g B B B N_B_c_204_n PM_SKY130_FD_SC_HD__NAND4B_2%B
x_PM_SKY130_FD_SC_HD__NAND4B_2%C N_C_M1010_g N_C_c_250_n N_C_M1004_g N_C_M1016_g
+ N_C_c_251_n N_C_M1014_g C C C N_C_c_253_n PM_SKY130_FD_SC_HD__NAND4B_2%C
x_PM_SKY130_FD_SC_HD__NAND4B_2%D N_D_M1008_g N_D_c_297_n N_D_M1001_g N_D_M1012_g
+ N_D_c_298_n N_D_M1005_g D D N_D_c_300_n PM_SKY130_FD_SC_HD__NAND4B_2%D
x_PM_SKY130_FD_SC_HD__NAND4B_2%VPWR N_VPWR_M1007_d N_VPWR_M1000_s N_VPWR_M1015_s
+ N_VPWR_M1013_d N_VPWR_M1016_d N_VPWR_M1012_d N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n VPWR N_VPWR_c_348_n
+ N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_337_n
+ PM_SKY130_FD_SC_HD__NAND4B_2%VPWR
x_PM_SKY130_FD_SC_HD__NAND4B_2%Y N_Y_M1002_s N_Y_M1000_d N_Y_M1011_s N_Y_M1010_s
+ N_Y_M1008_s N_Y_c_423_n N_Y_c_416_n N_Y_c_426_n N_Y_c_417_n N_Y_c_454_n
+ N_Y_c_418_n N_Y_c_459_n N_Y_c_419_n N_Y_c_420_n Y Y Y Y
+ PM_SKY130_FD_SC_HD__NAND4B_2%Y
x_PM_SKY130_FD_SC_HD__NAND4B_2%VGND N_VGND_M1017_d N_VGND_M1001_d N_VGND_c_498_n
+ N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n VGND N_VGND_c_502_n
+ N_VGND_c_503_n N_VGND_c_504_n N_VGND_c_505_n PM_SKY130_FD_SC_HD__NAND4B_2%VGND
x_PM_SKY130_FD_SC_HD__NAND4B_2%A_215_47# N_A_215_47#_M1002_d N_A_215_47#_M1003_d
+ N_A_215_47#_M1009_s N_A_215_47#_c_566_n N_A_215_47#_c_567_n
+ N_A_215_47#_c_576_n N_A_215_47#_c_568_n N_A_215_47#_c_569_n
+ PM_SKY130_FD_SC_HD__NAND4B_2%A_215_47#
x_PM_SKY130_FD_SC_HD__NAND4B_2%A_465_47# N_A_465_47#_M1006_d N_A_465_47#_M1004_d
+ N_A_465_47#_c_606_n PM_SKY130_FD_SC_HD__NAND4B_2%A_465_47#
x_PM_SKY130_FD_SC_HD__NAND4B_2%A_655_47# N_A_655_47#_M1004_s N_A_655_47#_M1014_s
+ N_A_655_47#_M1005_s N_A_655_47#_c_622_n N_A_655_47#_c_647_n
+ N_A_655_47#_c_623_n N_A_655_47#_c_624_n N_A_655_47#_c_625_n
+ PM_SKY130_FD_SC_HD__NAND4B_2%A_655_47#
cc_1 VNB N_A_N_M1017_g 0.0432803f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.0134299f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_86_n 0.037293f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_47#_c_113_n 0.0200369f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_5 VNB N_A_27_47#_c_114_n 0.01577f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_A_27_47#_c_115_n 0.0147647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_116_n 0.00359176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_117_n 6.77426e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_118_n 0.0230682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_119_n 0.0116462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_120_n 0.0509972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_201_n 0.0160098f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_B_c_202_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB B 0.00757421f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_15 VNB N_B_c_204_n 0.0483309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_C_c_250_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_17 VNB N_C_c_251_n 0.0168109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB C 0.00769179f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_19 VNB N_C_c_253_n 0.0401218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D_c_297_n 0.0168109f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_21 VNB N_D_c_298_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB D 0.00895653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_D_c_300_n 0.0622746f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.53
cc_24 VNB N_VPWR_c_337_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB Y 9.87696e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_498_n 0.0056135f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_27 VNB N_VGND_c_499_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_28 VNB N_VGND_c_500_n 0.0896918f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_501_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_30 VNB N_VGND_c_502_n 0.0143366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_503_n 0.0200298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_504_n 0.29037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_505_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_215_47#_c_566_n 0.00217944f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_35 VNB N_A_215_47#_c_567_n 0.0071501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_215_47#_c_568_n 0.00206682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_215_47#_c_569_n 0.00723412f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.53
cc_38 VNB N_A_465_47#_c_606_n 0.0103416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_655_47#_c_622_n 0.0086278f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_40 VNB N_A_655_47#_c_623_n 0.0121718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_655_47#_c_624_n 0.0182049f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.53
cc_42 VNB N_A_655_47#_c_625_n 0.00250338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_A_N_M1007_g 0.0725217f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_44 VPB A_N 0.01652f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_45 VPB N_A_N_c_86_n 0.0103072f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_46 VPB N_A_27_47#_M1000_g 0.0228659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_M1015_g 0.0178886f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.16
cc_48 VPB N_A_27_47#_c_123_n 0.0147827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_117_n 0.00711948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_125_n 0.0125758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_120_n 0.0134448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_B_M1011_g 0.0183716f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_53 VPB N_B_M1013_g 0.0250398f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_54 VPB N_B_c_204_n 0.0115682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_C_M1010_g 0.0250398f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_56 VPB N_C_M1016_g 0.0193602f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_57 VPB N_C_c_253_n 0.00822359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_D_M1008_g 0.0193602f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_59 VPB N_D_M1012_g 0.0258005f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_60 VPB N_D_c_300_n 0.0172717f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.53
cc_61 VPB N_VPWR_c_338_n 0.0117084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_339_n 0.00358794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_340_n 0.00617918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_341_n 0.004085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_342_n 0.0126404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_343_n 0.0449841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_344_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_345_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_346_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_347_n 0.00496849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_348_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_349_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_350_n 0.0143307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_351_n 0.0297812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_352_n 0.0122777f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_337_n 0.0435245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_Y_c_416_n 0.00412785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_Y_c_417_n 0.0106294f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_Y_c_418_n 0.00539385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_Y_c_419_n 0.00223196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_Y_c_420_n 0.00223196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB Y 9.38585e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB Y 0.00112774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 N_A_N_M1017_g N_A_27_47#_c_116_n 0.0112496f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_85 A_N N_A_27_47#_c_116_n 0.00553612f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_N_c_86_n N_A_27_47#_c_116_n 0.00227579f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_N_M1007_g N_A_27_47#_c_117_n 0.026127f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_88 A_N N_A_27_47#_c_117_n 0.0268282f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A_N_c_86_n N_A_27_47#_c_117_n 0.00227579f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_N_M1017_g N_A_27_47#_c_119_n 0.0165563f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_91 A_N N_A_27_47#_c_119_n 0.0174382f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A_N_c_86_n N_A_27_47#_c_119_n 0.00393367f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_N_M1007_g N_A_27_47#_c_125_n 0.016571f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_94 A_N N_A_27_47#_c_125_n 0.0134295f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_N_c_86_n N_A_27_47#_c_125_n 0.00241083f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_96 A_N N_A_27_47#_c_139_n 0.0132649f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_97 N_A_N_c_86_n N_A_27_47#_c_139_n 0.0062407f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_N_c_86_n N_A_27_47#_c_120_n 0.00654498f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_N_M1007_g N_VPWR_c_338_n 0.00626656f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_100 N_A_N_M1007_g N_VPWR_c_350_n 0.00339367f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_101 N_A_N_M1007_g N_VPWR_c_351_n 0.010062f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_102 N_A_N_M1007_g N_VPWR_c_337_n 0.00488264f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_103 N_A_N_M1017_g N_VGND_c_498_n 0.00944899f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_N_M1017_g N_VGND_c_502_n 0.00339367f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_N_M1017_g N_VGND_c_504_n 0.00489827f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_N_M1017_g N_A_215_47#_c_567_n 0.00438858f $X=0.47 $Y=0.445 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_114_n N_B_c_201_n 0.0230042f $X=1.83 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_27_47#_M1015_g N_B_M1011_g 0.0230042f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_120_n B 0.00193346f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_120_n N_B_c_204_n 0.0230042f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_125_n N_VPWR_M1007_d 9.71102e-19 $X=0.585 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_27_47#_M1000_g N_VPWR_c_338_n 8.89484e-19 $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_117_n N_VPWR_c_338_n 0.0214963f $X=0.585 $Y=1.915 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_118_n N_VPWR_c_338_n 0.0177704f $X=1.215 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_125_n N_VPWR_c_338_n 0.00842813f $X=0.585 $Y=2 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_120_n N_VPWR_c_338_n 0.0059184f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_27_47#_M1015_g N_VPWR_c_339_n 0.00146339f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_M1000_g N_VPWR_c_344_n 0.00541359f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_M1015_g N_VPWR_c_344_n 0.00541359f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_c_123_n N_VPWR_c_350_n 0.0169243f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_125_n N_VPWR_c_350_n 0.00246266f $X=0.585 $Y=2 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1000_g N_VPWR_c_351_n 0.00336547f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_125_n N_VPWR_c_351_n 0.00725006f $X=0.585 $Y=2 $X2=0 $Y2=0
cc_124 N_A_27_47#_M1007_s N_VPWR_c_337_n 0.0022756f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_M1000_g N_VPWR_c_337_n 0.0108251f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_27_47#_M1015_g N_VPWR_c_337_n 0.00952874f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_123_n N_VPWR_c_337_n 0.00960198f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_125_n N_VPWR_c_337_n 0.00490838f $X=0.585 $Y=2 $X2=0 $Y2=0
cc_129 N_A_27_47#_M1000_g N_Y_c_423_n 0.00901111f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_27_47#_M1015_g N_Y_c_423_n 0.00975139f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_27_47#_M1015_g N_Y_c_416_n 0.0157539f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_27_47#_M1015_g N_Y_c_426_n 6.1949e-19 $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_113_n Y 0.00322939f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_114_n Y 0.00237069f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_27_47#_M1000_g Y 0.0036711f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_27_47#_M1015_g Y 0.00105585f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_113_n Y 0.00266571f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1000_g Y 0.00296785f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_114_n Y 0.00332434f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1015_g Y 0.00311352f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_118_n Y 0.0130894f $X=1.215 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_120_n Y 0.0244855f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_119_n N_VGND_M1017_d 9.6948e-19 $X=0.585 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_144 N_A_27_47#_c_113_n N_VGND_c_498_n 0.00235149f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_118_n N_VGND_c_498_n 0.00565372f $X=1.215 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_119_n N_VGND_c_498_n 0.00721829f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_113_n N_VGND_c_500_n 0.00357877f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_114_n N_VGND_c_500_n 0.00357877f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_115_n N_VGND_c_502_n 0.0169243f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_119_n N_VGND_c_502_n 0.00247115f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_M1017_s N_VGND_c_504_n 0.0022756f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_113_n N_VGND_c_504_n 0.00655123f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_114_n N_VGND_c_504_n 0.0052923f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_115_n N_VGND_c_504_n 0.00960198f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_119_n N_VGND_c_504_n 0.00494211f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_113_n N_A_215_47#_c_567_n 4.72107e-19 $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_116_n N_A_215_47#_c_567_n 0.00457368f $X=0.585 $Y=1.075
+ $X2=0 $Y2=0
cc_158 N_A_27_47#_c_118_n N_A_215_47#_c_567_n 0.0199821f $X=1.215 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_119_n N_A_215_47#_c_567_n 0.00842813f $X=0.585 $Y=0.72 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_120_n N_A_215_47#_c_567_n 0.00598881f $X=1.83 $Y=1.16 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_113_n N_A_215_47#_c_576_n 0.0116213f $X=1.41 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_114_n N_A_215_47#_c_576_n 0.01333f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_118_n N_A_215_47#_c_576_n 0.00165197f $X=1.215 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_120_n N_A_215_47#_c_576_n 3.01257e-19 $X=1.83 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_114_n N_A_215_47#_c_568_n 7.34403e-19 $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_166 B C 0.0137573f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_167 N_B_c_204_n C 8.19518e-19 $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_168 B N_C_c_253_n 7.3417e-19 $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_169 N_B_c_204_n N_C_c_253_n 0.0100132f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B_M1011_g N_VPWR_c_339_n 0.00146448f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B_M1013_g N_VPWR_c_340_n 0.00334219f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_172 N_B_M1011_g N_VPWR_c_348_n 0.00541359f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B_M1013_g N_VPWR_c_348_n 0.00541359f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B_M1011_g N_VPWR_c_337_n 0.00952874f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_175 N_B_M1013_g N_VPWR_c_337_n 0.0108276f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B_M1011_g N_Y_c_423_n 6.1949e-19 $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B_M1011_g N_Y_c_416_n 0.0119784f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_178 B N_Y_c_416_n 0.021194f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_179 N_B_M1011_g N_Y_c_426_n 0.00975139f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B_M1013_g N_Y_c_426_n 0.0145598f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B_M1013_g N_Y_c_417_n 0.0147646f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_182 B N_Y_c_417_n 0.0348641f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_183 N_B_c_204_n N_Y_c_417_n 0.00681999f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_184 N_B_M1011_g N_Y_c_419_n 0.00149073f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_185 N_B_M1013_g N_Y_c_419_n 0.00149073f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_186 B N_Y_c_419_n 0.0266427f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_187 N_B_c_204_n N_Y_c_419_n 0.00222737f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_188 N_B_c_201_n Y 9.21687e-19 $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_189 B Y 0.0132337f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_190 N_B_c_204_n Y 0.00105183f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B_c_201_n N_VGND_c_500_n 0.00411651f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B_c_202_n N_VGND_c_500_n 0.00357877f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B_c_201_n N_VGND_c_504_n 0.00574374f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B_c_202_n N_VGND_c_504_n 0.00660224f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_195 B N_A_215_47#_c_568_n 0.00978542f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_196 N_B_c_201_n N_A_215_47#_c_569_n 0.0134979f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B_c_202_n N_A_215_47#_c_569_n 0.0113074f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_198 B N_A_215_47#_c_569_n 0.0681255f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_199 N_B_c_204_n N_A_215_47#_c_569_n 0.00935154f $X=2.865 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B_c_201_n N_A_465_47#_c_606_n 0.0028244f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B_c_202_n N_A_465_47#_c_606_n 0.0112708f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_202 B N_A_465_47#_c_606_n 0.00175186f $X=2.93 $Y=1.105 $X2=0 $Y2=0
cc_203 N_B_c_202_n N_A_655_47#_c_622_n 5.43931e-19 $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_204 N_C_M1016_g N_D_M1008_g 0.0210533f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_205 N_C_c_251_n N_D_c_297_n 0.00918758f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_206 C D 0.0167609f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_207 C N_D_c_300_n 0.00606758f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_208 N_C_c_253_n N_D_c_300_n 0.0239875f $X=4.03 $Y=1.16 $X2=0 $Y2=0
cc_209 N_C_M1010_g N_VPWR_c_340_n 0.0158485f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_210 N_C_M1016_g N_VPWR_c_341_n 0.00164968f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_211 N_C_M1010_g N_VPWR_c_346_n 0.00541359f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_212 N_C_M1016_g N_VPWR_c_346_n 0.00541359f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_213 N_C_M1010_g N_VPWR_c_337_n 0.0109543f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_214 N_C_M1016_g N_VPWR_c_337_n 0.0097341f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_215 N_C_M1010_g N_Y_c_417_n 0.0147646f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_216 C N_Y_c_417_n 0.0180842f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_217 N_C_M1010_g N_Y_c_454_n 0.0145598f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_218 N_C_M1016_g N_Y_c_454_n 0.0101674f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_219 N_C_M1016_g N_Y_c_418_n 0.0126115f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_220 C N_Y_c_418_n 0.0382251f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_221 N_C_c_253_n N_Y_c_418_n 0.00379745f $X=4.03 $Y=1.16 $X2=0 $Y2=0
cc_222 N_C_M1016_g N_Y_c_459_n 6.0188e-19 $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_223 N_C_M1010_g N_Y_c_420_n 0.00149073f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_224 N_C_M1016_g N_Y_c_420_n 0.00149073f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_225 C N_Y_c_420_n 0.0266427f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_226 N_C_c_253_n N_Y_c_420_n 0.00243558f $X=4.03 $Y=1.16 $X2=0 $Y2=0
cc_227 N_C_c_250_n N_VGND_c_500_n 0.00357877f $X=3.61 $Y=0.995 $X2=0 $Y2=0
cc_228 N_C_c_251_n N_VGND_c_500_n 0.00411651f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_229 N_C_c_250_n N_VGND_c_504_n 0.00660224f $X=3.61 $Y=0.995 $X2=0 $Y2=0
cc_230 N_C_c_251_n N_VGND_c_504_n 0.00590508f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_231 N_C_c_250_n N_A_215_47#_c_569_n 5.43931e-19 $X=3.61 $Y=0.995 $X2=0 $Y2=0
cc_232 N_C_c_250_n N_A_465_47#_c_606_n 0.0112708f $X=3.61 $Y=0.995 $X2=0 $Y2=0
cc_233 N_C_c_251_n N_A_465_47#_c_606_n 0.00285917f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_234 N_C_c_250_n N_A_655_47#_c_622_n 0.0113779f $X=3.61 $Y=0.995 $X2=0 $Y2=0
cc_235 N_C_c_251_n N_A_655_47#_c_622_n 0.0123515f $X=4.03 $Y=0.995 $X2=0 $Y2=0
cc_236 C N_A_655_47#_c_622_n 0.0589687f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_237 N_C_c_253_n N_A_655_47#_c_622_n 0.00516505f $X=4.03 $Y=1.16 $X2=0 $Y2=0
cc_238 C N_A_655_47#_c_625_n 0.0245883f $X=4.28 $Y=1.105 $X2=0 $Y2=0
cc_239 N_C_c_253_n N_A_655_47#_c_625_n 0.00127974f $X=4.03 $Y=1.16 $X2=0 $Y2=0
cc_240 N_D_M1008_g N_VPWR_c_341_n 0.00164968f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_241 N_D_M1012_g N_VPWR_c_343_n 0.0223289f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_242 D N_VPWR_c_343_n 0.0256479f $X=5.2 $Y=1.105 $X2=0 $Y2=0
cc_243 N_D_c_300_n N_VPWR_c_343_n 0.00883269f $X=4.96 $Y=1.16 $X2=0 $Y2=0
cc_244 N_D_M1008_g N_VPWR_c_349_n 0.00541359f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_245 N_D_M1012_g N_VPWR_c_349_n 0.00541359f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_246 N_D_M1008_g N_VPWR_c_337_n 0.0097341f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_247 N_D_M1012_g N_VPWR_c_337_n 0.0106821f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_248 N_D_M1008_g N_Y_c_454_n 6.0188e-19 $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_249 N_D_M1008_g N_Y_c_418_n 0.0175874f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_250 N_D_M1012_g N_Y_c_418_n 0.00725171f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_251 D N_Y_c_418_n 0.0198454f $X=5.2 $Y=1.105 $X2=0 $Y2=0
cc_252 N_D_c_300_n N_Y_c_418_n 0.00243558f $X=4.96 $Y=1.16 $X2=0 $Y2=0
cc_253 N_D_M1008_g N_Y_c_459_n 0.011789f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_254 N_D_M1012_g N_Y_c_459_n 0.0106465f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_255 N_D_c_297_n N_VGND_c_499_n 0.00268723f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_256 N_D_c_298_n N_VGND_c_499_n 0.00268723f $X=4.96 $Y=0.995 $X2=0 $Y2=0
cc_257 N_D_c_297_n N_VGND_c_500_n 0.00436487f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_258 N_D_c_298_n N_VGND_c_503_n 0.00422241f $X=4.96 $Y=0.995 $X2=0 $Y2=0
cc_259 N_D_c_297_n N_VGND_c_504_n 0.00609471f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_260 N_D_c_298_n N_VGND_c_504_n 0.00672659f $X=4.96 $Y=0.995 $X2=0 $Y2=0
cc_261 N_D_c_297_n N_A_655_47#_c_623_n 0.0126994f $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_262 N_D_c_298_n N_A_655_47#_c_623_n 0.0102289f $X=4.96 $Y=0.995 $X2=0 $Y2=0
cc_263 D N_A_655_47#_c_623_n 0.0547017f $X=5.2 $Y=1.105 $X2=0 $Y2=0
cc_264 N_D_c_300_n N_A_655_47#_c_623_n 0.0104862f $X=4.96 $Y=1.16 $X2=0 $Y2=0
cc_265 N_D_c_297_n N_A_655_47#_c_624_n 5.31244e-19 $X=4.54 $Y=0.995 $X2=0 $Y2=0
cc_266 N_D_c_298_n N_A_655_47#_c_624_n 0.00635814f $X=4.96 $Y=0.995 $X2=0 $Y2=0
cc_267 N_D_c_300_n N_A_655_47#_c_625_n 0.00119738f $X=4.96 $Y=1.16 $X2=0 $Y2=0
cc_268 N_VPWR_c_337_n N_Y_M1000_d 0.00215201f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_c_337_n N_Y_M1011_s 0.00215201f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_337_n N_Y_M1010_s 0.00215201f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_271 N_VPWR_c_337_n N_Y_M1008_s 0.00215201f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_272 N_VPWR_c_344_n N_Y_c_423_n 0.0189039f $X=1.955 $Y=2.72 $X2=0 $Y2=0
cc_273 N_VPWR_c_337_n N_Y_c_423_n 0.0122217f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_274 N_VPWR_M1015_s N_Y_c_416_n 0.00167154f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_275 N_VPWR_c_339_n N_Y_c_416_n 0.0129161f $X=2.04 $Y=2 $X2=0 $Y2=0
cc_276 N_VPWR_c_348_n N_Y_c_426_n 0.0189039f $X=2.795 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_337_n N_Y_c_426_n 0.0122217f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_M1013_d N_Y_c_417_n 0.0104725f $X=2.745 $Y=1.485 $X2=0 $Y2=0
cc_279 N_VPWR_c_340_n N_Y_c_417_n 0.0518301f $X=3.27 $Y=2 $X2=0 $Y2=0
cc_280 N_VPWR_c_346_n N_Y_c_454_n 0.0189039f $X=4.105 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_337_n N_Y_c_454_n 0.0122217f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_M1016_d N_Y_c_418_n 0.0026359f $X=4.055 $Y=1.485 $X2=0 $Y2=0
cc_283 N_VPWR_c_341_n N_Y_c_418_n 0.0203677f $X=4.225 $Y=2 $X2=0 $Y2=0
cc_284 N_VPWR_c_349_n N_Y_c_459_n 0.0189039f $X=5.035 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_337_n N_Y_c_459_n 0.0122217f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_c_338_n Y 0.0108296f $X=1.2 $Y=1.66 $X2=0 $Y2=0
cc_287 N_Y_M1002_s N_VGND_c_504_n 0.00216833f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_288 Y N_A_215_47#_c_567_n 0.00275701f $X=1.635 $Y=0.85 $X2=0 $Y2=0
cc_289 N_Y_M1002_s N_A_215_47#_c_576_n 0.00304479f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_290 Y N_A_215_47#_c_576_n 0.0160863f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_291 N_Y_c_416_n N_A_215_47#_c_568_n 0.00210886f $X=2.295 $Y=1.555 $X2=0 $Y2=0
cc_292 Y N_A_215_47#_c_568_n 0.0108762f $X=1.55 $Y=0.765 $X2=0 $Y2=0
cc_293 N_Y_c_417_n N_A_655_47#_c_622_n 0.00446358f $X=3.605 $Y=1.555 $X2=0 $Y2=0
cc_294 N_Y_c_418_n N_A_655_47#_c_623_n 0.00496247f $X=4.535 $Y=1.555 $X2=0 $Y2=0
cc_295 N_VGND_c_504_n N_A_215_47#_M1002_d 0.00209324f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_296 N_VGND_c_504_n N_A_215_47#_M1003_d 0.00235053f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_297 N_VGND_c_504_n N_A_215_47#_M1009_s 0.00210147f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_298 N_VGND_c_498_n N_A_215_47#_c_566_n 0.0171705f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_299 N_VGND_c_500_n N_A_215_47#_c_566_n 0.0173346f $X=4.665 $Y=0 $X2=0 $Y2=0
cc_300 N_VGND_c_504_n N_A_215_47#_c_566_n 0.00961661f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_c_500_n N_A_215_47#_c_576_n 0.0476962f $X=4.665 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_504_n N_A_215_47#_c_576_n 0.0301625f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_303 N_VGND_c_500_n N_A_215_47#_c_569_n 0.00250396f $X=4.665 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_504_n N_A_215_47#_c_569_n 0.00581016f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_504_n N_A_465_47#_M1006_d 0.00215227f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_306 N_VGND_c_504_n N_A_465_47#_M1004_d 0.00215227f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_500_n N_A_465_47#_c_606_n 0.0982292f $X=4.665 $Y=0 $X2=0 $Y2=0
cc_308 N_VGND_c_504_n N_A_465_47#_c_606_n 0.0613107f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_504_n N_A_655_47#_M1004_s 0.00210147f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_310 N_VGND_c_504_n N_A_655_47#_M1014_s 0.00321471f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_504_n N_A_655_47#_M1005_s 0.00209319f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_500_n N_A_655_47#_c_622_n 0.00250396f $X=4.665 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_504_n N_A_655_47#_c_622_n 0.00576854f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_500_n N_A_655_47#_c_647_n 0.0176675f $X=4.665 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_504_n N_A_655_47#_c_647_n 0.00992425f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_M1001_d N_A_655_47#_c_623_n 0.00162148f $X=4.615 $Y=0.235 $X2=0
+ $Y2=0
cc_317 N_VGND_c_499_n N_A_655_47#_c_623_n 0.0122675f $X=4.75 $Y=0.38 $X2=0 $Y2=0
cc_318 N_VGND_c_500_n N_A_655_47#_c_623_n 0.00253038f $X=4.665 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_503_n N_A_655_47#_c_623_n 0.00203746f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_504_n N_A_655_47#_c_623_n 0.00932974f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_503_n N_A_655_47#_c_624_n 0.0213324f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_504_n N_A_655_47#_c_624_n 0.0126042f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_504_n N_A_655_47#_c_625_n 0.00117665f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_324 N_A_215_47#_c_569_n N_A_465_47#_M1006_d 0.00162207f $X=2.88 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_325 N_A_215_47#_M1009_s N_A_465_47#_c_606_n 0.00479304f $X=2.745 $Y=0.235
+ $X2=0 $Y2=0
cc_326 N_A_215_47#_c_569_n N_A_465_47#_c_606_n 0.0410913f $X=2.88 $Y=0.72 $X2=0
+ $Y2=0
cc_327 N_A_215_47#_c_569_n N_A_655_47#_c_622_n 0.0231988f $X=2.88 $Y=0.72 $X2=0
+ $Y2=0
cc_328 N_A_465_47#_c_606_n N_A_655_47#_M1004_s 0.00501743f $X=3.82 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_329 N_A_465_47#_M1004_d N_A_655_47#_c_622_n 0.00162207f $X=3.685 $Y=0.235
+ $X2=0 $Y2=0
cc_330 N_A_465_47#_c_606_n N_A_655_47#_c_622_n 0.0410913f $X=3.82 $Y=0.38 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__fa_2.spice
* Created: Tue Sep  1 19:08:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__fa_2.pex.spice"
.subckt sky130_fd_sc_hd__fa_2  VNB VPB A B CIN VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_80_21#_M1008_g N_COUT_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_80_21#_M1014_g N_COUT_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.125626 AS=0.08775 PD=1.21495 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1004 A_294_47# N_A_M1004_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42 AD=0.06825
+ AS=0.0811738 PD=0.745 PS=0.785047 NRD=30.708 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1026 N_A_80_21#_M1026_d N_B_M1026_g A_294_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.06825 PD=0.69 PS=0.745 NRD=0 NRS=30.708 M=1 R=2.8 SA=75001.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1025 N_A_473_47#_M1025_d N_CIN_M1025_g N_A_80_21#_M1026_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_M1029_g N_A_473_47#_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1028 N_A_473_47#_M1028_d N_B_M1028_g N_VGND_M1029_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_A_829_47#_M1017_d N_B_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_CIN_M1015_g N_A_829_47#_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1021 N_A_829_47#_M1021_d N_A_M1021_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.0567 PD=0.715 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75003
+ A=0.063 P=1.14 MULT=1
MM1027 N_A_1086_47#_M1027_d N_A_80_21#_M1027_g N_A_829_47#_M1021_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0819 AS=0.06195 PD=0.81 PS=0.715 NRD=15.708 NRS=5.712 M=1
+ R=2.8 SA=75001.5 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1003 A_1194_47# N_CIN_M1003_g N_A_1086_47#_M1027_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=15.708 M=1 R=2.8 SA=75002
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 A_1266_47# N_B_M1006_g A_1194_47# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0441 PD=0.75 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8 SA=75002.4 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g A_1266_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0803495 AS=0.0693 PD=0.781121 PS=0.75 NRD=0 NRS=31.428 M=1 R=2.8
+ SA=75002.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1018 N_SUM_M1018_d N_A_1086_47#_M1018_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.65 AD=0.12675 AS=0.12435 PD=1.04 PS=1.20888 NRD=21.228 NRS=12.912 M=1
+ R=4.33333 SA=75002.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1031 N_SUM_M1018_d N_A_1086_47#_M1031_g N_VGND_M1031_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12675 AS=0.169 PD=1.04 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_80_21#_M1005_g N_COUT_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A_80_21#_M1019_g N_COUT_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.182362 AS=0.135 PD=1.62577 PS=1.27 NRD=6.8753 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1002 A_289_371# N_A_M1002_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=0.63
+ AD=0.092925 AS=0.114888 PD=0.925 PS=1.02423 NRD=28.9196 NRS=3.1126 M=1 R=4.2
+ SA=75001.1 SB=75001.9 A=0.0945 P=1.56 MULT=1
MM1013 N_A_80_21#_M1013_d N_B_M1013_g A_289_371# VPB PHIGHVT L=0.15 W=0.63
+ AD=0.102375 AS=0.092925 PD=0.955 PS=0.925 NRD=15.6221 NRS=28.9196 M=1 R=4.2
+ SA=75001.5 SB=75001.5 A=0.0945 P=1.56 MULT=1
MM1000 N_A_473_371#_M1000_d N_CIN_M1000_g N_A_80_21#_M1013_d VPB PHIGHVT L=0.15
+ W=0.63 AD=0.08505 AS=0.102375 PD=0.9 PS=0.955 NRD=0 NRS=0 M=1 R=4.2 SA=75002
+ SB=75001 A=0.0945 P=1.56 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_473_371#_M1000_d VPB PHIGHVT L=0.15 W=0.63
+ AD=0.08505 AS=0.08505 PD=0.9 PS=0.9 NRD=0 NRS=0 M=1 R=4.2 SA=75002.4
+ SB=75000.6 A=0.0945 P=1.56 MULT=1
MM1023 N_A_473_371#_M1023_d N_B_M1023_g N_VPWR_M1030_d VPB PHIGHVT L=0.15 W=0.63
+ AD=0.1638 AS=0.08505 PD=1.78 PS=0.9 NRD=0 NRS=0 M=1 R=4.2 SA=75002.8
+ SB=75000.2 A=0.0945 P=1.56 MULT=1
MM1024 N_A_829_369#_M1024_d N_B_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.8 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_CIN_M1016_g N_A_829_369#_M1024_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.0864 PD=0.91 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1012 N_A_829_369#_M1012_d N_A_M1012_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0944 AS=0.0864 PD=0.935 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1020 N_A_1086_47#_M1020_d N_A_80_21#_M1020_g N_A_829_369#_M1012_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.088 AS=0.0944 PD=0.915 PS=0.935 NRD=0 NRS=6.1464 M=1
+ R=4.26667 SA=75001.5 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1007 A_1171_369# N_CIN_M1007_g N_A_1086_47#_M1020_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.104441 AS=0.088 PD=0.972598 PS=0.915 NRD=33.293 NRS=0 M=1 R=4.26667
+ SA=75001.9 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1010 A_1266_371# N_B_M1010_g A_1171_369# VPB PHIGHVT L=0.15 W=0.63 AD=0.12285
+ AS=0.102809 PD=1.02 PS=0.957402 NRD=43.7734 NRS=33.8249 M=1 R=4.2 SA=75002.4
+ SB=75001.6 A=0.0945 P=1.56 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g A_1266_371# VPB PHIGHVT L=0.15 W=0.63
+ AD=0.114888 AS=0.12285 PD=1.02423 PS=1.02 NRD=14.0658 NRS=43.7734 M=1 R=4.2
+ SA=75002.9 SB=75001.1 A=0.0945 P=1.56 MULT=1
MM1001 N_VPWR_M1022_d N_A_1086_47#_M1001_g N_SUM_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.182362 AS=0.135 PD=1.62577 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_1086_47#_M1011_g N_SUM_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.8993 P=20.53
*
.include "sky130_fd_sc_hd__fa_2.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_hd__or2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
M1000 X a_219_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=4.057e+11p ps=4.04e+06u
M1001 VGND A a_219_297# VNB nshort w=420000u l=150000u
+  ad=5.1875e+11p pd=4.32e+06u as=1.134e+11p ps=1.38e+06u
M1002 a_219_297# a_27_53# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B_N a_27_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1004 X a_219_297# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1005 a_301_297# a_27_53# a_219_297# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u
M1006 VPWR A a_301_297# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_53# B_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
.ends


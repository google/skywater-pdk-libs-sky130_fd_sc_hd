* File: sky130_fd_sc_hd__clkbuf_4.spice.SKY130_FD_SC_HD__CLKBUF_4.pxi
* Created: Thu Aug 27 14:11:01 2020
* 
x_PM_SKY130_FD_SC_HD__CLKBUF_4%A N_A_M1003_g N_A_M1006_g A A N_A_c_57_n
+ PM_SKY130_FD_SC_HD__CLKBUF_4%A
x_PM_SKY130_FD_SC_HD__CLKBUF_4%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1006_s
+ N_A_27_47#_M1002_g N_A_27_47#_M1000_g N_A_27_47#_M1007_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1008_g N_A_27_47#_M1004_g N_A_27_47#_M1009_g N_A_27_47#_M1005_g
+ N_A_27_47#_c_98_n N_A_27_47#_c_106_n N_A_27_47#_c_117_n N_A_27_47#_c_107_n
+ N_A_27_47#_c_122_n N_A_27_47#_c_147_p N_A_27_47#_c_99_n N_A_27_47#_c_108_n
+ N_A_27_47#_c_100_n PM_SKY130_FD_SC_HD__CLKBUF_4%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKBUF_4%VPWR N_VPWR_M1006_d N_VPWR_M1007_s N_VPWR_M1009_s
+ N_VPWR_c_188_n N_VPWR_c_189_n N_VPWR_c_190_n N_VPWR_c_191_n VPWR
+ N_VPWR_c_192_n N_VPWR_c_193_n N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_196_n
+ N_VPWR_c_187_n PM_SKY130_FD_SC_HD__CLKBUF_4%VPWR
x_PM_SKY130_FD_SC_HD__CLKBUF_4%X N_X_M1000_d N_X_M1004_d N_X_M1002_d N_X_M1008_d
+ N_X_c_231_n N_X_c_273_n N_X_c_232_n N_X_c_233_n N_X_c_252_n N_X_c_256_n
+ N_X_c_234_n N_X_c_280_n X X X N_X_c_237_n PM_SKY130_FD_SC_HD__CLKBUF_4%X
x_PM_SKY130_FD_SC_HD__CLKBUF_4%VGND N_VGND_M1003_d N_VGND_M1001_s N_VGND_M1005_s
+ N_VGND_c_297_n N_VGND_c_298_n N_VGND_c_299_n N_VGND_c_300_n VGND
+ N_VGND_c_301_n N_VGND_c_302_n N_VGND_c_303_n N_VGND_c_304_n N_VGND_c_305_n
+ N_VGND_c_306_n PM_SKY130_FD_SC_HD__CLKBUF_4%VGND
cc_1 VNB N_A_M1003_g 0.0322943f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB A 0.00620969f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_3 VNB N_A_c_57_n 0.0251851f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_4 VNB N_A_27_47#_M1002_g 4.17371e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_5 VNB N_A_27_47#_M1000_g 0.0295782f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_6 VNB N_A_27_47#_M1007_g 4.55724e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_7 VNB N_A_27_47#_M1001_g 0.0276999f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_8 VNB N_A_27_47#_M1008_g 4.56723e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1004_g 0.0276748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1009_g 5.58244e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1005_g 0.0366072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_98_n 0.0330143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_99_n 0.0131987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_100_n 0.0707961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_187_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_X_c_231_n 6.31183e-19 $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_17 VNB N_X_c_232_n 0.00518223f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_18 VNB N_X_c_233_n 0.00217909f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.19
cc_19 VNB N_X_c_234_n 0.00204615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.0337654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_297_n 0.00475331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_298_n 0.00404131f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_23 VNB N_VGND_c_299_n 0.0120207f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.85
cc_24 VNB N_VGND_c_300_n 0.00474766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_301_n 0.0164986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_302_n 0.0175222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_303_n 0.0158977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_304_n 0.0052624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_305_n 0.0048778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_306_n 0.161822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_A_M1006_g 0.0229606f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_32 VPB A 0.00221579f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_33 VPB N_A_c_57_n 0.00536987f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_34 VPB N_A_27_47#_M1002_g 0.0198993f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_35 VPB N_A_27_47#_M1007_g 0.0197727f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_36 VPB N_A_27_47#_M1008_g 0.0197632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_M1009_g 0.0240996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_98_n 0.00904608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_106_n 0.0313553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_107_n 0.00175845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_108_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_188_n 0.0048939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_189_n 0.00398868f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_44 VPB N_VPWR_c_190_n 0.0121228f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.85
cc_45 VPB N_VPWR_c_191_n 0.00477568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_192_n 0.0172252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_193_n 0.0158982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_194_n 0.0160896f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_195_n 0.00593688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_196_n 0.00487698f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_187_n 0.0450154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB X 0.0058073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_X_c_237_n 0.0130264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 N_A_M1006_g N_A_27_47#_M1002_g 0.0228625f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_55 N_A_M1003_g N_A_27_47#_M1000_g 0.0183348f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_56 A N_A_27_47#_M1000_g 0.0050309f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_c_57_n N_A_27_47#_M1000_g 0.00287228f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_M1003_g N_A_27_47#_c_98_n 0.0101619f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_59 N_A_M1006_g N_A_27_47#_c_98_n 0.0059274f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_60 A N_A_27_47#_c_98_n 0.0429918f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_61 N_A_c_57_n N_A_27_47#_c_98_n 0.00797697f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_M1006_g N_A_27_47#_c_117_n 0.0139831f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_63 A N_A_27_47#_c_117_n 0.0251553f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_64 N_A_c_57_n N_A_27_47#_c_117_n 5.45329e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_A_27_47#_c_107_n 9.07197e-19 $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_66 A N_A_27_47#_c_107_n 0.00600199f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_67 A N_A_27_47#_c_122_n 0.0143279f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_68 A N_A_27_47#_c_100_n 0.00251756f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_69 N_A_c_57_n N_A_27_47#_c_100_n 0.0154138f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_M1006_g N_VPWR_c_188_n 0.00315548f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_M1006_g N_VPWR_c_192_n 0.00585385f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_M1006_g N_VPWR_c_187_n 0.0115761f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_X_c_231_n 7.63641e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_M1003_g N_X_c_233_n 2.1267e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_75 A N_X_c_233_n 0.00990658f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_VGND_c_297_n 0.00318753f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_77 A N_VGND_c_297_n 0.0152693f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_78 N_A_c_57_n N_VGND_c_297_n 3.07485e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_M1003_g N_VGND_c_301_n 0.00466641f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_80 A N_VGND_c_301_n 0.00176987f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_M1003_g N_VGND_c_306_n 0.00775648f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_82 A N_VGND_c_306_n 0.00378105f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_117_n N_VPWR_M1006_d 0.00585437f $X=0.945 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_27_47#_M1002_g N_VPWR_c_188_n 0.00174199f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_85 N_A_27_47#_c_117_n N_VPWR_c_188_n 0.0175734f $X=0.945 $Y=1.58 $X2=0 $Y2=0
cc_86 N_A_27_47#_M1007_g N_VPWR_c_189_n 0.00158973f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_87 N_A_27_47#_M1008_g N_VPWR_c_189_n 0.00161779f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_88 N_A_27_47#_M1009_g N_VPWR_c_191_n 0.00377306f $X=2.245 $Y=1.985 $X2=0
+ $Y2=0
cc_89 N_A_27_47#_c_106_n N_VPWR_c_192_n 0.0199493f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_90 N_A_27_47#_M1002_g N_VPWR_c_193_n 0.00585385f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_91 N_A_27_47#_M1007_g N_VPWR_c_193_n 0.00436487f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_M1008_g N_VPWR_c_194_n 0.00436487f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_M1009_g N_VPWR_c_194_n 0.00585385f $X=2.245 $Y=1.985 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_M1006_s N_VPWR_c_187_n 0.00230776f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_M1002_g N_VPWR_c_187_n 0.0106953f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_27_47#_M1007_g N_VPWR_c_187_n 0.00587239f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_M1008_g N_VPWR_c_187_n 0.00581455f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_M1009_g N_VPWR_c_187_n 0.0115843f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_106_n N_VPWR_c_187_n 0.0118616f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_117_n N_X_M1002_d 0.00266776f $X=0.945 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A_27_47#_M1000_g N_X_c_231_n 0.00655439f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A_27_47#_M1001_g N_X_c_231_n 0.00115565f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A_27_47#_M1001_g N_X_c_232_n 0.0122792f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_27_47#_M1004_g N_X_c_232_n 0.0122792f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_147_p N_X_c_232_n 0.054594f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_100_n N_X_c_232_n 0.0023301f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_107 N_A_27_47#_M1000_g N_X_c_233_n 0.00456754f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_122_n N_X_c_233_n 0.00901782f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_147_p N_X_c_233_n 0.0150434f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_100_n N_X_c_233_n 0.00240878f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_111 N_A_27_47#_M1007_g N_X_c_252_n 0.0134417f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_27_47#_M1008_g N_X_c_252_n 0.0120866f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_147_p N_X_c_252_n 0.0132831f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_100_n N_X_c_252_n 0.00167579f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_117_n N_X_c_256_n 0.00243987f $X=0.945 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_147_p N_X_c_256_n 0.00470582f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_100_n N_X_c_256_n 0.0017973f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_118 N_A_27_47#_M1004_g N_X_c_234_n 0.00114296f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A_27_47#_M1005_g N_X_c_234_n 0.00216977f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1008_g X 6.2445e-19 $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_27_47#_M1004_g X 6.0408e-19 $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1009_g X 0.00525161f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_27_47#_M1005_g X 0.018959f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_147_p X 0.0136122f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_100_n X 0.0174538f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_126 N_A_27_47#_M1008_g N_X_c_237_n 0.00226561f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1009_g N_X_c_237_n 0.0153884f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_147_p N_X_c_237_n 0.0128752f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_100_n N_X_c_237_n 0.00233619f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_130 N_A_27_47#_M1000_g N_VGND_c_297_n 0.00157173f $X=0.96 $Y=0.445 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_M1001_g N_VGND_c_298_n 0.00166998f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_M1004_g N_VGND_c_298_n 0.00159632f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_M1005_g N_VGND_c_300_n 0.00341661f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_99_n N_VGND_c_301_n 0.0186529f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_135 N_A_27_47#_M1000_g N_VGND_c_302_n 0.0055185f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A_27_47#_M1001_g N_VGND_c_302_n 0.00439206f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_M1004_g N_VGND_c_303_n 0.00439206f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_M1005_g N_VGND_c_303_n 0.00439206f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_M1003_s N_VGND_c_306_n 0.00262044f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_M1000_g N_VGND_c_306_n 0.00995296f $X=0.96 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_M1001_g N_VGND_c_306_n 0.00590932f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_M1004_g N_VGND_c_306_n 0.00592186f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_M1005_g N_VGND_c_306_n 0.0068734f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_99_n N_VGND_c_306_n 0.0113402f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_145 N_VPWR_c_187_n N_X_M1002_d 0.0028199f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_146 N_VPWR_c_187_n N_X_M1008_d 0.00246537f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_147 N_VPWR_c_193_n N_X_c_273_n 0.0148724f $X=1.475 $Y=2.72 $X2=0 $Y2=0
cc_148 N_VPWR_c_187_n N_X_c_273_n 0.00991615f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_149 N_VPWR_M1007_s N_X_c_252_n 0.00468845f $X=1.46 $Y=1.485 $X2=0 $Y2=0
cc_150 N_VPWR_c_189_n N_X_c_252_n 0.0129597f $X=1.6 $Y=2.34 $X2=0 $Y2=0
cc_151 N_VPWR_c_193_n N_X_c_252_n 0.00219745f $X=1.475 $Y=2.72 $X2=0 $Y2=0
cc_152 N_VPWR_c_194_n N_X_c_252_n 0.00223722f $X=2.335 $Y=2.72 $X2=0 $Y2=0
cc_153 N_VPWR_c_187_n N_X_c_252_n 0.00851676f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_c_194_n N_X_c_280_n 0.0149375f $X=2.335 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_187_n N_X_c_280_n 0.00993603f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_M1009_s N_X_c_237_n 0.00329253f $X=2.32 $Y=1.485 $X2=0 $Y2=0
cc_157 N_VPWR_c_191_n N_X_c_237_n 0.0188647f $X=2.46 $Y=1.93 $X2=0 $Y2=0
cc_158 N_X_c_232_n N_VGND_c_298_n 0.0162872f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_159 X N_VGND_c_299_n 6.74578e-19 $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_160 X N_VGND_c_300_n 0.0201078f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_161 N_X_c_231_n N_VGND_c_302_n 0.010662f $X=1.175 $Y=0.51 $X2=0 $Y2=0
cc_162 N_X_c_232_n N_VGND_c_302_n 0.00224999f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_163 N_X_c_232_n N_VGND_c_303_n 0.00461204f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_164 N_X_c_234_n N_VGND_c_303_n 0.0092385f $X=2.035 $Y=0.51 $X2=0 $Y2=0
cc_165 N_X_M1000_d N_VGND_c_306_n 0.0023797f $X=1.035 $Y=0.235 $X2=0 $Y2=0
cc_166 N_X_M1004_d N_VGND_c_306_n 0.00244557f $X=1.895 $Y=0.235 $X2=0 $Y2=0
cc_167 N_X_c_231_n N_VGND_c_306_n 0.0105577f $X=1.175 $Y=0.51 $X2=0 $Y2=0
cc_168 N_X_c_232_n N_VGND_c_306_n 0.0121304f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_169 N_X_c_234_n N_VGND_c_306_n 0.00930021f $X=2.035 $Y=0.51 $X2=0 $Y2=0
cc_170 X N_VGND_c_306_n 0.00223695f $X=2.445 $Y=0.765 $X2=0 $Y2=0

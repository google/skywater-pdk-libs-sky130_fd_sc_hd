* File: sky130_fd_sc_hd__dlclkp_1.pxi.spice
* Created: Thu Aug 27 14:16:18 2020
* 
x_PM_SKY130_FD_SC_HD__DLCLKP_1%CLK N_CLK_c_153_n N_CLK_c_142_n N_CLK_M1019_g
+ N_CLK_c_154_n N_CLK_M1008_g N_CLK_M1016_g N_CLK_M1013_g N_CLK_c_144_n
+ N_CLK_c_156_n CLK N_CLK_c_145_n N_CLK_c_146_n N_CLK_c_147_n N_CLK_c_148_n
+ N_CLK_c_149_n N_CLK_c_150_n N_CLK_c_151_n N_CLK_c_152_n
+ PM_SKY130_FD_SC_HD__DLCLKP_1%CLK
x_PM_SKY130_FD_SC_HD__DLCLKP_1%GATE N_GATE_c_277_n N_GATE_M1015_g N_GATE_c_278_n
+ N_GATE_M1017_g N_GATE_c_282_n GATE GATE GATE PM_SKY130_FD_SC_HD__DLCLKP_1%GATE
x_PM_SKY130_FD_SC_HD__DLCLKP_1%A_193_47# N_A_193_47#_M1010_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1005_g N_A_193_47#_M1014_g N_A_193_47#_c_322_n
+ N_A_193_47#_c_329_n N_A_193_47#_c_323_n N_A_193_47#_c_331_n
+ N_A_193_47#_c_324_n N_A_193_47#_c_325_n N_A_193_47#_c_332_n
+ N_A_193_47#_c_326_n PM_SKY130_FD_SC_HD__DLCLKP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__DLCLKP_1%A_27_47# N_A_27_47#_M1019_s N_A_27_47#_M1008_s
+ N_A_27_47#_c_415_n N_A_27_47#_M1010_g N_A_27_47#_c_416_n N_A_27_47#_M1000_g
+ N_A_27_47#_c_417_n N_A_27_47#_c_418_n N_A_27_47#_c_419_n N_A_27_47#_c_420_n
+ N_A_27_47#_M1009_g N_A_27_47#_c_422_n N_A_27_47#_c_423_n N_A_27_47#_M1002_g
+ N_A_27_47#_c_424_n N_A_27_47#_c_537_p N_A_27_47#_c_425_n N_A_27_47#_c_426_n
+ N_A_27_47#_c_434_n N_A_27_47#_c_435_n N_A_27_47#_c_436_n N_A_27_47#_c_427_n
+ N_A_27_47#_c_428_n N_A_27_47#_c_429_n PM_SKY130_FD_SC_HD__DLCLKP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__DLCLKP_1%A_642_307# N_A_642_307#_M1011_d
+ N_A_642_307#_M1018_s N_A_642_307#_M1003_g N_A_642_307#_M1004_g
+ N_A_642_307#_c_550_n N_A_642_307#_M1007_g N_A_642_307#_c_551_n
+ N_A_642_307#_c_552_n N_A_642_307#_M1001_g N_A_642_307#_c_560_n
+ N_A_642_307#_c_634_p N_A_642_307#_c_561_n N_A_642_307#_c_562_n
+ N_A_642_307#_c_553_n N_A_642_307#_c_554_n N_A_642_307#_c_555_n
+ N_A_642_307#_c_563_n PM_SKY130_FD_SC_HD__DLCLKP_1%A_642_307#
x_PM_SKY130_FD_SC_HD__DLCLKP_1%A_476_413# N_A_476_413#_M1009_d
+ N_A_476_413#_M1005_d N_A_476_413#_M1011_g N_A_476_413#_M1018_g
+ N_A_476_413#_c_678_n N_A_476_413#_c_671_n N_A_476_413#_c_666_n
+ N_A_476_413#_c_658_n N_A_476_413#_c_659_n N_A_476_413#_c_660_n
+ N_A_476_413#_c_661_n N_A_476_413#_c_662_n N_A_476_413#_c_663_n
+ N_A_476_413#_c_664_n PM_SKY130_FD_SC_HD__DLCLKP_1%A_476_413#
x_PM_SKY130_FD_SC_HD__DLCLKP_1%A_957_369# N_A_957_369#_M1001_s
+ N_A_957_369#_M1007_d N_A_957_369#_M1006_g N_A_957_369#_M1012_g
+ N_A_957_369#_c_747_n N_A_957_369#_c_760_n N_A_957_369#_c_748_n
+ N_A_957_369#_c_749_n N_A_957_369#_c_755_n N_A_957_369#_c_756_n
+ N_A_957_369#_c_750_n N_A_957_369#_c_751_n N_A_957_369#_c_758_n
+ N_A_957_369#_c_781_n N_A_957_369#_c_752_n N_A_957_369#_c_753_n
+ PM_SKY130_FD_SC_HD__DLCLKP_1%A_957_369#
x_PM_SKY130_FD_SC_HD__DLCLKP_1%VPWR N_VPWR_M1008_d N_VPWR_M1015_s N_VPWR_M1003_d
+ N_VPWR_M1018_d N_VPWR_M1013_d N_VPWR_c_827_n N_VPWR_c_828_n N_VPWR_c_829_n
+ N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_832_n VPWR N_VPWR_c_833_n
+ N_VPWR_c_834_n N_VPWR_c_835_n N_VPWR_c_836_n N_VPWR_c_837_n N_VPWR_c_826_n
+ N_VPWR_c_839_n N_VPWR_c_840_n N_VPWR_c_841_n N_VPWR_c_842_n N_VPWR_c_843_n
+ PM_SKY130_FD_SC_HD__DLCLKP_1%VPWR
x_PM_SKY130_FD_SC_HD__DLCLKP_1%GCLK N_GCLK_M1006_d N_GCLK_M1012_d N_GCLK_c_924_n
+ N_GCLK_c_922_n GCLK GCLK GCLK N_GCLK_c_926_n N_GCLK_c_923_n
+ PM_SKY130_FD_SC_HD__DLCLKP_1%GCLK
x_PM_SKY130_FD_SC_HD__DLCLKP_1%VGND N_VGND_M1019_d N_VGND_M1017_s N_VGND_M1004_d
+ N_VGND_M1016_d N_VGND_c_939_n N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n
+ VGND N_VGND_c_943_n N_VGND_c_944_n N_VGND_c_945_n N_VGND_c_946_n
+ N_VGND_c_947_n N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n
+ N_VGND_c_952_n PM_SKY130_FD_SC_HD__DLCLKP_1%VGND
cc_1 VNB N_CLK_c_142_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_M1016_g 0.0346763f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=0.445
cc_3 VNB N_CLK_c_144_n 0.0236526f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_4 VNB N_CLK_c_145_n 0.0512113f $X=-0.19 $Y=-0.24 $X2=5.15 $Y2=1.19
cc_5 VNB N_CLK_c_146_n 0.00982131f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_6 VNB N_CLK_c_147_n 0.0103308f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_7 VNB N_CLK_c_148_n 0.00277658f $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_8 VNB N_CLK_c_149_n 7.80019e-19 $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_9 VNB N_CLK_c_150_n 0.0198903f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_10 VNB N_CLK_c_151_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_11 VNB N_CLK_c_152_n 0.021223f $X=-0.19 $Y=-0.24 $X2=5.325 $Y2=1.27
cc_12 VNB N_GATE_c_277_n 0.0280986f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.88
cc_13 VNB N_GATE_c_278_n 0.0154714f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_14 VNB GATE 0.00988506f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=1.105
cc_15 VNB N_A_193_47#_M1014_g 0.0212024f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=0.445
cc_16 VNB N_A_193_47#_c_322_n 0.0159946f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=2.165
cc_17 VNB N_A_193_47#_c_323_n 0.00463956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_193_47#_c_324_n 0.00120332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_193_47#_c_325_n 0.0053269f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_20 VNB N_A_193_47#_c_326_n 0.0351829f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_21 VNB N_A_27_47#_c_415_n 0.014637f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_22 VNB N_A_27_47#_c_416_n 0.0125115f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=1.105
cc_23 VNB N_A_27_47#_c_417_n 0.0317905f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=2.165
cc_24 VNB N_A_27_47#_c_418_n 0.0267961f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_25 VNB N_A_27_47#_c_419_n 0.0761503f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_420_n 0.00988887f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_27 VNB N_A_27_47#_M1009_g 0.035085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_28 VNB N_A_27_47#_c_422_n 0.018035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_423_n 0.00453564f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_30 VNB N_A_27_47#_c_424_n 0.0052727f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_31 VNB N_A_27_47#_c_425_n 0.00177906f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_32 VNB N_A_27_47#_c_426_n 0.00553431f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_33 VNB N_A_27_47#_c_427_n 7.70731e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_428_n 0.00438392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_429_n 0.0241763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_642_307#_M1004_g 0.0460839f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=0.445
cc_37 VNB N_A_642_307#_c_550_n 0.0417074f $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=1.435
cc_38 VNB N_A_642_307#_c_551_n 0.027812f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_39 VNB N_A_642_307#_c_552_n 0.0174432f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_40 VNB N_A_642_307#_c_553_n 0.0041536f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_41 VNB N_A_642_307#_c_554_n 0.00390883f $X=-0.19 $Y=-0.24 $X2=5.325 $Y2=1.27
cc_42 VNB N_A_642_307#_c_555_n 0.00449335f $X=-0.19 $Y=-0.24 $X2=5.38 $Y2=1.435
cc_43 VNB N_A_476_413#_c_658_n 0.0037655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_476_413#_c_659_n 0.00267318f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_45 VNB N_A_476_413#_c_660_n 0.00317602f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_46 VNB N_A_476_413#_c_661_n 0.00694965f $X=-0.19 $Y=-0.24 $X2=0.38 $Y2=1.19
cc_47 VNB N_A_476_413#_c_662_n 0.026225f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_48 VNB N_A_476_413#_c_663_n 0.00436303f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_49 VNB N_A_476_413#_c_664_n 0.020237f $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_50 VNB N_A_957_369#_c_747_n 7.57877e-19 $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=1.435
cc_51 VNB N_A_957_369#_c_748_n 0.0122309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_957_369#_c_749_n 0.00325886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_53 VNB N_A_957_369#_c_750_n 0.00206875f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_54 VNB N_A_957_369#_c_751_n 0.0227277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_957_369#_c_752_n 6.10609e-19 $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_56 VNB N_A_957_369#_c_753_n 0.0193012f $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_57 VNB N_VPWR_c_826_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_GCLK_c_922_n 0.0304805f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_59 VNB N_GCLK_c_923_n 0.013586f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_60 VNB N_VGND_c_939_n 4.1623e-19 $X=-0.19 $Y=-0.24 $X2=5.495 $Y2=1.435
cc_61 VNB N_VGND_c_940_n 0.0107856f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_62 VNB N_VGND_c_941_n 0.00239192f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_63 VNB N_VGND_c_942_n 0.00472864f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_64 VNB N_VGND_c_943_n 0.0151256f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_65 VNB N_VGND_c_944_n 0.0155996f $X=-0.19 $Y=-0.24 $X2=5.295 $Y2=1.19
cc_66 VNB N_VGND_c_945_n 0.0570522f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_67 VNB N_VGND_c_946_n 0.042241f $X=-0.19 $Y=-0.24 $X2=5.325 $Y2=1.27
cc_68 VNB N_VGND_c_947_n 0.0184163f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_948_n 0.325204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_949_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_950_n 0.00439458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_951_n 0.00357019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_952_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VPB N_CLK_c_153_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_75 VPB N_CLK_c_154_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_76 VPB N_CLK_M1013_g 0.0379102f $X=-0.19 $Y=1.305 $X2=5.495 $Y2=2.165
cc_77 VPB N_CLK_c_156_n 0.0238508f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_78 VPB N_CLK_c_147_n 0.0156114f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_79 VPB N_CLK_c_148_n 3.91477e-19 $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_80 VPB N_CLK_c_149_n 0.00260386f $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_81 VPB N_CLK_c_150_n 0.0109496f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_82 VPB N_CLK_c_152_n 0.0175687f $X=-0.19 $Y=1.305 $X2=5.325 $Y2=1.27
cc_83 VPB N_GATE_c_277_n 0.0325214f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.88
cc_84 VPB N_GATE_M1015_g 0.0227685f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_85 VPB N_GATE_c_282_n 0.00990655f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_86 VPB GATE 0.0016051f $X=-0.19 $Y=1.305 $X2=5.495 $Y2=1.105
cc_87 VPB N_A_193_47#_M1005_g 0.0218483f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_88 VPB N_A_193_47#_c_322_n 0.0125206f $X=-0.19 $Y=1.305 $X2=5.495 $Y2=2.165
cc_89 VPB N_A_193_47#_c_329_n 0.0136055f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_90 VPB N_A_193_47#_c_323_n 0.00348173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_193_47#_c_331_n 0.0383239f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_92 VPB N_A_193_47#_c_332_n 0.00725072f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_27_47#_M1000_g 0.0415337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_47#_c_422_n 0.0178202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_47#_c_423_n 0.00326288f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_96 VPB N_A_27_47#_M1002_g 0.0482884f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.19
cc_97 VPB N_A_27_47#_c_434_n 0.00121249f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_98 VPB N_A_27_47#_c_435_n 0.00647616f $X=-0.19 $Y=1.305 $X2=5.325 $Y2=1.27
cc_99 VPB N_A_27_47#_c_436_n 0.00345702f $X=-0.19 $Y=1.305 $X2=5.38 $Y2=1.435
cc_100 VPB N_A_27_47#_c_427_n 0.00152564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_27_47#_c_429_n 0.0108287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_642_307#_M1003_g 0.023974f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_103 VPB N_A_642_307#_M1004_g 0.0152291f $X=-0.19 $Y=1.305 $X2=5.495 $Y2=0.445
cc_104 VPB N_A_642_307#_c_550_n 0.00479778f $X=-0.19 $Y=1.305 $X2=5.495
+ $Y2=1.435
cc_105 VPB N_A_642_307#_M1007_g 0.0431417f $X=-0.19 $Y=1.305 $X2=5.495 $Y2=2.165
cc_106 VPB N_A_642_307#_c_560_n 0.00440075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_642_307#_c_561_n 0.0015694f $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_108 VPB N_A_642_307#_c_562_n 0.00198847f $X=-0.19 $Y=1.305 $X2=0.242
+ $Y2=1.235
cc_109 VPB N_A_642_307#_c_563_n 0.0477574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_476_413#_M1018_g 0.023217f $X=-0.19 $Y=1.305 $X2=5.495 $Y2=0.445
cc_111 VPB N_A_476_413#_c_666_n 0.0086435f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_112 VPB N_A_476_413#_c_658_n 0.00294899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_476_413#_c_659_n 2.95714e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_114 VPB N_A_476_413#_c_661_n 0.00225196f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.19
cc_115 VPB N_A_476_413#_c_662_n 0.00644727f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_116 VPB N_A_957_369#_M1012_g 0.0217242f $X=-0.19 $Y=1.305 $X2=5.495 $Y2=0.445
cc_117 VPB N_A_957_369#_c_755_n 0.00314873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_957_369#_c_756_n 0.00629769f $X=-0.19 $Y=1.305 $X2=0.305
+ $Y2=1.665
cc_119 VPB N_A_957_369#_c_751_n 0.00478128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_957_369#_c_758_n 0.00121786f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.19
cc_121 VPB N_VPWR_c_827_n 0.00106176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_828_n 0.00540398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_829_n 0.00915038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_830_n 0.0175728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_831_n 0.00477366f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_126 VPB N_VPWR_c_832_n 0.0029422f $X=-0.19 $Y=1.305 $X2=5.295 $Y2=1.19
cc_127 VPB N_VPWR_c_833_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_128 VPB N_VPWR_c_834_n 0.0153955f $X=-0.19 $Y=1.305 $X2=5.325 $Y2=1.27
cc_129 VPB N_VPWR_c_835_n 0.0400543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_836_n 0.0278771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_837_n 0.0152176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_826_n 0.0587227f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_839_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_840_n 0.00557046f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_841_n 0.00574408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_842_n 0.00545601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_843_n 0.00549285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_GCLK_c_924_n 0.00502818f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_139 VPB N_GCLK_c_922_n 0.00893034f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_140 VPB N_GCLK_c_926_n 0.0318655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 N_CLK_c_145_n N_GATE_c_277_n 0.0167433f $X=5.15 $Y=1.19 $X2=-0.19
+ $Y2=-0.24
cc_142 N_CLK_c_145_n N_GATE_c_282_n 0.0157888f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_143 N_CLK_c_145_n GATE 0.024007f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_144 N_CLK_c_145_n N_A_193_47#_c_322_n 0.0314284f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_145 N_CLK_c_145_n N_A_193_47#_c_329_n 0.0143972f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_146 N_CLK_c_145_n N_A_193_47#_c_323_n 0.0226377f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_147 N_CLK_c_145_n N_A_193_47#_c_331_n 0.00405475f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_148 N_CLK_c_145_n N_A_193_47#_c_325_n 0.0254803f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_149 N_CLK_c_145_n N_A_193_47#_c_326_n 0.00789047f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_150 N_CLK_c_142_n N_A_27_47#_c_415_n 0.0101063f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_151 N_CLK_c_151_n N_A_27_47#_c_416_n 0.00406423f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_152 N_CLK_c_156_n N_A_27_47#_M1000_g 0.0256048f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_153 N_CLK_c_150_n N_A_27_47#_M1000_g 0.00439406f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_154 N_CLK_c_145_n N_A_27_47#_c_417_n 0.00590074f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_155 N_CLK_c_145_n N_A_27_47#_M1009_g 0.00145143f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_156 N_CLK_c_145_n N_A_27_47#_c_422_n 0.0179291f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_157 N_CLK_c_145_n N_A_27_47#_c_423_n 2.71279e-19 $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_158 N_CLK_c_144_n N_A_27_47#_c_424_n 0.0101063f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_159 N_CLK_c_142_n N_A_27_47#_c_425_n 0.00770412f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_160 N_CLK_c_144_n N_A_27_47#_c_425_n 0.00553647f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_161 N_CLK_c_145_n N_A_27_47#_c_425_n 0.00817564f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_162 N_CLK_c_146_n N_A_27_47#_c_425_n 0.00120578f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_163 N_CLK_c_144_n N_A_27_47#_c_426_n 0.0057713f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_164 N_CLK_c_146_n N_A_27_47#_c_426_n 0.00161409f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_165 N_CLK_c_147_n N_A_27_47#_c_426_n 0.0105869f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_166 N_CLK_c_150_n N_A_27_47#_c_426_n 3.38487e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_167 N_CLK_c_154_n N_A_27_47#_c_434_n 0.0107161f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_168 N_CLK_c_156_n N_A_27_47#_c_434_n 0.00220936f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_169 N_CLK_c_145_n N_A_27_47#_c_434_n 0.0067661f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_170 N_CLK_c_146_n N_A_27_47#_c_434_n 0.00108512f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_171 N_CLK_c_153_n N_A_27_47#_c_435_n 8.6683e-19 $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_172 N_CLK_c_156_n N_A_27_47#_c_435_n 0.00435948f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_173 N_CLK_c_154_n N_A_27_47#_c_436_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_174 N_CLK_c_156_n N_A_27_47#_c_436_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_175 N_CLK_c_146_n N_A_27_47#_c_436_n 0.00126485f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_176 N_CLK_c_147_n N_A_27_47#_c_436_n 0.0133866f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_177 N_CLK_c_150_n N_A_27_47#_c_436_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_178 N_CLK_c_145_n N_A_27_47#_c_427_n 0.0293907f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_179 N_CLK_c_146_n N_A_27_47#_c_427_n 0.00217711f $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_180 N_CLK_c_150_n N_A_27_47#_c_427_n 0.00320691f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_181 N_CLK_c_144_n N_A_27_47#_c_428_n 0.00227671f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_182 N_CLK_c_147_n N_A_27_47#_c_428_n 0.028836f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_183 N_CLK_c_151_n N_A_27_47#_c_428_n 0.00146736f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_184 N_CLK_c_145_n N_A_27_47#_c_429_n 0.0137802f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_185 N_CLK_c_146_n N_A_27_47#_c_429_n 4.33321e-19 $X=0.38 $Y=1.19 $X2=0 $Y2=0
cc_186 N_CLK_c_147_n N_A_27_47#_c_429_n 9.54145e-19 $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_187 N_CLK_c_150_n N_A_27_47#_c_429_n 0.0183177f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_188 N_CLK_M1016_g N_A_642_307#_c_550_n 0.00423242f $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_189 N_CLK_c_145_n N_A_642_307#_c_550_n 0.00512296f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_190 N_CLK_c_148_n N_A_642_307#_c_550_n 0.00133445f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_191 N_CLK_c_149_n N_A_642_307#_c_550_n 9.11216e-19 $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_192 N_CLK_c_152_n N_A_642_307#_c_550_n 0.00720036f $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_193 N_CLK_M1013_g N_A_642_307#_M1007_g 0.0172818f $X=5.495 $Y=2.165 $X2=0
+ $Y2=0
cc_194 N_CLK_c_149_n N_A_642_307#_M1007_g 4.07079e-19 $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_195 N_CLK_c_152_n N_A_642_307#_M1007_g 0.00292858f $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_196 N_CLK_c_145_n N_A_642_307#_c_551_n 0.0029373f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_197 N_CLK_c_152_n N_A_642_307#_c_551_n 0.00120126f $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_198 N_CLK_M1016_g N_A_642_307#_c_552_n 0.0480446f $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_199 N_CLK_c_145_n N_A_642_307#_c_560_n 0.00312808f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_200 N_CLK_c_149_n N_A_642_307#_c_561_n 0.00355136f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_201 N_CLK_c_152_n N_A_642_307#_c_561_n 4.24609e-19 $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_202 N_CLK_c_145_n N_A_642_307#_c_562_n 0.00829457f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_203 N_CLK_c_145_n N_A_642_307#_c_553_n 8.5633e-19 $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_204 N_CLK_M1016_g N_A_642_307#_c_554_n 4.56256e-19 $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_CLK_c_145_n N_A_642_307#_c_554_n 0.0505805f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_206 N_CLK_c_148_n N_A_642_307#_c_554_n 0.00263102f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_207 N_CLK_c_149_n N_A_642_307#_c_554_n 0.00449696f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_208 N_CLK_c_152_n N_A_642_307#_c_554_n 7.19579e-19 $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_209 N_CLK_c_145_n N_A_476_413#_c_671_n 0.00754428f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_210 N_CLK_c_145_n N_A_476_413#_c_658_n 0.0136361f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_211 N_CLK_c_145_n N_A_476_413#_c_659_n 0.0133794f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_212 N_CLK_c_145_n N_A_476_413#_c_661_n 0.0268066f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_213 N_CLK_c_145_n N_A_476_413#_c_662_n 0.00739349f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_214 N_CLK_c_145_n N_A_476_413#_c_663_n 0.0150785f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_215 N_CLK_c_152_n N_A_957_369#_M1012_g 0.0322481f $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_216 N_CLK_M1013_g N_A_957_369#_c_760_n 0.0109865f $X=5.495 $Y=2.165 $X2=0
+ $Y2=0
cc_217 N_CLK_M1016_g N_A_957_369#_c_748_n 0.0137901f $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_CLK_c_148_n N_A_957_369#_c_748_n 0.00873139f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_219 N_CLK_c_149_n N_A_957_369#_c_748_n 0.0206178f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_220 N_CLK_c_152_n N_A_957_369#_c_748_n 0.00153685f $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_221 N_CLK_c_145_n N_A_957_369#_c_749_n 0.0110704f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_222 N_CLK_c_148_n N_A_957_369#_c_749_n 2.81942e-19 $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_223 N_CLK_M1013_g N_A_957_369#_c_755_n 0.0154639f $X=5.495 $Y=2.165 $X2=0
+ $Y2=0
cc_224 N_CLK_c_148_n N_A_957_369#_c_755_n 5.69151e-19 $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_225 N_CLK_c_149_n N_A_957_369#_c_755_n 0.00778699f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_226 N_CLK_c_152_n N_A_957_369#_c_755_n 5.3256e-19 $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_227 N_CLK_c_145_n N_A_957_369#_c_756_n 0.00573426f $X=5.15 $Y=1.19 $X2=0
+ $Y2=0
cc_228 N_CLK_c_148_n N_A_957_369#_c_756_n 0.00268666f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_229 N_CLK_c_149_n N_A_957_369#_c_756_n 0.00704395f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_230 N_CLK_c_152_n N_A_957_369#_c_756_n 0.00106765f $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_231 N_CLK_M1016_g N_A_957_369#_c_750_n 0.0039753f $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_232 N_CLK_c_148_n N_A_957_369#_c_750_n 0.00245074f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_233 N_CLK_c_149_n N_A_957_369#_c_750_n 0.0179568f $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_234 N_CLK_M1016_g N_A_957_369#_c_751_n 0.0203801f $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_235 N_CLK_c_149_n N_A_957_369#_c_751_n 2.4238e-19 $X=5.295 $Y=1.19 $X2=0
+ $Y2=0
cc_236 N_CLK_M1013_g N_A_957_369#_c_758_n 0.0039753f $X=5.495 $Y=2.165 $X2=0
+ $Y2=0
cc_237 N_CLK_M1016_g N_A_957_369#_c_781_n 0.00211691f $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_238 N_CLK_c_145_n N_A_957_369#_c_781_n 0.0033383f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_239 N_CLK_c_152_n N_A_957_369#_c_752_n 0.0039753f $X=5.325 $Y=1.27 $X2=0
+ $Y2=0
cc_240 N_CLK_M1016_g N_A_957_369#_c_753_n 0.021487f $X=5.495 $Y=0.445 $X2=0
+ $Y2=0
cc_241 N_CLK_c_154_n N_VPWR_c_827_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_M1013_g N_VPWR_c_832_n 0.00324046f $X=5.495 $Y=2.165 $X2=0 $Y2=0
cc_243 N_CLK_c_154_n N_VPWR_c_833_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_244 N_CLK_M1013_g N_VPWR_c_836_n 0.00583607f $X=5.495 $Y=2.165 $X2=0 $Y2=0
cc_245 N_CLK_c_154_n N_VPWR_c_826_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_246 N_CLK_M1013_g N_VPWR_c_826_n 0.00691647f $X=5.495 $Y=2.165 $X2=0 $Y2=0
cc_247 N_CLK_c_142_n N_VGND_c_939_n 0.0082568f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_248 N_CLK_c_145_n N_VGND_c_940_n 0.0107999f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_249 N_CLK_c_145_n N_VGND_c_941_n 0.00164197f $X=5.15 $Y=1.19 $X2=0 $Y2=0
cc_250 N_CLK_M1016_g N_VGND_c_942_n 0.00518162f $X=5.495 $Y=0.445 $X2=0 $Y2=0
cc_251 N_CLK_c_142_n N_VGND_c_943_n 0.00337001f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_252 N_CLK_c_144_n N_VGND_c_943_n 4.4475e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_253 N_CLK_M1016_g N_VGND_c_946_n 0.00585385f $X=5.495 $Y=0.445 $X2=0 $Y2=0
cc_254 N_CLK_c_142_n N_VGND_c_948_n 0.00485988f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_255 N_CLK_M1016_g N_VGND_c_948_n 0.00617518f $X=5.495 $Y=0.445 $X2=0 $Y2=0
cc_256 N_GATE_M1015_g N_A_193_47#_M1005_g 0.020041f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_257 N_GATE_c_277_n N_A_193_47#_c_322_n 0.00825783f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_258 N_GATE_M1015_g N_A_193_47#_c_322_n 0.00442795f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_259 N_GATE_c_278_n N_A_193_47#_c_322_n 0.00417595f $X=1.905 $Y=1.09 $X2=0
+ $Y2=0
cc_260 N_GATE_c_282_n N_A_193_47#_c_322_n 0.0166772f $X=1.985 $Y=1.56 $X2=0
+ $Y2=0
cc_261 N_GATE_c_277_n N_A_193_47#_c_329_n 0.00267752f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_262 N_GATE_M1015_g N_A_193_47#_c_329_n 0.0136889f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_263 N_GATE_c_282_n N_A_193_47#_c_329_n 0.045043f $X=1.985 $Y=1.56 $X2=0 $Y2=0
cc_264 N_GATE_c_277_n N_A_193_47#_c_323_n 0.00155015f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_265 N_GATE_c_282_n N_A_193_47#_c_323_n 0.0183467f $X=1.985 $Y=1.56 $X2=0
+ $Y2=0
cc_266 GATE N_A_193_47#_c_323_n 0.0276354f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_267 N_GATE_c_277_n N_A_193_47#_c_331_n 0.020041f $X=1.83 $Y=1.685 $X2=0 $Y2=0
cc_268 N_GATE_c_282_n N_A_193_47#_c_331_n 8.60298e-19 $X=1.985 $Y=1.56 $X2=0
+ $Y2=0
cc_269 GATE N_A_193_47#_c_324_n 0.0116864f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_270 N_GATE_M1015_g N_A_193_47#_c_332_n 0.00359119f $X=1.83 $Y=2.165 $X2=0
+ $Y2=0
cc_271 N_GATE_c_278_n N_A_27_47#_c_418_n 0.00641991f $X=1.905 $Y=1.09 $X2=0
+ $Y2=0
cc_272 N_GATE_c_278_n N_A_27_47#_c_419_n 0.0104164f $X=1.905 $Y=1.09 $X2=0 $Y2=0
cc_273 GATE N_A_27_47#_c_419_n 0.00459101f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_274 N_GATE_c_277_n N_A_27_47#_M1009_g 0.00300861f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_275 N_GATE_c_278_n N_A_27_47#_M1009_g 0.0178241f $X=1.905 $Y=1.09 $X2=0 $Y2=0
cc_276 GATE N_A_27_47#_M1009_g 0.012688f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_277 N_GATE_c_277_n N_A_27_47#_c_429_n 0.00329527f $X=1.83 $Y=1.685 $X2=0
+ $Y2=0
cc_278 GATE N_A_476_413#_c_671_n 0.00530459f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_279 N_GATE_M1015_g N_VPWR_c_828_n 0.0140188f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_280 N_GATE_M1015_g N_VPWR_c_835_n 0.00259464f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_281 N_GATE_M1015_g N_VPWR_c_826_n 0.00340558f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_282 N_GATE_c_277_n N_VGND_c_940_n 0.00394422f $X=1.83 $Y=1.685 $X2=0 $Y2=0
cc_283 N_GATE_c_278_n N_VGND_c_940_n 0.00122676f $X=1.905 $Y=1.09 $X2=0 $Y2=0
cc_284 N_GATE_c_282_n N_VGND_c_940_n 0.00393477f $X=1.985 $Y=1.56 $X2=0 $Y2=0
cc_285 GATE N_VGND_c_940_n 0.0164199f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_286 GATE N_VGND_c_945_n 0.0076037f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_287 N_GATE_c_278_n N_VGND_c_948_n 9.32477e-19 $X=1.905 $Y=1.09 $X2=0 $Y2=0
cc_288 GATE N_VGND_c_948_n 0.00629773f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_289 GATE A_396_119# 0.0135437f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_290 N_A_193_47#_c_322_n N_A_27_47#_c_415_n 8.4897e-19 $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_291 N_A_193_47#_c_322_n N_A_27_47#_c_416_n 0.0184126f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_292 N_A_193_47#_c_332_n N_A_27_47#_M1000_g 2.19569e-19 $X=1.1 $Y=1.96 $X2=0
+ $Y2=0
cc_293 N_A_193_47#_c_322_n N_A_27_47#_c_417_n 0.0167691f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_294 N_A_193_47#_c_322_n N_A_27_47#_c_418_n 0.0042868f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_295 N_A_193_47#_M1014_g N_A_27_47#_c_419_n 0.0109825f $X=3.18 $Y=0.43 $X2=0
+ $Y2=0
cc_296 N_A_193_47#_c_323_n N_A_27_47#_M1009_g 0.00780067f $X=2.475 $Y=1.74 $X2=0
+ $Y2=0
cc_297 N_A_193_47#_c_324_n N_A_27_47#_M1009_g 0.00948518f $X=2.59 $Y=0.9 $X2=0
+ $Y2=0
cc_298 N_A_193_47#_c_326_n N_A_27_47#_M1009_g 0.00927066f $X=3.18 $Y=0.9 $X2=0
+ $Y2=0
cc_299 N_A_193_47#_c_323_n N_A_27_47#_c_422_n 0.00566797f $X=2.475 $Y=1.74 $X2=0
+ $Y2=0
cc_300 N_A_193_47#_c_325_n N_A_27_47#_c_422_n 0.00887274f $X=3.055 $Y=0.9 $X2=0
+ $Y2=0
cc_301 N_A_193_47#_c_326_n N_A_27_47#_c_422_n 0.00778651f $X=3.18 $Y=0.9 $X2=0
+ $Y2=0
cc_302 N_A_193_47#_c_323_n N_A_27_47#_c_423_n 0.00402836f $X=2.475 $Y=1.74 $X2=0
+ $Y2=0
cc_303 N_A_193_47#_c_331_n N_A_27_47#_c_423_n 0.01702f $X=2.475 $Y=1.74 $X2=0
+ $Y2=0
cc_304 N_A_193_47#_M1005_g N_A_27_47#_M1002_g 0.0178331f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_305 N_A_193_47#_c_329_n N_A_27_47#_M1002_g 0.00167159f $X=2.39 $Y=1.94 $X2=0
+ $Y2=0
cc_306 N_A_193_47#_c_323_n N_A_27_47#_M1002_g 0.00500062f $X=2.475 $Y=1.74 $X2=0
+ $Y2=0
cc_307 N_A_193_47#_c_331_n N_A_27_47#_M1002_g 0.0165844f $X=2.475 $Y=1.74 $X2=0
+ $Y2=0
cc_308 N_A_193_47#_c_322_n N_A_27_47#_c_425_n 0.00863104f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_309 N_A_193_47#_c_322_n N_A_27_47#_c_434_n 0.0013042f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_310 N_A_193_47#_c_322_n N_A_27_47#_c_435_n 0.0250776f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_311 N_A_193_47#_c_322_n N_A_27_47#_c_427_n 0.0232864f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_312 N_A_193_47#_c_322_n N_A_27_47#_c_428_n 0.0166222f $X=1.1 $Y=0.425 $X2=0
+ $Y2=0
cc_313 N_A_193_47#_M1014_g N_A_642_307#_M1004_g 0.0349903f $X=3.18 $Y=0.43 $X2=0
+ $Y2=0
cc_314 N_A_193_47#_c_326_n N_A_642_307#_c_563_n 8.61266e-19 $X=3.18 $Y=0.9 $X2=0
+ $Y2=0
cc_315 N_A_193_47#_M1005_g N_A_476_413#_c_678_n 0.00290984f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_316 N_A_193_47#_c_329_n N_A_476_413#_c_678_n 0.00700812f $X=2.39 $Y=1.94
+ $X2=0 $Y2=0
cc_317 N_A_193_47#_c_331_n N_A_476_413#_c_678_n 0.00202018f $X=2.475 $Y=1.74
+ $X2=0 $Y2=0
cc_318 N_A_193_47#_M1014_g N_A_476_413#_c_671_n 0.00947094f $X=3.18 $Y=0.43
+ $X2=0 $Y2=0
cc_319 N_A_193_47#_c_325_n N_A_476_413#_c_671_n 0.0177012f $X=3.055 $Y=0.9 $X2=0
+ $Y2=0
cc_320 N_A_193_47#_c_326_n N_A_476_413#_c_671_n 0.0044688f $X=3.18 $Y=0.9 $X2=0
+ $Y2=0
cc_321 N_A_193_47#_c_329_n N_A_476_413#_c_666_n 0.00700895f $X=2.39 $Y=1.94
+ $X2=0 $Y2=0
cc_322 N_A_193_47#_c_323_n N_A_476_413#_c_666_n 0.0187722f $X=2.475 $Y=1.74
+ $X2=0 $Y2=0
cc_323 N_A_193_47#_c_326_n N_A_476_413#_c_658_n 4.27554e-19 $X=3.18 $Y=0.9 $X2=0
+ $Y2=0
cc_324 N_A_193_47#_c_323_n N_A_476_413#_c_659_n 0.00509542f $X=2.475 $Y=1.74
+ $X2=0 $Y2=0
cc_325 N_A_193_47#_c_325_n N_A_476_413#_c_659_n 0.010612f $X=3.055 $Y=0.9 $X2=0
+ $Y2=0
cc_326 N_A_193_47#_c_326_n N_A_476_413#_c_659_n 0.00425627f $X=3.18 $Y=0.9 $X2=0
+ $Y2=0
cc_327 N_A_193_47#_M1014_g N_A_476_413#_c_660_n 0.00454479f $X=3.18 $Y=0.43
+ $X2=0 $Y2=0
cc_328 N_A_193_47#_c_325_n N_A_476_413#_c_660_n 0.00805965f $X=3.055 $Y=0.9
+ $X2=0 $Y2=0
cc_329 N_A_193_47#_c_326_n N_A_476_413#_c_663_n 9.61131e-19 $X=3.18 $Y=0.9 $X2=0
+ $Y2=0
cc_330 N_A_193_47#_c_329_n N_VPWR_M1015_s 0.00507355f $X=2.39 $Y=1.94 $X2=0
+ $Y2=0
cc_331 N_A_193_47#_c_332_n N_VPWR_c_827_n 0.0127357f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_332 N_A_193_47#_M1005_g N_VPWR_c_828_n 0.00221309f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_333 N_A_193_47#_c_329_n N_VPWR_c_828_n 0.0235582f $X=2.39 $Y=1.94 $X2=0 $Y2=0
cc_334 N_A_193_47#_c_332_n N_VPWR_c_828_n 0.0189906f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_335 N_A_193_47#_c_329_n N_VPWR_c_834_n 0.002731f $X=2.39 $Y=1.94 $X2=0 $Y2=0
cc_336 N_A_193_47#_c_332_n N_VPWR_c_834_n 0.016699f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_337 N_A_193_47#_M1005_g N_VPWR_c_835_n 0.00433717f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_338 N_A_193_47#_c_329_n N_VPWR_c_835_n 0.00976688f $X=2.39 $Y=1.94 $X2=0
+ $Y2=0
cc_339 N_A_193_47#_M1005_g N_VPWR_c_826_n 0.00664549f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_340 N_A_193_47#_c_329_n N_VPWR_c_826_n 0.0232398f $X=2.39 $Y=1.94 $X2=0 $Y2=0
cc_341 N_A_193_47#_c_332_n N_VPWR_c_826_n 0.00973235f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_342 N_A_193_47#_c_329_n A_381_369# 0.00559323f $X=2.39 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_343 N_A_193_47#_c_322_n N_VGND_c_940_n 0.0464822f $X=1.1 $Y=0.425 $X2=0 $Y2=0
cc_344 N_A_193_47#_c_322_n N_VGND_c_944_n 0.0177915f $X=1.1 $Y=0.425 $X2=0 $Y2=0
cc_345 N_A_193_47#_M1014_g N_VGND_c_945_n 0.00384492f $X=3.18 $Y=0.43 $X2=0
+ $Y2=0
cc_346 N_A_193_47#_M1010_d N_VGND_c_948_n 0.00381667f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_347 N_A_193_47#_M1014_g N_VGND_c_948_n 0.00616835f $X=3.18 $Y=0.43 $X2=0
+ $Y2=0
cc_348 N_A_193_47#_c_322_n N_VGND_c_948_n 0.0101048f $X=1.1 $Y=0.425 $X2=0 $Y2=0
cc_349 N_A_193_47#_c_324_n N_VGND_c_948_n 0.00692839f $X=2.59 $Y=0.9 $X2=0 $Y2=0
cc_350 N_A_193_47#_c_325_n N_VGND_c_948_n 0.00776489f $X=3.055 $Y=0.9 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_422_n N_A_642_307#_M1004_g 0.00385724f $X=2.85 $Y=1.32 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_M1002_g N_A_642_307#_c_563_n 0.0656786f $X=2.925 $Y=2.275
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_M1002_g N_A_476_413#_c_678_n 0.0146203f $X=2.925 $Y=2.275
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_M1009_g N_A_476_413#_c_671_n 0.00218822f $X=2.455 $Y=0.54
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_422_n N_A_476_413#_c_666_n 0.00957693f $X=2.85 $Y=1.32 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_M1009_g N_A_476_413#_c_659_n 3.86069e-19 $X=2.455 $Y=0.54
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_c_422_n N_A_476_413#_c_659_n 0.00151673f $X=2.85 $Y=1.32 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_434_n N_VPWR_M1008_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_359 N_A_27_47#_M1000_g N_VPWR_c_827_n 0.00940337f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_434_n N_VPWR_c_827_n 0.0155904f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_361 N_A_27_47#_c_436_n N_VPWR_c_827_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_362 N_A_27_47#_M1000_g N_VPWR_c_828_n 0.00181768f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_434_n N_VPWR_c_833_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_364 N_A_27_47#_c_436_n N_VPWR_c_833_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_365 N_A_27_47#_M1000_g N_VPWR_c_834_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_M1002_g N_VPWR_c_835_n 0.00366111f $X=2.925 $Y=2.275 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_M1000_g N_VPWR_c_826_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_M1002_g N_VPWR_c_826_n 0.00560345f $X=2.925 $Y=2.275 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_434_n N_VPWR_c_826_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_370 N_A_27_47#_c_436_n N_VPWR_c_826_n 0.00646745f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_371 N_A_27_47#_c_425_n N_VGND_M1019_d 0.00169549f $X=0.61 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_372 N_A_27_47#_c_415_n N_VGND_c_939_n 0.00727594f $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_373 N_A_27_47#_c_420_n N_VGND_c_939_n 6.19779e-19 $X=1.45 $Y=0.18 $X2=0 $Y2=0
cc_374 N_A_27_47#_c_425_n N_VGND_c_939_n 0.0149823f $X=0.61 $Y=0.7 $X2=0 $Y2=0
cc_375 N_A_27_47#_c_427_n N_VGND_c_939_n 0.00122968f $X=0.755 $Y=1.225 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_429_n N_VGND_c_939_n 5.68744e-19 $X=0.89 $Y=1.225 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_415_n N_VGND_c_940_n 3.97733e-19 $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_378 N_A_27_47#_c_418_n N_VGND_c_940_n 0.00934292f $X=1.375 $Y=0.73 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_419_n N_VGND_c_940_n 0.0229858f $X=2.38 $Y=0.18 $X2=0 $Y2=0
cc_380 N_A_27_47#_M1009_g N_VGND_c_940_n 0.00327004f $X=2.455 $Y=0.54 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_537_p N_VGND_c_943_n 0.0110394f $X=0.26 $Y=0.425 $X2=0 $Y2=0
cc_382 N_A_27_47#_c_425_n N_VGND_c_943_n 0.00255672f $X=0.61 $Y=0.7 $X2=0 $Y2=0
cc_383 N_A_27_47#_c_415_n N_VGND_c_944_n 0.0046653f $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_384 N_A_27_47#_c_417_n N_VGND_c_944_n 3.66494e-19 $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_385 N_A_27_47#_c_420_n N_VGND_c_944_n 0.00698559f $X=1.45 $Y=0.18 $X2=0 $Y2=0
cc_386 N_A_27_47#_c_419_n N_VGND_c_945_n 0.023604f $X=2.38 $Y=0.18 $X2=0 $Y2=0
cc_387 N_A_27_47#_M1019_s N_VGND_c_948_n 0.00367415f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_415_n N_VGND_c_948_n 0.00805453f $X=0.89 $Y=0.73 $X2=0 $Y2=0
cc_389 N_A_27_47#_c_419_n N_VGND_c_948_n 0.0302007f $X=2.38 $Y=0.18 $X2=0 $Y2=0
cc_390 N_A_27_47#_c_420_n N_VGND_c_948_n 0.0100087f $X=1.45 $Y=0.18 $X2=0 $Y2=0
cc_391 N_A_27_47#_c_537_p N_VGND_c_948_n 0.00641103f $X=0.26 $Y=0.425 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_425_n N_VGND_c_948_n 0.00557795f $X=0.61 $Y=0.7 $X2=0 $Y2=0
cc_393 N_A_642_307#_M1004_g N_A_476_413#_M1018_g 0.0106889f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_394 N_A_642_307#_M1007_g N_A_476_413#_M1018_g 0.0322927f $X=4.71 $Y=2.165
+ $X2=0 $Y2=0
cc_395 N_A_642_307#_c_561_n N_A_476_413#_M1018_g 0.00358342f $X=4.527 $Y=1.535
+ $X2=0 $Y2=0
cc_396 N_A_642_307#_c_562_n N_A_476_413#_M1018_g 0.0184612f $X=4.025 $Y=1.755
+ $X2=0 $Y2=0
cc_397 N_A_642_307#_M1003_g N_A_476_413#_c_678_n 0.00338501f $X=3.285 $Y=2.275
+ $X2=0 $Y2=0
cc_398 N_A_642_307#_M1004_g N_A_476_413#_c_671_n 0.0074137f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_399 N_A_642_307#_M1003_g N_A_476_413#_c_666_n 0.0140667f $X=3.285 $Y=2.275
+ $X2=0 $Y2=0
cc_400 N_A_642_307#_M1004_g N_A_476_413#_c_666_n 0.00390654f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_401 N_A_642_307#_c_560_n N_A_476_413#_c_666_n 0.0214954f $X=3.91 $Y=1.7 $X2=0
+ $Y2=0
cc_402 N_A_642_307#_c_563_n N_A_476_413#_c_666_n 0.00742928f $X=3.655 $Y=1.7
+ $X2=0 $Y2=0
cc_403 N_A_642_307#_c_560_n N_A_476_413#_c_658_n 0.00714741f $X=3.91 $Y=1.7
+ $X2=0 $Y2=0
cc_404 N_A_642_307#_c_563_n N_A_476_413#_c_658_n 0.0101207f $X=3.655 $Y=1.7
+ $X2=0 $Y2=0
cc_405 N_A_642_307#_M1004_g N_A_476_413#_c_660_n 0.0134126f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_406 N_A_642_307#_c_555_n N_A_476_413#_c_660_n 0.00996062f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_407 N_A_642_307#_M1004_g N_A_476_413#_c_661_n 0.00326591f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_408 N_A_642_307#_c_550_n N_A_476_413#_c_661_n 3.09008e-19 $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_409 N_A_642_307#_c_560_n N_A_476_413#_c_661_n 0.0117588f $X=3.91 $Y=1.7 $X2=0
+ $Y2=0
cc_410 N_A_642_307#_c_562_n N_A_476_413#_c_661_n 0.0148361f $X=4.025 $Y=1.755
+ $X2=0 $Y2=0
cc_411 N_A_642_307#_c_554_n N_A_476_413#_c_661_n 0.0256428f $X=4.655 $Y=1.16
+ $X2=0 $Y2=0
cc_412 N_A_642_307#_M1004_g N_A_476_413#_c_662_n 0.0195941f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_413 N_A_642_307#_c_550_n N_A_476_413#_c_662_n 0.021275f $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_414 N_A_642_307#_c_562_n N_A_476_413#_c_662_n 0.00463369f $X=4.025 $Y=1.755
+ $X2=0 $Y2=0
cc_415 N_A_642_307#_c_554_n N_A_476_413#_c_662_n 0.00358342f $X=4.655 $Y=1.16
+ $X2=0 $Y2=0
cc_416 N_A_642_307#_M1004_g N_A_476_413#_c_663_n 0.0122771f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_642_307#_c_560_n N_A_476_413#_c_663_n 0.0104303f $X=3.91 $Y=1.7 $X2=0
+ $Y2=0
cc_418 N_A_642_307#_c_563_n N_A_476_413#_c_663_n 5.70452e-19 $X=3.655 $Y=1.7
+ $X2=0 $Y2=0
cc_419 N_A_642_307#_M1004_g N_A_476_413#_c_664_n 0.0185609f $X=3.655 $Y=0.445
+ $X2=0 $Y2=0
cc_420 N_A_642_307#_c_550_n N_A_476_413#_c_664_n 0.00652245f $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_421 N_A_642_307#_c_555_n N_A_476_413#_c_664_n 0.00621473f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_422 N_A_642_307#_c_551_n N_A_957_369#_c_747_n 0.0043908f $X=5.06 $Y=0.805
+ $X2=0 $Y2=0
cc_423 N_A_642_307#_c_552_n N_A_957_369#_c_747_n 0.00371139f $X=5.135 $Y=0.73
+ $X2=0 $Y2=0
cc_424 N_A_642_307#_c_555_n N_A_957_369#_c_747_n 0.00661846f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_425 N_A_642_307#_M1007_g N_A_957_369#_c_760_n 0.00795417f $X=4.71 $Y=2.165
+ $X2=0 $Y2=0
cc_426 N_A_642_307#_c_551_n N_A_957_369#_c_748_n 0.00338363f $X=5.06 $Y=0.805
+ $X2=0 $Y2=0
cc_427 N_A_642_307#_c_550_n N_A_957_369#_c_749_n 7.22329e-19 $X=4.71 $Y=1.325
+ $X2=0 $Y2=0
cc_428 N_A_642_307#_c_551_n N_A_957_369#_c_749_n 0.00753447f $X=5.06 $Y=0.805
+ $X2=0 $Y2=0
cc_429 N_A_642_307#_c_555_n N_A_957_369#_c_749_n 0.00824229f $X=4.542 $Y=0.995
+ $X2=0 $Y2=0
cc_430 N_A_642_307#_M1007_g N_A_957_369#_c_756_n 0.00281757f $X=4.71 $Y=2.165
+ $X2=0 $Y2=0
cc_431 N_A_642_307#_c_562_n N_A_957_369#_c_756_n 0.00677764f $X=4.025 $Y=1.755
+ $X2=0 $Y2=0
cc_432 N_A_642_307#_c_551_n N_A_957_369#_c_781_n 0.00372863f $X=5.06 $Y=0.805
+ $X2=0 $Y2=0
cc_433 N_A_642_307#_c_552_n N_A_957_369#_c_781_n 0.00812233f $X=5.135 $Y=0.73
+ $X2=0 $Y2=0
cc_434 N_A_642_307#_c_553_n N_A_957_369#_c_781_n 0.0194395f $X=4.405 $Y=0.45
+ $X2=0 $Y2=0
cc_435 N_A_642_307#_c_562_n N_VPWR_M1018_d 0.00213578f $X=4.025 $Y=1.755 $X2=0
+ $Y2=0
cc_436 N_A_642_307#_M1003_g N_VPWR_c_829_n 0.00467052f $X=3.285 $Y=2.275 $X2=0
+ $Y2=0
cc_437 N_A_642_307#_c_560_n N_VPWR_c_829_n 0.0144253f $X=3.91 $Y=1.7 $X2=0 $Y2=0
cc_438 N_A_642_307#_c_634_p N_VPWR_c_829_n 0.0199633f $X=4.025 $Y=2.27 $X2=0
+ $Y2=0
cc_439 N_A_642_307#_c_563_n N_VPWR_c_829_n 0.00709979f $X=3.655 $Y=1.7 $X2=0
+ $Y2=0
cc_440 N_A_642_307#_c_634_p N_VPWR_c_830_n 0.0121002f $X=4.025 $Y=2.27 $X2=0
+ $Y2=0
cc_441 N_A_642_307#_M1007_g N_VPWR_c_831_n 0.00338987f $X=4.71 $Y=2.165 $X2=0
+ $Y2=0
cc_442 N_A_642_307#_c_562_n N_VPWR_c_831_n 0.0198055f $X=4.025 $Y=1.755 $X2=0
+ $Y2=0
cc_443 N_A_642_307#_M1003_g N_VPWR_c_835_n 0.00563437f $X=3.285 $Y=2.275 $X2=0
+ $Y2=0
cc_444 N_A_642_307#_M1007_g N_VPWR_c_836_n 0.00585385f $X=4.71 $Y=2.165 $X2=0
+ $Y2=0
cc_445 N_A_642_307#_M1018_s N_VPWR_c_826_n 0.00340182f $X=3.89 $Y=1.485 $X2=0
+ $Y2=0
cc_446 N_A_642_307#_M1003_g N_VPWR_c_826_n 0.0112135f $X=3.285 $Y=2.275 $X2=0
+ $Y2=0
cc_447 N_A_642_307#_M1007_g N_VPWR_c_826_n 0.0115396f $X=4.71 $Y=2.165 $X2=0
+ $Y2=0
cc_448 N_A_642_307#_c_560_n N_VPWR_c_826_n 0.00859146f $X=3.91 $Y=1.7 $X2=0
+ $Y2=0
cc_449 N_A_642_307#_c_634_p N_VPWR_c_826_n 0.00827281f $X=4.025 $Y=2.27 $X2=0
+ $Y2=0
cc_450 N_A_642_307#_c_563_n N_VPWR_c_826_n 0.00167685f $X=3.655 $Y=1.7 $X2=0
+ $Y2=0
cc_451 N_A_642_307#_M1004_g N_VGND_c_941_n 0.00749145f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_642_307#_M1004_g N_VGND_c_945_n 0.00391009f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_453 N_A_642_307#_c_550_n N_VGND_c_946_n 0.00398989f $X=4.71 $Y=1.325 $X2=0
+ $Y2=0
cc_454 N_A_642_307#_c_551_n N_VGND_c_946_n 3.02019e-19 $X=5.06 $Y=0.805 $X2=0
+ $Y2=0
cc_455 N_A_642_307#_c_552_n N_VGND_c_946_n 0.00447211f $X=5.135 $Y=0.73 $X2=0
+ $Y2=0
cc_456 N_A_642_307#_c_553_n N_VGND_c_946_n 0.0179446f $X=4.405 $Y=0.45 $X2=0
+ $Y2=0
cc_457 N_A_642_307#_M1011_d N_VGND_c_948_n 0.00387172f $X=4.27 $Y=0.235 $X2=0
+ $Y2=0
cc_458 N_A_642_307#_M1004_g N_VGND_c_948_n 0.00602379f $X=3.655 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_A_642_307#_c_550_n N_VGND_c_948_n 0.00516342f $X=4.71 $Y=1.325 $X2=0
+ $Y2=0
cc_460 N_A_642_307#_c_552_n N_VGND_c_948_n 0.00684735f $X=5.135 $Y=0.73 $X2=0
+ $Y2=0
cc_461 N_A_642_307#_c_553_n N_VGND_c_948_n 0.00992144f $X=4.405 $Y=0.45 $X2=0
+ $Y2=0
cc_462 N_A_476_413#_c_678_n N_VPWR_c_828_n 0.00474258f $X=3.055 $Y=2.34 $X2=0
+ $Y2=0
cc_463 N_A_476_413#_M1018_g N_VPWR_c_829_n 0.00237885f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_464 N_A_476_413#_M1018_g N_VPWR_c_830_n 0.00583607f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_465 N_A_476_413#_M1018_g N_VPWR_c_831_n 0.00222005f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_466 N_A_476_413#_c_678_n N_VPWR_c_835_n 0.0344605f $X=3.055 $Y=2.34 $X2=0
+ $Y2=0
cc_467 N_A_476_413#_M1005_d N_VPWR_c_826_n 0.00425502f $X=2.38 $Y=2.065 $X2=0
+ $Y2=0
cc_468 N_A_476_413#_M1018_g N_VPWR_c_826_n 0.0121029f $X=4.235 $Y=1.985 $X2=0
+ $Y2=0
cc_469 N_A_476_413#_c_678_n N_VPWR_c_826_n 0.0267056f $X=3.055 $Y=2.34 $X2=0
+ $Y2=0
cc_470 N_A_476_413#_c_678_n A_600_413# 0.00102341f $X=3.055 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_471 N_A_476_413#_c_671_n N_VGND_c_941_n 0.0137306f $X=3.555 $Y=0.475 $X2=0
+ $Y2=0
cc_472 N_A_476_413#_c_660_n N_VGND_c_941_n 0.00358434f $X=3.64 $Y=0.995 $X2=0
+ $Y2=0
cc_473 N_A_476_413#_c_661_n N_VGND_c_941_n 0.00829692f $X=4.09 $Y=1.16 $X2=0
+ $Y2=0
cc_474 N_A_476_413#_c_662_n N_VGND_c_941_n 0.00311808f $X=4.09 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_A_476_413#_c_664_n N_VGND_c_941_n 0.0099666f $X=4.132 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_A_476_413#_c_671_n N_VGND_c_945_n 0.0293579f $X=3.555 $Y=0.475 $X2=0
+ $Y2=0
cc_477 N_A_476_413#_c_664_n N_VGND_c_946_n 0.00486043f $X=4.132 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_476_413#_M1009_d N_VGND_c_948_n 0.00392318f $X=2.53 $Y=0.33 $X2=0
+ $Y2=0
cc_479 N_A_476_413#_c_671_n N_VGND_c_948_n 0.0306841f $X=3.555 $Y=0.475 $X2=0
+ $Y2=0
cc_480 N_A_476_413#_c_664_n N_VGND_c_948_n 0.00965187f $X=4.132 $Y=0.995 $X2=0
+ $Y2=0
cc_481 N_A_476_413#_c_671_n A_651_47# 0.00632435f $X=3.555 $Y=0.475 $X2=-0.19
+ $Y2=-0.24
cc_482 N_A_957_369#_c_755_n N_VPWR_M1013_d 0.00653118f $X=5.75 $Y=1.81 $X2=0
+ $Y2=0
cc_483 N_A_957_369#_c_758_n N_VPWR_M1013_d 0.00279081f $X=5.835 $Y=1.725 $X2=0
+ $Y2=0
cc_484 N_A_957_369#_M1012_g N_VPWR_c_832_n 0.00981345f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_A_957_369#_c_760_n N_VPWR_c_832_n 0.0217852f $X=5.17 $Y=2 $X2=0 $Y2=0
cc_486 N_A_957_369#_c_755_n N_VPWR_c_832_n 0.0147141f $X=5.75 $Y=1.81 $X2=0
+ $Y2=0
cc_487 N_A_957_369#_c_760_n N_VPWR_c_836_n 0.0230652f $X=5.17 $Y=2 $X2=0 $Y2=0
cc_488 N_A_957_369#_M1012_g N_VPWR_c_837_n 0.00486043f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_489 N_A_957_369#_M1007_d N_VPWR_c_826_n 0.013359f $X=4.785 $Y=1.845 $X2=0
+ $Y2=0
cc_490 N_A_957_369#_M1012_g N_VPWR_c_826_n 0.00915314f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_491 N_A_957_369#_c_760_n N_VPWR_c_826_n 0.0126319f $X=5.17 $Y=2 $X2=0 $Y2=0
cc_492 N_A_957_369#_c_755_n N_VPWR_c_826_n 0.00847738f $X=5.75 $Y=1.81 $X2=0
+ $Y2=0
cc_493 N_A_957_369#_M1012_g N_GCLK_c_922_n 0.00340846f $X=5.97 $Y=1.985 $X2=0
+ $Y2=0
cc_494 N_A_957_369#_c_748_n N_GCLK_c_922_n 0.0135077f $X=5.75 $Y=0.85 $X2=0
+ $Y2=0
cc_495 N_A_957_369#_c_750_n N_GCLK_c_922_n 0.0287817f $X=5.915 $Y=1.16 $X2=0
+ $Y2=0
cc_496 N_A_957_369#_c_751_n N_GCLK_c_922_n 0.00754825f $X=5.915 $Y=1.16 $X2=0
+ $Y2=0
cc_497 N_A_957_369#_c_758_n N_GCLK_c_922_n 0.00911561f $X=5.835 $Y=1.725 $X2=0
+ $Y2=0
cc_498 N_A_957_369#_c_753_n N_GCLK_c_922_n 0.0104416f $X=5.915 $Y=0.995 $X2=0
+ $Y2=0
cc_499 N_A_957_369#_c_748_n N_VGND_M1016_d 0.0024638f $X=5.75 $Y=0.85 $X2=0
+ $Y2=0
cc_500 N_A_957_369#_c_748_n N_VGND_c_942_n 0.0110864f $X=5.75 $Y=0.85 $X2=0
+ $Y2=0
cc_501 N_A_957_369#_c_751_n N_VGND_c_942_n 2.76169e-19 $X=5.915 $Y=1.16 $X2=0
+ $Y2=0
cc_502 N_A_957_369#_c_781_n N_VGND_c_942_n 0.00788856f $X=4.925 $Y=0.455 $X2=0
+ $Y2=0
cc_503 N_A_957_369#_c_753_n N_VGND_c_942_n 0.00274164f $X=5.915 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_957_369#_c_781_n N_VGND_c_946_n 0.0158526f $X=4.925 $Y=0.455 $X2=0
+ $Y2=0
cc_505 N_A_957_369#_c_753_n N_VGND_c_947_n 0.00585385f $X=5.915 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_A_957_369#_M1001_s N_VGND_c_948_n 0.00258814f $X=4.8 $Y=0.235 $X2=0
+ $Y2=0
cc_507 N_A_957_369#_c_748_n N_VGND_c_948_n 0.0238999f $X=5.75 $Y=0.85 $X2=0
+ $Y2=0
cc_508 N_A_957_369#_c_781_n N_VGND_c_948_n 0.0113132f $X=4.925 $Y=0.455 $X2=0
+ $Y2=0
cc_509 N_A_957_369#_c_753_n N_VGND_c_948_n 0.00846015f $X=5.915 $Y=0.995 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_826_n A_381_369# 0.00410346f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_511 N_VPWR_c_826_n A_600_413# 0.00170467f $X=6.21 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_512 N_VPWR_c_826_n N_GCLK_M1012_d 0.00365806f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_513 N_VPWR_c_837_n N_GCLK_c_926_n 0.0170871f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_514 N_VPWR_c_826_n N_GCLK_c_926_n 0.0100807f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_515 N_GCLK_c_923_n N_VGND_c_947_n 0.018533f $X=6.262 $Y=0.425 $X2=0 $Y2=0
cc_516 N_GCLK_M1006_d N_VGND_c_948_n 0.00240587f $X=6.045 $Y=0.235 $X2=0 $Y2=0
cc_517 N_GCLK_c_923_n N_VGND_c_948_n 0.0113482f $X=6.262 $Y=0.425 $X2=0 $Y2=0
cc_518 N_VGND_c_948_n A_651_47# 0.00282601f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24
cc_519 N_VGND_c_948_n A_1042_47# 0.00285576f $X=6.21 $Y=0 $X2=-0.19 $Y2=-0.24

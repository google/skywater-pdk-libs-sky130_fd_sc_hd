* File: sky130_fd_sc_hd__xnor3_4.spice
* Created: Thu Aug 27 14:49:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__xnor3_4.spice.pex"
.subckt sky130_fd_sc_hd__xnor3_4  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_101_21#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_101_21#_M1015_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.08775 PD=0.93 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1015_d N_A_101_21#_M1022_g N_X_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.08775 PD=0.93 PS=0.92 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1027_d N_A_101_21#_M1027_g N_X_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.141542 AS=0.08775 PD=1.25748 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1016 N_A_492_93#_M1016_d N_C_M1016_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1785 AS=0.0914579 PD=1.69 PS=0.812523 NRD=39.996 NRS=46.5 M=1 R=2.8
+ SA=75002 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1024 N_A_101_21#_M1024_d N_C_M1024_g N_A_631_49#_M1024_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=0.936 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1020 N_A_607_325#_M1020_d N_A_492_93#_M1020_g N_A_101_21#_M1024_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.224 AS=0.0928 PD=1.98 PS=0.93 NRD=12.18 NRS=0.936 M=1
+ R=4.26667 SA=75000.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1003 N_A_1011_297#_M1003_d N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.16515 AS=0.1885 PD=1.82 PS=1.88 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_607_325#_M1007_d N_B_M1007_g N_A_1117_297#_M1007_s VNB NSHORT L=0.15
+ W=0.64 AD=0.219834 AS=0.16275 PD=1.5034 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1021 N_A_1382_49#_M1021_d N_A_1011_297#_M1021_g N_A_607_325#_M1007_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.152666 AS=0.144266 PD=1.0183 PS=0.986604 NRD=88.14
+ NRS=94.284 M=1 R=2.8 SA=75000.9 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1023 N_A_631_49#_M1023_d N_B_M1023_g N_A_1382_49#_M1021_d VNB NSHORT L=0.15
+ W=0.64 AD=0.145368 AS=0.232634 PD=1.13548 PS=1.5517 NRD=0.936 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_1117_297#_M1006_d N_A_1011_297#_M1006_g N_A_631_49#_M1023_d VNB
+ NSHORT L=0.15 W=0.6 AD=0.106452 AS=0.136282 PD=0.958065 PS=1.06452 NRD=15
+ NRS=32.988 M=1 R=4 SA=75001.9 SB=75001.1 A=0.09 P=1.5 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_1117_297#_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.113548 PD=0.91 PS=1.02194 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_1382_49#_M1009_d N_A_1117_297#_M1009_g N_VGND_M1004_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0864 PD=1.85 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_101_21#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_101_21#_M1002_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.135 PD=1.3 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1002_d N_A_101_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.135 PD=1.3 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_A_101_21#_M1014_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.206098 AS=0.135 PD=1.66463 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1025 N_A_492_93#_M1025_d N_C_M1025_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1792 AS=0.131902 PD=1.84 PS=1.06537 NRD=0 NRS=46.492 M=1 R=4.26667
+ SA=75002 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_A_101_21#_M1011_d N_C_M1011_g N_A_607_325#_M1011_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.15295 AS=0.273 PD=1.315 PS=2.33 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1026 N_A_631_49#_M1026_d N_A_492_93#_M1026_g N_A_101_21#_M1011_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.32235 AS=0.15295 PD=2.45 PS=1.315 NRD=23.443 NRS=15.2281
+ M=1 R=5.6 SA=75000.6 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1000 N_A_1011_297#_M1000_d N_B_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.25655 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1018 N_A_631_49#_M1018_d N_B_M1018_g N_A_1117_297#_M1018_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.275951 AS=0.3528 PD=1.64027 PS=2.52 NRD=45.7237 NRS=36.3465 M=1
+ R=5.6 SA=75000.3 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1019 N_A_1382_49#_M1019_d N_A_1011_297#_M1019_g N_A_631_49#_M1018_d VPB
+ PHIGHVT L=0.15 W=0.64 AD=0.246 AS=0.210249 PD=1.525 PS=1.24973 NRD=138.511
+ NRS=40.0107 M=1 R=4.26667 SA=75001.1 SB=75002 A=0.096 P=1.58 MULT=1
MM1013 N_A_607_325#_M1013_d N_B_M1013_g N_A_1382_49#_M1019_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.126097 AS=0.246 PD=1.04216 PS=1.525 NRD=43.7143 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_1117_297#_M1008_d N_A_1011_297#_M1008_g N_A_607_325#_M1013_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.156587 AS=0.165503 PD=1.23717 PS=1.36784
+ NRD=30.8108 NRS=0 M=1 R=5.6 SA=75001.6 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g N_A_1117_297#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.186413 PD=1.27 PS=1.47283 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_A_1382_49#_M1012_d N_A_1117_297#_M1012_g N_VPWR_M1017_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.285 AS=0.135 PD=2.57 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=16.1142 P=23.29
*
.include "sky130_fd_sc_hd__xnor3_4.spice.SKY130_FD_SC_HD__XNOR3_4.pxi"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.075000 5.395000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.350000 1.075000 4.680000 1.445000 ;
        RECT 4.350000 1.445000 5.735000 1.615000 ;
        RECT 5.565000 1.075000 6.355000 1.275000 ;
        RECT 5.565000 1.275000 5.735000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.075000 3.680000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.420000 1.075000 2.955000 1.445000 ;
        RECT 2.420000 1.445000 4.180000 1.615000 ;
        RECT 3.850000 1.075000 4.180000 1.445000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.770000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.730000 1.615000 ;
        RECT 0.600000 0.265000 0.930000 0.725000 ;
        RECT 0.640000 1.615000 0.890000 2.465000 ;
        RECT 1.440000 0.255000 1.770000 0.725000 ;
        RECT 1.480000 1.615000 1.730000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.220000  1.825000 0.470000 2.635000 ;
      RECT 0.260000  0.085000 0.430000 0.555000 ;
      RECT 0.540000  1.075000 2.230000 1.275000 ;
      RECT 1.060000  1.795000 1.310000 2.635000 ;
      RECT 1.100000  0.085000 1.270000 0.555000 ;
      RECT 1.900000  1.275000 2.230000 1.785000 ;
      RECT 1.900000  1.785000 3.930000 1.955000 ;
      RECT 1.900000  2.125000 2.150000 2.635000 ;
      RECT 1.940000  0.085000 2.630000 0.555000 ;
      RECT 1.940000  0.735000 5.310000 0.905000 ;
      RECT 1.940000  0.905000 2.230000 1.075000 ;
      RECT 2.420000  2.125000 2.670000 2.295000 ;
      RECT 2.420000  2.295000 4.430000 2.465000 ;
      RECT 2.800000  0.255000 3.970000 0.475000 ;
      RECT 2.840000  1.955000 3.090000 2.125000 ;
      RECT 3.170000  0.645000 3.605000 0.735000 ;
      RECT 3.260000  2.125000 3.510000 2.295000 ;
      RECT 3.680000  1.955000 3.930000 2.125000 ;
      RECT 4.100000  1.785000 6.110000 1.955000 ;
      RECT 4.100000  1.955000 4.430000 2.295000 ;
      RECT 4.185000  0.085000 4.355000 0.555000 ;
      RECT 4.560000  0.255000 5.730000 0.475000 ;
      RECT 4.600000  2.125000 4.850000 2.635000 ;
      RECT 4.935000  0.645000 5.310000 0.735000 ;
      RECT 5.020000  1.955000 5.270000 2.465000 ;
      RECT 5.440000  2.125000 5.690000 2.635000 ;
      RECT 5.480000  0.475000 5.730000 0.895000 ;
      RECT 5.900000  0.085000 6.070000 0.895000 ;
      RECT 5.905000  1.455000 6.110000 1.785000 ;
      RECT 5.905000  1.955000 6.110000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__a22o_4
END LIBRARY

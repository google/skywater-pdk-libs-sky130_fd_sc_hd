* File: sky130_fd_sc_hd__dfbbn_1.spice
* Created: Tue Sep  1 19:02:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dfbbn_1.pex.spice"
.subckt sky130_fd_sc_hd__dfbbn_1  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_CLK_N_M1033_g N_A_27_47#_M1033_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_193_47#_M1013_d N_A_27_47#_M1013_g N_VGND_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_381_47#_M1002_d N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.1092 PD=0.802308 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1026 N_A_473_413#_M1026_d N_A_193_47#_M1026_g N_A_381_47#_M1002_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0675 AS=0.0609231 PD=0.735 PS=0.687692 NRD=14.988
+ NRS=16.656 M=1 R=2.4 SA=75000.7 SB=75002.7 A=0.054 P=1.02 MULT=1
MM1038 A_581_47# N_A_27_47#_M1038_g N_A_473_413#_M1026_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0618923 AS=0.0675 PD=0.692308 PS=0.735 NRD=38.964 NRS=16.656 M=1
+ R=2.4 SA=75001.2 SB=75002.1 A=0.054 P=1.02 MULT=1
MM1007 N_VGND_M1007_d N_A_647_21#_M1007_g A_581_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0722077 PD=0.84 PS=0.807692 NRD=41.424 NRS=33.396 M=1 R=2.8
+ SA=75001.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_791_47#_M1016_d N_SET_B_M1016_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0771453 AS=0.0882 PD=0.768679 PS=0.84 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1035 N_A_647_21#_M1035_d N_A_473_413#_M1035_g N_A_791_47#_M1016_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0864 AS=0.117555 PD=0.91 PS=1.17132 NRD=0 NRS=10.308 M=1
+ R=4.26667 SA=75001.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1031 N_A_791_47#_M1031_d N_A_941_21#_M1031_g N_A_647_21#_M1035_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1019 A_1159_47# N_A_647_21#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.64
+ AD=0.14848 AS=0.1664 PD=1.3952 PS=1.8 NRD=33.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1001 N_A_1256_413#_M1001_d N_A_27_47#_M1001_g A_1159_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0486 AS=0.08352 PD=0.63 PS=0.7848 NRD=0 NRS=58.992 M=1 R=2.4
+ SA=75000.8 SB=75002.5 A=0.054 P=1.02 MULT=1
MM1036 A_1363_47# N_A_193_47#_M1036_g N_A_1256_413#_M1001_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0486 PD=0.687692 PS=0.63 NRD=38.076 NRS=0 M=1 R=2.4
+ SA=75001.2 SB=75002.1 A=0.054 P=1.02 MULT=1
MM1020 N_VGND_M1020_d N_A_1415_315#_M1020_g A_1363_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0710769 PD=0.755 PS=0.802308 NRD=17.136 NRS=32.628 M=1 R=2.8
+ SA=75001.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_1555_47#_M1009_d N_SET_B_M1009_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0866943 AS=0.07035 PD=0.816226 PS=0.755 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1025 N_A_1415_315#_M1025_d N_A_1256_413#_M1025_g N_A_1555_47#_M1009_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.0864 AS=0.132106 PD=0.91 PS=1.24377 NRD=0 NRS=21.552
+ M=1 R=4.26667 SA=75001.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1032 N_A_1555_47#_M1032_d N_A_941_21#_M1032_g N_A_1415_315#_M1025_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_RESET_B_M1015_g N_A_941_21#_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_Q_N_M1030_d N_A_1415_315#_M1030_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_1415_315#_M1010_g N_A_2136_47#_M1010_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=14.28 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1027 N_Q_M1027_d N_A_2136_47#_M1027_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_CLK_N_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_381_47#_M1017_d N_D_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0651 AS=0.1092 PD=0.73 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75007
+ A=0.063 P=1.14 MULT=1
MM1021 N_A_473_413#_M1021_d N_A_27_47#_M1021_g N_A_381_47#_M1017_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.0651 PD=0.69 PS=0.73 NRD=0 NRS=16.4101 M=1 R=2.8
+ SA=75000.6 SB=75006.5 A=0.063 P=1.14 MULT=1
MM1014 A_557_413# N_A_193_47#_M1014_g N_A_473_413#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0945 AS=0.0567 PD=0.87 PS=0.69 NRD=79.7259 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75006.1 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_647_21#_M1023_g A_557_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0945 PD=0.8 PS=0.87 NRD=21.0987 NRS=79.7259 M=1 R=2.8
+ SA=75001.7 SB=75005.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_647_21#_M1004_d N_SET_B_M1004_g N_VPWR_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.098 AS=0.0798 PD=0.82 PS=0.8 NRD=53.9386 NRS=25.7873 M=1 R=2.8
+ SA=75002.2 SB=75005 A=0.063 P=1.14 MULT=1
MM1024 A_891_329# N_A_473_413#_M1024_g N_A_647_21#_M1004_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1134 AS=0.196 PD=1.11 PS=1.64 NRD=18.7544 NRS=0 M=1 R=5.6
+ SA=75001.5 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_A_941_21#_M1018_g A_891_329# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2247 AS=0.1134 PD=1.375 PS=1.11 NRD=5.8509 NRS=18.7544 M=1 R=5.6
+ SA=75001.9 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1028 A_1112_329# N_A_647_21#_M1028_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2324 AS=0.2247 PD=1.88 PS=1.375 NRD=51.9686 NRS=53.9386 M=1 R=5.6
+ SA=75002.6 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1034 N_A_1256_413#_M1034_d N_A_193_47#_M1034_g A_1112_329# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.1162 PD=0.69 PS=0.94 NRD=0 NRS=103.957 M=1 R=2.8
+ SA=75004.6 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1022 A_1340_413# N_A_27_47#_M1022_g N_A_1256_413#_M1034_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07875 AS=0.0567 PD=0.795 PS=0.69 NRD=62.1338 NRS=0 M=1 R=2.8
+ SA=75005 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1415_315#_M1008_g A_1340_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09555 AS=0.07875 PD=0.875 PS=0.795 NRD=56.2829 NRS=62.1338 M=1
+ R=2.8 SA=75005.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1012 N_A_1415_315#_M1012_d N_SET_B_M1012_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0882 AS=0.09555 PD=0.813333 PS=0.875 NRD=25.7873 NRS=25.7873 M=1
+ R=2.8 SA=75006.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_1672_329# N_A_1256_413#_M1003_g N_A_1415_315#_M1012_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.0882 AS=0.1764 PD=1.05 PS=1.62667 NRD=11.7215 NRS=10.5395
+ M=1 R=5.6 SA=75003.4 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_A_941_21#_M1005_g A_1672_329# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2184 AS=0.0882 PD=2.2 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75003.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1029 N_VPWR_M1029_d N_RESET_B_M1029_g N_A_941_21#_M1029_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.120117 AS=0.1696 PD=1.04195 PS=1.81 NRD=40.8381 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1039 N_Q_N_M1039_d N_A_1415_315#_M1039_g N_VPWR_M1029_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.187683 PD=2.52 PS=1.62805 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_1415_315#_M1006_g N_A_2136_47#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.116293 AS=0.1664 PD=1.03415 PS=1.8 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1037 N_Q_M1037_d N_A_2136_47#_M1037_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.181707 PD=2.52 PS=1.61585 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.8057 P=27.89
c_256 VPB 0 1.39343e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dfbbn_1.pxi.spice"
*
.ends
*
*

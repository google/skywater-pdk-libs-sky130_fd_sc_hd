* File: sky130_fd_sc_hd__mux2_8.spice.SKY130_FD_SC_HD__MUX2_8.pxi
* Created: Thu Aug 27 14:27:48 2020
* 
x_PM_SKY130_FD_SC_HD__MUX2_8%A_79_21# N_A_79_21#_M1022_d N_A_79_21#_M1015_s
+ N_A_79_21#_M1001_s N_A_79_21#_M1016_s N_A_79_21#_c_130_n N_A_79_21#_M1009_g
+ N_A_79_21#_M1000_g N_A_79_21#_c_131_n N_A_79_21#_M1013_g N_A_79_21#_M1002_g
+ N_A_79_21#_c_132_n N_A_79_21#_M1014_g N_A_79_21#_M1003_g N_A_79_21#_c_133_n
+ N_A_79_21#_M1017_g N_A_79_21#_M1004_g N_A_79_21#_c_134_n N_A_79_21#_M1021_g
+ N_A_79_21#_M1019_g N_A_79_21#_c_135_n N_A_79_21#_M1026_g N_A_79_21#_M1024_g
+ N_A_79_21#_c_136_n N_A_79_21#_M1027_g N_A_79_21#_M1029_g N_A_79_21#_c_137_n
+ N_A_79_21#_M1031_g N_A_79_21#_M1030_g N_A_79_21#_c_292_p N_A_79_21#_c_138_n
+ N_A_79_21#_c_139_n N_A_79_21#_c_164_p N_A_79_21#_c_339_p N_A_79_21#_c_246_p
+ N_A_79_21#_c_158_p N_A_79_21#_c_196_p N_A_79_21#_c_140_n N_A_79_21#_c_141_n
+ N_A_79_21#_c_142_n N_A_79_21#_c_143_n N_A_79_21#_c_144_n N_A_79_21#_c_145_n
+ N_A_79_21#_c_146_n PM_SKY130_FD_SC_HD__MUX2_8%A_79_21#
x_PM_SKY130_FD_SC_HD__MUX2_8%S N_S_M1005_g N_S_M1010_g N_S_c_400_n N_S_M1011_g
+ N_S_M1033_g N_S_M1023_g N_S_M1012_g N_S_c_411_n N_S_c_401_n N_S_c_436_n
+ N_S_c_439_n N_S_c_440_n N_S_c_402_n N_S_c_403_n N_S_c_415_n N_S_c_416_n S
+ N_S_c_404_n N_S_c_405_n N_S_c_406_n N_S_c_407_n PM_SKY130_FD_SC_HD__MUX2_8%S
x_PM_SKY130_FD_SC_HD__MUX2_8%A1 N_A1_c_560_n N_A1_M1022_g N_A1_c_561_n
+ N_A1_M1032_g N_A1_c_566_n N_A1_M1016_g N_A1_c_567_n N_A1_M1025_g N_A1_c_562_n
+ N_A1_c_563_n A1 N_A1_c_568_n N_A1_c_564_n N_A1_c_607_n
+ PM_SKY130_FD_SC_HD__MUX2_8%A1
x_PM_SKY130_FD_SC_HD__MUX2_8%A0 N_A0_c_659_n N_A0_M1001_g N_A0_c_660_n
+ N_A0_M1020_g N_A0_c_652_n N_A0_M1015_g N_A0_c_653_n N_A0_M1018_g N_A0_c_654_n
+ N_A0_c_676_n N_A0_c_655_n N_A0_c_682_n N_A0_c_656_n N_A0_c_657_n A0
+ N_A0_c_658_n N_A0_c_691_n A0 N_A0_c_692_n PM_SKY130_FD_SC_HD__MUX2_8%A0
x_PM_SKY130_FD_SC_HD__MUX2_8%A_1259_199# N_A_1259_199#_M1023_d
+ N_A_1259_199#_M1012_d N_A_1259_199#_M1006_g N_A_1259_199#_M1007_g
+ N_A_1259_199#_M1028_g N_A_1259_199#_M1008_g N_A_1259_199#_c_777_n
+ N_A_1259_199#_c_770_n N_A_1259_199#_c_786_n N_A_1259_199#_c_789_n
+ N_A_1259_199#_c_771_n N_A_1259_199#_c_772_n N_A_1259_199#_c_790_n
+ N_A_1259_199#_c_824_n N_A_1259_199#_c_895_p N_A_1259_199#_c_828_n
+ N_A_1259_199#_c_791_n N_A_1259_199#_c_905_p N_A_1259_199#_c_832_n
+ N_A_1259_199#_c_881_p N_A_1259_199#_c_835_n N_A_1259_199#_c_773_n
+ N_A_1259_199#_c_774_n PM_SKY130_FD_SC_HD__MUX2_8%A_1259_199#
x_PM_SKY130_FD_SC_HD__MUX2_8%VPWR N_VPWR_M1000_s N_VPWR_M1002_s N_VPWR_M1004_s
+ N_VPWR_M1024_s N_VPWR_M1030_s N_VPWR_M1033_s N_VPWR_M1008_s N_VPWR_c_914_n
+ N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_917_n N_VPWR_c_918_n N_VPWR_c_919_n
+ N_VPWR_c_920_n N_VPWR_c_921_n N_VPWR_c_922_n N_VPWR_c_923_n N_VPWR_c_924_n
+ N_VPWR_c_925_n N_VPWR_c_926_n N_VPWR_c_927_n VPWR N_VPWR_c_928_n
+ N_VPWR_c_929_n N_VPWR_c_930_n N_VPWR_c_931_n N_VPWR_c_913_n N_VPWR_c_933_n
+ N_VPWR_c_934_n N_VPWR_c_935_n PM_SKY130_FD_SC_HD__MUX2_8%VPWR
x_PM_SKY130_FD_SC_HD__MUX2_8%X N_X_M1009_s N_X_M1014_s N_X_M1021_s N_X_M1027_s
+ N_X_M1000_d N_X_M1003_d N_X_M1019_d N_X_M1029_d N_X_c_1120_p N_X_c_1092_n
+ N_X_c_1048_n N_X_c_1052_n N_X_c_1113_p N_X_c_1096_n N_X_c_1056_n N_X_c_1060_n
+ N_X_c_1116_p N_X_c_1100_n N_X_c_1064_n N_X_c_1068_n N_X_c_1119_p N_X_c_1104_n
+ N_X_c_1072_n N_X_c_1073_n N_X_c_1074_n N_X_c_1076_n N_X_c_1078_n N_X_c_1080_n
+ X PM_SKY130_FD_SC_HD__MUX2_8%X
x_PM_SKY130_FD_SC_HD__MUX2_8%A_792_297# N_A_792_297#_M1010_d
+ N_A_792_297#_M1020_d N_A_792_297#_c_1136_n
+ PM_SKY130_FD_SC_HD__MUX2_8%A_792_297#
x_PM_SKY130_FD_SC_HD__MUX2_8%A_1302_297# N_A_1302_297#_M1007_d
+ N_A_1302_297#_M1025_d N_A_1302_297#_c_1149_n
+ PM_SKY130_FD_SC_HD__MUX2_8%A_1302_297#
x_PM_SKY130_FD_SC_HD__MUX2_8%VGND N_VGND_M1009_d N_VGND_M1013_d N_VGND_M1017_d
+ N_VGND_M1026_d N_VGND_M1031_d N_VGND_M1011_s N_VGND_M1028_s N_VGND_c_1163_n
+ N_VGND_c_1164_n N_VGND_c_1165_n N_VGND_c_1166_n N_VGND_c_1167_n
+ N_VGND_c_1168_n N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n
+ N_VGND_c_1172_n N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n
+ N_VGND_c_1176_n VGND N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n
+ N_VGND_c_1180_n N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n
+ N_VGND_c_1184_n PM_SKY130_FD_SC_HD__MUX2_8%VGND
x_PM_SKY130_FD_SC_HD__MUX2_8%A_792_47# N_A_792_47#_M1005_d N_A_792_47#_M1032_s
+ N_A_792_47#_c_1318_n PM_SKY130_FD_SC_HD__MUX2_8%A_792_47#
x_PM_SKY130_FD_SC_HD__MUX2_8%A_1302_47# N_A_1302_47#_M1006_d
+ N_A_1302_47#_M1018_d N_A_1302_47#_c_1339_n
+ PM_SKY130_FD_SC_HD__MUX2_8%A_1302_47#
cc_1 VNB N_A_79_21#_c_130_n 0.0210549f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_131_n 0.0157281f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_132_n 0.0157715f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_133_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_134_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=0.995
cc_6 VNB N_A_79_21#_c_135_n 0.0157781f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.995
cc_7 VNB N_A_79_21#_c_136_n 0.0157701f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.995
cc_8 VNB N_A_79_21#_c_137_n 0.0158368f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.995
cc_9 VNB N_A_79_21#_c_138_n 0.00153202f $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=1.075
cc_10 VNB N_A_79_21#_c_139_n 3.30931e-19 $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=1.835
cc_11 VNB N_A_79_21#_c_140_n 9.74472e-19 $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=1.16
cc_12 VNB N_A_79_21#_c_141_n 0.00907575f $X=-0.19 $Y=-0.24 $X2=7.44 $Y2=0.85
cc_13 VNB N_A_79_21#_c_142_n 0.00110822f $X=-0.19 $Y=-0.24 $X2=4.98 $Y2=0.85
cc_14 VNB N_A_79_21#_c_143_n 0.00435351f $X=-0.19 $Y=-0.24 $X2=7.585 $Y2=0.85
cc_15 VNB N_A_79_21#_c_144_n 0.138486f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.17
cc_16 VNB N_A_79_21#_c_145_n 0.00109173f $X=-0.19 $Y=-0.24 $X2=4.835 $Y2=0.72
cc_17 VNB N_A_79_21#_c_146_n 0.00164881f $X=-0.19 $Y=-0.24 $X2=7.585 $Y2=0.72
cc_18 VNB N_S_c_400_n 0.021459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_S_c_401_n 0.0232313f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_20 VNB N_S_c_402_n 0.00364594f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_21 VNB N_S_c_403_n 0.019578f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_22 VNB N_S_c_404_n 0.017751f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=0.56
cc_23 VNB N_S_c_405_n 0.0294018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_S_c_406_n 0.0144623f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.995
cc_25 VNB N_S_c_407_n 0.0226348f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.56
cc_26 VNB N_A1_c_560_n 0.0151572f $X=-0.19 $Y=-0.24 $X2=4.405 $Y2=0.235
cc_27 VNB N_A1_c_561_n 0.0518982f $X=-0.19 $Y=-0.24 $X2=7.925 $Y2=1.485
cc_28 VNB N_A1_c_562_n 0.0109137f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_29 VNB N_A1_c_563_n 0.00217219f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_30 VNB N_A1_c_564_n 0.0584715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A0_c_652_n 0.0160263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A0_c_653_n 0.0183348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A0_c_654_n 0.00232214f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_34 VNB N_A0_c_655_n 0.00253547f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_35 VNB N_A0_c_656_n 0.00397678f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.345
cc_36 VNB N_A0_c_657_n 0.0365893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A0_c_658_n 0.0442265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_1259_199#_c_770_n 0.025781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_39 VNB N_A_1259_199#_c_771_n 0.00123525f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_40 VNB N_A_1259_199#_c_772_n 0.0243306f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_41 VNB N_A_1259_199#_c_773_n 0.0186241f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.345
cc_42 VNB N_A_1259_199#_c_774_n 0.023078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VPWR_c_913_n 0.402575f $X=-0.19 $Y=-0.24 $X2=7.5 $Y2=0.72
cc_44 VNB X 0.00203507f $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=0.805
cc_45 VNB N_VGND_c_1163_n 0.0102396f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_46 VNB N_VGND_c_1164_n 0.0133383f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_47 VNB N_VGND_c_1165_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_48 VNB N_VGND_c_1166_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_49 VNB N_VGND_c_1167_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_50 VNB N_VGND_c_1168_n 0.00267136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1169_n 0.00280471f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.345
cc_52 VNB N_VGND_c_1170_n 0.00280526f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.995
cc_53 VNB N_VGND_c_1171_n 0.011083f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.345
cc_54 VNB N_VGND_c_1172_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.985
cc_55 VNB N_VGND_c_1173_n 0.0109642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1174_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.995
cc_57 VNB N_VGND_c_1175_n 0.0118467f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.56
cc_58 VNB N_VGND_c_1176_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.345
cc_59 VNB N_VGND_c_1177_n 0.0117274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1178_n 0.0561984f $X=-0.19 $Y=-0.24 $X2=3.19 $Y2=1.16
cc_61 VNB N_VGND_c_1179_n 0.0634881f $X=-0.19 $Y=-0.24 $X2=4.54 $Y2=0.72
cc_62 VNB N_VGND_c_1180_n 0.0152743f $X=-0.19 $Y=-0.24 $X2=7.28 $Y2=0.72
cc_63 VNB N_VGND_c_1181_n 0.450172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1182_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=4.835 $Y2=0.85
cc_65 VNB N_VGND_c_1183_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=7.585 $Y2=0.85
cc_66 VNB N_VGND_c_1184_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.17
cc_67 VPB N_A_79_21#_M1000_g 0.0234477f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_68 VPB N_A_79_21#_M1002_g 0.0172197f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_69 VPB N_A_79_21#_M1003_g 0.0172704f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_70 VPB N_A_79_21#_M1004_g 0.0172788f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_71 VPB N_A_79_21#_M1019_g 0.0172788f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_72 VPB N_A_79_21#_M1024_g 0.0172788f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.985
cc_73 VPB N_A_79_21#_M1029_g 0.0172686f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.985
cc_74 VPB N_A_79_21#_M1030_g 0.0172791f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_75 VPB N_A_79_21#_c_139_n 0.00108569f $X=-0.19 $Y=1.305 $X2=3.54 $Y2=1.835
cc_76 VPB N_A_79_21#_c_144_n 0.0320798f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.17
cc_77 VPB N_S_M1010_g 0.0230132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_S_M1033_g 0.0179902f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_79 VPB N_S_M1012_g 0.0237648f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_80 VPB N_S_c_411_n 0.0064904f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_81 VPB N_S_c_401_n 0.00460543f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_82 VPB N_S_c_402_n 0.00318057f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_83 VPB N_S_c_403_n 0.0046518f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_84 VPB N_S_c_415_n 0.0284264f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_85 VPB N_S_c_416_n 0.00137559f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_86 VPB S 0.0130498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_S_c_405_n 0.00644343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_S_c_406_n 0.00494387f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=0.995
cc_89 VPB N_A1_c_561_n 0.0170701f $X=-0.19 $Y=1.305 $X2=7.925 $Y2=1.485
cc_90 VPB N_A1_c_566_n 0.0187456f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A1_c_567_n 0.0141974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A1_c_568_n 0.00157676f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_93 VPB N_A1_c_564_n 0.0154578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A0_c_659_n 0.0191084f $X=-0.19 $Y=1.305 $X2=4.405 $Y2=0.235
cc_95 VPB N_A0_c_660_n 0.0143405f $X=-0.19 $Y=1.305 $X2=7.925 $Y2=1.485
cc_96 VPB N_A0_c_656_n 0.0012601f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.345
cc_97 VPB N_A0_c_657_n 0.0176671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A0_c_658_n 0.0153869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_1259_199#_M1007_g 0.0231172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_1259_199#_M1008_g 0.0189568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_1259_199#_c_777_n 0.00612163f $X=-0.19 $Y=1.305 $X2=0.89
+ $Y2=1.345
cc_102 VPB N_A_1259_199#_c_770_n 0.00623332f $X=-0.19 $Y=1.305 $X2=0.89
+ $Y2=1.985
cc_103 VPB N_A_1259_199#_c_771_n 0.00121743f $X=-0.19 $Y=1.305 $X2=1.31
+ $Y2=1.985
cc_104 VPB N_A_1259_199#_c_772_n 0.00547927f $X=-0.19 $Y=1.305 $X2=1.31
+ $Y2=1.985
cc_105 VPB N_VPWR_c_914_n 0.0102469f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_106 VPB N_VPWR_c_915_n 0.026632f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_107 VPB N_VPWR_c_916_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_108 VPB N_VPWR_c_917_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_109 VPB N_VPWR_c_918_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_110 VPB N_VPWR_c_919_n 0.00267136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_920_n 0.00468906f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.345
cc_112 VPB N_VPWR_c_921_n 0.00276587f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=0.995
cc_113 VPB N_VPWR_c_922_n 0.0124915f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.345
cc_114 VPB N_VPWR_c_923_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.985
cc_115 VPB N_VPWR_c_924_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_925_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=0.995
cc_117 VPB N_VPWR_c_926_n 0.0124915f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=0.56
cc_118 VPB N_VPWR_c_927_n 0.00507168f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.345
cc_119 VPB N_VPWR_c_928_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_929_n 0.0545962f $X=-0.19 $Y=1.305 $X2=3.19 $Y2=1.16
cc_121 VPB N_VPWR_c_930_n 0.0614592f $X=-0.19 $Y=1.305 $X2=4.54 $Y2=0.72
cc_122 VPB N_VPWR_c_931_n 0.0151407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_913_n 0.0477524f $X=-0.19 $Y=1.305 $X2=7.5 $Y2=0.72
cc_124 VPB N_VPWR_c_933_n 0.00436868f $X=-0.19 $Y=1.305 $X2=4.98 $Y2=0.85
cc_125 VPB N_VPWR_c_934_n 0.0032427f $X=-0.19 $Y=1.305 $X2=4.835 $Y2=0.85
cc_126 VPB N_VPWR_c_935_n 0.00507168f $X=-0.19 $Y=1.305 $X2=7.585 $Y2=0.85
cc_127 VPB X 0.00259518f $X=-0.19 $Y=1.305 $X2=3.54 $Y2=0.805
cc_128 N_A_79_21#_c_139_n N_S_M1010_g 0.004594f $X=3.54 $Y=1.835 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_158_p N_S_M1010_g 0.0144f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_144_n N_S_M1010_g 0.0352929f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_141_n N_S_c_400_n 0.00333325f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_158_p N_S_M1033_g 0.0120327f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_138_n N_S_c_411_n 0.00568393f $X=3.54 $Y=1.075 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_139_n N_S_c_411_n 0.0179481f $X=3.54 $Y=1.835 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_164_p N_S_c_411_n 0.0111255f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_140_n N_S_c_411_n 0.013341f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_144_n N_S_c_411_n 6.87836e-19 $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_138_n N_S_c_401_n 5.08741e-19 $X=3.54 $Y=1.075 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_139_n N_S_c_401_n 5.08741e-19 $X=3.54 $Y=1.835 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_164_p N_S_c_401_n 0.00230473f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_158_p N_S_c_401_n 8.37305e-19 $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_140_n N_S_c_401_n 0.00124809f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_144_n N_S_c_401_n 0.0154128f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_144 N_A_79_21#_M1001_s N_S_c_436_n 0.00306754f $X=5.185 $Y=1.485 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_158_p N_S_c_436_n 0.0994837f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_145_n N_S_c_436_n 0.00244587f $X=4.835 $Y=0.72 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_158_p N_S_c_439_n 0.0114121f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_158_p N_S_c_440_n 0.0215806f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_141_n N_S_c_402_n 0.00296505f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_150 N_A_79_21#_c_158_p N_S_c_403_n 8.96773e-19 $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_141_n N_S_c_403_n 8.26873e-19 $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_158_p N_S_c_415_n 0.0261278f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_158_p N_S_c_416_n 0.00207706f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_137_n N_S_c_404_n 0.0201714f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_138_n N_S_c_404_n 0.00392431f $X=3.54 $Y=1.075 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_164_p N_S_c_404_n 0.0121866f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_164_p N_A1_c_560_n 0.00865779f $X=4.75 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_79_21#_c_142_n N_A1_c_560_n 6.97795e-19 $X=4.98 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_79_21#_c_145_n N_A1_c_560_n 0.00100061f $X=4.835 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_79_21#_c_164_p N_A1_c_561_n 0.00758604f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_161 N_A_79_21#_c_142_n N_A1_c_561_n 0.00416495f $X=4.98 $Y=0.85 $X2=0 $Y2=0
cc_162 N_A_79_21#_c_145_n N_A1_c_561_n 0.011863f $X=4.835 $Y=0.72 $X2=0 $Y2=0
cc_163 N_A_79_21#_c_158_p N_A1_c_566_n 0.0108654f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_164 N_A_79_21#_c_158_p N_A1_c_567_n 0.00365224f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_164_p N_A1_c_562_n 0.00666166f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_158_p N_A1_c_562_n 3.3156e-19 $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_196_p N_A1_c_562_n 0.00221421f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_141_n N_A1_c_562_n 0.196389f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_142_n N_A1_c_562_n 0.027636f $X=4.98 $Y=0.85 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_143_n N_A1_c_562_n 0.02766f $X=7.585 $Y=0.85 $X2=0 $Y2=0
cc_171 N_A_79_21#_c_145_n N_A1_c_562_n 8.74703e-19 $X=4.835 $Y=0.72 $X2=0 $Y2=0
cc_172 N_A_79_21#_c_146_n N_A1_c_562_n 8.48533e-19 $X=7.585 $Y=0.72 $X2=0 $Y2=0
cc_173 N_A_79_21#_c_164_p N_A1_c_563_n 0.00542467f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_174 N_A_79_21#_c_164_p N_A1_c_568_n 0.0092174f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_175 N_A_79_21#_c_158_p N_A0_c_659_n 0.0108768f $X=8.06 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_79_21#_c_158_p N_A0_c_660_n 0.0087706f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_177 N_A_79_21#_c_196_p N_A0_c_652_n 0.00263491f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_178 N_A_79_21#_c_141_n N_A0_c_652_n 0.00392968f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_179 N_A_79_21#_c_146_n N_A0_c_652_n 3.8728e-19 $X=7.585 $Y=0.72 $X2=0 $Y2=0
cc_180 N_A_79_21#_c_196_p N_A0_c_653_n 0.0046877f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_181 N_A_79_21#_c_141_n N_A0_c_653_n 4.5949e-19 $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_182 N_A_79_21#_c_143_n N_A0_c_653_n 7.55118e-19 $X=7.585 $Y=0.85 $X2=0 $Y2=0
cc_183 N_A_79_21#_c_146_n N_A0_c_653_n 0.0106473f $X=7.585 $Y=0.72 $X2=0 $Y2=0
cc_184 N_A_79_21#_c_141_n N_A0_c_654_n 0.00933542f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_185 N_A_79_21#_c_142_n N_A0_c_654_n 0.00185586f $X=4.98 $Y=0.85 $X2=0 $Y2=0
cc_186 N_A_79_21#_c_145_n N_A0_c_654_n 0.00536876f $X=4.835 $Y=0.72 $X2=0 $Y2=0
cc_187 N_A_79_21#_c_196_p N_A0_c_676_n 0.0103375f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_188 N_A_79_21#_c_141_n N_A0_c_676_n 0.0362184f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_189 N_A_79_21#_c_143_n N_A0_c_676_n 2.04554e-19 $X=7.585 $Y=0.85 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_141_n N_A0_c_655_n 0.0103849f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_143_n N_A0_c_655_n 0.00118928f $X=7.585 $Y=0.85 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_146_n N_A0_c_655_n 0.00155989f $X=7.585 $Y=0.72 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_141_n N_A0_c_682_n 0.00474837f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_194 N_A_79_21#_c_142_n N_A0_c_682_n 0.00136313f $X=4.98 $Y=0.85 $X2=0 $Y2=0
cc_195 N_A_79_21#_c_145_n N_A0_c_682_n 0.0093695f $X=4.835 $Y=0.72 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_196_p N_A0_c_656_n 0.00373756f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_197 N_A_79_21#_c_141_n N_A0_c_656_n 0.00338508f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_198 N_A_79_21#_c_196_p N_A0_c_657_n 0.00315413f $X=7.5 $Y=0.72 $X2=0 $Y2=0
cc_199 N_A_79_21#_c_141_n N_A0_c_657_n 0.0015376f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_200 N_A_79_21#_c_143_n N_A0_c_657_n 0.00102189f $X=7.585 $Y=0.85 $X2=0 $Y2=0
cc_201 N_A_79_21#_c_141_n N_A0_c_658_n 0.00805385f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_202 N_A_79_21#_c_141_n N_A0_c_691_n 0.0173495f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_203 N_A_79_21#_c_141_n N_A0_c_692_n 0.00667593f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_204 N_A_79_21#_c_158_p N_A_1259_199#_M1007_g 0.014182f $X=8.06 $Y=1.92 $X2=0
+ $Y2=0
cc_205 N_A_79_21#_c_158_p N_A_1259_199#_M1008_g 4.80266e-19 $X=8.06 $Y=1.92
+ $X2=0 $Y2=0
cc_206 N_A_79_21#_c_141_n N_A_1259_199#_c_777_n 0.00128493f $X=7.44 $Y=0.85
+ $X2=0 $Y2=0
cc_207 N_A_79_21#_c_158_p N_A_1259_199#_c_770_n 9.07657e-19 $X=8.06 $Y=1.92
+ $X2=0 $Y2=0
cc_208 N_A_79_21#_c_141_n N_A_1259_199#_c_770_n 0.0027076f $X=7.44 $Y=0.85 $X2=0
+ $Y2=0
cc_209 N_A_79_21#_M1016_s N_A_1259_199#_c_786_n 0.00240193f $X=7.925 $Y=1.485
+ $X2=0 $Y2=0
cc_210 N_A_79_21#_c_158_p N_A_1259_199#_c_786_n 0.0983108f $X=8.06 $Y=1.92 $X2=0
+ $Y2=0
cc_211 N_A_79_21#_c_146_n N_A_1259_199#_c_786_n 0.00278871f $X=7.585 $Y=0.72
+ $X2=0 $Y2=0
cc_212 N_A_79_21#_c_158_p N_A_1259_199#_c_789_n 0.0105851f $X=8.06 $Y=1.92 $X2=0
+ $Y2=0
cc_213 N_A_79_21#_c_158_p N_A_1259_199#_c_790_n 0.00266034f $X=8.06 $Y=1.92
+ $X2=0 $Y2=0
cc_214 N_A_79_21#_c_158_p N_A_1259_199#_c_791_n 0.0033398f $X=8.06 $Y=1.92 $X2=0
+ $Y2=0
cc_215 N_A_79_21#_c_141_n N_A_1259_199#_c_773_n 0.0026463f $X=7.44 $Y=0.85 $X2=0
+ $Y2=0
cc_216 N_A_79_21#_c_139_n N_VPWR_M1030_s 0.00349139f $X=3.54 $Y=1.835 $X2=0
+ $Y2=0
cc_217 N_A_79_21#_c_246_p N_VPWR_M1030_s 0.00104554f $X=3.625 $Y=1.92 $X2=0
+ $Y2=0
cc_218 N_A_79_21#_c_158_p N_VPWR_M1030_s 0.00621781f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_219 N_A_79_21#_c_158_p N_VPWR_M1033_s 0.00573688f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_220 N_A_79_21#_M1000_g N_VPWR_c_915_n 0.0123531f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_79_21#_M1002_g N_VPWR_c_915_n 6.0928e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A_79_21#_M1000_g N_VPWR_c_916_n 6.0901e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_79_21#_M1002_g N_VPWR_c_916_n 0.0101939f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_79_21#_M1003_g N_VPWR_c_916_n 0.0101939f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_79_21#_M1004_g N_VPWR_c_916_n 6.0901e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A_79_21#_M1003_g N_VPWR_c_917_n 6.0901e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_79_21#_M1004_g N_VPWR_c_917_n 0.0101939f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_79_21#_M1019_g N_VPWR_c_917_n 0.0101939f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A_79_21#_M1024_g N_VPWR_c_917_n 6.0901e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A_79_21#_M1019_g N_VPWR_c_918_n 6.0901e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A_79_21#_M1024_g N_VPWR_c_918_n 0.0101939f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A_79_21#_M1029_g N_VPWR_c_918_n 0.0101939f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A_79_21#_M1030_g N_VPWR_c_918_n 6.0901e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_79_21#_M1029_g N_VPWR_c_919_n 5.08801e-19 $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_79_21#_M1030_g N_VPWR_c_919_n 0.00671377f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_c_246_p N_VPWR_c_919_n 0.00660099f $X=3.625 $Y=1.92 $X2=0
+ $Y2=0
cc_237 N_A_79_21#_c_158_p N_VPWR_c_919_n 0.00706171f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_238 N_A_79_21#_c_158_p N_VPWR_c_920_n 0.0122669f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_239 N_A_79_21#_M1003_g N_VPWR_c_922_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_79_21#_M1004_g N_VPWR_c_922_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A_79_21#_M1019_g N_VPWR_c_924_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A_79_21#_M1024_g N_VPWR_c_924_n 0.0046653f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_79_21#_M1029_g N_VPWR_c_926_n 0.0046653f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A_79_21#_M1030_g N_VPWR_c_926_n 0.0046653f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_79_21#_M1000_g N_VPWR_c_928_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A_79_21#_M1002_g N_VPWR_c_928_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_79_21#_c_158_p N_VPWR_c_929_n 0.00420597f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_248 N_A_79_21#_c_158_p N_VPWR_c_930_n 0.00294412f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_249 N_A_79_21#_M1001_s N_VPWR_c_913_n 0.00219239f $X=5.185 $Y=1.485 $X2=0
+ $Y2=0
cc_250 N_A_79_21#_M1016_s N_VPWR_c_913_n 0.00219239f $X=7.925 $Y=1.485 $X2=0
+ $Y2=0
cc_251 N_A_79_21#_M1000_g N_VPWR_c_913_n 0.00789179f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_252 N_A_79_21#_M1002_g N_VPWR_c_913_n 0.00789179f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_253 N_A_79_21#_M1003_g N_VPWR_c_913_n 0.00789179f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_254 N_A_79_21#_M1004_g N_VPWR_c_913_n 0.00789179f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_255 N_A_79_21#_M1019_g N_VPWR_c_913_n 0.00789179f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_79_21#_M1024_g N_VPWR_c_913_n 0.00789179f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_A_79_21#_M1029_g N_VPWR_c_913_n 0.00789179f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_A_79_21#_M1030_g N_VPWR_c_913_n 0.00789179f $X=3.41 $Y=1.985 $X2=0
+ $Y2=0
cc_259 N_A_79_21#_c_246_p N_VPWR_c_913_n 8.86197e-19 $X=3.625 $Y=1.92 $X2=0
+ $Y2=0
cc_260 N_A_79_21#_c_158_p N_VPWR_c_913_n 0.0234588f $X=8.06 $Y=1.92 $X2=0 $Y2=0
cc_261 N_A_79_21#_c_131_n N_X_c_1048_n 0.0140058f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A_79_21#_c_132_n N_X_c_1048_n 0.0117424f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_79_21#_c_292_p N_X_c_1048_n 0.0180804f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_79_21#_c_144_n N_X_c_1048_n 0.00209469f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_265 N_A_79_21#_M1002_g N_X_c_1052_n 0.0165948f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A_79_21#_M1003_g N_X_c_1052_n 0.014911f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A_79_21#_c_292_p N_X_c_1052_n 0.0154322f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_79_21#_c_144_n N_X_c_1052_n 0.00204956f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_269 N_A_79_21#_c_133_n N_X_c_1056_n 0.0117865f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_79_21#_c_134_n N_X_c_1056_n 0.0120311f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_79_21#_c_292_p N_X_c_1056_n 0.026745f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_79_21#_c_144_n N_X_c_1056_n 0.00209469f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_273 N_A_79_21#_M1004_g N_X_c_1060_n 0.0149551f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A_79_21#_M1019_g N_X_c_1060_n 0.0149551f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A_79_21#_c_292_p N_X_c_1060_n 0.0228035f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_79_21#_c_144_n N_X_c_1060_n 0.00204956f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_277 N_A_79_21#_c_135_n N_X_c_1064_n 0.0119869f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_79_21#_c_136_n N_X_c_1064_n 0.011364f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A_79_21#_c_292_p N_X_c_1064_n 0.035502f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_79_21#_c_144_n N_X_c_1064_n 0.00427415f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_281 N_A_79_21#_M1024_g N_X_c_1068_n 0.014911f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A_79_21#_M1029_g N_X_c_1068_n 0.0144787f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A_79_21#_c_292_p N_X_c_1068_n 0.0304885f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_79_21#_c_144_n N_X_c_1068_n 0.00422654f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_285 N_A_79_21#_c_131_n N_X_c_1072_n 0.00146775f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_79_21#_M1002_g N_X_c_1073_n 0.00146775f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A_79_21#_c_292_p N_X_c_1074_n 0.00875702f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_79_21#_c_144_n N_X_c_1074_n 0.00217946f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_289 N_A_79_21#_c_292_p N_X_c_1076_n 0.00768502f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_79_21#_c_144_n N_X_c_1076_n 0.00217698f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_291 N_A_79_21#_c_292_p N_X_c_1078_n 0.00881067f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_79_21#_c_144_n N_X_c_1078_n 0.00218592f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_293 N_A_79_21#_c_292_p N_X_c_1080_n 0.00768502f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_79_21#_c_144_n N_X_c_1080_n 0.00217698f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_295 N_A_79_21#_c_130_n X 0.00306467f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A_79_21#_M1000_g X 0.00385866f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A_79_21#_c_131_n X 0.00328117f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A_79_21#_M1002_g X 0.00412925f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A_79_21#_c_292_p X 0.0130288f $X=3.455 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_79_21#_c_144_n X 0.036294f $X=3.41 $Y=1.17 $X2=0 $Y2=0
cc_301 N_A_79_21#_c_158_p N_A_792_297#_M1010_d 0.0278488f $X=8.06 $Y=1.92
+ $X2=-0.19 $Y2=-0.24
cc_302 N_A_79_21#_c_158_p N_A_792_297#_M1020_d 0.00338684f $X=8.06 $Y=1.92 $X2=0
+ $Y2=0
cc_303 N_A_79_21#_M1001_s N_A_792_297#_c_1136_n 0.00357033f $X=5.185 $Y=1.485
+ $X2=0 $Y2=0
cc_304 N_A_79_21#_c_158_p N_A_792_297#_c_1136_n 0.0780283f $X=8.06 $Y=1.92 $X2=0
+ $Y2=0
cc_305 N_A_79_21#_c_158_p N_A_1302_297#_M1007_d 0.0331645f $X=8.06 $Y=1.92
+ $X2=-0.19 $Y2=-0.24
cc_306 N_A_79_21#_M1016_s N_A_1302_297#_c_1149_n 0.00357033f $X=7.925 $Y=1.485
+ $X2=0 $Y2=0
cc_307 N_A_79_21#_c_158_p N_A_1302_297#_c_1149_n 0.0746945f $X=8.06 $Y=1.92
+ $X2=0 $Y2=0
cc_308 N_A_79_21#_c_138_n N_VGND_M1031_d 9.25699e-19 $X=3.54 $Y=1.075 $X2=0
+ $Y2=0
cc_309 N_A_79_21#_c_164_p N_VGND_M1031_d 0.00593339f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_310 N_A_79_21#_c_339_p N_VGND_M1031_d 8.83574e-19 $X=3.625 $Y=0.72 $X2=0
+ $Y2=0
cc_311 N_A_79_21#_c_130_n N_VGND_c_1164_n 0.00877218f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_312 N_A_79_21#_c_131_n N_VGND_c_1164_n 5.0911e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_A_79_21#_c_130_n N_VGND_c_1165_n 5.08801e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_79_21#_c_131_n N_VGND_c_1165_n 0.00664421f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_315 N_A_79_21#_c_132_n N_VGND_c_1165_n 0.00692315f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_79_21#_c_133_n N_VGND_c_1165_n 5.8955e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_79_21#_c_132_n N_VGND_c_1166_n 5.8955e-19 $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_318 N_A_79_21#_c_133_n N_VGND_c_1166_n 0.00692315f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_319 N_A_79_21#_c_134_n N_VGND_c_1166_n 0.00664421f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_A_79_21#_c_135_n N_VGND_c_1166_n 5.08801e-19 $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_A_79_21#_c_134_n N_VGND_c_1167_n 5.08801e-19 $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_322 N_A_79_21#_c_135_n N_VGND_c_1167_n 0.00664421f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_79_21#_c_136_n N_VGND_c_1167_n 0.00692315f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_79_21#_c_137_n N_VGND_c_1167_n 5.8955e-19 $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_A_79_21#_c_136_n N_VGND_c_1168_n 5.8955e-19 $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_A_79_21#_c_137_n N_VGND_c_1168_n 0.00689993f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_79_21#_c_164_p N_VGND_c_1168_n 0.0097332f $X=4.75 $Y=0.72 $X2=0 $Y2=0
cc_328 N_A_79_21#_c_339_p N_VGND_c_1168_n 0.00924733f $X=3.625 $Y=0.72 $X2=0
+ $Y2=0
cc_329 N_A_79_21#_c_141_n N_VGND_c_1169_n 0.00128242f $X=7.44 $Y=0.85 $X2=0
+ $Y2=0
cc_330 N_A_79_21#_c_132_n N_VGND_c_1171_n 0.00339367f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_331 N_A_79_21#_c_133_n N_VGND_c_1171_n 0.00339367f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_A_79_21#_c_134_n N_VGND_c_1173_n 0.00339367f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_333 N_A_79_21#_c_135_n N_VGND_c_1173_n 0.00339367f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_79_21#_c_136_n N_VGND_c_1175_n 0.00339367f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_A_79_21#_c_137_n N_VGND_c_1175_n 0.0046653f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_A_79_21#_c_130_n N_VGND_c_1177_n 0.0046653f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_337 N_A_79_21#_c_131_n N_VGND_c_1177_n 0.00339367f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A_79_21#_c_164_p N_VGND_c_1178_n 0.00260755f $X=4.75 $Y=0.72 $X2=0
+ $Y2=0
cc_339 N_A_79_21#_M1022_d N_VGND_c_1181_n 0.00219239f $X=4.405 $Y=0.235 $X2=0
+ $Y2=0
cc_340 N_A_79_21#_M1015_s N_VGND_c_1181_n 0.00179951f $X=7.145 $Y=0.235 $X2=0
+ $Y2=0
cc_341 N_A_79_21#_c_130_n N_VGND_c_1181_n 0.00789179f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_342 N_A_79_21#_c_131_n N_VGND_c_1181_n 0.00394406f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A_79_21#_c_132_n N_VGND_c_1181_n 0.00398704f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A_79_21#_c_133_n N_VGND_c_1181_n 0.00398704f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A_79_21#_c_134_n N_VGND_c_1181_n 0.00394406f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_79_21#_c_135_n N_VGND_c_1181_n 0.00394406f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_347 N_A_79_21#_c_136_n N_VGND_c_1181_n 0.00398704f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_348 N_A_79_21#_c_137_n N_VGND_c_1181_n 0.00796766f $X=3.41 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_79_21#_c_164_p N_VGND_c_1181_n 0.00620673f $X=4.75 $Y=0.72 $X2=0
+ $Y2=0
cc_350 N_A_79_21#_c_339_p N_VGND_c_1181_n 8.3983e-19 $X=3.625 $Y=0.72 $X2=0
+ $Y2=0
cc_351 N_A_79_21#_c_141_n N_VGND_c_1181_n 0.112877f $X=7.44 $Y=0.85 $X2=0 $Y2=0
cc_352 N_A_79_21#_c_142_n N_VGND_c_1181_n 0.0146685f $X=4.98 $Y=0.85 $X2=0 $Y2=0
cc_353 N_A_79_21#_c_143_n N_VGND_c_1181_n 0.0146781f $X=7.585 $Y=0.85 $X2=0
+ $Y2=0
cc_354 N_A_79_21#_c_164_p N_A_792_47#_M1005_d 0.00864706f $X=4.75 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_355 N_A_79_21#_c_141_n N_A_792_47#_M1032_s 0.00213562f $X=7.44 $Y=0.85 $X2=0
+ $Y2=0
cc_356 N_A_79_21#_c_142_n N_A_792_47#_M1032_s 8.49639e-19 $X=4.98 $Y=0.85 $X2=0
+ $Y2=0
cc_357 N_A_79_21#_c_145_n N_A_792_47#_M1032_s 0.00268397f $X=4.835 $Y=0.72 $X2=0
+ $Y2=0
cc_358 N_A_79_21#_M1022_d N_A_792_47#_c_1318_n 0.00314285f $X=4.405 $Y=0.235
+ $X2=0 $Y2=0
cc_359 N_A_79_21#_c_164_p N_A_792_47#_c_1318_n 0.0372551f $X=4.75 $Y=0.72 $X2=0
+ $Y2=0
cc_360 N_A_79_21#_c_141_n N_A_792_47#_c_1318_n 0.00376946f $X=7.44 $Y=0.85 $X2=0
+ $Y2=0
cc_361 N_A_79_21#_c_142_n N_A_792_47#_c_1318_n 0.00240796f $X=4.98 $Y=0.85 $X2=0
+ $Y2=0
cc_362 N_A_79_21#_c_145_n N_A_792_47#_c_1318_n 0.00706558f $X=4.835 $Y=0.72
+ $X2=0 $Y2=0
cc_363 N_A_79_21#_c_141_n N_A_1302_47#_M1006_d 8.05638e-19 $X=7.44 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_364 N_A_79_21#_c_143_n N_A_1302_47#_M1018_d 0.0064111f $X=7.585 $Y=0.85 $X2=0
+ $Y2=0
cc_365 N_A_79_21#_c_146_n N_A_1302_47#_M1018_d 0.00669004f $X=7.585 $Y=0.72
+ $X2=0 $Y2=0
cc_366 N_A_79_21#_M1015_s N_A_1302_47#_c_1339_n 0.00306531f $X=7.145 $Y=0.235
+ $X2=0 $Y2=0
cc_367 N_A_79_21#_c_196_p N_A_1302_47#_c_1339_n 0.0167969f $X=7.5 $Y=0.72 $X2=0
+ $Y2=0
cc_368 N_A_79_21#_c_141_n N_A_1302_47#_c_1339_n 0.00450758f $X=7.44 $Y=0.85
+ $X2=0 $Y2=0
cc_369 N_A_79_21#_c_143_n N_A_1302_47#_c_1339_n 0.00241219f $X=7.585 $Y=0.85
+ $X2=0 $Y2=0
cc_370 N_A_79_21#_c_146_n N_A_1302_47#_c_1339_n 0.00710927f $X=7.585 $Y=0.72
+ $X2=0 $Y2=0
cc_371 N_S_c_404_n N_A1_c_560_n 0.0249248f $X=3.882 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_372 N_S_c_411_n N_A1_c_561_n 0.00100109f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_373 N_S_c_401_n N_A1_c_561_n 0.0189371f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_374 N_S_c_436_n N_A1_c_561_n 0.0164287f $X=5.67 $Y=1.58 $X2=0 $Y2=0
cc_375 N_S_c_415_n N_A1_c_566_n 0.00222909f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_376 N_S_c_415_n N_A1_c_567_n 0.0045181f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_377 N_S_c_436_n N_A1_c_562_n 0.0346191f $X=5.67 $Y=1.58 $X2=0 $Y2=0
cc_378 N_S_c_402_n N_A1_c_562_n 0.0187893f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_379 N_S_c_403_n N_A1_c_562_n 0.00108868f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_380 N_S_c_415_n N_A1_c_562_n 0.16206f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_381 N_S_c_416_n N_A1_c_562_n 0.0255809f $X=5.9 $Y=1.53 $X2=0 $Y2=0
cc_382 N_S_c_411_n N_A1_c_563_n 0.00681217f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_383 N_S_c_401_n N_A1_c_563_n 0.00400245f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_384 N_S_c_436_n N_A1_c_563_n 0.00618462f $X=5.67 $Y=1.58 $X2=0 $Y2=0
cc_385 N_S_c_415_n A1 0.0265308f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_386 N_S_c_411_n N_A1_c_568_n 0.0102456f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_387 N_S_c_401_n N_A1_c_568_n 0.00132404f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_388 N_S_c_436_n N_A1_c_568_n 0.0121998f $X=5.67 $Y=1.58 $X2=0 $Y2=0
cc_389 N_S_c_415_n N_A1_c_564_n 0.00154717f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_390 N_S_c_415_n N_A1_c_607_n 0.00258524f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_391 N_S_c_436_n N_A0_c_659_n 0.0127182f $X=5.67 $Y=1.58 $X2=-0.19 $Y2=-0.24
cc_392 N_S_c_436_n N_A0_c_660_n 0.0106341f $X=5.67 $Y=1.58 $X2=0 $Y2=0
cc_393 N_S_c_416_n N_A0_c_660_n 0.00151681f $X=5.9 $Y=1.53 $X2=0 $Y2=0
cc_394 N_S_c_400_n N_A0_c_654_n 0.00327471f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_395 N_S_c_436_n N_A0_c_654_n 0.010462f $X=5.67 $Y=1.58 $X2=0 $Y2=0
cc_396 N_S_c_402_n N_A0_c_654_n 0.0139256f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_397 N_S_c_403_n N_A0_c_654_n 3.12617e-19 $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_398 N_S_c_400_n N_A0_c_676_n 0.00855755f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_399 N_S_c_403_n N_A0_c_676_n 0.00143275f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_400 N_S_c_415_n N_A0_c_656_n 0.00215282f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_401 N_S_c_415_n N_A0_c_657_n 0.00774887f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_402 N_S_M1033_g N_A0_c_658_n 0.046573f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_403 N_S_c_436_n N_A0_c_658_n 0.00260029f $X=5.67 $Y=1.58 $X2=0 $Y2=0
cc_404 N_S_c_402_n N_A0_c_658_n 0.00728079f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_405 N_S_c_403_n N_A0_c_658_n 0.0217853f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_406 N_S_c_402_n N_A0_c_691_n 0.0221807f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_407 N_S_c_400_n N_A0_c_692_n 0.0135864f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_408 N_S_c_403_n N_A0_c_692_n 3.43952e-19 $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_409 S N_A_1259_199#_M1012_d 0.00363235f $X=9.34 $Y=1.445 $X2=0 $Y2=0
cc_410 N_S_c_406_n N_A_1259_199#_M1012_d 0.00383138f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_411 N_S_M1033_g N_A_1259_199#_M1007_g 0.0418025f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_412 N_S_c_440_n N_A_1259_199#_M1007_g 2.38734e-19 $X=5.852 $Y=1.495 $X2=0
+ $Y2=0
cc_413 N_S_c_402_n N_A_1259_199#_M1007_g 6.32827e-19 $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_414 N_S_M1012_g N_A_1259_199#_M1008_g 0.0361345f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_415 N_S_c_415_n N_A_1259_199#_M1008_g 0.00312552f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_416 N_S_c_406_n N_A_1259_199#_M1008_g 3.79247e-19 $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_417 N_S_M1033_g N_A_1259_199#_c_777_n 5.59831e-19 $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_S_c_402_n N_A_1259_199#_c_777_n 0.0209681f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_419 N_S_c_403_n N_A_1259_199#_c_777_n 0.00107715f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_420 N_S_c_415_n N_A_1259_199#_c_777_n 0.0049194f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_421 N_S_c_416_n N_A_1259_199#_c_777_n 2.46737e-19 $X=5.9 $Y=1.53 $X2=0 $Y2=0
cc_422 N_S_c_402_n N_A_1259_199#_c_770_n 0.0011199f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_423 N_S_c_403_n N_A_1259_199#_c_770_n 0.0215254f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_424 N_S_c_415_n N_A_1259_199#_c_770_n 0.00259714f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_425 N_S_c_415_n N_A_1259_199#_c_786_n 0.0905481f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_426 N_S_M1033_g N_A_1259_199#_c_789_n 2.42036e-19 $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_427 N_S_c_440_n N_A_1259_199#_c_789_n 0.00215289f $X=5.852 $Y=1.495 $X2=0
+ $Y2=0
cc_428 N_S_c_415_n N_A_1259_199#_c_789_n 0.00569808f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_429 N_S_c_416_n N_A_1259_199#_c_789_n 2.89971e-19 $X=5.9 $Y=1.53 $X2=0 $Y2=0
cc_430 N_S_M1012_g N_A_1259_199#_c_771_n 0.00112998f $X=9.19 $Y=1.985 $X2=0
+ $Y2=0
cc_431 N_S_c_415_n N_A_1259_199#_c_771_n 0.00868653f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_432 S N_A_1259_199#_c_771_n 2.75926e-19 $X=9.34 $Y=1.445 $X2=0 $Y2=0
cc_433 N_S_c_405_n N_A_1259_199#_c_771_n 0.00113668f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_434 N_S_c_406_n N_A_1259_199#_c_771_n 0.0192071f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_435 N_S_c_407_n N_A_1259_199#_c_771_n 0.0034322f $X=9.275 $Y=0.995 $X2=0
+ $Y2=0
cc_436 N_S_c_415_n N_A_1259_199#_c_772_n 0.00125669f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_437 N_S_c_405_n N_A_1259_199#_c_772_n 0.020416f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_438 N_S_c_406_n N_A_1259_199#_c_772_n 9.97845e-19 $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_439 N_S_M1012_g N_A_1259_199#_c_790_n 0.00341949f $X=9.19 $Y=1.985 $X2=0
+ $Y2=0
cc_440 S N_A_1259_199#_c_824_n 7.47844e-19 $X=9.34 $Y=1.445 $X2=0 $Y2=0
cc_441 N_S_c_405_n N_A_1259_199#_c_824_n 8.95436e-19 $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_442 N_S_c_406_n N_A_1259_199#_c_824_n 0.0189058f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_443 N_S_c_407_n N_A_1259_199#_c_824_n 0.0160113f $X=9.275 $Y=0.995 $X2=0
+ $Y2=0
cc_444 N_S_M1012_g N_A_1259_199#_c_828_n 0.0105158f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_445 N_S_c_415_n N_A_1259_199#_c_828_n 0.0138667f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_446 S N_A_1259_199#_c_828_n 9.16562e-19 $X=9.34 $Y=1.445 $X2=0 $Y2=0
cc_447 N_S_c_406_n N_A_1259_199#_c_828_n 0.00236949f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_448 S N_A_1259_199#_c_832_n 0.00497232f $X=9.34 $Y=1.445 $X2=0 $Y2=0
cc_449 N_S_c_405_n N_A_1259_199#_c_832_n 4.92502e-19 $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_450 N_S_c_406_n N_A_1259_199#_c_832_n 0.0111382f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_451 N_S_M1012_g N_A_1259_199#_c_835_n 0.00200433f $X=9.19 $Y=1.985 $X2=0
+ $Y2=0
cc_452 N_S_c_415_n N_A_1259_199#_c_835_n 0.012197f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_453 S N_A_1259_199#_c_835_n 0.00140336f $X=9.34 $Y=1.445 $X2=0 $Y2=0
cc_454 N_S_c_406_n N_A_1259_199#_c_835_n 0.00362486f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_455 N_S_c_400_n N_A_1259_199#_c_773_n 0.0267415f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_456 N_S_c_407_n N_A_1259_199#_c_774_n 0.0231835f $X=9.275 $Y=0.995 $X2=0
+ $Y2=0
cc_457 N_S_c_415_n N_VPWR_M1033_s 0.00304429f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_458 N_S_c_415_n N_VPWR_M1008_s 0.00244334f $X=9.28 $Y=1.53 $X2=0 $Y2=0
cc_459 N_S_M1010_g N_VPWR_c_919_n 0.00310635f $X=3.885 $Y=1.985 $X2=0 $Y2=0
cc_460 N_S_M1033_g N_VPWR_c_920_n 0.00278284f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_461 N_S_M1012_g N_VPWR_c_921_n 0.00839292f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_462 N_S_M1010_g N_VPWR_c_929_n 0.00434141f $X=3.885 $Y=1.985 $X2=0 $Y2=0
cc_463 N_S_M1033_g N_VPWR_c_929_n 0.00422411f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_464 N_S_M1012_g N_VPWR_c_931_n 0.00339367f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_465 N_S_M1010_g N_VPWR_c_913_n 0.00722426f $X=3.885 $Y=1.985 $X2=0 $Y2=0
cc_466 N_S_M1033_g N_VPWR_c_913_n 0.00591461f $X=5.95 $Y=1.985 $X2=0 $Y2=0
cc_467 N_S_M1012_g N_VPWR_c_913_n 0.00489827f $X=9.19 $Y=1.985 $X2=0 $Y2=0
cc_468 N_S_c_436_n N_A_792_297#_M1010_d 0.030937f $X=5.67 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_469 N_S_c_440_n N_A_792_297#_M1020_d 0.00163f $X=5.852 $Y=1.495 $X2=0 $Y2=0
cc_470 N_S_M1010_g N_A_792_297#_c_1136_n 0.00148617f $X=3.885 $Y=1.985 $X2=0
+ $Y2=0
cc_471 N_S_M1033_g N_A_792_297#_c_1136_n 0.00256562f $X=5.95 $Y=1.985 $X2=0
+ $Y2=0
cc_472 N_S_c_404_n N_VGND_c_1168_n 0.00310635f $X=3.882 $Y=0.995 $X2=0 $Y2=0
cc_473 N_S_c_400_n N_VGND_c_1169_n 0.00423719f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_474 N_S_c_407_n N_VGND_c_1170_n 0.00971505f $X=9.275 $Y=0.995 $X2=0 $Y2=0
cc_475 N_S_c_400_n N_VGND_c_1178_n 0.00422995f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_476 N_S_c_404_n N_VGND_c_1178_n 0.00423128f $X=3.882 $Y=0.995 $X2=0 $Y2=0
cc_477 N_S_c_407_n N_VGND_c_1180_n 0.00340533f $X=9.275 $Y=0.995 $X2=0 $Y2=0
cc_478 N_S_c_400_n N_VGND_c_1181_n 0.00699162f $X=5.95 $Y=0.995 $X2=0 $Y2=0
cc_479 N_S_c_404_n N_VGND_c_1181_n 0.00579719f $X=3.882 $Y=0.995 $X2=0 $Y2=0
cc_480 N_S_c_407_n N_VGND_c_1181_n 0.00499747f $X=9.275 $Y=0.995 $X2=0 $Y2=0
cc_481 N_S_c_404_n N_A_792_47#_c_1318_n 0.00148617f $X=3.882 $Y=0.995 $X2=0
+ $Y2=0
cc_482 N_A1_c_561_n N_A0_c_654_n 0.00443549f $X=4.75 $Y=0.96 $X2=0 $Y2=0
cc_483 N_A1_c_562_n N_A0_c_654_n 0.0131387f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_484 N_A1_c_562_n N_A0_c_676_n 0.00317988f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_485 N_A1_c_561_n N_A0_c_682_n 0.00465662f $X=4.75 $Y=0.96 $X2=0 $Y2=0
cc_486 N_A1_c_562_n N_A0_c_656_n 0.020072f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_487 N_A1_c_564_n N_A0_c_656_n 0.00144174f $X=8.27 $Y=1.202 $X2=0 $Y2=0
cc_488 N_A1_c_562_n N_A0_c_657_n 0.00658252f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_489 A1 N_A0_c_657_n 4.6869e-19 $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_490 N_A1_c_564_n N_A0_c_657_n 0.0239569f $X=8.27 $Y=1.202 $X2=0 $Y2=0
cc_491 N_A1_c_607_n N_A0_c_657_n 0.00234591f $X=8.045 $Y=1.19 $X2=0 $Y2=0
cc_492 N_A1_c_561_n N_A0_c_658_n 0.0237812f $X=4.75 $Y=0.96 $X2=0 $Y2=0
cc_493 N_A1_c_562_n N_A0_c_658_n 0.00806863f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_494 N_A1_c_563_n N_A0_c_658_n 3.81565e-19 $X=4.52 $Y=1.19 $X2=0 $Y2=0
cc_495 N_A1_c_568_n N_A0_c_658_n 0.00170161f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_496 N_A1_c_562_n N_A0_c_691_n 0.00208806f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_497 N_A1_c_567_n N_A_1259_199#_M1008_g 0.0305877f $X=8.27 $Y=1.41 $X2=0 $Y2=0
cc_498 N_A1_c_562_n N_A_1259_199#_c_777_n 0.0114043f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_499 N_A1_c_562_n N_A_1259_199#_c_770_n 0.00301167f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_500 N_A1_c_566_n N_A_1259_199#_c_786_n 0.0138558f $X=7.85 $Y=1.41 $X2=0 $Y2=0
cc_501 N_A1_c_567_n N_A_1259_199#_c_786_n 0.0125443f $X=8.27 $Y=1.41 $X2=0 $Y2=0
cc_502 N_A1_c_562_n N_A_1259_199#_c_786_n 0.00760558f $X=7.9 $Y=1.19 $X2=0 $Y2=0
cc_503 A1 N_A_1259_199#_c_786_n 8.31423e-19 $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_504 N_A1_c_564_n N_A_1259_199#_c_786_n 0.00229962f $X=8.27 $Y=1.202 $X2=0
+ $Y2=0
cc_505 N_A1_c_607_n N_A_1259_199#_c_786_n 0.0169278f $X=8.045 $Y=1.19 $X2=0
+ $Y2=0
cc_506 A1 N_A_1259_199#_c_771_n 0.00119888f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_507 N_A1_c_564_n N_A_1259_199#_c_771_n 0.00241497f $X=8.27 $Y=1.202 $X2=0
+ $Y2=0
cc_508 N_A1_c_607_n N_A_1259_199#_c_771_n 0.00945118f $X=8.045 $Y=1.19 $X2=0
+ $Y2=0
cc_509 N_A1_c_564_n N_A_1259_199#_c_772_n 0.0305877f $X=8.27 $Y=1.202 $X2=0
+ $Y2=0
cc_510 N_A1_c_607_n N_A_1259_199#_c_772_n 0.00109146f $X=8.045 $Y=1.19 $X2=0
+ $Y2=0
cc_511 N_A1_c_567_n N_A_1259_199#_c_790_n 0.00118897f $X=8.27 $Y=1.41 $X2=0
+ $Y2=0
cc_512 N_A1_c_567_n N_A_1259_199#_c_791_n 7.19151e-19 $X=8.27 $Y=1.41 $X2=0
+ $Y2=0
cc_513 N_A1_c_566_n N_VPWR_c_930_n 0.00366111f $X=7.85 $Y=1.41 $X2=0 $Y2=0
cc_514 N_A1_c_567_n N_VPWR_c_930_n 0.00366111f $X=8.27 $Y=1.41 $X2=0 $Y2=0
cc_515 N_A1_c_566_n N_VPWR_c_913_n 0.00665614f $X=7.85 $Y=1.41 $X2=0 $Y2=0
cc_516 N_A1_c_567_n N_VPWR_c_913_n 0.00526729f $X=8.27 $Y=1.41 $X2=0 $Y2=0
cc_517 N_A1_c_566_n N_A_1302_297#_c_1149_n 0.012448f $X=7.85 $Y=1.41 $X2=0 $Y2=0
cc_518 N_A1_c_567_n N_A_1302_297#_c_1149_n 0.00957594f $X=8.27 $Y=1.41 $X2=0
+ $Y2=0
cc_519 N_A1_c_560_n N_VGND_c_1178_n 0.00366111f $X=4.33 $Y=0.96 $X2=0 $Y2=0
cc_520 N_A1_c_561_n N_VGND_c_1178_n 0.00366111f $X=4.75 $Y=0.96 $X2=0 $Y2=0
cc_521 N_A1_c_560_n N_VGND_c_1181_n 0.00532774f $X=4.33 $Y=0.96 $X2=0 $Y2=0
cc_522 N_A1_c_561_n N_VGND_c_1181_n 0.00646315f $X=4.75 $Y=0.96 $X2=0 $Y2=0
cc_523 N_A1_c_560_n N_A_792_47#_c_1318_n 0.00788636f $X=4.33 $Y=0.96 $X2=0 $Y2=0
cc_524 N_A1_c_561_n N_A_792_47#_c_1318_n 0.00783096f $X=4.75 $Y=0.96 $X2=0 $Y2=0
cc_525 N_A1_c_564_n N_A_1302_47#_c_1339_n 0.00256393f $X=8.27 $Y=1.202 $X2=0
+ $Y2=0
cc_526 N_A0_c_676_n N_A_1259_199#_c_777_n 0.0100535f $X=6.725 $Y=0.73 $X2=0
+ $Y2=0
cc_527 N_A0_c_656_n N_A_1259_199#_c_777_n 0.0140592f $X=6.81 $Y=1.16 $X2=0 $Y2=0
cc_528 N_A0_c_657_n N_A_1259_199#_c_777_n 7.08588e-19 $X=7.11 $Y=1.16 $X2=0
+ $Y2=0
cc_529 N_A0_c_676_n N_A_1259_199#_c_770_n 0.00501517f $X=6.725 $Y=0.73 $X2=0
+ $Y2=0
cc_530 N_A0_c_656_n N_A_1259_199#_c_770_n 0.0021229f $X=6.81 $Y=1.16 $X2=0 $Y2=0
cc_531 N_A0_c_657_n N_A_1259_199#_c_770_n 0.0119823f $X=7.11 $Y=1.16 $X2=0 $Y2=0
cc_532 N_A0_c_656_n N_A_1259_199#_c_786_n 0.0216019f $X=6.81 $Y=1.16 $X2=0 $Y2=0
cc_533 N_A0_c_657_n N_A_1259_199#_c_786_n 0.0155054f $X=7.11 $Y=1.16 $X2=0 $Y2=0
cc_534 N_A0_c_652_n N_A_1259_199#_c_773_n 0.0206856f $X=7.07 $Y=0.96 $X2=0 $Y2=0
cc_535 N_A0_c_676_n N_A_1259_199#_c_773_n 0.0116237f $X=6.725 $Y=0.73 $X2=0
+ $Y2=0
cc_536 N_A0_c_655_n N_A_1259_199#_c_773_n 0.0032974f $X=6.81 $Y=0.995 $X2=0
+ $Y2=0
cc_537 N_A0_c_692_n N_A_1259_199#_c_773_n 5.86574e-19 $X=5.89 $Y=0.62 $X2=0
+ $Y2=0
cc_538 N_A0_c_659_n N_VPWR_c_929_n 0.00366111f $X=5.11 $Y=1.41 $X2=0 $Y2=0
cc_539 N_A0_c_660_n N_VPWR_c_929_n 0.00366111f $X=5.53 $Y=1.41 $X2=0 $Y2=0
cc_540 N_A0_c_659_n N_VPWR_c_913_n 0.00665614f $X=5.11 $Y=1.41 $X2=0 $Y2=0
cc_541 N_A0_c_660_n N_VPWR_c_913_n 0.00526729f $X=5.53 $Y=1.41 $X2=0 $Y2=0
cc_542 N_A0_c_659_n N_A_792_297#_c_1136_n 0.012448f $X=5.11 $Y=1.41 $X2=0 $Y2=0
cc_543 N_A0_c_660_n N_A_792_297#_c_1136_n 0.00835778f $X=5.53 $Y=1.41 $X2=0
+ $Y2=0
cc_544 N_A0_c_676_n N_VGND_M1011_s 0.00603121f $X=6.725 $Y=0.73 $X2=0 $Y2=0
cc_545 N_A0_c_652_n N_VGND_c_1169_n 0.00114889f $X=7.07 $Y=0.96 $X2=0 $Y2=0
cc_546 N_A0_c_676_n N_VGND_c_1169_n 0.016507f $X=6.725 $Y=0.73 $X2=0 $Y2=0
cc_547 N_A0_c_676_n N_VGND_c_1178_n 0.00247619f $X=6.725 $Y=0.73 $X2=0 $Y2=0
cc_548 N_A0_c_682_n N_VGND_c_1178_n 0.00385827f $X=5.35 $Y=0.62 $X2=0 $Y2=0
cc_549 N_A0_c_691_n N_VGND_c_1178_n 0.0163503f $X=5.695 $Y=0.62 $X2=0 $Y2=0
cc_550 N_A0_c_652_n N_VGND_c_1179_n 0.00366111f $X=7.07 $Y=0.96 $X2=0 $Y2=0
cc_551 N_A0_c_653_n N_VGND_c_1179_n 0.00366111f $X=7.49 $Y=0.96 $X2=0 $Y2=0
cc_552 N_A0_c_676_n N_VGND_c_1179_n 0.00258949f $X=6.725 $Y=0.73 $X2=0 $Y2=0
cc_553 N_A0_c_652_n N_VGND_c_1181_n 0.00570745f $X=7.07 $Y=0.96 $X2=0 $Y2=0
cc_554 N_A0_c_653_n N_VGND_c_1181_n 0.00646071f $X=7.49 $Y=0.96 $X2=0 $Y2=0
cc_555 N_A0_c_676_n N_VGND_c_1181_n 0.00495678f $X=6.725 $Y=0.73 $X2=0 $Y2=0
cc_556 N_A0_c_682_n N_VGND_c_1181_n 0.00247927f $X=5.35 $Y=0.62 $X2=0 $Y2=0
cc_557 N_A0_c_691_n N_VGND_c_1181_n 0.0084779f $X=5.695 $Y=0.62 $X2=0 $Y2=0
cc_558 N_A0_c_654_n N_A_792_47#_M1032_s 0.00142043f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_559 N_A0_c_682_n N_A_792_47#_M1032_s 0.0102597f $X=5.35 $Y=0.62 $X2=0 $Y2=0
cc_560 N_A0_c_691_n N_A_792_47#_M1032_s 0.0175284f $X=5.695 $Y=0.62 $X2=0 $Y2=0
cc_561 N_A0_c_692_n N_A_792_47#_M1032_s 0.0022425f $X=5.89 $Y=0.62 $X2=0 $Y2=0
cc_562 N_A0_c_682_n N_A_792_47#_c_1318_n 0.00333203f $X=5.35 $Y=0.62 $X2=0 $Y2=0
cc_563 N_A0_c_658_n N_A_792_47#_c_1318_n 0.00256393f $X=5.53 $Y=1.202 $X2=0
+ $Y2=0
cc_564 N_A0_c_676_n N_A_1302_47#_M1006_d 0.00969025f $X=6.725 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_565 N_A0_c_655_n N_A_1302_47#_M1006_d 0.0019707f $X=6.81 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_566 N_A0_c_652_n N_A_1302_47#_c_1339_n 0.0118435f $X=7.07 $Y=0.96 $X2=0 $Y2=0
cc_567 N_A0_c_653_n N_A_1302_47#_c_1339_n 0.00782822f $X=7.49 $Y=0.96 $X2=0
+ $Y2=0
cc_568 N_A0_c_676_n N_A_1302_47#_c_1339_n 0.0203831f $X=6.725 $Y=0.73 $X2=0
+ $Y2=0
cc_569 N_A0_c_656_n N_A_1302_47#_c_1339_n 0.00241368f $X=6.81 $Y=1.16 $X2=0
+ $Y2=0
cc_570 N_A_1259_199#_c_790_n N_VPWR_M1008_s 0.00303355f $X=8.77 $Y=1.915 $X2=0
+ $Y2=0
cc_571 N_A_1259_199#_c_828_n N_VPWR_M1008_s 0.00470892f $X=9.315 $Y=2 $X2=0
+ $Y2=0
cc_572 N_A_1259_199#_c_791_n N_VPWR_M1008_s 3.40655e-19 $X=8.855 $Y=2 $X2=0
+ $Y2=0
cc_573 N_A_1259_199#_c_835_n N_VPWR_M1008_s 0.00162349f $X=8.77 $Y=1.58 $X2=0
+ $Y2=0
cc_574 N_A_1259_199#_M1007_g N_VPWR_c_920_n 0.00691784f $X=6.435 $Y=1.985 $X2=0
+ $Y2=0
cc_575 N_A_1259_199#_M1008_g N_VPWR_c_921_n 0.00417809f $X=8.69 $Y=1.985 $X2=0
+ $Y2=0
cc_576 N_A_1259_199#_c_828_n N_VPWR_c_921_n 0.0174856f $X=9.315 $Y=2 $X2=0 $Y2=0
cc_577 N_A_1259_199#_c_791_n N_VPWR_c_921_n 0.00274045f $X=8.855 $Y=2 $X2=0
+ $Y2=0
cc_578 N_A_1259_199#_M1007_g N_VPWR_c_930_n 0.00422411f $X=6.435 $Y=1.985 $X2=0
+ $Y2=0
cc_579 N_A_1259_199#_M1008_g N_VPWR_c_930_n 0.00455963f $X=8.69 $Y=1.985 $X2=0
+ $Y2=0
cc_580 N_A_1259_199#_c_791_n N_VPWR_c_930_n 0.00190971f $X=8.855 $Y=2 $X2=0
+ $Y2=0
cc_581 N_A_1259_199#_c_828_n N_VPWR_c_931_n 0.00243651f $X=9.315 $Y=2 $X2=0
+ $Y2=0
cc_582 N_A_1259_199#_c_881_p N_VPWR_c_931_n 0.0115924f $X=9.4 $Y=2.3 $X2=0 $Y2=0
cc_583 N_A_1259_199#_M1012_d N_VPWR_c_913_n 0.00368727f $X=9.265 $Y=1.485 $X2=0
+ $Y2=0
cc_584 N_A_1259_199#_M1007_g N_VPWR_c_913_n 0.00738741f $X=6.435 $Y=1.985 $X2=0
+ $Y2=0
cc_585 N_A_1259_199#_M1008_g N_VPWR_c_913_n 0.00715673f $X=8.69 $Y=1.985 $X2=0
+ $Y2=0
cc_586 N_A_1259_199#_c_828_n N_VPWR_c_913_n 0.00546438f $X=9.315 $Y=2 $X2=0
+ $Y2=0
cc_587 N_A_1259_199#_c_791_n N_VPWR_c_913_n 0.00369058f $X=8.855 $Y=2 $X2=0
+ $Y2=0
cc_588 N_A_1259_199#_c_881_p N_VPWR_c_913_n 0.00646745f $X=9.4 $Y=2.3 $X2=0
+ $Y2=0
cc_589 N_A_1259_199#_c_786_n N_A_1302_297#_M1007_d 0.0345215f $X=8.685 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_590 N_A_1259_199#_c_786_n N_A_1302_297#_M1025_d 0.00573593f $X=8.685 $Y=1.58
+ $X2=0 $Y2=0
cc_591 N_A_1259_199#_M1007_g N_A_1302_297#_c_1149_n 0.00282243f $X=6.435
+ $Y=1.985 $X2=0 $Y2=0
cc_592 N_A_1259_199#_M1008_g N_A_1302_297#_c_1149_n 0.00286794f $X=8.69 $Y=1.985
+ $X2=0 $Y2=0
cc_593 N_A_1259_199#_c_786_n N_A_1302_297#_c_1149_n 0.00808849f $X=8.685 $Y=1.58
+ $X2=0 $Y2=0
cc_594 N_A_1259_199#_c_771_n N_VGND_M1028_s 7.32946e-19 $X=8.77 $Y=1.16 $X2=0
+ $Y2=0
cc_595 N_A_1259_199#_c_824_n N_VGND_M1028_s 0.00852769f $X=9.315 $Y=0.73 $X2=0
+ $Y2=0
cc_596 N_A_1259_199#_c_895_p N_VGND_M1028_s 3.60207e-19 $X=8.855 $Y=0.73 $X2=0
+ $Y2=0
cc_597 N_A_1259_199#_c_773_n N_VGND_c_1169_n 0.00846933f $X=6.462 $Y=0.995 $X2=0
+ $Y2=0
cc_598 N_A_1259_199#_c_772_n N_VGND_c_1170_n 2.25622e-19 $X=8.77 $Y=1.16 $X2=0
+ $Y2=0
cc_599 N_A_1259_199#_c_824_n N_VGND_c_1170_n 0.0166668f $X=9.315 $Y=0.73 $X2=0
+ $Y2=0
cc_600 N_A_1259_199#_c_895_p N_VGND_c_1170_n 0.00264959f $X=8.855 $Y=0.73 $X2=0
+ $Y2=0
cc_601 N_A_1259_199#_c_774_n N_VGND_c_1170_n 0.00417809f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_602 N_A_1259_199#_c_895_p N_VGND_c_1179_n 0.00187308f $X=8.855 $Y=0.73 $X2=0
+ $Y2=0
cc_603 N_A_1259_199#_c_773_n N_VGND_c_1179_n 0.00340533f $X=6.462 $Y=0.995 $X2=0
+ $Y2=0
cc_604 N_A_1259_199#_c_774_n N_VGND_c_1179_n 0.00500603f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_605 N_A_1259_199#_c_824_n N_VGND_c_1180_n 0.00237932f $X=9.315 $Y=0.73 $X2=0
+ $Y2=0
cc_606 N_A_1259_199#_c_905_p N_VGND_c_1180_n 0.00905679f $X=9.4 $Y=0.46 $X2=0
+ $Y2=0
cc_607 N_A_1259_199#_M1023_d N_VGND_c_1181_n 0.00372073f $X=9.265 $Y=0.235 $X2=0
+ $Y2=0
cc_608 N_A_1259_199#_c_824_n N_VGND_c_1181_n 0.00547535f $X=9.315 $Y=0.73 $X2=0
+ $Y2=0
cc_609 N_A_1259_199#_c_895_p N_VGND_c_1181_n 0.00367222f $X=8.855 $Y=0.73 $X2=0
+ $Y2=0
cc_610 N_A_1259_199#_c_905_p N_VGND_c_1181_n 0.00629232f $X=9.4 $Y=0.46 $X2=0
+ $Y2=0
cc_611 N_A_1259_199#_c_773_n N_VGND_c_1181_n 0.00426385f $X=6.462 $Y=0.995 $X2=0
+ $Y2=0
cc_612 N_A_1259_199#_c_774_n N_VGND_c_1181_n 0.00966499f $X=8.76 $Y=0.995 $X2=0
+ $Y2=0
cc_613 N_A_1259_199#_c_773_n N_A_1302_47#_c_1339_n 0.00179047f $X=6.462 $Y=0.995
+ $X2=0 $Y2=0
cc_614 N_VPWR_c_913_n N_X_M1000_d 0.00562358f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_615 N_VPWR_c_913_n N_X_M1003_d 0.00562358f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_616 N_VPWR_c_913_n N_X_M1019_d 0.00562358f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_617 N_VPWR_c_913_n N_X_M1029_d 0.00562358f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_618 N_VPWR_c_928_n N_X_c_1092_n 0.0113958f $X=0.935 $Y=2.72 $X2=0 $Y2=0
cc_619 N_VPWR_c_913_n N_X_c_1092_n 0.00646998f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_620 N_VPWR_M1002_s N_X_c_1052_n 0.00362893f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_621 N_VPWR_c_916_n N_X_c_1052_n 0.0170259f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_622 N_VPWR_c_922_n N_X_c_1096_n 0.0113958f $X=1.775 $Y=2.72 $X2=0 $Y2=0
cc_623 N_VPWR_c_913_n N_X_c_1096_n 0.00646998f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_624 N_VPWR_M1004_s N_X_c_1060_n 0.00362893f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_625 N_VPWR_c_917_n N_X_c_1060_n 0.0170259f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_626 N_VPWR_c_924_n N_X_c_1100_n 0.0113958f $X=2.615 $Y=2.72 $X2=0 $Y2=0
cc_627 N_VPWR_c_913_n N_X_c_1100_n 0.00646998f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_628 N_VPWR_M1024_s N_X_c_1068_n 0.00362893f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_629 N_VPWR_c_918_n N_X_c_1068_n 0.0170259f $X=2.78 $Y=2 $X2=0 $Y2=0
cc_630 N_VPWR_c_926_n N_X_c_1104_n 0.0113958f $X=3.455 $Y=2.72 $X2=0 $Y2=0
cc_631 N_VPWR_c_913_n N_X_c_1104_n 0.00646998f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_632 N_VPWR_c_913_n N_A_792_297#_M1010_d 0.00884105f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_633 N_VPWR_c_913_n N_A_792_297#_M1020_d 0.00214367f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_634 N_VPWR_c_929_n N_A_792_297#_c_1136_n 0.0904622f $X=6.075 $Y=2.72 $X2=0
+ $Y2=0
cc_635 N_VPWR_c_913_n N_A_792_297#_c_1136_n 0.0691003f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_636 N_VPWR_c_913_n N_A_1302_297#_M1007_d 0.0104158f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_637 N_VPWR_c_913_n N_A_1302_297#_M1025_d 0.00217615f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_638 N_VPWR_c_920_n N_A_1302_297#_c_1149_n 0.0102747f $X=6.16 $Y=2.34 $X2=0
+ $Y2=0
cc_639 N_VPWR_c_930_n N_A_1302_297#_c_1149_n 0.10129f $X=8.815 $Y=2.72 $X2=0
+ $Y2=0
cc_640 N_VPWR_c_913_n N_A_1302_297#_c_1149_n 0.076797f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_641 N_X_c_1048_n N_VGND_M1013_d 0.00337587f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_642 N_X_c_1056_n N_VGND_M1017_d 0.00337587f $X=2.275 $Y=0.72 $X2=0 $Y2=0
cc_643 N_X_c_1064_n N_VGND_M1026_d 0.00337587f $X=3.115 $Y=0.72 $X2=0 $Y2=0
cc_644 N_X_c_1048_n N_VGND_c_1165_n 0.0159625f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_645 N_X_c_1056_n N_VGND_c_1166_n 0.0159625f $X=2.275 $Y=0.72 $X2=0 $Y2=0
cc_646 N_X_c_1064_n N_VGND_c_1167_n 0.0159625f $X=3.115 $Y=0.72 $X2=0 $Y2=0
cc_647 N_X_c_1048_n N_VGND_c_1171_n 0.00243651f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_648 N_X_c_1113_p N_VGND_c_1171_n 0.00888874f $X=1.52 $Y=0.46 $X2=0 $Y2=0
cc_649 N_X_c_1056_n N_VGND_c_1171_n 0.00243651f $X=2.275 $Y=0.72 $X2=0 $Y2=0
cc_650 N_X_c_1056_n N_VGND_c_1173_n 0.00244309f $X=2.275 $Y=0.72 $X2=0 $Y2=0
cc_651 N_X_c_1116_p N_VGND_c_1173_n 0.0112274f $X=2.36 $Y=0.42 $X2=0 $Y2=0
cc_652 N_X_c_1064_n N_VGND_c_1173_n 0.00244309f $X=3.115 $Y=0.72 $X2=0 $Y2=0
cc_653 N_X_c_1064_n N_VGND_c_1175_n 0.00243651f $X=3.115 $Y=0.72 $X2=0 $Y2=0
cc_654 N_X_c_1119_p N_VGND_c_1175_n 0.00888874f $X=3.2 $Y=0.46 $X2=0 $Y2=0
cc_655 N_X_c_1120_p N_VGND_c_1177_n 0.0113958f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_656 N_X_c_1048_n N_VGND_c_1177_n 0.00194726f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_657 N_X_M1009_s N_VGND_c_1181_n 0.00405782f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_658 N_X_M1014_s N_VGND_c_1181_n 0.00253139f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_659 N_X_M1021_s N_VGND_c_1181_n 0.00249348f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_660 N_X_M1027_s N_VGND_c_1181_n 0.00412751f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_661 N_X_c_1120_p N_VGND_c_1181_n 0.00646998f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_662 N_X_c_1048_n N_VGND_c_1181_n 0.00848151f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_663 N_X_c_1113_p N_VGND_c_1181_n 0.00628881f $X=1.52 $Y=0.46 $X2=0 $Y2=0
cc_664 N_X_c_1056_n N_VGND_c_1181_n 0.00987412f $X=2.275 $Y=0.72 $X2=0 $Y2=0
cc_665 N_X_c_1116_p N_VGND_c_1181_n 0.00643448f $X=2.36 $Y=0.42 $X2=0 $Y2=0
cc_666 N_X_c_1064_n N_VGND_c_1181_n 0.00987412f $X=3.115 $Y=0.72 $X2=0 $Y2=0
cc_667 N_X_c_1119_p N_VGND_c_1181_n 0.00628881f $X=3.2 $Y=0.46 $X2=0 $Y2=0
cc_668 N_X_c_1072_n N_VGND_c_1181_n 0.00148162f $X=0.705 $Y=0.72 $X2=0 $Y2=0
cc_669 N_VGND_c_1181_n N_A_792_47#_M1005_d 0.00237915f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_670 N_VGND_c_1181_n N_A_792_47#_M1032_s 0.00809734f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_671 N_VGND_c_1178_n N_A_792_47#_c_1318_n 0.0523253f $X=6.06 $Y=0 $X2=0 $Y2=0
cc_672 N_VGND_c_1181_n N_A_792_47#_c_1318_n 0.0324524f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_673 N_VGND_c_1181_n N_A_1302_47#_M1006_d 0.00339599f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_674 N_VGND_c_1181_n N_A_1302_47#_M1018_d 0.034326f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_675 N_VGND_c_1169_n N_A_1302_47#_c_1339_n 0.012994f $X=6.225 $Y=0.38 $X2=0
+ $Y2=0
cc_676 N_VGND_c_1179_n N_A_1302_47#_c_1339_n 0.0596907f $X=8.815 $Y=0 $X2=0
+ $Y2=0
cc_677 N_VGND_c_1181_n N_A_1302_47#_c_1339_n 0.023152f $X=9.43 $Y=0 $X2=0 $Y2=0

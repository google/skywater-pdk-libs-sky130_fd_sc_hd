* File: sky130_fd_sc_hd__a211o_2.spice
* Created: Thu Aug 27 13:59:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a211o_2.spice.pex"
.subckt sky130_fd_sc_hd__a211o_2  VNB VPB A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1010 N_X_M1010_d N_A_79_21#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.169 PD=0.93 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1010_d N_A_79_21#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.199875 PD=0.93 PS=1.265 NRD=0.456 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1001 A_348_47# N_A2_M1001_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65 AD=0.13325
+ AS=0.199875 PD=1.06 PS=1.265 NRD=27.684 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1008 N_A_79_21#_M1008_d N_A1_M1008_g A_348_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.13325 PD=1.005 PS=1.06 NRD=0 NRS=27.684 M=1 R=4.33333
+ SA=75001.9 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_A_79_21#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.115375 PD=0.98 PS=1.005 NRD=4.608 NRS=13.836 M=1 R=4.33333
+ SA=75002.4 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_A_79_21#_M1006_d N_C1_M1006_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=4.608 M=1 R=4.33333 SA=75002.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_79_21#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_79_21#_M1005_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_299_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.26 PD=1.39 PS=2.52 NRD=11.8003 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_299_297#_M1003_d N_A1_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.195 PD=1.33 PS=1.39 NRD=8.8453 NRS=9.8303 M=1 R=6.66667
+ SA=75000.7 SB=75001 A=0.15 P=2.3 MULT=1
MM1009 A_585_297# N_B1_M1009_g N_A_299_297#_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.165 PD=1.21 PS=1.33 NRD=9.8303 NRS=0.9653 M=1 R=6.66667
+ SA=75001.2 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1000 N_A_79_21#_M1000_d N_C1_M1000_g A_585_297# VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75001.6 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__a211o_2.spice.SKY130_FD_SC_HD__A211O_2.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdfsbp_1.pex.spice
* Created: Tue Sep  1 19:30:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%SCD 1 2 3 5 6 8 11 13 14
r35 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r36 14 19 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.53
+ $X2=0.215 $Y2=1.16
r37 13 19 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=0.215 $Y=0.85
+ $X2=0.215 $Y2=1.16
r38 9 11 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.32 $Y=1.695
+ $X2=0.47 $Y2=1.695
r39 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=1.695
r40 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=2.165
r41 3 18 87.8413 $w=2.62e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r42 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r43 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.32 $Y=1.62 $X2=0.32
+ $Y2=1.695
r44 1 18 39.0894 $w=2.62e-07 $l=1.68464e-07 $layer=POLY_cond $X=0.32 $Y=1.325
+ $X2=0.327 $Y2=1.16
r45 1 2 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.32 $Y=1.325
+ $X2=0.32 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%SCE 3 5 7 11 15 17 19 20 26 33 34
c103 26 0 1.07953e-19 $X=2.53 $Y=1.19
c104 7 0 1.67072e-19 $X=0.89 $Y=2.165
r105 33 36 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.557 $Y=1.16
+ $X2=2.557 $Y2=1.325
r106 33 35 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.557 $Y=1.16
+ $X2=2.557 $Y2=0.995
r107 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=1.16 $X2=2.535 $Y2=1.16
r108 26 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r109 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.19
+ $X2=0.695 $Y2=1.19
r110 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r111 19 20 1.91213 $w=1.4e-07 $l=1.545e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.84 $Y2=1.19
r112 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.74
+ $Y=1.25 $X2=0.74 $Y2=1.25
r113 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.19
+ $X2=0.695 $Y2=1.19
r114 15 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.64 $Y=0.445
+ $X2=2.64 $Y2=0.995
r115 11 36 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.61 $Y=2.165
+ $X2=2.61 $Y2=1.325
r116 5 30 38.5818 $w=3.27e-07 $l=2.11069e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.785 $Y2=1.25
r117 5 7 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.89 $Y2=2.165
r118 1 30 38.5818 $w=3.27e-07 $l=1.86145e-07 $layer=POLY_cond $X=0.83 $Y=1.085
+ $X2=0.785 $Y2=1.25
r119 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.83 $Y=1.085 $X2=0.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%D 1 3 6 8 9 13
c42 13 0 1.62439e-19 $X=1.25 $Y=0.93
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=0.93 $X2=1.25 $Y2=0.93
r44 9 14 24.6952 $w=2.78e-07 $l=6e-07 $layer=LI1_cond $X=1.195 $Y=1.53 $X2=1.195
+ $Y2=0.93
r45 8 14 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=1.195 $Y=0.85 $X2=1.195
+ $Y2=0.93
r46 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.095
+ $X2=1.25 $Y2=0.93
r47 4 6 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.25 $Y=1.095 $X2=1.25
+ $Y2=2.165
r48 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=0.765
+ $X2=1.25 $Y2=0.93
r49 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.25 $Y=0.765 $X2=1.25
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_319_21# 1 2 9 13 18 19 20 22 32 34
c73 19 0 1.59069e-19 $X=1.95 $Y=1.16
r74 32 34 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=2.395 $Y=1.927
+ $X2=2.4 $Y2=1.927
r75 20 22 12.4283 $w=2.53e-07 $l=2.75e-07 $layer=LI1_cond $X=2.387 $Y=0.715
+ $X2=2.387 $Y2=0.44
r76 19 36 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=1.95 $Y=1.16
+ $X2=1.67 $Y2=1.16
r77 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.16 $X2=1.95 $Y2=1.16
r78 16 32 13.2805 $w=3.13e-07 $l=3.63e-07 $layer=LI1_cond $X=2.032 $Y=1.927
+ $X2=2.395 $Y2=1.927
r79 16 18 20.9848 $w=3.33e-07 $l=6.1e-07 $layer=LI1_cond $X=2.032 $Y=1.77
+ $X2=2.032 $Y2=1.16
r80 15 20 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=2.032 $Y=0.81
+ $X2=2.387 $Y2=0.81
r81 15 18 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.032 $Y=0.905
+ $X2=2.032 $Y2=1.16
r82 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.325
+ $X2=1.67 $Y2=1.16
r83 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.67 $Y=1.325
+ $X2=1.67 $Y2=2.165
r84 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=0.995
+ $X2=1.67 $Y2=1.16
r85 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.67 $Y=0.995 $X2=1.67
+ $Y2=0.445
r86 2 34 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.845 $X2=2.4 $Y2=1.99
r87 1 22 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.235 $X2=2.43 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%CLK 7 8 10 13 15 16 17 18 19 20 26 28
c78 20 0 9.44719e-20 $X=3.45 $Y=1.19
c79 13 0 1.07242e-19 $X=3.58 $Y=0.805
r80 34 41 7.22265 $w=1.8e-07 $l=2.68e-07 $layer=LI1_cond $X=2.995 $Y=1.59
+ $X2=2.995 $Y2=1.322
r81 30 41 0.156496 $w=5.33e-07 $l=7e-09 $layer=LI1_cond $X=3.002 $Y=1.322
+ $X2=2.995 $Y2=1.322
r82 26 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.42
r83 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.09
r84 20 30 9.56863 $w=5.33e-07 $l=4.28e-07 $layer=LI1_cond $X=3.43 $Y=1.322
+ $X2=3.002 $Y2=1.322
r85 20 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.255 $X2=3.43 $Y2=1.255
r86 19 34 17.2525 $w=1.78e-07 $l=2.8e-07 $layer=LI1_cond $X=2.995 $Y=1.87
+ $X2=2.995 $Y2=1.59
r87 18 41 0.111783 $w=5.33e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=1.322
+ $X2=2.995 $Y2=1.322
r88 17 30 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.002 $Y=0.85
+ $X2=3.002 $Y2=1.055
r89 15 16 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.52 $Y=1.62
+ $X2=3.52 $Y2=1.77
r90 15 29 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.49 $Y=1.62 $X2=3.49
+ $Y2=1.42
r91 11 13 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.49 $Y=0.805 $X2=3.58
+ $Y2=0.805
r92 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.58 $Y=0.73 $X2=3.58
+ $Y2=0.805
r93 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.58 $Y=0.73 $X2=3.58
+ $Y2=0.445
r94 7 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.55 $Y=2.165
+ $X2=3.55 $Y2=1.77
r95 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.88 $X2=3.49
+ $Y2=0.805
r96 1 28 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.49 $Y=0.88 $X2=3.49
+ $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_643_369# 1 2 9 13 15 16 18 20 23 27 31 33
+ 36 40 42 43 44 45 47 49 50 54 55 56 57 60 61 63 64 65 66 67 76 80 83 84
c295 84 0 1.78722e-19 $X=5.33 $Y=1.74
c296 80 0 3.22574e-20 $X=3.917 $Y=1.09
c297 76 0 2.00397e-19 $X=7.59 $Y=1.87
c298 66 0 1.66008e-19 $X=7.445 $Y=1.87
c299 64 0 1.42859e-19 $X=5.145 $Y=1.87
c300 61 0 6.90487e-20 $X=8.9 $Y=1.08
r301 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=1.74 $X2=5.33 $Y2=1.74
r302 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=1.87
+ $X2=7.59 $Y2=1.87
r303 73 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r304 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=1.87
+ $X2=3.91 $Y2=1.87
r305 67 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r306 66 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=7.59 $Y2=1.87
r307 66 67 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=5.435 $Y2=1.87
r308 65 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=1.87
+ $X2=3.91 $Y2=1.87
r309 64 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r310 64 65 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=4.055 $Y2=1.87
r311 63 77 6.37042 $w=4.58e-07 $l=2.45e-07 $layer=LI1_cond $X=7.835 $Y=1.725
+ $X2=7.59 $Y2=1.725
r312 61 90 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=8.897 $Y=1.08
+ $X2=8.897 $Y2=0.915
r313 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.9
+ $Y=1.08 $X2=8.9 $Y2=1.08
r314 58 60 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=8.925 $Y=0.895
+ $X2=8.925 $Y2=1.08
r315 56 58 6.85974 $w=2e-07 $l=1.57242e-07 $layer=LI1_cond $X=8.81 $Y=0.795
+ $X2=8.925 $Y2=0.895
r316 56 57 44.6409 $w=1.98e-07 $l=8.05e-07 $layer=LI1_cond $X=8.81 $Y=0.795
+ $X2=8.005 $Y2=0.795
r317 55 88 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.92 $Y=1.16
+ $X2=7.92 $Y2=1.325
r318 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.92
+ $Y=1.16 $X2=7.92 $Y2=1.16
r319 52 63 8.89075 $w=4.6e-07 $l=2.69165e-07 $layer=LI1_cond $X=7.92 $Y=1.495
+ $X2=7.835 $Y2=1.725
r320 52 54 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.92 $Y=1.495
+ $X2=7.92 $Y2=1.16
r321 51 57 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.92 $Y=0.895
+ $X2=8.005 $Y2=0.795
r322 51 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.92 $Y=0.895
+ $X2=7.92 $Y2=1.16
r323 50 81 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.917 $Y=1.255
+ $X2=3.917 $Y2=1.42
r324 50 80 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.917 $Y=1.255
+ $X2=3.917 $Y2=1.09
r325 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.91
+ $Y=1.255 $X2=3.91 $Y2=1.255
r326 47 70 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=3.865 $Y=1.775
+ $X2=3.865 $Y2=1.865
r327 47 49 23.0489 $w=2.58e-07 $l=5.2e-07 $layer=LI1_cond $X=3.865 $Y=1.775
+ $X2=3.865 $Y2=1.255
r328 46 49 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.865 $Y=0.885
+ $X2=3.865 $Y2=1.255
r329 44 46 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.865 $Y2=0.885
r330 44 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.455 $Y2=0.8
r331 42 70 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.735 $Y=1.865
+ $X2=3.865 $Y2=1.865
r332 42 43 19.101 $w=1.78e-07 $l=3.1e-07 $layer=LI1_cond $X=3.735 $Y=1.865
+ $X2=3.425 $Y2=1.865
r333 38 45 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.362 $Y=0.715
+ $X2=3.455 $Y2=0.8
r334 38 40 16.4865 $w=1.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.362 $Y=0.715
+ $X2=3.362 $Y2=0.44
r335 34 43 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.34 $Y=1.955
+ $X2=3.425 $Y2=1.865
r336 34 36 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.34 $Y=1.955
+ $X2=3.34 $Y2=2.16
r337 31 90 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=8.96 $Y=0.445 $X2=8.96
+ $Y2=0.915
r338 27 88 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.86 $Y=2.065
+ $X2=7.86 $Y2=1.325
r339 21 83 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.33 $Y=1.905
+ $X2=5.33 $Y2=1.74
r340 21 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.33 $Y=1.905
+ $X2=5.33 $Y2=2.275
r341 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.94 $Y=0.73
+ $X2=4.94 $Y2=0.445
r342 17 33 5.30422 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=4.075 $Y=0.805
+ $X2=3.992 $Y2=0.805
r343 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.94 $Y2=0.73
r344 16 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.075 $Y2=0.805
r345 13 33 20.4101 $w=1.5e-07 $l=7.88987e-08 $layer=POLY_cond $X=4 $Y=0.73
+ $X2=3.992 $Y2=0.805
r346 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4 $Y=0.73 $X2=4
+ $Y2=0.445
r347 11 33 20.4101 $w=1.5e-07 $l=7.84219e-08 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=3.992 $Y2=0.805
r348 11 80 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=3.985 $Y2=1.09
r349 9 81 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.97 $Y=2.165
+ $X2=3.97 $Y2=1.42
r350 2 36 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.845 $X2=3.34 $Y2=2.16
r351 1 40 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.37 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_809_369# 1 2 8 9 11 13 16 20 22 24 28 35
+ 36 39 42 43 46 49 50 57 66
c182 66 0 8.01298e-20 $X=4.327 $Y=1.09
c183 50 0 9.95379e-21 $X=8.51 $Y=1.19
c184 46 0 3.47594e-20 $X=4.37 $Y=1.19
c185 22 0 5.6211e-20 $X=8.485 $Y=1.905
c186 16 0 9.48056e-20 $X=5.36 $Y=0.445
c187 9 0 1.42859e-19 $X=5.285 $Y=1.165
c188 8 0 1.78722e-19 $X=4.615 $Y=1.84
r189 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.505
+ $Y=1.74 $X2=8.505 $Y2=1.74
r190 56 57 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.615 $Y=1.255
+ $X2=4.69 $Y2=1.255
r191 53 56 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.405 $Y=1.255
+ $X2=4.615 $Y2=1.255
r192 50 60 27.5584 $w=2.28e-07 $l=5.5e-07 $layer=LI1_cond $X=8.48 $Y=1.19
+ $X2=8.48 $Y2=1.74
r193 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=1.19
+ $X2=8.51 $Y2=1.19
r194 46 67 8.46186 $w=3.23e-07 $l=2.3e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.42
r195 46 66 6.15528 $w=3.23e-07 $l=1e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.09
r196 46 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.255 $X2=4.405 $Y2=1.255
r197 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=1.19
+ $X2=4.37 $Y2=1.19
r198 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=1.19
+ $X2=4.37 $Y2=1.19
r199 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=8.51 $Y2=1.19
r200 42 43 4.76484 $w=1.4e-07 $l=3.85e-06 $layer=MET1_cond $X=8.365 $Y=1.19
+ $X2=4.515 $Y2=1.19
r201 41 66 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.25 $Y=0.585
+ $X2=4.25 $Y2=1.09
r202 39 41 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=4.222 $Y=0.42
+ $X2=4.222 $Y2=0.585
r203 36 67 29.9635 $w=2.73e-07 $l=7.15e-07 $layer=LI1_cond $X=4.302 $Y=2.135
+ $X2=4.302 $Y2=1.42
r204 35 36 6.01906 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.267 $Y=2.3
+ $X2=4.267 $Y2=2.135
r205 26 28 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=4.615 $Y=1.915
+ $X2=4.91 $Y2=1.915
r206 22 59 38.5406 $w=3.17e-07 $l=1.80748e-07 $layer=POLY_cond $X=8.485 $Y=1.905
+ $X2=8.452 $Y2=1.74
r207 22 24 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.485 $Y=1.905
+ $X2=8.485 $Y2=2.275
r208 18 59 38.5406 $w=3.17e-07 $l=2.13787e-07 $layer=POLY_cond $X=8.34 $Y=1.575
+ $X2=8.452 $Y2=1.74
r209 18 20 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=8.34 $Y=1.575
+ $X2=8.34 $Y2=0.555
r210 14 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.36 $Y=1.09
+ $X2=5.36 $Y2=0.445
r211 11 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.91 $Y=1.99
+ $X2=4.91 $Y2=1.915
r212 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.91 $Y=1.99
+ $X2=4.91 $Y2=2.275
r213 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.285 $Y=1.165
+ $X2=5.36 $Y2=1.09
r214 9 57 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.285 $Y=1.165
+ $X2=4.69 $Y2=1.165
r215 8 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.615 $Y=1.84
+ $X2=4.615 $Y2=1.915
r216 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.615 $Y=1.42
+ $X2=4.615 $Y2=1.255
r217 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.615 $Y=1.42
+ $X2=4.615 $Y2=1.84
r218 2 35 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.845 $X2=4.18 $Y2=2.3
r219 1 39 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.235 $X2=4.21 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_1129_21# 1 2 9 15 19 20 22 24 25 28 32 34
+ 38 44
c97 34 0 4.26244e-20 $X=5.792 $Y=0.72
c98 22 0 4.90363e-20 $X=6.275 $Y=0.72
c99 20 0 5.68782e-20 $X=6.01 $Y=1.74
r100 42 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.84 $Y=1.065
+ $X2=5.84 $Y2=1.575
r101 38 42 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=1.065
r102 38 41 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=0.795
r103 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.81
+ $Y=0.93 $X2=5.81 $Y2=0.93
r104 34 37 6.63049 $w=3.63e-07 $l=2.1e-07 $layer=LI1_cond $X=5.792 $Y=0.72
+ $X2=5.792 $Y2=0.93
r105 30 32 9.64836 $w=2.13e-07 $l=1.8e-07 $layer=LI1_cond $X=6.657 $Y=2.105
+ $X2=6.657 $Y2=2.285
r106 26 28 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=0.635
+ $X2=6.405 $Y2=0.51
r107 24 30 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.55 $Y=2.02
+ $X2=6.657 $Y2=2.105
r108 24 25 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.55 $Y=2.02
+ $X2=6.095 $Y2=2.02
r109 23 34 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=5.975 $Y=0.72
+ $X2=5.792 $Y2=0.72
r110 22 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.275 $Y=0.72
+ $X2=6.405 $Y2=0.635
r111 22 23 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.275 $Y=0.72
+ $X2=5.975 $Y2=0.72
r112 20 45 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.74
+ $X2=5.955 $Y2=1.905
r113 20 44 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.74
+ $X2=5.955 $Y2=1.575
r114 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.01
+ $Y=1.74 $X2=6.01 $Y2=1.74
r115 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.01 $Y=1.935
+ $X2=6.095 $Y2=2.02
r116 17 19 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.01 $Y=1.935
+ $X2=6.01 $Y2=1.74
r117 15 45 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.84 $Y=2.275
+ $X2=5.84 $Y2=1.905
r118 9 41 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.72 $Y=0.445
+ $X2=5.72 $Y2=0.795
r119 2 32 600 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_PDIFF $count=1 $X=6.505
+ $Y=2.065 $X2=6.66 $Y2=2.285
r120 1 28 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.325
+ $Y=0.235 $X2=6.45 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_997_413# 1 2 7 9 12 13 15 18 21 25 29 31
+ 36 38 46 47 49 50 51 55
c152 21 0 1.34667e-19 $X=7.495 $Y=2.065
c153 12 0 4.26244e-20 $X=6.44 $Y=1.095
c154 7 0 1.66008e-19 $X=6.43 $Y=1.365
r155 50 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.44 $Y=1.16
+ $X2=7.44 $Y2=1.325
r156 50 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.44 $Y=1.16
+ $X2=7.44 $Y2=0.995
r157 49 51 4.87734 $w=3.48e-07 $l=1.4e-07 $layer=LI1_cond $X=7.44 $Y=1.15
+ $X2=7.3 $Y2=1.15
r158 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.44
+ $Y=1.16 $X2=7.44 $Y2=1.16
r159 47 51 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=6.435 $Y=1.125
+ $X2=7.3 $Y2=1.125
r160 44 47 3.29018 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.35 $Y=1.185
+ $X2=6.435 $Y2=1.185
r161 44 46 6.95306 $w=4.18e-07 $l=1e-07 $layer=LI1_cond $X=6.35 $Y=1.185
+ $X2=6.25 $Y2=1.185
r162 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.35
+ $Y=1.23 $X2=6.35 $Y2=1.23
r163 38 42 6.20468 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=1.31
+ $X2=5.67 $Y2=1.31
r164 38 46 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.755 $Y=1.31
+ $X2=6.25 $Y2=1.31
r165 35 42 0.18542 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=1.395
+ $X2=5.67 $Y2=1.31
r166 35 36 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.67 $Y=1.395
+ $X2=5.67 $Y2=2.135
r167 31 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.585 $Y=2.3
+ $X2=5.67 $Y2=2.135
r168 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.585 $Y=2.3
+ $X2=5.12 $Y2=2.3
r169 27 42 35.1923 $w=1.56e-07 $l=4.5e-07 $layer=LI1_cond $X=5.22 $Y=1.31
+ $X2=5.67 $Y2=1.31
r170 27 29 21.0845 $w=4.38e-07 $l=8.05e-07 $layer=LI1_cond $X=5.22 $Y=1.225
+ $X2=5.22 $Y2=0.42
r171 23 25 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=6.44 $Y=0.805
+ $X2=6.66 $Y2=0.805
r172 21 56 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.495 $Y=2.065
+ $X2=7.495 $Y2=1.325
r173 18 55 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.495 $Y=0.555
+ $X2=7.495 $Y2=0.995
r174 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.66 $Y=0.73
+ $X2=6.66 $Y2=0.805
r175 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.66 $Y=0.73
+ $X2=6.66 $Y2=0.445
r176 12 45 34.1986 $w=3.29e-07 $l=1.74284e-07 $layer=POLY_cond $X=6.44 $Y=1.095
+ $X2=6.35 $Y2=1.23
r177 11 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.44 $Y=0.88
+ $X2=6.44 $Y2=0.805
r178 11 12 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.44 $Y=0.88
+ $X2=6.44 $Y2=1.095
r179 7 45 34.1986 $w=3.29e-07 $l=1.70367e-07 $layer=POLY_cond $X=6.43 $Y=1.365
+ $X2=6.35 $Y2=1.23
r180 7 9 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=6.43 $Y=1.365
+ $X2=6.43 $Y2=2.275
r181 2 33 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=2.065 $X2=5.12 $Y2=2.3
r182 1 29 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%SET_B 5 9 11 13 16 20 25 27 31 32 34 36 37
+ 43 44 48 50
c147 37 0 1.34667e-19 $X=6.87 $Y=1.53
c148 34 0 4.62344e-20 $X=6.725 $Y=1.53
c149 25 0 1.33399e-19 $X=9.9 $Y=1.835
c150 9 0 4.90363e-20 $X=7.02 $Y=0.445
c151 5 0 1.54163e-19 $X=6.915 $Y=2.275
r152 48 51 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.852 $Y=1.68
+ $X2=6.852 $Y2=1.845
r153 48 50 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.852 $Y=1.68
+ $X2=6.852 $Y2=1.515
r154 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.68 $X2=6.85 $Y2=1.68
r155 44 59 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=8.997 $Y=1.53
+ $X2=8.997 $Y2=1.625
r156 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=1.53
+ $X2=8.97 $Y2=1.53
r157 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.87 $Y=1.53
+ $X2=6.725 $Y2=1.53
r158 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.825 $Y=1.53
+ $X2=8.97 $Y2=1.53
r159 36 37 2.41955 $w=1.4e-07 $l=1.955e-06 $layer=MET1_cond $X=8.825 $Y=1.53
+ $X2=6.87 $Y2=1.53
r160 34 49 4.60977 $w=3.73e-07 $l=1.5e-07 $layer=LI1_cond $X=6.827 $Y=1.53
+ $X2=6.827 $Y2=1.68
r161 34 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.725 $Y=1.53
+ $X2=6.725 $Y2=1.53
r162 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.9
+ $Y=1.61 $X2=9.9 $Y2=1.61
r163 29 59 1.42499 $w=2e-07 $l=1.13e-07 $layer=LI1_cond $X=9.11 $Y=1.625
+ $X2=8.997 $Y2=1.625
r164 29 31 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=9.11 $Y=1.625
+ $X2=9.9 $Y2=1.625
r165 27 32 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=9.9 $Y=1.58 $X2=9.9
+ $Y2=1.61
r166 27 28 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=9.9 $Y=1.58
+ $X2=9.9 $Y2=1.445
r167 25 32 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=9.9 $Y=1.835
+ $X2=9.9 $Y2=1.61
r168 22 25 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=9.57 $Y=1.91
+ $X2=9.9 $Y2=1.91
r169 18 20 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=6.915 $Y=1.29
+ $X2=7.02 $Y2=1.29
r170 16 28 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=9.96 $Y=0.445
+ $X2=9.96 $Y2=1.445
r171 11 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.57 $Y=1.985
+ $X2=9.57 $Y2=1.91
r172 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.57 $Y=1.985
+ $X2=9.57 $Y2=2.275
r173 7 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.02 $Y=1.215
+ $X2=7.02 $Y2=1.29
r174 7 9 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.02 $Y=1.215 $X2=7.02
+ $Y2=0.445
r175 5 51 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.915 $Y=2.275
+ $X2=6.915 $Y2=1.845
r176 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.915 $Y=1.365
+ $X2=6.915 $Y2=1.29
r177 1 50 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.915 $Y=1.365
+ $X2=6.915 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_1770_295# 1 2 9 11 12 15 18 21 22 24 25
+ 28 31 35 37
c101 25 0 6.90487e-20 $X=9.465 $Y=1.27
c102 15 0 1.2016e-19 $X=9.32 $Y=0.445
c103 9 0 9.95379e-21 $X=8.925 $Y=2.275
r104 33 35 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=10.725 $Y=0.397
+ $X2=10.805 $Y2=0.397
r105 31 37 4.14756 $w=2.2e-07 $l=1.03078e-07 $layer=LI1_cond $X=10.805 $Y=1.185
+ $X2=10.765 $Y2=1.27
r106 30 35 3.4259 $w=1.8e-07 $l=1.43e-07 $layer=LI1_cond $X=10.805 $Y=0.54
+ $X2=10.805 $Y2=0.397
r107 30 31 39.7424 $w=1.78e-07 $l=6.45e-07 $layer=LI1_cond $X=10.805 $Y=0.54
+ $X2=10.805 $Y2=1.185
r108 26 37 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=10.765 $Y=1.355
+ $X2=10.765 $Y2=1.27
r109 26 28 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=10.765 $Y=1.355
+ $X2=10.765 $Y2=2.285
r110 24 37 2.28545 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.635 $Y=1.27
+ $X2=10.765 $Y2=1.27
r111 24 25 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=10.635 $Y=1.27
+ $X2=9.465 $Y2=1.27
r112 22 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.38 $Y=1.02
+ $X2=9.38 $Y2=1.185
r113 22 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.38 $Y=1.02
+ $X2=9.38 $Y2=0.855
r114 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.38
+ $Y=1.02 $X2=9.38 $Y2=1.02
r115 19 25 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=9.377 $Y=1.185
+ $X2=9.465 $Y2=1.27
r116 19 21 10.4571 $w=1.73e-07 $l=1.65e-07 $layer=LI1_cond $X=9.377 $Y=1.185
+ $X2=9.377 $Y2=1.02
r117 18 40 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.32 $Y=1.475
+ $X2=9.32 $Y2=1.185
r118 15 39 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.32 $Y=0.445
+ $X2=9.32 $Y2=0.855
r119 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.245 $Y=1.55
+ $X2=9.32 $Y2=1.475
r120 11 12 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=9.245 $Y=1.55
+ $X2=9 $Y2=1.55
r121 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.925 $Y=1.625
+ $X2=9 $Y2=1.55
r122 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=8.925 $Y=1.625
+ $X2=8.925 $Y2=2.275
r123 2 28 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=10.585
+ $Y=2.065 $X2=10.72 $Y2=2.285
r124 1 33 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.235 $X2=10.725 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_1587_329# 1 2 3 12 16 17 19 21 24 26 30
+ 34 37 38 39 40 44 48 51 54 56 58 59 61 65 66 68 72 76
c168 68 0 1.41057e-19 $X=8.85 $Y=1.98
c169 65 0 1.93782e-19 $X=10.38 $Y=1.69
c170 56 0 1.2016e-19 $X=9.825 $Y=0.93
r171 77 78 27.5977 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=10.417 $Y=1.16
+ $X2=10.417 $Y2=1.325
r172 66 78 61.9472 $w=3.4e-07 $l=3.65e-07 $layer=POLY_cond $X=10.415 $Y=1.69
+ $X2=10.415 $Y2=1.325
r173 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.38
+ $Y=1.69 $X2=10.38 $Y2=1.69
r174 63 65 10.7387 $w=2.18e-07 $l=2.05e-07 $layer=LI1_cond $X=10.355 $Y=1.895
+ $X2=10.355 $Y2=1.69
r175 62 72 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=9.91 $Y=1.98
+ $X2=9.802 $Y2=1.98
r176 61 63 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=10.245 $Y=1.98
+ $X2=10.355 $Y2=1.895
r177 61 62 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.245 $Y=1.98
+ $X2=9.91 $Y2=1.98
r178 59 77 38.4695 $w=3.45e-07 $l=2.3e-07 $layer=POLY_cond $X=10.417 $Y=0.93
+ $X2=10.417 $Y2=1.16
r179 59 76 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=10.417 $Y=0.93
+ $X2=10.417 $Y2=0.765
r180 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.38
+ $Y=0.93 $X2=10.38 $Y2=0.93
r181 56 58 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=9.825 $Y=0.93
+ $X2=10.38 $Y2=0.93
r182 52 72 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=9.802 $Y=2.065
+ $X2=9.802 $Y2=1.98
r183 52 54 11.7924 $w=2.13e-07 $l=2.2e-07 $layer=LI1_cond $X=9.802 $Y=2.065
+ $X2=9.802 $Y2=2.285
r184 51 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.74 $Y=0.845
+ $X2=9.825 $Y2=0.93
r185 50 51 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.74 $Y=0.445
+ $X2=9.74 $Y2=0.845
r186 49 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=1.98
+ $X2=8.85 $Y2=1.98
r187 48 72 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=9.695 $Y=1.98
+ $X2=9.802 $Y2=1.98
r188 48 49 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=9.695 $Y=1.98
+ $X2=8.935 $Y2=1.98
r189 44 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.655 $Y=0.36
+ $X2=9.74 $Y2=0.445
r190 44 46 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=9.655 $Y=0.36
+ $X2=8.575 $Y2=0.36
r191 40 68 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=8.85 $Y=2.292
+ $X2=8.85 $Y2=1.98
r192 40 42 18.9207 $w=3.33e-07 $l=5.5e-07 $layer=LI1_cond $X=8.765 $Y=2.292
+ $X2=8.215 $Y2=2.292
r193 36 66 2.54577 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=10.415 $Y=1.705
+ $X2=10.415 $Y2=1.69
r194 36 37 47.1551 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=10.415 $Y=1.705
+ $X2=10.415 $Y2=1.875
r195 32 39 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.395 $Y=1.325
+ $X2=12.395 $Y2=1.16
r196 32 34 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=12.395 $Y=1.325
+ $X2=12.395 $Y2=2.095
r197 28 39 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.395 $Y=0.995
+ $X2=12.395 $Y2=1.16
r198 28 30 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=12.395 $Y=0.995
+ $X2=12.395 $Y2=0.445
r199 27 38 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.53 $Y=1.16
+ $X2=11.455 $Y2=1.16
r200 26 39 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.32 $Y=1.16
+ $X2=12.395 $Y2=1.16
r201 26 27 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=12.32 $Y=1.16
+ $X2=11.53 $Y2=1.16
r202 22 38 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.455 $Y=1.325
+ $X2=11.455 $Y2=1.16
r203 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.455 $Y=1.325
+ $X2=11.455 $Y2=1.985
r204 19 38 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.455 $Y=0.995
+ $X2=11.455 $Y2=1.16
r205 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.455 $Y=0.995
+ $X2=11.455 $Y2=0.56
r206 18 77 3.89586 $w=3.3e-07 $l=1.73e-07 $layer=POLY_cond $X=10.59 $Y=1.16
+ $X2=10.417 $Y2=1.16
r207 17 38 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.38 $Y=1.16
+ $X2=11.455 $Y2=1.16
r208 17 18 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=11.38 $Y=1.16
+ $X2=10.59 $Y2=1.16
r209 16 76 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.515 $Y=0.445
+ $X2=10.515 $Y2=0.765
r210 12 37 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.51 $Y=2.275
+ $X2=10.51 $Y2=1.875
r211 3 54 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=2.065 $X2=9.78 $Y2=2.285
r212 2 42 600 $w=1.7e-07 $l=7.72415e-07 $layer=licon1_PDIFF $count=1 $X=7.935
+ $Y=1.645 $X2=8.215 $Y2=2.29
r213 1 46 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=8.415
+ $Y=0.235 $X2=8.575 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_2412_47# 1 2 9 12 16 20 24 25 27 29
r47 25 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=12.815 $Y=1.16
+ $X2=12.815 $Y2=1.325
r48 25 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=12.815 $Y=1.16
+ $X2=12.815 $Y2=0.995
r49 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.815
+ $Y=1.16 $X2=12.815 $Y2=1.16
r50 22 27 0.221902 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=12.27 $Y=1.16
+ $X2=12.165 $Y2=1.16
r51 22 24 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=12.27 $Y=1.16
+ $X2=12.815 $Y2=1.16
r52 18 27 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=12.165 $Y=1.325
+ $X2=12.165 $Y2=1.16
r53 18 20 31.9524 $w=2.08e-07 $l=6.05e-07 $layer=LI1_cond $X=12.165 $Y=1.325
+ $X2=12.165 $Y2=1.93
r54 14 27 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=12.165 $Y=0.995
+ $X2=12.165 $Y2=1.16
r55 14 16 29.3117 $w=2.08e-07 $l=5.55e-07 $layer=LI1_cond $X=12.165 $Y=0.995
+ $X2=12.165 $Y2=0.44
r56 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.87 $Y=1.985
+ $X2=12.87 $Y2=1.325
r57 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.87 $Y=0.56
+ $X2=12.87 $Y2=0.995
r58 2 20 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=12.06
+ $Y=1.775 $X2=12.185 $Y2=1.93
r59 1 16 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=12.06
+ $Y=0.235 $X2=12.185 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_27_369# 1 2 7 10 11 13 14 16
r48 14 16 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=1.105 $Y=2.36
+ $X2=1.88 $Y2=2.36
r49 13 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.02 $Y=2.255
+ $X2=1.105 $Y2=2.36
r50 12 13 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.02 $Y=2.025
+ $X2=1.02 $Y2=2.255
r51 10 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.935 $Y=1.935
+ $X2=1.02 $Y2=2.025
r52 10 11 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=0.935 $Y=1.935
+ $X2=0.345 $Y2=1.935
r53 7 11 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.345 $Y2=1.935
r54 7 9 2.11154 $w=2.6e-07 $l=4.5e-08 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.215 $Y2=2.07
r55 2 16 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=1.845 $X2=1.88 $Y2=2.34
r56 1 9 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 58 62 65 66 68 69 70 72 81 93 101 106 113 114 117 120 124 128 130 133 136 139
+ 143
c200 114 0 1.05431e-19 $X=13.11 $Y=2.72
c201 34 0 2.10013e-20 $X=2.82 $Y=2.34
r202 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r203 137 140 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.65 $Y2=2.72
r204 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r205 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r206 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r207 126 128 14.2822 $w=6.78e-07 $l=3.7e-07 $layer=LI1_cond $X=7.59 $Y=2.465
+ $X2=7.96 $Y2=2.465
r208 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r209 123 126 7.38754 $w=6.78e-07 $l=4.2e-07 $layer=LI1_cond $X=7.17 $Y=2.465
+ $X2=7.59 $Y2=2.465
r210 123 124 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=2.465
+ $X2=7.005 $Y2=2.465
r211 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r212 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r213 114 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=12.65 $Y2=2.72
r214 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r215 111 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.745 $Y=2.72
+ $X2=12.66 $Y2=2.72
r216 111 113 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.745 $Y=2.72
+ $X2=13.11 $Y2=2.72
r217 110 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r218 110 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=10.35 $Y2=2.72
r219 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r220 107 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.465 $Y=2.72
+ $X2=10.3 $Y2=2.72
r221 107 109 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.465 $Y=2.72
+ $X2=10.81 $Y2=2.72
r222 106 136 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.12 $Y=2.72
+ $X2=11.225 $Y2=2.72
r223 106 109 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.12 $Y=2.72
+ $X2=10.81 $Y2=2.72
r224 105 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r225 105 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r226 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r227 102 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.525 $Y=2.72
+ $X2=9.36 $Y2=2.72
r228 102 104 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.525 $Y=2.72
+ $X2=9.89 $Y2=2.72
r229 101 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.135 $Y=2.72
+ $X2=10.3 $Y2=2.72
r230 101 104 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=10.135 $Y=2.72
+ $X2=9.89 $Y2=2.72
r231 100 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r232 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r233 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r234 97 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r235 96 99 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r236 96 128 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=7.96 $Y2=2.72
r237 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r238 93 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.195 $Y=2.72
+ $X2=9.36 $Y2=2.72
r239 93 99 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.195 $Y=2.72
+ $X2=8.97 $Y2=2.72
r240 92 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r241 91 124 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=7.005 $Y2=2.72
r242 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r243 88 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r244 88 121 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r245 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r246 85 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=3.76 $Y2=2.72
r247 85 87 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r248 84 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r249 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r250 81 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.76 $Y2=2.72
r251 81 83 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.45 $Y2=2.72
r252 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r253 80 118 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=0.69 $Y2=2.72
r254 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r255 77 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.64 $Y2=2.72
r256 77 79 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=2.53 $Y2=2.72
r257 74 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r258 72 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.64 $Y2=2.72
r259 72 74 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r260 70 118 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r261 70 143 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r262 68 87 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=5.75 $Y2=2.72
r263 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=6.11 $Y2=2.72
r264 67 91 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.67 $Y2=2.72
r265 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.11 $Y2=2.72
r266 65 79 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r267 65 66 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.86 $Y2=2.72
r268 64 83 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.03 $Y=2.72
+ $X2=3.45 $Y2=2.72
r269 64 66 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.03 $Y=2.72
+ $X2=2.86 $Y2=2.72
r270 60 139 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.66 $Y=2.635
+ $X2=12.66 $Y2=2.72
r271 60 62 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=12.66 $Y=2.635
+ $X2=12.66 $Y2=1.9
r272 59 136 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.33 $Y=2.72
+ $X2=11.225 $Y2=2.72
r273 58 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.575 $Y=2.72
+ $X2=12.66 $Y2=2.72
r274 58 59 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=12.575 $Y=2.72
+ $X2=11.33 $Y2=2.72
r275 54 57 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=11.225 $Y=1.66
+ $X2=11.225 $Y2=2.34
r276 52 136 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=11.225 $Y=2.635
+ $X2=11.225 $Y2=2.72
r277 52 57 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=11.225 $Y=2.635
+ $X2=11.225 $Y2=2.34
r278 48 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.3 $Y=2.635
+ $X2=10.3 $Y2=2.72
r279 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.3 $Y=2.635
+ $X2=10.3 $Y2=2.34
r280 44 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.36 $Y=2.635
+ $X2=9.36 $Y2=2.72
r281 44 46 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.36 $Y=2.635
+ $X2=9.36 $Y2=2.36
r282 40 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.11 $Y=2.635
+ $X2=6.11 $Y2=2.72
r283 40 42 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.11 $Y=2.635
+ $X2=6.11 $Y2=2.36
r284 36 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=2.635
+ $X2=3.76 $Y2=2.72
r285 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.76 $Y=2.635
+ $X2=3.76 $Y2=2.36
r286 32 66 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=2.635
+ $X2=2.86 $Y2=2.72
r287 32 34 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.86 $Y=2.635
+ $X2=2.86 $Y2=2.34
r288 28 117 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=2.635
+ $X2=0.64 $Y2=2.72
r289 28 30 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.64 $Y=2.635
+ $X2=0.64 $Y2=2.36
r290 9 62 300 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=2 $X=12.47
+ $Y=1.775 $X2=12.66 $Y2=1.9
r291 8 57 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=11.12
+ $Y=1.485 $X2=11.245 $Y2=2.34
r292 8 54 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=11.12
+ $Y=1.485 $X2=11.245 $Y2=1.66
r293 7 50 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=10.175
+ $Y=2.065 $X2=10.3 $Y2=2.34
r294 6 46 600 $w=1.7e-07 $l=4.85592e-07 $layer=licon1_PDIFF $count=1 $X=9
+ $Y=2.065 $X2=9.36 $Y2=2.36
r295 5 123 600 $w=1.7e-07 $l=3.74333e-07 $layer=licon1_PDIFF $count=1 $X=6.99
+ $Y=2.065 $X2=7.17 $Y2=2.36
r296 4 42 600 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_PDIFF $count=1 $X=5.915
+ $Y=2.065 $X2=6.11 $Y2=2.36
r297 3 38 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.845 $X2=3.76 $Y2=2.36
r298 2 34 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.845 $X2=2.82 $Y2=2.34
r299 1 30 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%A_181_47# 1 2 3 4 13 19 21 23 26 31 33 35
+ 36 37 40 43
c139 43 0 3.47594e-20 $X=4.83 $Y=1.53
c140 37 0 1.59069e-19 $X=1.755 $Y=1.53
c141 33 0 1.62439e-19 $X=1.6 $Y=0.705
c142 31 0 1.67072e-19 $X=1.6 $Y=1.87
c143 19 0 9.48056e-20 $X=4.73 $Y=0.42
r144 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.53
+ $X2=4.83 $Y2=1.53
r145 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.53
+ $X2=1.61 $Y2=1.53
r146 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.53
+ $X2=1.61 $Y2=1.53
r147 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.53
+ $X2=4.83 $Y2=1.53
r148 36 37 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=4.685 $Y=1.53
+ $X2=1.755 $Y2=1.53
r149 33 40 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=1.6 $Y=0.705
+ $X2=1.6 $Y2=1.53
r150 33 34 14.2801 $w=2.6e-07 $l=3.14929e-07 $layer=LI1_cond $X=1.6 $Y=0.705
+ $X2=1.537 $Y2=0.42
r151 31 40 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=1.6 $Y=1.87 $X2=1.6
+ $Y2=1.53
r152 28 31 7.57428 $w=2.03e-07 $l=1.4e-07 $layer=LI1_cond $X=1.46 $Y=1.972
+ $X2=1.6 $Y2=1.972
r153 26 44 5.45986 $w=2.62e-07 $l=9.31128e-08 $layer=LI1_cond $X=4.745 $Y=1.445
+ $X2=4.762 $Y2=1.53
r154 26 35 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.745 $Y=1.445
+ $X2=4.745 $Y2=0.92
r155 21 44 4.30723 $w=2.62e-07 $l=1.03899e-07 $layer=LI1_cond $X=4.72 $Y=1.615
+ $X2=4.762 $Y2=1.53
r156 21 23 35.8829 $w=2.18e-07 $l=6.85e-07 $layer=LI1_cond $X=4.72 $Y=1.615
+ $X2=4.72 $Y2=2.3
r157 17 35 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=4.667 $Y=0.758
+ $X2=4.667 $Y2=0.92
r158 17 19 11.9854 $w=3.23e-07 $l=3.38e-07 $layer=LI1_cond $X=4.667 $Y=0.758
+ $X2=4.667 $Y2=0.42
r159 13 34 0.25943 $w=2.8e-07 $l=1.57e-07 $layer=LI1_cond $X=1.38 $Y=0.42
+ $X2=1.537 $Y2=0.42
r160 13 15 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.38 $Y=0.42
+ $X2=1.04 $Y2=0.42
r161 4 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=4.575
+ $Y=2.065 $X2=4.7 $Y2=2.3
r162 3 28 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=1.845 $X2=1.46 $Y2=1.97
r163 2 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.605
+ $Y=0.235 $X2=4.73 $Y2=0.42
r164 1 15 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=0.905
+ $Y=0.235 $X2=1.04 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%Q_N 1 2 7 8 9 10 11 12 20
r18 12 37 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=11.665 $Y=2.21
+ $X2=11.665 $Y2=2.335
r19 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.665 $Y=1.87
+ $X2=11.665 $Y2=2.21
r20 11 31 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=11.665 $Y=1.87
+ $X2=11.665 $Y2=1.655
r21 10 31 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=11.665 $Y=1.53
+ $X2=11.665 $Y2=1.655
r22 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.665 $Y=1.19
+ $X2=11.665 $Y2=1.53
r23 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.665 $Y=0.85
+ $X2=11.665 $Y2=1.19
r24 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.665 $Y=0.51
+ $X2=11.665 $Y2=0.85
r25 7 20 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=11.665 $Y=0.51
+ $X2=11.665 $Y2=0.38
r26 2 37 400 $w=1.7e-07 $l=9.15014e-07 $layer=licon1_PDIFF $count=1 $X=11.53
+ $Y=1.485 $X2=11.665 $Y2=2.335
r27 2 31 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=11.53
+ $Y=1.485 $X2=11.665 $Y2=1.655
r28 1 20 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=11.53
+ $Y=0.235 $X2=11.665 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%Q 1 2 7 8 9 10 11 12 23 30 46
r22 46 47 3.56481 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=13.085 $Y=1.53
+ $X2=13.085 $Y2=1.495
r23 35 50 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=13.085 $Y=1.665
+ $X2=13.085 $Y2=1.66
r24 30 44 1.49877 $w=1.83e-07 $l=2.5e-08 $layer=LI1_cond $X=13.162 $Y=0.85
+ $X2=13.162 $Y2=0.825
r25 12 41 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=13.085 $Y=2.21
+ $X2=13.085 $Y2=2.34
r26 11 12 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=13.085 $Y=1.87
+ $X2=13.085 $Y2=2.21
r27 11 35 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=13.085 $Y=1.87
+ $X2=13.085 $Y2=1.665
r28 10 50 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=13.085 $Y=1.555
+ $X2=13.085 $Y2=1.66
r29 10 46 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=13.085 $Y=1.555
+ $X2=13.085 $Y2=1.53
r30 10 47 1.49877 $w=1.83e-07 $l=2.5e-08 $layer=LI1_cond $X=13.162 $Y=1.47
+ $X2=13.162 $Y2=1.495
r31 9 10 16.7862 $w=1.83e-07 $l=2.8e-07 $layer=LI1_cond $X=13.162 $Y=1.19
+ $X2=13.162 $Y2=1.47
r32 8 44 3.39533 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=13.085 $Y=0.795
+ $X2=13.085 $Y2=0.825
r33 8 21 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=13.085 $Y=0.795
+ $X2=13.085 $Y2=0.655
r34 8 9 18.5848 $w=1.83e-07 $l=3.1e-07 $layer=LI1_cond $X=13.162 $Y=0.88
+ $X2=13.162 $Y2=1.19
r35 8 30 1.79853 $w=1.83e-07 $l=3e-08 $layer=LI1_cond $X=13.162 $Y=0.88
+ $X2=13.162 $Y2=0.85
r36 7 21 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=13.085 $Y=0.51
+ $X2=13.085 $Y2=0.655
r37 7 23 3.72849 $w=3.38e-07 $l=1.1e-07 $layer=LI1_cond $X=13.085 $Y=0.51
+ $X2=13.085 $Y2=0.4
r38 2 50 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=12.945
+ $Y=1.485 $X2=13.08 $Y2=1.66
r39 2 41 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.945
+ $Y=1.485 $X2=13.08 $Y2=2.34
r40 1 23 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=12.945
+ $Y=0.235 $X2=13.08 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSBP_1%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 57 58 60 61 63 64 65 77 81 95 99 106 107 113 125 131 133 136 140
c186 107 0 2.71124e-20 $X=13.11 $Y=0
c187 38 0 4.12131e-20 $X=2.85 $Y=0.38
r188 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r189 133 134 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r190 129 131 10.5001 $w=8.88e-07 $l=4e-08 $layer=LI1_cond $X=7.59 $Y=0.36
+ $X2=7.63 $Y2=0.36
r191 129 130 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r192 127 129 4.93483 $w=8.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.23 $Y=0.36
+ $X2=7.59 $Y2=0.36
r193 124 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r194 123 127 1.37079 $w=8.88e-07 $l=1e-07 $layer=LI1_cond $X=7.13 $Y=0.36
+ $X2=7.23 $Y2=0.36
r195 123 125 15.3664 $w=8.88e-07 $l=3.95e-07 $layer=LI1_cond $X=7.13 $Y=0.36
+ $X2=6.735 $Y2=0.36
r196 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r197 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r198 110 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r199 107 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=12.65 $Y2=0
r200 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r201 104 136 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=12.745 $Y=0
+ $X2=12.642 $Y2=0
r202 104 106 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.745 $Y=0
+ $X2=13.11 $Y2=0
r203 103 137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=12.65 $Y2=0
r204 103 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.27 $Y2=0
r205 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r206 100 133 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.33 $Y=0
+ $X2=11.225 $Y2=0
r207 100 102 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=11.33 $Y=0
+ $X2=12.19 $Y2=0
r208 99 136 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=12.54 $Y=0
+ $X2=12.642 $Y2=0
r209 99 102 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.54 $Y=0
+ $X2=12.19 $Y2=0
r210 98 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r211 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r212 95 133 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.12 $Y=0
+ $X2=11.225 $Y2=0
r213 95 97 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.12 $Y=0
+ $X2=10.81 $Y2=0
r214 94 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r215 94 130 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=7.59 $Y2=0
r216 93 131 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=7.63 $Y2=0
r217 93 94 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r218 90 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r219 90 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=5.75 $Y2=0
r220 89 125 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=6.735 $Y2=0
r221 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r222 87 89 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.67 $Y2=0
r223 85 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r224 85 114 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=3.91 $Y2=0
r225 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r226 82 113 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.94 $Y=0
+ $X2=3.785 $Y2=0
r227 82 84 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.94 $Y=0 $X2=5.29
+ $Y2=0
r228 81 120 9.37134 $w=4.83e-07 $l=3.8e-07 $layer=LI1_cond $X=5.852 $Y=0
+ $X2=5.852 $Y2=0.38
r229 81 87 6.96588 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=5.852 $Y=0
+ $X2=6.095 $Y2=0
r230 81 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r231 81 84 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.29
+ $Y2=0
r232 80 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r233 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r234 77 113 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.63 $Y=0
+ $X2=3.785 $Y2=0
r235 77 79 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.63 $Y=0 $X2=3.45
+ $Y2=0
r236 76 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r237 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r238 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r239 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r240 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r241 69 72 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r242 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r243 67 110 5.44567 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r244 67 69 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.69
+ $Y2=0
r245 65 70 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r246 65 140 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r247 63 93 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.22 $Y=0 $X2=9.89
+ $Y2=0
r248 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.22 $Y=0
+ $X2=10.305 $Y2=0
r249 62 97 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.39 $Y=0
+ $X2=10.81 $Y2=0
r250 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=0
+ $X2=10.305 $Y2=0
r251 60 75 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.53
+ $Y2=0
r252 60 61 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.86
+ $Y2=0
r253 59 79 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.45
+ $Y2=0
r254 59 61 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.86
+ $Y2=0
r255 57 72 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=1.61 $Y2=0
r256 57 58 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.915
+ $Y2=0
r257 56 75 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.53 $Y2=0
r258 56 58 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.915
+ $Y2=0
r259 52 136 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=12.642 $Y=0.085
+ $X2=12.642 $Y2=0
r260 52 54 18.6652 $w=2.03e-07 $l=3.45e-07 $layer=LI1_cond $X=12.642 $Y=0.085
+ $X2=12.642 $Y2=0.43
r261 48 133 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=11.225 $Y=0.085
+ $X2=11.225 $Y2=0
r262 48 50 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=11.225 $Y=0.085
+ $X2=11.225 $Y2=0.38
r263 44 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=0.085
+ $X2=10.305 $Y2=0
r264 44 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.305 $Y=0.085
+ $X2=10.305 $Y2=0.36
r265 40 113 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0
r266 40 42 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.785 $Y=0.085
+ $X2=3.785 $Y2=0.36
r267 36 61 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r268 36 38 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.38
r269 32 58 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=0.085
+ $X2=1.915 $Y2=0
r270 32 34 18.1768 $w=1.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.915 $Y=0.085
+ $X2=1.915 $Y2=0.38
r271 28 110 2.88167 $w=3.95e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.282 $Y=0.085
+ $X2=0.24 $Y2=0
r272 28 30 10.0656 $w=3.93e-07 $l=3.45e-07 $layer=LI1_cond $X=0.282 $Y=0.085
+ $X2=0.282 $Y2=0.43
r273 9 54 182 $w=1.7e-07 $l=2.73998e-07 $layer=licon1_NDIFF $count=1 $X=12.47
+ $Y=0.235 $X2=12.66 $Y2=0.43
r274 8 50 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=11.12
+ $Y=0.235 $X2=11.245 $Y2=0.38
r275 7 46 182 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_NDIFF $count=1 $X=10.035
+ $Y=0.235 $X2=10.305 $Y2=0.36
r276 6 127 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.095
+ $Y=0.235 $X2=7.23 $Y2=0.36
r277 5 120 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.235 $X2=5.93 $Y2=0.38
r278 4 42 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.235 $X2=3.79 $Y2=0.36
r279 3 38 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.85 $Y2=0.38
r280 2 34 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=1.745
+ $Y=0.235 $X2=1.91 $Y2=0.38
r281 1 30 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends


* File: sky130_fd_sc_hd__a41oi_4.spice.pex
* Created: Thu Aug 27 14:06:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A41OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 34 50 51
r79 49 50 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r80 47 49 2.98452 $w=3.23e-07 $l=2e-08 $layer=POLY_cond $X=1.29 $Y=1.16 $X2=1.31
+ $Y2=1.16
r81 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.29
+ $Y=1.16 $X2=1.29 $Y2=1.16
r82 45 47 59.6904 $w=3.23e-07 $l=4e-07 $layer=POLY_cond $X=0.89 $Y=1.16 $X2=1.29
+ $Y2=1.16
r83 44 45 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r84 42 44 29.8452 $w=3.23e-07 $l=2e-07 $layer=POLY_cond $X=0.27 $Y=1.16 $X2=0.47
+ $Y2=1.16
r85 34 48 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.61 $Y=1.19 $X2=1.29
+ $Y2=1.19
r86 33 48 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.15 $Y=1.19
+ $X2=1.29 $Y2=1.19
r87 32 33 23.0489 $w=2.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=1.19
+ $X2=1.15 $Y2=1.19
r88 32 57 18.2888 $w=2.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.69 $Y=1.19
+ $X2=0.325 $Y2=1.19
r89 30 31 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=0.215 $Y=1.53
+ $X2=0.215 $Y2=1.87
r90 30 51 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=0.215 $Y=1.53
+ $X2=0.215 $Y2=1.305
r91 29 51 3.48622 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=0.215 $Y=1.19
+ $X2=0.215 $Y2=1.305
r92 29 57 3.33465 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.215 $Y=1.19
+ $X2=0.325 $Y2=1.19
r93 29 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r94 25 50 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r95 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r96 22 50 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r97 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r98 18 49 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r99 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r100 15 49 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r101 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r102 11 45 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r103 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r104 8 45 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r105 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r106 4 44 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r107 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r108 1 44 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r109 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A1 3 5 7 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 47 48
r72 46 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4 $Y=1.16 $X2=4.06
+ $Y2=1.16
r73 46 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4 $Y=1.16
+ $X2=4 $Y2=1.16
r74 44 46 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.64 $Y=1.16 $X2=4
+ $Y2=1.16
r75 43 44 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.22 $Y=1.16
+ $X2=3.64 $Y2=1.16
r76 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.8 $Y=1.16 $X2=3.22
+ $Y2=1.16
r77 40 42 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.64 $Y=1.16 $X2=2.8
+ $Y2=1.16
r78 40 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.64
+ $Y=1.16 $X2=2.64 $Y2=1.16
r79 37 40 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.46 $Y=1.16 $X2=2.64
+ $Y2=1.16
r80 32 47 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.885 $Y=1.16 $X2=4
+ $Y2=1.16
r81 31 32 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=3.425 $Y=1.16
+ $X2=3.885 $Y2=1.16
r82 30 31 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.965 $Y=1.16
+ $X2=3.425 $Y2=1.16
r83 30 41 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=1.16
+ $X2=2.64 $Y2=1.16
r84 29 41 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.505 $Y=1.16
+ $X2=2.64 $Y2=1.16
r85 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.325
+ $X2=4.06 $Y2=1.16
r86 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.06 $Y=1.325
+ $X2=4.06 $Y2=1.985
r87 22 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=0.995
+ $X2=4.06 $Y2=1.16
r88 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.06 $Y=0.995
+ $X2=4.06 $Y2=0.56
r89 18 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.325
+ $X2=3.64 $Y2=1.16
r90 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.64 $Y=1.325
+ $X2=3.64 $Y2=1.985
r91 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=0.995
+ $X2=3.64 $Y2=1.16
r92 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.64 $Y=0.995
+ $X2=3.64 $Y2=0.56
r93 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.325
+ $X2=3.22 $Y2=1.16
r94 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.22 $Y=1.325
+ $X2=3.22 $Y2=1.985
r95 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=0.995
+ $X2=3.22 $Y2=1.16
r96 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.22 $Y=0.995
+ $X2=3.22 $Y2=0.56
r97 5 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=0.995 $X2=2.8
+ $Y2=1.16
r98 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.8 $Y=0.995 $X2=2.8
+ $Y2=0.56
r99 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.325
+ $X2=2.46 $Y2=1.16
r100 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.46 $Y=1.325
+ $X2=2.46 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 38
r72 49 50 13.2725 $w=3.45e-07 $l=9.5e-08 $layer=POLY_cond $X=5.32 $Y=1.17
+ $X2=5.415 $Y2=1.17
r73 48 49 45.4058 $w=3.45e-07 $l=3.25e-07 $layer=POLY_cond $X=4.995 $Y=1.17
+ $X2=5.32 $Y2=1.17
r74 47 48 13.2725 $w=3.45e-07 $l=9.5e-08 $layer=POLY_cond $X=4.9 $Y=1.17
+ $X2=4.995 $Y2=1.17
r75 45 47 15.3681 $w=3.45e-07 $l=1.1e-07 $layer=POLY_cond $X=4.79 $Y=1.17
+ $X2=4.9 $Y2=1.17
r76 43 45 30.0377 $w=3.45e-07 $l=2.15e-07 $layer=POLY_cond $X=4.575 $Y=1.17
+ $X2=4.79 $Y2=1.17
r77 42 43 13.2725 $w=3.45e-07 $l=9.5e-08 $layer=POLY_cond $X=4.48 $Y=1.17
+ $X2=4.575 $Y2=1.17
r78 38 40 57.7042 $w=3.35e-07 $l=3.35e-07 $layer=POLY_cond $X=5.815 $Y=1.177
+ $X2=6.15 $Y2=1.177
r79 33 40 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.15
+ $Y=1.16 $X2=6.15 $Y2=1.16
r80 32 33 22.4459 $w=2.08e-07 $l=4.25e-07 $layer=LI1_cond $X=5.725 $Y=1.18
+ $X2=6.15 $Y2=1.18
r81 31 32 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=5.265 $Y=1.18
+ $X2=5.725 $Y2=1.18
r82 30 31 25.0866 $w=2.08e-07 $l=4.75e-07 $layer=LI1_cond $X=4.79 $Y=1.18
+ $X2=5.265 $Y2=1.18
r83 30 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.79
+ $Y=1.16 $X2=4.79 $Y2=1.16
r84 29 40 2.58377 $w=3.35e-07 $l=1.5e-08 $layer=POLY_cond $X=6.165 $Y=1.177
+ $X2=6.15 $Y2=1.177
r85 25 29 32.3722 $w=3.35e-07 $l=2.02049e-07 $layer=POLY_cond $X=6.24 $Y=1.345
+ $X2=6.165 $Y2=1.177
r86 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.24 $Y=1.345
+ $X2=6.24 $Y2=1.985
r87 22 38 10.4783 $w=3.45e-07 $l=7.84219e-08 $layer=POLY_cond $X=5.74 $Y=1.17
+ $X2=5.815 $Y2=1.177
r88 22 50 45.4058 $w=3.45e-07 $l=3.25e-07 $layer=POLY_cond $X=5.74 $Y=1.17
+ $X2=5.415 $Y2=1.17
r89 22 24 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.74 $Y=1.01 $X2=5.74
+ $Y2=0.56
r90 18 50 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.415 $Y=1.345
+ $X2=5.415 $Y2=1.17
r91 18 20 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.415 $Y=1.345
+ $X2=5.415 $Y2=1.985
r92 15 49 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=1.17
r93 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=0.56
r94 11 48 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.995 $Y=1.345
+ $X2=4.995 $Y2=1.17
r95 11 13 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.995 $Y=1.345
+ $X2=4.995 $Y2=1.985
r96 8 47 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.9 $Y=0.995 $X2=4.9
+ $Y2=1.17
r97 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.9 $Y=0.995 $X2=4.9
+ $Y2=0.56
r98 4 43 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.575 $Y=1.345
+ $X2=4.575 $Y2=1.17
r99 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.575 $Y=1.345
+ $X2=4.575 $Y2=1.985
r100 1 42 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.48 $Y=0.995
+ $X2=4.48 $Y2=1.17
r101 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.48 $Y=0.995
+ $X2=4.48 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 43
r65 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.79
+ $Y=1.16 $X2=7.79 $Y2=1.16
r66 40 42 37.7217 $w=3.45e-07 $l=2.7e-07 $layer=POLY_cond $X=7.52 $Y=1.17
+ $X2=7.79 $Y2=1.17
r67 39 40 58.6783 $w=3.45e-07 $l=4.2e-07 $layer=POLY_cond $X=7.1 $Y=1.17
+ $X2=7.52 $Y2=1.17
r68 37 39 46.1043 $w=3.45e-07 $l=3.3e-07 $layer=POLY_cond $X=6.77 $Y=1.17
+ $X2=7.1 $Y2=1.17
r69 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.77
+ $Y=1.16 $X2=6.77 $Y2=1.16
r70 35 37 12.5739 $w=3.45e-07 $l=9e-08 $layer=POLY_cond $X=6.68 $Y=1.17 $X2=6.77
+ $Y2=1.17
r71 31 43 10.5 $w=2.23e-07 $l=2.05e-07 $layer=LI1_cond $X=7.585 $Y=1.187
+ $X2=7.79 $Y2=1.187
r72 30 31 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=7.125 $Y=1.187
+ $X2=7.585 $Y2=1.187
r73 30 38 18.183 $w=2.23e-07 $l=3.55e-07 $layer=LI1_cond $X=7.125 $Y=1.187
+ $X2=6.77 $Y2=1.187
r74 29 38 5.37807 $w=2.23e-07 $l=1.05e-07 $layer=LI1_cond $X=6.665 $Y=1.187
+ $X2=6.77 $Y2=1.187
r75 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.94 $Y=1.345
+ $X2=7.94 $Y2=1.985
r76 22 25 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.94 $Y=1.17
+ $X2=7.94 $Y2=1.345
r77 22 42 20.9565 $w=3.45e-07 $l=1.5e-07 $layer=POLY_cond $X=7.94 $Y=1.17
+ $X2=7.79 $Y2=1.17
r78 22 24 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.94 $Y=1.01 $X2=7.94
+ $Y2=0.56
r79 18 40 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.52 $Y=1.345
+ $X2=7.52 $Y2=1.17
r80 18 20 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.52 $Y=1.345
+ $X2=7.52 $Y2=1.985
r81 15 40 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.52 $Y=0.995
+ $X2=7.52 $Y2=1.17
r82 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.52 $Y=0.995
+ $X2=7.52 $Y2=0.56
r83 11 39 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.1 $Y=1.345
+ $X2=7.1 $Y2=1.17
r84 11 13 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.1 $Y=1.345 $X2=7.1
+ $Y2=1.985
r85 8 39 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.1 $Y=0.995 $X2=7.1
+ $Y2=1.17
r86 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995 $X2=7.1
+ $Y2=0.56
r87 4 35 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.68 $Y=1.345
+ $X2=6.68 $Y2=1.17
r88 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.68 $Y=1.345 $X2=6.68
+ $Y2=1.985
r89 1 35 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.68 $Y=0.995
+ $X2=6.68 $Y2=1.17
r90 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.68 $Y=0.995 $X2=6.68
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A4 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 43
c67 1 0 1.25206e-19 $X=8.36 $Y=0.995
r68 43 45 28.3529 $w=3.23e-07 $l=1.9e-07 $layer=POLY_cond $X=9.62 $Y=1.16
+ $X2=9.81 $Y2=1.16
r69 42 43 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=9.2 $Y=1.16
+ $X2=9.62 $Y2=1.16
r70 41 42 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=8.78 $Y=1.16
+ $X2=9.2 $Y2=1.16
r71 39 41 49.2446 $w=3.23e-07 $l=3.3e-07 $layer=POLY_cond $X=8.45 $Y=1.16
+ $X2=8.78 $Y2=1.16
r72 37 39 13.4303 $w=3.23e-07 $l=9e-08 $layer=POLY_cond $X=8.36 $Y=1.16 $X2=8.45
+ $Y2=1.16
r73 32 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.81
+ $Y=1.16 $X2=9.81 $Y2=1.16
r74 31 32 20.8293 $w=2.03e-07 $l=3.85e-07 $layer=LI1_cond $X=9.425 $Y=1.177
+ $X2=9.81 $Y2=1.177
r75 30 31 24.8869 $w=2.03e-07 $l=4.6e-07 $layer=LI1_cond $X=8.965 $Y=1.177
+ $X2=9.425 $Y2=1.177
r76 29 30 27.8625 $w=2.03e-07 $l=5.15e-07 $layer=LI1_cond $X=8.45 $Y=1.177
+ $X2=8.965 $Y2=1.177
r77 29 39 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.45
+ $Y=1.16 $X2=8.45 $Y2=1.16
r78 25 43 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.62 $Y=1.325
+ $X2=9.62 $Y2=1.16
r79 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.62 $Y=1.325
+ $X2=9.62 $Y2=1.985
r80 22 43 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.62 $Y=0.995
+ $X2=9.62 $Y2=1.16
r81 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.62 $Y=0.995
+ $X2=9.62 $Y2=0.56
r82 18 42 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.2 $Y=1.325
+ $X2=9.2 $Y2=1.16
r83 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.2 $Y=1.325 $X2=9.2
+ $Y2=1.985
r84 15 42 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.2 $Y=0.995
+ $X2=9.2 $Y2=1.16
r85 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.2 $Y=0.995 $X2=9.2
+ $Y2=0.56
r86 11 41 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.78 $Y=1.325
+ $X2=8.78 $Y2=1.16
r87 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.78 $Y=1.325
+ $X2=8.78 $Y2=1.985
r88 8 41 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.78 $Y=0.995
+ $X2=8.78 $Y2=1.16
r89 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.78 $Y=0.995
+ $X2=8.78 $Y2=0.56
r90 4 37 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.36 $Y=1.325
+ $X2=8.36 $Y2=1.16
r91 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.36 $Y=1.325 $X2=8.36
+ $Y2=1.985
r92 1 37 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.36 $Y=0.995
+ $X2=8.36 $Y2=1.16
r93 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.36 $Y=0.995 $X2=8.36
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A_27_297# 1 2 3 4 5 6 7 8 9 10 11 34 41 42
+ 43 48 50 51 54 56 60 62 66 68 72 74 78 80 84 86 90 95 96 98 100
r119 88 90 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.86 $Y=1.745
+ $X2=9.86 $Y2=1.96
r120 87 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.075 $Y=1.66
+ $X2=8.99 $Y2=1.66
r121 86 88 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.775 $Y=1.66
+ $X2=9.86 $Y2=1.745
r122 86 87 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.775 $Y=1.66
+ $X2=9.075 $Y2=1.66
r123 82 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=1.745
+ $X2=8.99 $Y2=1.66
r124 82 84 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.99 $Y=1.745
+ $X2=8.99 $Y2=1.96
r125 81 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.235 $Y=1.66
+ $X2=8.15 $Y2=1.66
r126 80 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=1.66
+ $X2=8.99 $Y2=1.66
r127 80 81 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.905 $Y=1.66
+ $X2=8.235 $Y2=1.66
r128 76 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.15 $Y=1.745
+ $X2=8.15 $Y2=1.66
r129 76 78 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.15 $Y=1.745
+ $X2=8.15 $Y2=1.96
r130 75 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=1.66
+ $X2=7.31 $Y2=1.66
r131 74 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.065 $Y=1.66
+ $X2=8.15 $Y2=1.66
r132 74 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.065 $Y=1.66
+ $X2=7.395 $Y2=1.66
r133 70 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=1.745
+ $X2=7.31 $Y2=1.66
r134 70 72 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.31 $Y=1.745
+ $X2=7.31 $Y2=1.96
r135 69 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.66
+ $X2=6.47 $Y2=1.66
r136 68 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=1.66
+ $X2=7.31 $Y2=1.66
r137 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.225 $Y=1.66
+ $X2=6.555 $Y2=1.66
r138 64 97 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=1.745
+ $X2=6.47 $Y2=1.66
r139 64 66 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.47 $Y=1.745
+ $X2=6.47 $Y2=1.96
r140 63 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=1.66
+ $X2=5.205 $Y2=1.66
r141 62 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=1.66
+ $X2=6.47 $Y2=1.66
r142 62 63 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=6.385 $Y=1.66
+ $X2=5.29 $Y2=1.66
r143 58 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=1.745
+ $X2=5.205 $Y2=1.66
r144 58 60 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.205 $Y=1.745
+ $X2=5.205 $Y2=1.96
r145 57 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=1.66
+ $X2=4.27 $Y2=1.66
r146 56 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=1.66
+ $X2=5.205 $Y2=1.66
r147 56 57 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.12 $Y=1.66
+ $X2=4.355 $Y2=1.66
r148 52 95 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=1.745
+ $X2=4.27 $Y2=1.66
r149 52 54 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.27 $Y=1.745
+ $X2=4.27 $Y2=2.26
r150 50 95 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=1.66
+ $X2=4.27 $Y2=1.66
r151 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.185 $Y=1.66
+ $X2=3.515 $Y2=1.66
r152 46 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=2.075
+ $X2=3.43 $Y2=1.99
r153 46 48 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.43 $Y=2.075
+ $X2=3.43 $Y2=2.3
r154 45 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=1.905
+ $X2=3.43 $Y2=1.99
r155 44 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=1.745
+ $X2=3.515 $Y2=1.66
r156 44 45 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.43 $Y=1.745
+ $X2=3.43 $Y2=1.905
r157 42 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=1.99
+ $X2=3.43 $Y2=1.99
r158 42 43 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.345 $Y=1.99
+ $X2=2.335 $Y2=1.99
r159 41 93 3.40825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.25 $Y=2.255
+ $X2=2.25 $Y2=2.36
r160 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=2.075
+ $X2=2.335 $Y2=1.99
r161 40 41 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=2.075
+ $X2=2.25 $Y2=2.255
r162 36 39 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.26 $Y=2.34
+ $X2=1.1 $Y2=2.34
r163 34 93 3.40825 $w=1.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.165 $Y=2.34
+ $X2=2.25 $Y2=2.36
r164 34 39 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=2.165 $Y=2.34
+ $X2=1.1 $Y2=2.34
r165 11 90 300 $w=1.7e-07 $l=5.51362e-07 $layer=licon1_PDIFF $count=2 $X=9.695
+ $Y=1.485 $X2=9.86 $Y2=1.96
r166 10 84 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.855
+ $Y=1.485 $X2=8.99 $Y2=1.96
r167 9 78 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.015
+ $Y=1.485 $X2=8.15 $Y2=1.96
r168 8 72 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.175
+ $Y=1.485 $X2=7.31 $Y2=1.96
r169 7 66 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=6.315
+ $Y=1.485 $X2=6.47 $Y2=1.96
r170 6 60 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.07
+ $Y=1.485 $X2=5.205 $Y2=1.96
r171 5 54 600 $w=1.7e-07 $l=8.39792e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.27 $Y2=2.26
r172 4 48 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.485 $X2=3.43 $Y2=2.3
r173 3 93 600 $w=1.7e-07 $l=1.01336e-06 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=2.25 $Y2=2.3
r174 2 39 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r175 1 36 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%Y 1 2 3 4 5 6 23 25 26 27 33 35 37 40 42 43
+ 44 45 46 54 56 66
r90 63 66 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.01 $Y=0.72
+ $X2=3.85 $Y2=0.72
r91 53 56 2.35727 $w=2.18e-07 $l=4.5e-08 $layer=LI1_cond $X=2.045 $Y=0.805
+ $X2=2.045 $Y2=0.85
r92 46 54 3.18091 $w=2.2e-07 $l=9.5e-08 $layer=LI1_cond $X=2.045 $Y=1.59
+ $X2=2.045 $Y2=1.495
r93 46 54 1.30959 $w=2.18e-07 $l=2.5e-08 $layer=LI1_cond $X=2.045 $Y=1.47
+ $X2=2.045 $Y2=1.495
r94 45 46 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=2.045 $Y=1.19
+ $X2=2.045 $Y2=1.47
r95 44 53 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.72
+ $X2=2.045 $Y2=0.805
r96 44 63 45.5907 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=2.155 $Y=0.72
+ $X2=3.01 $Y2=0.72
r97 44 45 16.7628 $w=2.18e-07 $l=3.2e-07 $layer=LI1_cond $X=2.045 $Y=0.87
+ $X2=2.045 $Y2=1.19
r98 44 56 1.04768 $w=2.18e-07 $l=2e-08 $layer=LI1_cond $X=2.045 $Y=0.87
+ $X2=2.045 $Y2=0.85
r99 38 42 8.35856 $w=1.8e-07 $l=1.82384e-07 $layer=LI1_cond $X=1.685 $Y=1.59
+ $X2=1.517 $Y2=1.62
r100 37 46 3.68316 $w=1.9e-07 $l=1.1e-07 $layer=LI1_cond $X=1.935 $Y=1.59
+ $X2=2.045 $Y2=1.59
r101 37 38 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.935 $Y=1.59
+ $X2=1.685 $Y2=1.59
r102 36 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.72
+ $X2=1.52 $Y2=0.72
r103 35 44 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.935 $Y=0.72
+ $X2=2.045 $Y2=0.72
r104 35 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.935 $Y=0.72
+ $X2=1.605 $Y2=0.72
r105 31 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.635
+ $X2=1.52 $Y2=0.72
r106 31 33 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.52 $Y=0.635
+ $X2=1.52 $Y2=0.46
r107 28 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.66
+ $X2=0.68 $Y2=1.66
r108 27 42 8.35856 $w=1.8e-07 $l=1.85927e-07 $layer=LI1_cond $X=1.35 $Y=1.66
+ $X2=1.517 $Y2=1.62
r109 27 28 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.35 $Y=1.66
+ $X2=0.845 $Y2=1.66
r110 25 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=1.52 $Y2=0.72
r111 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=0.765 $Y2=0.72
r112 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.765 $Y2=0.72
r113 21 23 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.68 $Y2=0.42
r114 6 42 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r115 5 40 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r116 4 66 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.715
+ $Y=0.235 $X2=3.85 $Y2=0.72
r117 3 63 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.235 $X2=3.01 $Y2=0.72
r118 2 33 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.46
r119 1 23 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 41 45 49 53
+ 55 56 57 64 69 74 83 88 95 96 101 107 109 112 115 118 121 124
r150 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r151 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r152 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r153 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r155 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r156 106 107 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=2.53
+ $X2=3.175 $Y2=2.53
r157 103 106 0.434938 $w=5.48e-07 $l=2e-08 $layer=LI1_cond $X=2.99 $Y=2.53
+ $X2=3.01 $Y2=2.53
r158 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r159 100 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r160 99 103 10.0036 $w=5.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=2.53
+ $X2=2.99 $Y2=2.53
r161 99 101 6.78742 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=2.53 $Y=2.53
+ $X2=2.505 $Y2=2.53
r162 99 100 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r163 96 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r164 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r165 93 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.575 $Y=2.72
+ $X2=9.41 $Y2=2.72
r166 93 95 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.575 $Y=2.72
+ $X2=9.89 $Y2=2.72
r167 92 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r168 92 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r169 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r170 89 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.735 $Y=2.72
+ $X2=8.57 $Y2=2.72
r171 89 91 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.735 $Y=2.72
+ $X2=8.97 $Y2=2.72
r172 88 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.245 $Y=2.72
+ $X2=9.41 $Y2=2.72
r173 88 91 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.245 $Y=2.72
+ $X2=8.97 $Y2=2.72
r174 87 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r175 87 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r176 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r177 84 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.895 $Y=2.72
+ $X2=7.73 $Y2=2.72
r178 84 86 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.895 $Y=2.72
+ $X2=8.05 $Y2=2.72
r179 83 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=2.72
+ $X2=8.57 $Y2=2.72
r180 83 86 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.405 $Y=2.72
+ $X2=8.05 $Y2=2.72
r181 82 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r182 82 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r183 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r184 79 115 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=6.165 $Y=2.72
+ $X2=5.83 $Y2=2.72
r185 79 81 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.165 $Y=2.72
+ $X2=6.67 $Y2=2.72
r186 78 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r187 78 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r188 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r189 75 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=4.785 $Y2=2.72
r190 75 77 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=5.29 $Y2=2.72
r191 74 115 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.83 $Y2=2.72
r192 74 77 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.29 $Y2=2.72
r193 73 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r194 73 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r195 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r196 70 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.85 $Y2=2.72
r197 70 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.37 $Y2=2.72
r198 69 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.785 $Y2=2.72
r199 69 72 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.37 $Y2=2.72
r200 68 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r201 68 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r202 67 107 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.175 $Y2=2.72
r203 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r204 64 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.85 $Y2=2.72
r205 64 67 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.45 $Y2=2.72
r206 61 101 148.422 $w=1.68e-07 $l=2.275e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.505 $Y2=2.72
r207 57 100 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r208 57 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r209 55 81 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.725 $Y=2.72
+ $X2=6.67 $Y2=2.72
r210 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=2.72
+ $X2=6.89 $Y2=2.72
r211 51 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.41 $Y=2.635
+ $X2=9.41 $Y2=2.72
r212 51 53 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=9.41 $Y=2.635
+ $X2=9.41 $Y2=2
r213 47 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.57 $Y=2.635
+ $X2=8.57 $Y2=2.72
r214 47 49 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=8.57 $Y=2.635
+ $X2=8.57 $Y2=2
r215 43 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.73 $Y=2.635
+ $X2=7.73 $Y2=2.72
r216 43 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.73 $Y=2.635
+ $X2=7.73 $Y2=2.34
r217 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=2.72
+ $X2=6.89 $Y2=2.72
r218 41 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.565 $Y=2.72
+ $X2=7.73 $Y2=2.72
r219 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.565 $Y=2.72
+ $X2=7.055 $Y2=2.72
r220 37 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=2.635
+ $X2=6.89 $Y2=2.72
r221 37 39 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.89 $Y=2.635
+ $X2=6.89 $Y2=2
r222 33 115 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=2.635
+ $X2=5.83 $Y2=2.72
r223 33 35 11.336 $w=6.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.83 $Y=2.635
+ $X2=5.83 $Y2=2
r224 29 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.635
+ $X2=4.785 $Y2=2.72
r225 29 31 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.785 $Y=2.635
+ $X2=4.785 $Y2=2
r226 25 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2.72
r227 25 27 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2
r228 8 53 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.275
+ $Y=1.485 $X2=9.41 $Y2=2
r229 7 49 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.435
+ $Y=1.485 $X2=8.57 $Y2=2
r230 6 45 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.595
+ $Y=1.485 $X2=7.73 $Y2=2.34
r231 5 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.755
+ $Y=1.485 $X2=6.89 $Y2=2
r232 4 35 150 $w=1.7e-07 $l=7.2655e-07 $layer=licon1_PDIFF $count=4 $X=5.49
+ $Y=1.485 $X2=6 $Y2=2
r233 3 31 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.65
+ $Y=1.485 $X2=4.785 $Y2=2
r234 2 27 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.715
+ $Y=1.485 $X2=3.85 $Y2=2
r235 1 106 300 $w=1.7e-07 $l=1.06637e-06 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.485 $X2=3.01 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 60 61 67 70 73 76
r136 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r137 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r138 70 71 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r139 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r140 61 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0 $X2=9.43
+ $Y2=0
r141 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r142 58 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.575 $Y=0 $X2=9.41
+ $Y2=0
r143 58 60 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.575 $Y=0
+ $X2=9.89 $Y2=0
r144 57 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.43
+ $Y2=0
r145 57 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=8.51
+ $Y2=0
r146 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r147 54 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.735 $Y=0 $X2=8.57
+ $Y2=0
r148 54 56 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.735 $Y=0
+ $X2=8.97 $Y2=0
r149 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.245 $Y=0 $X2=9.41
+ $Y2=0
r150 53 56 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.245 $Y=0
+ $X2=8.97 $Y2=0
r151 52 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.51
+ $Y2=0
r152 52 71 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=8.05 $Y=0 $X2=2.07
+ $Y2=0
r153 51 52 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r154 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=1.94
+ $Y2=0
r155 49 51 387.856 $w=1.68e-07 $l=5.945e-06 $layer=LI1_cond $X=2.105 $Y=0
+ $X2=8.05 $Y2=0
r156 48 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=0 $X2=8.57
+ $Y2=0
r157 48 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.405 $Y=0
+ $X2=8.05 $Y2=0
r158 47 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r159 47 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r160 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r161 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r162 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r163 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.94
+ $Y2=0
r164 43 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.61 $Y2=0
r165 42 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r166 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r167 39 64 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r168 39 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r169 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r170 38 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r171 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r172 36 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r173 32 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.41 $Y=0.085
+ $X2=9.41 $Y2=0
r174 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.41 $Y=0.085
+ $X2=9.41 $Y2=0.38
r175 28 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.57 $Y=0.085
+ $X2=8.57 $Y2=0
r176 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.57 $Y=0.085
+ $X2=8.57 $Y2=0.38
r177 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r178 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.38
r179 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r180 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r181 16 64 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r182 16 18 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r183 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=9.275
+ $Y=0.235 $X2=9.41 $Y2=0.38
r184 4 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.435
+ $Y=0.235 $X2=8.57 $Y2=0.38
r185 3 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r186 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r187 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A_493_47# 1 2 3 4 5 26
r30 24 26 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.11 $Y=0.38
+ $X2=5.95 $Y2=0.38
r31 22 24 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.27 $Y=0.38
+ $X2=5.11 $Y2=0.38
r32 20 22 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.43 $Y=0.38
+ $X2=4.27 $Y2=0.38
r33 17 20 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.59 $Y=0.38
+ $X2=3.43 $Y2=0.38
r34 5 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.38
r35 4 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.235 $X2=5.11 $Y2=0.38
r36 3 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.135
+ $Y=0.235 $X2=4.27 $Y2=0.38
r37 2 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.295
+ $Y=0.235 $X2=3.43 $Y2=0.38
r38 1 17 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.59 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A_911_47# 1 2 3 4 21
c31 21 0 1.25206e-19 $X=7.73 $Y=0.72
r32 19 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.89 $Y=0.72
+ $X2=7.73 $Y2=0.72
r33 17 19 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=5.53 $Y=0.72
+ $X2=6.89 $Y2=0.72
r34 14 17 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.69 $Y=0.72
+ $X2=5.53 $Y2=0.72
r35 4 21 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=7.595
+ $Y=0.235 $X2=7.73 $Y2=0.72
r36 3 19 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.755
+ $Y=0.235 $X2=6.89 $Y2=0.72
r37 2 17 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.53 $Y2=0.72
r38 1 14 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.555
+ $Y=0.235 $X2=4.69 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_4%A_1269_47# 1 2 3 4 5 16 22 24 28 30 34 38
r45 32 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.83 $Y=0.635
+ $X2=9.83 $Y2=0.42
r46 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.075 $Y=0.72
+ $X2=8.99 $Y2=0.72
r47 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.745 $Y=0.72
+ $X2=9.83 $Y2=0.635
r48 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.745 $Y=0.72
+ $X2=9.075 $Y2=0.72
r49 26 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=0.635
+ $X2=8.99 $Y2=0.72
r50 26 28 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.99 $Y=0.635
+ $X2=8.99 $Y2=0.42
r51 24 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=0.72
+ $X2=8.99 $Y2=0.72
r52 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.905 $Y=0.72
+ $X2=8.235 $Y2=0.72
r53 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.15 $Y=0.635
+ $X2=8.235 $Y2=0.72
r54 22 37 3.40825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.15 $Y=0.465
+ $X2=8.15 $Y2=0.36
r55 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.15 $Y=0.465
+ $X2=8.15 $Y2=0.635
r56 18 21 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.47 $Y=0.38
+ $X2=7.31 $Y2=0.38
r57 16 37 3.40825 $w=1.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=8.065 $Y=0.38
+ $X2=8.15 $Y2=0.36
r58 16 21 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.065 $Y=0.38
+ $X2=7.31 $Y2=0.38
r59 5 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.695
+ $Y=0.235 $X2=9.83 $Y2=0.42
r60 4 28 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.855
+ $Y=0.235 $X2=8.99 $Y2=0.42
r61 3 37 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.015
+ $Y=0.235 $X2=8.15 $Y2=0.42
r62 2 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.31 $Y2=0.38
r63 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.345
+ $Y=0.235 $X2=6.47 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o2111ai_4.spice
* Created: Thu Aug 27 14:34:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2111ai_4.spice.pex"
.subckt sky130_fd_sc_hd__o2111ai_4  VNB VPB D1 C1 B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1016 N_A_27_47#_M1016_d N_D1_M1016_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1020 N_A_27_47#_M1020_d N_D1_M1020_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1023 N_A_27_47#_M1020_d N_D1_M1023_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1039 N_A_27_47#_M1039_d N_D1_M1039_g N_Y_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1021 N_A_445_47#_M1021_d N_C1_M1021_g N_A_27_47#_M1039_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1026 N_A_445_47#_M1021_d N_C1_M1026_g N_A_27_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1032 N_A_445_47#_M1032_d N_C1_M1032_g N_A_27_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1033 N_A_445_47#_M1032_d N_C1_M1033_g N_A_27_47#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_A_445_47#_M1014_d N_B1_M1014_g N_A_803_47#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1017 N_A_445_47#_M1014_d N_B1_M1017_g N_A_803_47#_M1017_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1022 N_A_445_47#_M1022_d N_B1_M1022_g N_A_803_47#_M1017_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1027 N_A_445_47#_M1022_d N_B1_M1027_g N_A_803_47#_M1027_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.095875 PD=0.92 PS=0.945 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75001.4 SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1024 N_A_803_47#_M1027_s N_A2_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.08775 PD=0.945 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1028 N_A_803_47#_M1028_d N_A2_M1028_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.08775 PD=0.94 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1029 N_A_803_47#_M1028_d N_A2_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.08775 PD=0.94 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1031 N_A_803_47#_M1031_d N_A2_M1031_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.08775 PD=0.945 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75003.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_803_47#_M1031_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.095875 PD=0.92 PS=0.945 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1005_d N_A1_M1006_g N_A_803_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A1_M1012_g N_A_803_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1012_d N_A1_M1018_g N_A_803_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.18525 PD=0.92 PS=1.87 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_D1_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75006.7 A=0.15
+ P=2.3 MULT=1
MM1009 N_VPWR_M1003_d N_D1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75006.3
+ A=0.15 P=2.3 MULT=1
MM1025 N_VPWR_M1025_d N_D1_M1025_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75005.9 A=0.15
+ P=2.3 MULT=1
MM1036 N_VPWR_M1025_d N_D1_M1036_g N_Y_M1036_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75005.4
+ A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_C1_M1001_g N_Y_M1036_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75005 A=0.15
+ P=2.3 MULT=1
MM1010 N_VPWR_M1001_d N_C1_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75004.6
+ A=0.15 P=2.3 MULT=1
MM1030 N_VPWR_M1030_d N_C1_M1030_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7 SB=75004.2
+ A=0.15 P=2.3 MULT=1
MM1037 N_VPWR_M1030_d N_C1_M1037_g N_Y_M1037_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.2375 PD=1.27 PS=1.475 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1 SB=75003.8
+ A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_Y_M1037_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.2375 PD=1.27 PS=1.475 NRD=0 NRS=39.4 M=1 R=6.66667 SA=75003.7 SB=75003.1
+ A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1007_d N_B1_M1013_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.2 SB=75002.7
+ A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_B1_M1015_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.6 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1038 N_VPWR_M1015_d N_B1_M1038_g N_Y_M1038_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.1475 PD=1.27 PS=1.295 NRD=0 NRS=0 M=1 R=6.66667 SA=75005 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1002 N_Y_M1038_s N_A2_M1002_g N_A_1163_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1475 AS=0.135 PD=1.295 PS=1.27 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75005.5
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1008 N_Y_M1008_d N_A2_M1008_g N_A_1163_297#_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.9
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1011 N_Y_M1008_d N_A2_M1011_g N_A_1163_297#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.3
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1034 N_Y_M1034_d N_A2_M1034_g N_A_1163_297#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.25335 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_1163_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.25285 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_1163_297#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1004_d N_A1_M1019_g N_A_1163_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1035 N_VPWR_M1035_d N_A1_M1035_g N_A_1163_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_67 VNB 0 1.11453e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__o2111ai_4.spice.SKY130_FD_SC_HD__O2111AI_4.pxi"
*
.ends
*
*

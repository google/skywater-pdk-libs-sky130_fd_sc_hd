* File: sky130_fd_sc_hd__o2111a_4.pxi.spice
* Created: Tue Sep  1 19:20:03 2020
* 
x_PM_SKY130_FD_SC_HD__O2111A_4%D1 N_D1_c_122_n N_D1_M1009_g N_D1_M1002_g
+ N_D1_c_123_n N_D1_M1024_g N_D1_M1015_g D1 D1 PM_SKY130_FD_SC_HD__O2111A_4%D1
x_PM_SKY130_FD_SC_HD__O2111A_4%C1 N_C1_c_162_n N_C1_M1011_g N_C1_M1000_g
+ N_C1_M1014_g N_C1_M1003_g N_C1_c_164_n N_C1_c_165_n N_C1_c_179_n C1 C1
+ N_C1_c_166_n N_C1_c_221_p N_C1_c_167_n PM_SKY130_FD_SC_HD__O2111A_4%C1
x_PM_SKY130_FD_SC_HD__O2111A_4%B1 N_B1_M1020_g N_B1_M1016_g N_B1_M1012_g
+ N_B1_M1022_g B1 N_B1_c_251_n PM_SKY130_FD_SC_HD__O2111A_4%B1
x_PM_SKY130_FD_SC_HD__O2111A_4%A2 N_A2_M1008_g N_A2_c_294_n N_A2_M1018_g
+ N_A2_c_295_n N_A2_M1026_g N_A2_M1021_g N_A2_c_315_p N_A2_c_302_n N_A2_c_297_n
+ A2 A2 N_A2_c_299_n N_A2_c_337_p PM_SKY130_FD_SC_HD__O2111A_4%A2
x_PM_SKY130_FD_SC_HD__O2111A_4%A1 N_A1_c_381_n N_A1_M1004_g N_A1_c_377_n
+ N_A1_M1001_g N_A1_c_382_n N_A1_M1019_g N_A1_c_378_n N_A1_M1005_g A1
+ N_A1_c_380_n PM_SKY130_FD_SC_HD__O2111A_4%A1
x_PM_SKY130_FD_SC_HD__O2111A_4%A_27_297# N_A_27_297#_M1009_s N_A_27_297#_M1002_d
+ N_A_27_297#_M1015_d N_A_27_297#_M1016_s N_A_27_297#_M1003_s
+ N_A_27_297#_M1026_d N_A_27_297#_M1006_g N_A_27_297#_M1007_g
+ N_A_27_297#_M1013_g N_A_27_297#_M1010_g N_A_27_297#_M1025_g
+ N_A_27_297#_M1017_g N_A_27_297#_M1027_g N_A_27_297#_M1023_g
+ N_A_27_297#_c_437_n N_A_27_297#_c_444_n N_A_27_297#_c_461_n
+ N_A_27_297#_c_438_n N_A_27_297#_c_465_n N_A_27_297#_c_478_n
+ N_A_27_297#_c_439_n N_A_27_297#_c_440_n N_A_27_297#_c_431_n
+ N_A_27_297#_c_441_n N_A_27_297#_c_520_p N_A_27_297#_c_466_n
+ N_A_27_297#_c_467_n N_A_27_297#_c_470_n N_A_27_297#_c_442_n
+ N_A_27_297#_c_432_n PM_SKY130_FD_SC_HD__O2111A_4%A_27_297#
x_PM_SKY130_FD_SC_HD__O2111A_4%VPWR N_VPWR_M1002_s N_VPWR_M1000_d N_VPWR_M1022_d
+ N_VPWR_M1004_s N_VPWR_M1007_s N_VPWR_M1010_s N_VPWR_M1023_s N_VPWR_c_598_n
+ N_VPWR_c_599_n N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n N_VPWR_c_603_n
+ N_VPWR_c_604_n N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n N_VPWR_c_608_n
+ N_VPWR_c_609_n VPWR N_VPWR_c_610_n N_VPWR_c_611_n N_VPWR_c_612_n
+ N_VPWR_c_613_n N_VPWR_c_614_n N_VPWR_c_615_n N_VPWR_c_616_n N_VPWR_c_617_n
+ N_VPWR_c_618_n N_VPWR_c_597_n PM_SKY130_FD_SC_HD__O2111A_4%VPWR
x_PM_SKY130_FD_SC_HD__O2111A_4%X N_X_M1006_d N_X_M1025_d N_X_M1007_d N_X_M1017_d
+ N_X_c_738_n N_X_c_763_n N_X_c_739_n N_X_c_743_n N_X_c_746_n N_X_c_750_n
+ N_X_c_782_p N_X_c_767_n N_X_c_752_n N_X_c_753_n N_X_c_754_n N_X_c_756_n X X X
+ N_X_c_735_n N_X_c_737_n PM_SKY130_FD_SC_HD__O2111A_4%X
x_PM_SKY130_FD_SC_HD__O2111A_4%A_27_47# N_A_27_47#_M1009_d N_A_27_47#_M1024_d
+ N_A_27_47#_M1014_s N_A_27_47#_c_791_n N_A_27_47#_c_792_n
+ PM_SKY130_FD_SC_HD__O2111A_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O2111A_4%A_361_47# N_A_361_47#_M1020_d N_A_361_47#_M1018_s
+ N_A_361_47#_M1005_s N_A_361_47#_c_821_n N_A_361_47#_c_857_p
+ N_A_361_47#_c_836_n N_A_361_47#_c_822_n N_A_361_47#_c_854_p
+ N_A_361_47#_c_823_n PM_SKY130_FD_SC_HD__O2111A_4%A_361_47#
x_PM_SKY130_FD_SC_HD__O2111A_4%VGND N_VGND_M1018_d N_VGND_M1001_d N_VGND_M1021_d
+ N_VGND_M1013_s N_VGND_M1027_s N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n
+ N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n
+ N_VGND_c_879_n N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n VGND
+ N_VGND_c_883_n N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n
+ PM_SKY130_FD_SC_HD__O2111A_4%VGND
cc_1 VNB N_D1_c_122_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_D1_c_123_n 0.0611703f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_3 VNB N_D1_M1024_g 0.0171276f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_4 VNB N_D1_M1015_g 4.05031e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_5 VNB D1 0.00204204f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_C1_c_162_n 0.0164838f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_7 VNB N_C1_M1014_g 0.0221101f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_8 VNB N_C1_c_164_n 0.00365621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C1_c_165_n 0.0207255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_C1_c_166_n 0.0285962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_C1_c_167_n 0.00194425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_M1020_g 0.0177028f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_B1_M1016_g 4.05412e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B1_M1012_g 0.0170795f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_M1022_g 4.26256e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_c_251_n 0.0301236f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_17 VNB N_A2_M1008_g 4.28981e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_18 VNB N_A2_c_294_n 0.0187383f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_19 VNB N_A2_c_295_n 0.031896f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_20 VNB N_A2_M1021_g 0.0207111f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_21 VNB N_A2_c_297_n 0.00338548f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_22 VNB A2 0.00371495f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_23 VNB N_A2_c_299_n 0.0400877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A1_c_377_n 0.0158468f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_25 VNB N_A1_c_378_n 0.0160662f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_26 VNB A1 0.0017762f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_27 VNB N_A1_c_380_n 0.0427275f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_28 VNB N_A_27_297#_M1006_g 0.0203289f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_29 VNB N_A_27_297#_M1007_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_30 VNB N_A_27_297#_M1013_g 0.0185737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_297#_M1010_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_297#_M1025_g 0.0177469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_297#_M1017_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_297#_M1027_g 0.0201822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_297#_M1023_g 4.85024e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_27_297#_c_431_n 0.00338475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_27_297#_c_432_n 0.0786941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_597_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB X 0.0227943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_X_c_735_n 0.00765935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_27_47#_c_791_n 0.00400317f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_42 VNB N_A_27_47#_c_792_n 0.0233894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_361_47#_c_821_n 0.0163832f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_44 VNB N_A_361_47#_c_822_n 0.0023793f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_45 VNB N_A_361_47#_c_823_n 0.0025711f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_46 VNB N_VGND_c_871_n 0.00539026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_872_n 3.35563e-19 $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_48 VNB N_VGND_c_873_n 0.00474897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_874_n 0.00257633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_875_n 0.0105642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_876_n 0.0146805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_877_n 0.0729641f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_878_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_879_n 0.0120314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_880_n 0.00489469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_881_n 0.0170488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_882_n 0.00506925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_883_n 0.0217032f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_884_n 0.0118058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_885_n 0.00452805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_886_n 0.354649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VPB N_D1_M1002_g 0.0209706f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_63 VPB N_D1_c_123_n 0.0101638f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.025
cc_64 VPB N_D1_M1015_g 0.0188363f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_65 VPB D1 0.0128458f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_66 VPB N_C1_M1000_g 0.0172688f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_C1_M1003_g 0.0207856f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_C1_c_164_n 0.00302148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_C1_c_165_n 0.00428608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB C1 0.0037219f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_71 VPB N_C1_c_166_n 0.00500449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_C1_c_167_n 0.00258653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B1_M1016_g 0.0197688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B1_M1022_g 0.0195553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB B1 0.00249609f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_76 VPB N_A2_M1008_g 0.0223544f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_77 VPB N_A2_c_295_n 0.0271263f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.025
cc_78 VPB N_A2_c_302_n 0.00255463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A2_c_297_n 0.00256985f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_80 VPB A2 0.00189249f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_81 VPB A2 0.00160609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A1_c_381_n 0.0143411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_83 VPB N_A1_c_382_n 0.0149555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB A1 0.00215977f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_85 VPB N_A1_c_380_n 0.0132751f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_86 VPB N_A_27_297#_M1007_g 0.0221269f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_87 VPB N_A_27_297#_M1010_g 0.0191857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_27_297#_M1017_g 0.0192606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_27_297#_M1023_g 0.0221659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_27_297#_c_437_n 0.017641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_27_297#_c_438_n 0.00852169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_27_297#_c_439_n 0.0122513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_27_297#_c_440_n 0.00339654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_297#_c_441_n 0.00846493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_297#_c_442_n 0.00724245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_598_n 4.03531e-19 $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_97 VPB N_VPWR_c_599_n 0.00367883f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.53
cc_98 VPB N_VPWR_c_600_n 4.06069e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_601_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_602_n 0.00623686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_603_n 3.05427e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_604_n 0.0100112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_605_n 0.0282835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_606_n 0.0134295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_607_n 0.00429685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_608_n 0.013458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_609_n 0.00436611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_610_n 0.0146402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_611_n 0.030314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_612_n 0.0283851f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_613_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_614_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_615_n 0.00436611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_616_n 0.00436584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_617_n 0.0052688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_618_n 0.00423552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_597_n 0.0467425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB X 0.00947675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_X_c_737_n 0.00785406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 N_D1_M1024_g N_C1_c_162_n 0.0270204f $X=0.89 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_121 N_D1_M1015_g N_C1_M1000_g 0.0260359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_122 N_D1_M1024_g N_C1_c_164_n 0.00348438f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_123 N_D1_M1024_g N_C1_c_165_n 0.0214191f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_124 N_D1_M1015_g N_C1_c_179_n 0.00135261f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_125 D1 N_A_27_297#_M1002_d 0.00396794f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_126 N_D1_c_122_n N_A_27_297#_c_444_n 0.0109603f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_127 N_D1_M1002_g N_A_27_297#_c_444_n 0.0171771f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_128 N_D1_c_123_n N_A_27_297#_c_444_n 0.021035f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_129 N_D1_M1024_g N_A_27_297#_c_444_n 0.00933244f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_130 N_D1_M1015_g N_A_27_297#_c_444_n 0.0146909f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_131 D1 N_A_27_297#_c_444_n 0.0417872f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_132 N_D1_M1002_g N_A_27_297#_c_438_n 0.0133175f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_133 N_D1_c_123_n N_A_27_297#_c_438_n 8.48834e-19 $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_134 N_D1_M1015_g N_A_27_297#_c_438_n 0.0124758f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_135 D1 N_A_27_297#_c_438_n 0.018644f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_136 N_D1_M1002_g N_VPWR_c_598_n 0.00922823f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_137 N_D1_M1015_g N_VPWR_c_598_n 0.00758592f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_138 N_D1_M1015_g N_VPWR_c_606_n 0.00348296f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_139 N_D1_M1002_g N_VPWR_c_610_n 0.00348296f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_140 N_D1_M1002_g N_VPWR_c_597_n 0.0050535f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_141 N_D1_M1015_g N_VPWR_c_597_n 0.0041265f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_142 N_D1_c_122_n N_A_27_47#_c_791_n 0.0130183f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_143 N_D1_c_123_n N_A_27_47#_c_791_n 2.99382e-19 $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_144 N_D1_M1024_g N_A_27_47#_c_791_n 0.0124787f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_145 N_D1_c_123_n N_A_27_47#_c_792_n 0.00168825f $X=0.89 $Y=1.025 $X2=0 $Y2=0
cc_146 D1 N_A_27_47#_c_792_n 0.0187382f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_147 N_D1_c_122_n N_VGND_c_877_n 0.00357877f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_148 N_D1_M1024_g N_VGND_c_877_n 0.00357877f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_149 N_D1_c_122_n N_VGND_c_886_n 0.00617937f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_150 N_D1_M1024_g N_VGND_c_886_n 0.00525237f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_151 N_C1_c_162_n N_B1_M1020_g 0.0441466f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_152 N_C1_c_164_n N_B1_M1020_g 0.00146486f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_153 N_C1_c_165_n N_B1_M1020_g 0.0213318f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_154 N_C1_M1000_g N_B1_M1016_g 0.0459625f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_155 N_C1_c_164_n N_B1_M1016_g 0.00317217f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_156 C1 N_B1_M1016_g 0.013063f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_157 N_C1_M1014_g N_B1_M1012_g 0.0392465f $X=2.51 $Y=0.56 $X2=0 $Y2=0
cc_158 C1 N_B1_M1022_g 0.0137869f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_159 N_C1_c_166_n N_B1_M1022_g 0.0466515f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_160 N_C1_c_164_n B1 0.00955418f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_161 N_C1_c_165_n B1 7.02332e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_162 C1 B1 0.0282665f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_163 N_C1_c_166_n B1 8.19412e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_164 N_C1_c_167_n B1 0.0147269f $X=2.552 $Y=1.197 $X2=0 $Y2=0
cc_165 C1 N_B1_c_251_n 5.93738e-19 $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_166 N_C1_c_166_n N_B1_c_251_n 0.0392465f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_167 N_C1_c_167_n N_B1_c_251_n 8.56423e-19 $X=2.552 $Y=1.197 $X2=0 $Y2=0
cc_168 N_C1_M1003_g N_A2_M1008_g 0.0124528f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_169 C1 N_A2_M1008_g 0.00111062f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_170 N_C1_c_166_n N_A2_M1008_g 2.3171e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_171 N_C1_c_166_n A2 3.24534e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_172 N_C1_c_167_n A2 0.0117826f $X=2.552 $Y=1.197 $X2=0 $Y2=0
cc_173 C1 A2 0.00454775f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_174 N_C1_M1014_g N_A2_c_299_n 0.00159065f $X=2.51 $Y=0.56 $X2=0 $Y2=0
cc_175 N_C1_c_166_n N_A2_c_299_n 0.0117048f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_176 N_C1_c_167_n N_A2_c_299_n 4.19817e-19 $X=2.552 $Y=1.197 $X2=0 $Y2=0
cc_177 N_C1_c_179_n N_A_27_297#_M1015_d 0.00215164f $X=1.395 $Y=1.575 $X2=0
+ $Y2=0
cc_178 C1 N_A_27_297#_M1016_s 0.00312144f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_179 N_C1_c_162_n N_A_27_297#_c_444_n 0.00172638f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_180 N_C1_M1000_g N_A_27_297#_c_444_n 0.00104684f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_181 N_C1_c_164_n N_A_27_297#_c_444_n 0.0256978f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_182 N_C1_c_165_n N_A_27_297#_c_444_n 3.42171e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_183 N_C1_c_179_n N_A_27_297#_c_444_n 0.00934241f $X=1.395 $Y=1.575 $X2=0
+ $Y2=0
cc_184 N_C1_M1000_g N_A_27_297#_c_461_n 0.0101581f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_185 N_C1_c_179_n N_A_27_297#_c_461_n 0.0113935f $X=1.395 $Y=1.575 $X2=0 $Y2=0
cc_186 C1 N_A_27_297#_c_461_n 0.0208319f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_187 N_C1_c_179_n N_A_27_297#_c_438_n 0.00246268f $X=1.395 $Y=1.575 $X2=0
+ $Y2=0
cc_188 N_C1_M1000_g N_A_27_297#_c_465_n 5.52189e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_189 C1 N_A_27_297#_c_466_n 0.013379f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_190 N_C1_M1003_g N_A_27_297#_c_467_n 0.0132218f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_191 C1 N_A_27_297#_c_467_n 0.0215453f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_192 N_C1_c_221_p N_A_27_297#_c_467_n 0.0113061f $X=2.552 $Y=1.49 $X2=0 $Y2=0
cc_193 N_C1_c_166_n N_A_27_297#_c_470_n 8.75972e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_194 N_C1_c_167_n N_A_27_297#_c_470_n 0.00529866f $X=2.552 $Y=1.197 $X2=0
+ $Y2=0
cc_195 C1 N_VPWR_M1000_d 0.00750015f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_196 C1 N_VPWR_M1022_d 0.00472172f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_197 N_C1_M1000_g N_VPWR_c_598_n 5.51123e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_198 N_C1_M1000_g N_VPWR_c_599_n 0.0014971f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_199 N_C1_M1003_g N_VPWR_c_600_n 0.00922086f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_200 N_C1_M1000_g N_VPWR_c_606_n 0.00436487f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_201 N_C1_M1003_g N_VPWR_c_611_n 0.00348405f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_202 N_C1_M1000_g N_VPWR_c_597_n 0.00582874f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_203 N_C1_M1003_g N_VPWR_c_597_n 0.00475565f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_204 N_C1_c_162_n N_A_27_47#_c_791_n 0.0108385f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_205 N_C1_M1014_g N_A_27_47#_c_791_n 0.00859109f $X=2.51 $Y=0.56 $X2=0 $Y2=0
cc_206 N_C1_c_164_n N_A_27_47#_c_791_n 0.00687433f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_207 N_C1_c_165_n N_A_27_47#_c_791_n 9.06076e-19 $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_208 N_C1_c_162_n N_A_361_47#_c_821_n 0.00124376f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_209 N_C1_M1014_g N_A_361_47#_c_821_n 0.0151132f $X=2.51 $Y=0.56 $X2=0 $Y2=0
cc_210 C1 N_A_361_47#_c_821_n 0.00530528f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_211 N_C1_c_166_n N_A_361_47#_c_821_n 0.00560355f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_212 N_C1_c_167_n N_A_361_47#_c_821_n 0.0241185f $X=2.552 $Y=1.197 $X2=0 $Y2=0
cc_213 N_C1_M1014_g N_VGND_c_871_n 0.00222873f $X=2.51 $Y=0.56 $X2=0 $Y2=0
cc_214 N_C1_c_162_n N_VGND_c_877_n 0.00357877f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_215 N_C1_M1014_g N_VGND_c_877_n 0.00357877f $X=2.51 $Y=0.56 $X2=0 $Y2=0
cc_216 N_C1_c_162_n N_VGND_c_886_n 0.00528062f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_217 N_C1_M1014_g N_VGND_c_886_n 0.00641668f $X=2.51 $Y=0.56 $X2=0 $Y2=0
cc_218 N_B1_M1016_g N_A_27_297#_c_461_n 0.00961342f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B1_M1016_g N_A_27_297#_c_465_n 0.00642869f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_220 N_B1_M1016_g N_A_27_297#_c_466_n 0.00232001f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B1_M1022_g N_A_27_297#_c_467_n 0.0118623f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_222 N_B1_M1016_g N_VPWR_c_599_n 0.00145759f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B1_M1016_g N_VPWR_c_600_n 4.71778e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_224 N_B1_M1022_g N_VPWR_c_600_n 0.00758755f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_225 N_B1_M1016_g N_VPWR_c_608_n 0.0043275f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B1_M1022_g N_VPWR_c_608_n 0.00348405f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_227 N_B1_M1016_g N_VPWR_c_597_n 0.00578153f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_228 N_B1_M1022_g N_VPWR_c_597_n 0.00410128f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B1_M1020_g N_A_27_47#_c_791_n 0.0138856f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_230 N_B1_M1012_g N_A_27_47#_c_791_n 0.0112735f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_231 N_B1_M1020_g N_A_361_47#_c_821_n 0.00858956f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_232 N_B1_M1012_g N_A_361_47#_c_821_n 0.00960749f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_233 B1 N_A_361_47#_c_821_n 0.0253424f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_234 N_B1_c_251_n N_A_361_47#_c_821_n 0.00204539f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B1_M1020_g N_VGND_c_877_n 0.00357877f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_236 N_B1_M1012_g N_VGND_c_877_n 0.00357877f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B1_M1020_g N_VGND_c_886_n 0.0052923f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B1_M1012_g N_VGND_c_886_n 0.00512949f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_239 N_A2_c_315_p N_A1_c_381_n 0.0115024f $X=4.655 $Y=1.575 $X2=-0.19
+ $Y2=-0.24
cc_240 N_A2_c_294_n N_A1_c_377_n 0.00810501f $X=3.485 $Y=0.96 $X2=0 $Y2=0
cc_241 N_A2_c_315_p N_A1_c_382_n 0.0109024f $X=4.655 $Y=1.575 $X2=0 $Y2=0
cc_242 N_A2_M1021_g N_A1_c_378_n 0.010422f $X=4.89 $Y=0.56 $X2=0 $Y2=0
cc_243 N_A2_c_295_n A1 0.00123191f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_244 N_A2_c_315_p A1 0.035393f $X=4.655 $Y=1.575 $X2=0 $Y2=0
cc_245 N_A2_c_297_n A1 0.0201128f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_246 A2 A1 0.0123597f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_247 N_A2_c_299_n A1 2.1194e-19 $X=3.33 $Y=1.127 $X2=0 $Y2=0
cc_248 N_A2_M1008_g N_A1_c_380_n 0.0606277f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A2_c_295_n N_A1_c_380_n 0.0586377f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_250 N_A2_c_315_p N_A1_c_380_n 0.00377231f $X=4.655 $Y=1.575 $X2=0 $Y2=0
cc_251 N_A2_c_302_n N_A1_c_380_n 0.00102205f $X=4.74 $Y=1.49 $X2=0 $Y2=0
cc_252 N_A2_c_297_n N_A1_c_380_n 2.31305e-19 $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_253 A2 N_A1_c_380_n 0.00239931f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_254 A2 N_A1_c_380_n 0.00444041f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_255 N_A2_c_299_n N_A1_c_380_n 0.0141055f $X=3.33 $Y=1.127 $X2=0 $Y2=0
cc_256 N_A2_c_315_p N_A_27_297#_M1026_d 0.00340393f $X=4.655 $Y=1.575 $X2=0
+ $Y2=0
cc_257 N_A2_M1021_g N_A_27_297#_M1006_g 0.0192248f $X=4.89 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A2_M1008_g N_A_27_297#_c_478_n 0.00875403f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A2_c_295_n N_A_27_297#_c_478_n 0.0105985f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_260 N_A2_c_315_p N_A_27_297#_c_478_n 0.0621529f $X=4.655 $Y=1.575 $X2=0 $Y2=0
cc_261 N_A2_c_337_p N_A_27_297#_c_478_n 0.0186062f $X=3.452 $Y=1.49 $X2=0 $Y2=0
cc_262 N_A2_c_295_n N_A_27_297#_c_440_n 0.00462588f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_263 N_A2_c_315_p N_A_27_297#_c_440_n 0.0057166f $X=4.655 $Y=1.575 $X2=0 $Y2=0
cc_264 N_A2_c_302_n N_A_27_297#_c_440_n 0.00558653f $X=4.74 $Y=1.49 $X2=0 $Y2=0
cc_265 N_A2_c_295_n N_A_27_297#_c_431_n 0.00120986f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_266 N_A2_c_297_n N_A_27_297#_c_431_n 0.0110718f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A2_M1008_g N_A_27_297#_c_470_n 0.00996693f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_268 A2 N_A_27_297#_c_470_n 0.00487856f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_269 N_A2_c_299_n N_A_27_297#_c_470_n 6.31812e-19 $X=3.33 $Y=1.127 $X2=0 $Y2=0
cc_270 N_A2_c_295_n N_A_27_297#_c_442_n 0.00100085f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_271 N_A2_c_297_n N_A_27_297#_c_442_n 0.00613873f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A2_c_295_n N_A_27_297#_c_432_n 0.00770175f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_273 N_A2_c_297_n N_A_27_297#_c_432_n 2.58369e-19 $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A2_c_315_p N_VPWR_M1004_s 0.00349895f $X=4.655 $Y=1.575 $X2=0 $Y2=0
cc_275 N_A2_M1008_g N_VPWR_c_601_n 0.00195655f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A2_c_295_n N_VPWR_c_601_n 0.00189899f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_277 N_A2_c_295_n N_VPWR_c_602_n 0.00284653f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_278 N_A2_M1008_g N_VPWR_c_611_n 0.00420765f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A2_c_295_n N_VPWR_c_612_n 0.00436487f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_280 N_A2_M1008_g N_VPWR_c_597_n 0.00656811f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A2_c_295_n N_VPWR_c_597_n 0.00758582f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_282 N_A2_c_315_p A_681_297# 6.74115e-19 $X=4.655 $Y=1.575 $X2=-0.19 $Y2=-0.24
cc_283 N_A2_c_337_p A_681_297# 0.00151284f $X=3.452 $Y=1.49 $X2=-0.19 $Y2=-0.24
cc_284 N_A2_c_315_p A_852_297# 0.00560096f $X=4.655 $Y=1.575 $X2=-0.19 $Y2=-0.24
cc_285 N_A2_c_294_n N_A_361_47#_c_821_n 0.0140636f $X=3.485 $Y=0.96 $X2=0 $Y2=0
cc_286 A2 N_A_361_47#_c_821_n 0.0294096f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_287 N_A2_c_299_n N_A_361_47#_c_821_n 0.00749007f $X=3.33 $Y=1.127 $X2=0 $Y2=0
cc_288 N_A2_c_315_p N_A_361_47#_c_836_n 0.00144847f $X=4.655 $Y=1.575 $X2=0
+ $Y2=0
cc_289 N_A2_c_295_n N_A_361_47#_c_822_n 0.00478161f $X=4.69 $Y=1.405 $X2=0 $Y2=0
cc_290 N_A2_c_315_p N_A_361_47#_c_822_n 0.00283979f $X=4.655 $Y=1.575 $X2=0
+ $Y2=0
cc_291 N_A2_c_297_n N_A_361_47#_c_822_n 0.00881652f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A2_c_315_p N_A_361_47#_c_823_n 0.00534062f $X=4.655 $Y=1.575 $X2=0
+ $Y2=0
cc_293 N_A2_c_294_n N_VGND_c_871_n 0.00808217f $X=3.485 $Y=0.96 $X2=0 $Y2=0
cc_294 N_A2_c_294_n N_VGND_c_872_n 5.04642e-19 $X=3.485 $Y=0.96 $X2=0 $Y2=0
cc_295 N_A2_M1021_g N_VGND_c_872_n 5.55765e-19 $X=4.89 $Y=0.56 $X2=0 $Y2=0
cc_296 N_A2_M1021_g N_VGND_c_873_n 0.00302344f $X=4.89 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A2_c_294_n N_VGND_c_879_n 0.00341689f $X=3.485 $Y=0.96 $X2=0 $Y2=0
cc_298 N_A2_M1021_g N_VGND_c_881_n 0.00585385f $X=4.89 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A2_c_294_n N_VGND_c_886_n 0.00411698f $X=3.485 $Y=0.96 $X2=0 $Y2=0
cc_300 N_A2_M1021_g N_VGND_c_886_n 0.0112386f $X=4.89 $Y=0.56 $X2=0 $Y2=0
cc_301 N_A1_c_381_n N_A_27_297#_c_478_n 0.0120202f $X=3.755 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A1_c_382_n N_A_27_297#_c_478_n 0.0124666f $X=4.185 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A1_c_381_n N_A_27_297#_c_470_n 0.00169493f $X=3.755 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A1_c_381_n N_VPWR_c_601_n 0.0104101f $X=3.755 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A1_c_382_n N_VPWR_c_601_n 0.0110905f $X=4.185 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A1_c_381_n N_VPWR_c_611_n 0.00362954f $X=3.755 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A1_c_382_n N_VPWR_c_612_n 0.00362954f $X=4.185 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A1_c_381_n N_VPWR_c_597_n 0.0043358f $X=3.755 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A1_c_382_n N_VPWR_c_597_n 0.00452531f $X=4.185 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A1_c_377_n N_A_361_47#_c_836_n 0.0113936f $X=3.95 $Y=0.985 $X2=0 $Y2=0
cc_311 N_A1_c_378_n N_A_361_47#_c_836_n 0.0108187f $X=4.37 $Y=0.985 $X2=0 $Y2=0
cc_312 A1 N_A_361_47#_c_836_n 0.0340921f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_313 N_A1_c_380_n N_A_361_47#_c_836_n 0.00261576f $X=4.185 $Y=1.197 $X2=0
+ $Y2=0
cc_314 N_A1_c_380_n N_A_361_47#_c_823_n 0.00364018f $X=4.185 $Y=1.197 $X2=0
+ $Y2=0
cc_315 N_A1_c_377_n N_VGND_c_871_n 5.0237e-19 $X=3.95 $Y=0.985 $X2=0 $Y2=0
cc_316 N_A1_c_377_n N_VGND_c_872_n 0.00698067f $X=3.95 $Y=0.985 $X2=0 $Y2=0
cc_317 N_A1_c_378_n N_VGND_c_872_n 0.00961104f $X=4.37 $Y=0.985 $X2=0 $Y2=0
cc_318 N_A1_c_377_n N_VGND_c_879_n 0.00341689f $X=3.95 $Y=0.985 $X2=0 $Y2=0
cc_319 N_A1_c_378_n N_VGND_c_881_n 0.0022755f $X=4.37 $Y=0.985 $X2=0 $Y2=0
cc_320 N_A1_c_377_n N_VGND_c_886_n 0.00411698f $X=3.95 $Y=0.985 $X2=0 $Y2=0
cc_321 N_A1_c_378_n N_VGND_c_886_n 0.00313008f $X=4.37 $Y=0.985 $X2=0 $Y2=0
cc_322 N_A_27_297#_c_438_n N_VPWR_M1002_s 0.00168211f $X=1.23 $Y=1.917 $X2=-0.19
+ $Y2=-0.24
cc_323 N_A_27_297#_c_461_n N_VPWR_M1000_d 0.00324921f $X=1.795 $Y=1.917 $X2=0
+ $Y2=0
cc_324 N_A_27_297#_c_467_n N_VPWR_M1022_d 0.00324921f $X=2.695 $Y=2.147 $X2=0
+ $Y2=0
cc_325 N_A_27_297#_c_478_n N_VPWR_M1004_s 0.00333567f $X=4.775 $Y=1.917 $X2=0
+ $Y2=0
cc_326 N_A_27_297#_c_439_n N_VPWR_M1007_s 0.0071628f $X=5.38 $Y=1.915 $X2=0
+ $Y2=0
cc_327 N_A_27_297#_c_440_n N_VPWR_M1007_s 0.00791766f $X=5.465 $Y=1.83 $X2=0
+ $Y2=0
cc_328 N_A_27_297#_c_438_n N_VPWR_c_598_n 0.0180684f $X=1.23 $Y=1.917 $X2=0
+ $Y2=0
cc_329 N_A_27_297#_c_461_n N_VPWR_c_599_n 0.0122019f $X=1.795 $Y=1.917 $X2=0
+ $Y2=0
cc_330 N_A_27_297#_c_467_n N_VPWR_c_600_n 0.0163661f $X=2.695 $Y=2.147 $X2=0
+ $Y2=0
cc_331 N_A_27_297#_c_478_n N_VPWR_c_601_n 0.0160033f $X=4.775 $Y=1.917 $X2=0
+ $Y2=0
cc_332 N_A_27_297#_c_470_n N_VPWR_c_601_n 0.008955f $X=3.285 $Y=2.147 $X2=0
+ $Y2=0
cc_333 N_A_27_297#_M1007_g N_VPWR_c_602_n 0.00969206f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_334 N_A_27_297#_M1010_g N_VPWR_c_602_n 5.34447e-19 $X=6.05 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_27_297#_c_439_n N_VPWR_c_602_n 0.0207369f $X=5.38 $Y=1.915 $X2=0
+ $Y2=0
cc_336 N_A_27_297#_c_442_n N_VPWR_c_602_n 0.0234191f $X=4.9 $Y=1.96 $X2=0 $Y2=0
cc_337 N_A_27_297#_M1007_g N_VPWR_c_603_n 6.32056e-19 $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A_27_297#_M1010_g N_VPWR_c_603_n 0.0110282f $X=6.05 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A_27_297#_M1017_g N_VPWR_c_603_n 0.0102125f $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_27_297#_M1023_g N_VPWR_c_603_n 6.24225e-19 $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_27_297#_M1017_g N_VPWR_c_605_n 6.24498e-19 $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_27_297#_M1023_g N_VPWR_c_605_n 0.011324f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_343 N_A_27_297#_c_461_n N_VPWR_c_606_n 0.00220126f $X=1.795 $Y=1.917 $X2=0
+ $Y2=0
cc_344 N_A_27_297#_c_438_n N_VPWR_c_606_n 0.00166354f $X=1.23 $Y=1.917 $X2=0
+ $Y2=0
cc_345 N_A_27_297#_c_520_p N_VPWR_c_606_n 0.0129375f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_346 N_A_27_297#_c_461_n N_VPWR_c_608_n 0.00214376f $X=1.795 $Y=1.917 $X2=0
+ $Y2=0
cc_347 N_A_27_297#_c_465_n N_VPWR_c_608_n 0.0137286f $X=1.94 $Y=2.3 $X2=0 $Y2=0
cc_348 N_A_27_297#_c_467_n N_VPWR_c_608_n 0.0020345f $X=2.695 $Y=2.147 $X2=0
+ $Y2=0
cc_349 N_A_27_297#_c_437_n N_VPWR_c_610_n 0.0175447f $X=0.217 $Y=2.005 $X2=0
+ $Y2=0
cc_350 N_A_27_297#_c_438_n N_VPWR_c_610_n 0.00164067f $X=1.23 $Y=1.917 $X2=0
+ $Y2=0
cc_351 N_A_27_297#_c_478_n N_VPWR_c_611_n 0.00663483f $X=4.775 $Y=1.917 $X2=0
+ $Y2=0
cc_352 N_A_27_297#_c_467_n N_VPWR_c_611_n 0.0020345f $X=2.695 $Y=2.147 $X2=0
+ $Y2=0
cc_353 N_A_27_297#_c_470_n N_VPWR_c_611_n 0.0387224f $X=3.285 $Y=2.147 $X2=0
+ $Y2=0
cc_354 N_A_27_297#_c_478_n N_VPWR_c_612_n 0.00830426f $X=4.775 $Y=1.917 $X2=0
+ $Y2=0
cc_355 N_A_27_297#_c_439_n N_VPWR_c_612_n 0.00275452f $X=5.38 $Y=1.915 $X2=0
+ $Y2=0
cc_356 N_A_27_297#_c_442_n N_VPWR_c_612_n 0.0185484f $X=4.9 $Y=1.96 $X2=0 $Y2=0
cc_357 N_A_27_297#_M1007_g N_VPWR_c_613_n 0.0046653f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_358 N_A_27_297#_M1010_g N_VPWR_c_613_n 0.0046653f $X=6.05 $Y=1.985 $X2=0
+ $Y2=0
cc_359 N_A_27_297#_M1017_g N_VPWR_c_614_n 0.00505556f $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_360 N_A_27_297#_M1023_g N_VPWR_c_614_n 0.00505556f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_361 N_A_27_297#_M1002_d N_VPWR_c_597_n 0.00382897f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_362 N_A_27_297#_M1015_d N_VPWR_c_597_n 0.00384765f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_363 N_A_27_297#_M1016_s N_VPWR_c_597_n 0.00238028f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_364 N_A_27_297#_M1003_s N_VPWR_c_597_n 0.00516104f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_M1026_d N_VPWR_c_597_n 0.00212856f $X=4.765 $Y=1.485 $X2=0
+ $Y2=0
cc_366 N_A_27_297#_M1007_g N_VPWR_c_597_n 0.00789179f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_M1010_g N_VPWR_c_597_n 0.00789179f $X=6.05 $Y=1.985 $X2=0
+ $Y2=0
cc_368 N_A_27_297#_M1017_g N_VPWR_c_597_n 0.00850607f $X=6.47 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_M1023_g N_VPWR_c_597_n 0.00850607f $X=6.89 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_437_n N_VPWR_c_597_n 0.00972398f $X=0.217 $Y=2.005 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_461_n N_VPWR_c_597_n 0.00834033f $X=1.795 $Y=1.917 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_438_n N_VPWR_c_597_n 0.0066751f $X=1.23 $Y=1.917 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_465_n N_VPWR_c_597_n 0.00865145f $X=1.94 $Y=2.3 $X2=0 $Y2=0
cc_374 N_A_27_297#_c_478_n N_VPWR_c_597_n 0.0296029f $X=4.775 $Y=1.917 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_c_439_n N_VPWR_c_597_n 0.00605575f $X=5.38 $Y=1.915 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_c_520_p N_VPWR_c_597_n 0.00818828f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_377 N_A_27_297#_c_467_n N_VPWR_c_597_n 0.0090937f $X=2.695 $Y=2.147 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_c_470_n N_VPWR_c_597_n 0.022459f $X=3.285 $Y=2.147 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_c_442_n N_VPWR_c_597_n 0.0110612f $X=4.9 $Y=1.96 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_478_n A_681_297# 0.00473472f $X=4.775 $Y=1.917 $X2=-0.19
+ $Y2=-0.24
cc_381 N_A_27_297#_c_478_n A_852_297# 0.0070666f $X=4.775 $Y=1.917 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_27_297#_M1006_g N_X_c_738_n 0.00664399f $X=5.485 $Y=0.56 $X2=0 $Y2=0
cc_383 N_A_27_297#_M1013_g N_X_c_739_n 0.0123127f $X=5.99 $Y=0.56 $X2=0 $Y2=0
cc_384 N_A_27_297#_M1025_g N_X_c_739_n 0.012149f $X=6.425 $Y=0.56 $X2=0 $Y2=0
cc_385 N_A_27_297#_c_441_n N_X_c_739_n 0.0341798f $X=6.595 $Y=1.16 $X2=0 $Y2=0
cc_386 N_A_27_297#_c_432_n N_X_c_739_n 0.0026299f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A_27_297#_M1006_g N_X_c_743_n 0.0053072f $X=5.485 $Y=0.56 $X2=0 $Y2=0
cc_388 N_A_27_297#_c_441_n N_X_c_743_n 0.0146869f $X=6.595 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_27_297#_c_432_n N_X_c_743_n 0.00476923f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A_27_297#_M1010_g N_X_c_746_n 0.0136163f $X=6.05 $Y=1.985 $X2=0 $Y2=0
cc_391 N_A_27_297#_M1017_g N_X_c_746_n 0.0143544f $X=6.47 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A_27_297#_c_441_n N_X_c_746_n 0.0400225f $X=6.595 $Y=1.16 $X2=0 $Y2=0
cc_393 N_A_27_297#_c_432_n N_X_c_746_n 5.8591e-19 $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_394 N_A_27_297#_c_441_n N_X_c_750_n 0.0135068f $X=6.595 $Y=1.16 $X2=0 $Y2=0
cc_395 N_A_27_297#_c_432_n N_X_c_750_n 6.59861e-19 $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_396 N_A_27_297#_M1027_g N_X_c_752_n 0.0153866f $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_397 N_A_27_297#_M1023_g N_X_c_753_n 0.0178458f $X=6.89 $Y=1.985 $X2=0 $Y2=0
cc_398 N_A_27_297#_c_441_n N_X_c_754_n 0.0129079f $X=6.595 $Y=1.16 $X2=0 $Y2=0
cc_399 N_A_27_297#_c_432_n N_X_c_754_n 0.00288743f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_400 N_A_27_297#_c_441_n N_X_c_756_n 0.0137025f $X=6.595 $Y=1.16 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_432_n N_X_c_756_n 6.64183e-19 $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_402 N_A_27_297#_M1027_g X 0.00648664f $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_403 N_A_27_297#_c_441_n X 0.0153604f $X=6.595 $Y=1.16 $X2=0 $Y2=0
cc_404 N_A_27_297#_c_432_n X 0.0172713f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_405 N_A_27_297#_M1009_s N_A_27_47#_c_791_n 0.00305588f $X=0.545 $Y=0.235
+ $X2=0 $Y2=0
cc_406 N_A_27_297#_c_444_n N_A_27_47#_c_791_n 0.0176071f $X=0.68 $Y=0.76 $X2=0
+ $Y2=0
cc_407 N_A_27_297#_M1006_g N_VGND_c_873_n 0.00632033f $X=5.485 $Y=0.56 $X2=0
+ $Y2=0
cc_408 N_A_27_297#_M1013_g N_VGND_c_874_n 0.00310297f $X=5.99 $Y=0.56 $X2=0
+ $Y2=0
cc_409 N_A_27_297#_M1025_g N_VGND_c_874_n 0.00685754f $X=6.425 $Y=0.56 $X2=0
+ $Y2=0
cc_410 N_A_27_297#_M1027_g N_VGND_c_874_n 5.12898e-19 $X=6.87 $Y=0.56 $X2=0
+ $Y2=0
cc_411 N_A_27_297#_M1025_g N_VGND_c_876_n 5.22966e-19 $X=6.425 $Y=0.56 $X2=0
+ $Y2=0
cc_412 N_A_27_297#_M1027_g N_VGND_c_876_n 0.00851608f $X=6.87 $Y=0.56 $X2=0
+ $Y2=0
cc_413 N_A_27_297#_M1006_g N_VGND_c_883_n 0.00585385f $X=5.485 $Y=0.56 $X2=0
+ $Y2=0
cc_414 N_A_27_297#_M1013_g N_VGND_c_883_n 0.00433717f $X=5.99 $Y=0.56 $X2=0
+ $Y2=0
cc_415 N_A_27_297#_M1025_g N_VGND_c_884_n 0.00360664f $X=6.425 $Y=0.56 $X2=0
+ $Y2=0
cc_416 N_A_27_297#_M1027_g N_VGND_c_884_n 0.00346207f $X=6.87 $Y=0.56 $X2=0
+ $Y2=0
cc_417 N_A_27_297#_M1009_s N_VGND_c_886_n 0.00216833f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_418 N_A_27_297#_M1006_g N_VGND_c_886_n 0.0114418f $X=5.485 $Y=0.56 $X2=0
+ $Y2=0
cc_419 N_A_27_297#_M1013_g N_VGND_c_886_n 0.00596108f $X=5.99 $Y=0.56 $X2=0
+ $Y2=0
cc_420 N_A_27_297#_M1025_g N_VGND_c_886_n 0.00427414f $X=6.425 $Y=0.56 $X2=0
+ $Y2=0
cc_421 N_A_27_297#_M1027_g N_VGND_c_886_n 0.0041266f $X=6.87 $Y=0.56 $X2=0 $Y2=0
cc_422 N_VPWR_c_597_n A_681_297# 0.00353442f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_423 N_VPWR_c_597_n A_852_297# 0.00456261f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_424 N_VPWR_c_597_n N_X_M1007_d 0.00562358f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_425 N_VPWR_c_597_n N_X_M1017_d 0.00492927f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_426 N_VPWR_c_613_n N_X_c_763_n 0.0113958f $X=6.095 $Y=2.72 $X2=0 $Y2=0
cc_427 N_VPWR_c_597_n N_X_c_763_n 0.00646998f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_M1010_s N_X_c_746_n 0.00313971f $X=6.125 $Y=1.485 $X2=0 $Y2=0
cc_429 N_VPWR_c_603_n N_X_c_746_n 0.0162641f $X=6.26 $Y=2 $X2=0 $Y2=0
cc_430 N_VPWR_c_614_n N_X_c_767_n 0.0121054f $X=6.945 $Y=2.72 $X2=0 $Y2=0
cc_431 N_VPWR_c_597_n N_X_c_767_n 0.00724021f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_432 N_VPWR_c_605_n N_X_c_753_n 0.00140521f $X=7.1 $Y=2 $X2=0 $Y2=0
cc_433 N_VPWR_M1023_s N_X_c_737_n 0.00299921f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_434 N_VPWR_c_605_n N_X_c_737_n 0.0224255f $X=7.1 $Y=2 $X2=0 $Y2=0
cc_435 N_X_c_739_n N_VGND_M1013_s 0.00348735f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_436 X N_VGND_M1027_s 3.26185e-19 $X=7.045 $Y=0.765 $X2=0 $Y2=0
cc_437 N_X_c_735_n N_VGND_M1027_s 0.00330652f $X=7.14 $Y=0.865 $X2=0 $Y2=0
cc_438 N_X_c_738_n N_VGND_c_873_n 0.0130652f $X=5.78 $Y=0.42 $X2=0 $Y2=0
cc_439 N_X_c_739_n N_VGND_c_874_n 0.0149821f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_440 N_X_c_752_n N_VGND_c_876_n 0.00219925f $X=7.005 $Y=0.78 $X2=0 $Y2=0
cc_441 N_X_c_735_n N_VGND_c_876_n 0.023242f $X=7.14 $Y=0.865 $X2=0 $Y2=0
cc_442 N_X_c_738_n N_VGND_c_883_n 0.0150088f $X=5.78 $Y=0.42 $X2=0 $Y2=0
cc_443 N_X_c_739_n N_VGND_c_883_n 0.00255372f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_444 N_X_c_739_n N_VGND_c_884_n 0.00215462f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_445 N_X_c_782_p N_VGND_c_884_n 0.0132304f $X=6.64 $Y=0.42 $X2=0 $Y2=0
cc_446 N_X_c_752_n N_VGND_c_884_n 0.00212504f $X=7.005 $Y=0.78 $X2=0 $Y2=0
cc_447 N_X_M1006_d N_VGND_c_886_n 0.00617019f $X=5.56 $Y=0.235 $X2=0 $Y2=0
cc_448 N_X_M1025_d N_VGND_c_886_n 0.0027576f $X=6.5 $Y=0.235 $X2=0 $Y2=0
cc_449 N_X_c_738_n N_VGND_c_886_n 0.00856376f $X=5.78 $Y=0.42 $X2=0 $Y2=0
cc_450 N_X_c_739_n N_VGND_c_886_n 0.00971708f $X=6.545 $Y=0.78 $X2=0 $Y2=0
cc_451 N_X_c_782_p N_VGND_c_886_n 0.00760369f $X=6.64 $Y=0.42 $X2=0 $Y2=0
cc_452 N_X_c_752_n N_VGND_c_886_n 0.00432648f $X=7.005 $Y=0.78 $X2=0 $Y2=0
cc_453 N_X_c_735_n N_VGND_c_886_n 0.00122142f $X=7.14 $Y=0.865 $X2=0 $Y2=0
cc_454 N_A_27_47#_c_791_n A_445_47# 0.00753415f $X=2.72 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_455 N_A_27_47#_c_791_n N_A_361_47#_M1020_d 0.0030596f $X=2.72 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_456 N_A_27_47#_M1014_s N_A_361_47#_c_821_n 0.00565317f $X=2.585 $Y=0.235
+ $X2=0 $Y2=0
cc_457 N_A_27_47#_c_791_n N_A_361_47#_c_821_n 0.065996f $X=2.72 $Y=0.38 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_791_n A_277_47# 0.00194265f $X=2.72 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_459 N_A_27_47#_c_791_n N_VGND_c_871_n 0.0201689f $X=2.72 $Y=0.38 $X2=0 $Y2=0
cc_460 N_A_27_47#_c_791_n N_VGND_c_877_n 0.14622f $X=2.72 $Y=0.38 $X2=0 $Y2=0
cc_461 N_A_27_47#_c_792_n N_VGND_c_877_n 0.0168179f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_462 N_A_27_47#_M1009_d N_VGND_c_886_n 0.00209324f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_M1024_d N_VGND_c_886_n 0.00215227f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_M1014_s N_VGND_c_886_n 0.00209344f $X=2.585 $Y=0.235 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_791_n N_VGND_c_886_n 0.0928998f $X=2.72 $Y=0.38 $X2=0 $Y2=0
cc_466 N_A_27_47#_c_792_n N_VGND_c_886_n 0.00939253f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_467 A_445_47# N_VGND_c_886_n 0.00216833f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_468 N_A_361_47#_c_821_n A_277_47# 0.00293715f $X=3.61 $Y=0.77 $X2=-0.19
+ $Y2=-0.24
cc_469 N_A_361_47#_c_821_n N_VGND_M1018_d 0.0048535f $X=3.61 $Y=0.77 $X2=-0.19
+ $Y2=-0.24
cc_470 N_A_361_47#_c_836_n N_VGND_M1001_d 0.00313435f $X=4.535 $Y=0.77 $X2=0
+ $Y2=0
cc_471 N_A_361_47#_c_821_n N_VGND_c_871_n 0.0211503f $X=3.61 $Y=0.77 $X2=0 $Y2=0
cc_472 N_A_361_47#_c_836_n N_VGND_c_872_n 0.0193182f $X=4.535 $Y=0.77 $X2=0
+ $Y2=0
cc_473 N_A_361_47#_c_854_p N_VGND_c_872_n 0.0176835f $X=4.63 $Y=0.42 $X2=0 $Y2=0
cc_474 N_A_361_47#_c_821_n N_VGND_c_877_n 0.0030357f $X=3.61 $Y=0.77 $X2=0 $Y2=0
cc_475 N_A_361_47#_c_821_n N_VGND_c_879_n 0.00235985f $X=3.61 $Y=0.77 $X2=0
+ $Y2=0
cc_476 N_A_361_47#_c_857_p N_VGND_c_879_n 0.0144814f $X=3.74 $Y=0.42 $X2=0 $Y2=0
cc_477 N_A_361_47#_c_836_n N_VGND_c_879_n 0.00235985f $X=4.535 $Y=0.77 $X2=0
+ $Y2=0
cc_478 N_A_361_47#_c_836_n N_VGND_c_881_n 0.00234422f $X=4.535 $Y=0.77 $X2=0
+ $Y2=0
cc_479 N_A_361_47#_c_854_p N_VGND_c_881_n 0.0168014f $X=4.63 $Y=0.42 $X2=0 $Y2=0
cc_480 N_A_361_47#_M1020_d N_VGND_c_886_n 0.00216833f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_481 N_A_361_47#_M1018_s N_VGND_c_886_n 0.00288323f $X=3.56 $Y=0.235 $X2=0
+ $Y2=0
cc_482 N_A_361_47#_M1005_s N_VGND_c_886_n 0.00402052f $X=4.445 $Y=0.235 $X2=0
+ $Y2=0
cc_483 N_A_361_47#_c_821_n N_VGND_c_886_n 0.0127334f $X=3.61 $Y=0.77 $X2=0 $Y2=0
cc_484 N_A_361_47#_c_857_p N_VGND_c_886_n 0.00818659f $X=3.74 $Y=0.42 $X2=0
+ $Y2=0
cc_485 N_A_361_47#_c_836_n N_VGND_c_886_n 0.0101303f $X=4.535 $Y=0.77 $X2=0
+ $Y2=0
cc_486 N_A_361_47#_c_854_p N_VGND_c_886_n 0.00991615f $X=4.63 $Y=0.42 $X2=0
+ $Y2=0
cc_487 A_277_47# N_VGND_c_886_n 0.00168648f $X=2.225 $Y=0.235 $X2=0 $Y2=0

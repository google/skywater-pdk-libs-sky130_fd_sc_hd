* File: sky130_fd_sc_hd__a222oi_1.pex.spice
* Created: Thu Aug 27 14:02:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A222OI_1%C1 3 6 8 11 12 13 16
r30 11 14 46.6684 $w=4.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.325 $Y=1.165
+ $X2=0.325 $Y2=1.33
r31 11 13 46.6684 $w=4.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.325 $Y=1.165
+ $X2=0.325 $Y2=1
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.38
+ $Y=1.165 $X2=0.38 $Y2=1.165
r33 8 12 5.12197 $w=3.13e-07 $l=1.4e-07 $layer=LI1_cond $X=0.24 $Y=1.157
+ $X2=0.38 $Y2=1.157
r34 8 16 0.548782 $w=3.13e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=1.157
+ $X2=0.225 $Y2=1.157
r35 6 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.33
r36 3 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.47 $Y=0.555
+ $X2=0.47 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%C2 3 6 8 11 13
c34 6 0 1.04686e-19 $X=0.89 $Y=1.985
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.165
+ $X2=0.89 $Y2=1
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.165 $X2=0.89 $Y2=1.165
r37 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.33
+ $X2=0.89 $Y2=1.165
r38 4 6 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.33 $X2=0.89
+ $Y2=1.985
r39 3 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.83 $Y=0.555
+ $X2=0.83 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%B2 3 6 8 11 13
r35 11 14 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.165
+ $X2=1.81 $Y2=1.33
r36 11 13 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.165
+ $X2=1.81 $Y2=1
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.165 $X2=1.82 $Y2=1.165
r38 6 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=1.89 $Y=1.985
+ $X2=1.89 $Y2=1.33
r39 3 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.89 $Y=0.555
+ $X2=1.89 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%B1 3 6 8 11 13
c33 11 0 2.04008e-19 $X=2.31 $Y=1.165
c34 8 0 6.28217e-20 $X=2.31 $Y=1.175
c35 6 0 8.31507e-20 $X=2.31 $Y=1.985
r36 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.165
+ $X2=2.31 $Y2=1
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.165 $X2=2.31 $Y2=1.165
r38 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.33
+ $X2=2.31 $Y2=1.165
r39 4 6 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.31 $Y=1.33 $X2=2.31
+ $Y2=1.985
r40 3 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.25 $Y=0.555
+ $X2=2.25 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%A1 3 6 8 11 13
r32 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.165
+ $X2=2.79 $Y2=1.33
r33 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.165
+ $X2=2.79 $Y2=1
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.165 $X2=2.79 $Y2=1.165
r35 6 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.73 $Y=1.985
+ $X2=2.73 $Y2=1.33
r36 3 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.73 $Y=0.555
+ $X2=2.73 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%A2 3 6 8 11 13
c25 6 0 1.97589e-19 $X=3.21 $Y=1.985
r26 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.165
+ $X2=3.27 $Y2=1.33
r27 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.165
+ $X2=3.27 $Y2=1
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.165 $X2=3.27 $Y2=1.165
r29 6 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=3.21 $Y=1.985
+ $X2=3.21 $Y2=1.33
r30 3 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.21 $Y=0.555
+ $X2=3.21 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%Y 1 2 3 4 15 17 19 20 21 24 25 29 34 35 38
+ 41 42 48
c78 42 0 6.9407e-20 $X=1.255 $Y=1.09
c79 17 0 1.04686e-19 $X=0.22 $Y=1.68
r80 45 48 2.20245 $w=2.23e-07 $l=4.3e-08 $layer=LI1_cond $X=1.367 $Y=1.218
+ $X2=1.367 $Y2=1.175
r81 42 50 5.3766 $w=2.23e-07 $l=9.1e-08 $layer=LI1_cond $X=1.367 $Y=1.239
+ $X2=1.367 $Y2=1.33
r82 42 45 1.07561 $w=2.23e-07 $l=2.1e-08 $layer=LI1_cond $X=1.367 $Y=1.239
+ $X2=1.367 $Y2=1.218
r83 42 48 1.07561 $w=2.23e-07 $l=2.1e-08 $layer=LI1_cond $X=1.367 $Y=1.154
+ $X2=1.367 $Y2=1.175
r84 40 42 17.3635 $w=2.23e-07 $l=3.39e-07 $layer=LI1_cond $X=1.367 $Y=0.815
+ $X2=1.367 $Y2=1.154
r85 40 41 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.367 $Y=0.815
+ $X2=1.367 $Y2=0.73
r86 38 39 12.4068 $w=2.36e-07 $l=2.4e-07 $layer=LI1_cond $X=1.1 $Y=1.665
+ $X2=1.34 $Y2=1.665
r87 34 35 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.34
+ $X2=0.26 $Y2=2.255
r88 27 29 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.48 $Y=0.645
+ $X2=2.48 $Y2=0.38
r89 26 41 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.48 $Y=0.73
+ $X2=1.367 $Y2=0.73
r90 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.315 $Y=0.73
+ $X2=2.48 $Y2=0.645
r91 25 26 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.315 $Y=0.73
+ $X2=1.48 $Y2=0.73
r92 24 39 2.65936 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=1.5 $X2=1.34
+ $Y2=1.665
r93 24 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.34 $Y=1.5 $X2=1.34
+ $Y2=1.33
r94 22 32 3.92174 $w=1.7e-07 $l=1.66493e-07 $layer=LI1_cond $X=0.425 $Y=1.585
+ $X2=0.26 $Y2=1.582
r95 21 38 5.36806 $w=2.36e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.015 $Y=1.585
+ $X2=1.1 $Y2=1.665
r96 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.015 $Y=1.585
+ $X2=0.425 $Y2=1.585
r97 19 41 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.255 $Y=0.73
+ $X2=1.367 $Y2=0.73
r98 19 20 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.255 $Y=0.73
+ $X2=0.425 $Y2=0.73
r99 17 32 3.22143 $w=2.5e-07 $l=1.16293e-07 $layer=LI1_cond $X=0.22 $Y=1.68
+ $X2=0.26 $Y2=1.582
r100 17 35 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=0.22 $Y=1.68
+ $X2=0.22 $Y2=2.255
r101 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.645
+ $X2=0.425 $Y2=0.73
r102 13 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.26 $Y=0.645
+ $X2=0.26 $Y2=0.38
r103 4 38 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.665
r104 3 34 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r105 3 32 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
r106 2 29 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.235 $X2=2.48 $Y2=0.38
r107 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%A_109_297# 1 2 8 9 12 17
r26 10 15 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.38
+ $X2=0.68 $Y2=2.38
r27 9 17 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.015 $Y=2.38
+ $X2=2.1 $Y2=2.3
r28 9 10 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.015 $Y=2.38
+ $X2=0.765 $Y2=2.38
r29 8 15 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.295 $X2=0.68
+ $Y2=2.38
r30 7 12 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.68 $Y=2.075
+ $X2=0.68 $Y2=1.96
r31 7 8 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.68 $Y=2.075 $X2=0.68
+ $Y2=2.295
r32 2 17 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.485 $X2=2.1 $Y2=2.3
r33 1 15 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.3
r34 1 12 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%A_311_297# 1 2 3 10 14 16 19 25 26 33 37 38
+ 41
c48 26 0 8.31507e-20 $X=1.93 $Y=1.74
c49 16 0 1.97589e-19 $X=2.48 $Y=1.825
c50 14 0 1.97423e-19 $X=2.355 $Y=1.74
r51 41 42 3.54783 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=2.34
+ $X2=3.425 $Y2=2.255
r52 37 38 10.7092 $w=2.33e-07 $l=2e-07 $layer=LI1_cond $X=3.42 $Y=1.617 $X2=3.22
+ $Y2=1.617
r53 33 34 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.34
+ $X2=2.52 $Y2=2.255
r54 30 31 3.57655 $w=3.07e-07 $l=9e-08 $layer=LI1_cond $X=2.52 $Y=1.65 $X2=2.52
+ $Y2=1.74
r55 28 30 2.58306 $w=3.07e-07 $l=6.5e-08 $layer=LI1_cond $X=2.52 $Y=1.585
+ $X2=2.52 $Y2=1.65
r56 26 27 12.8025 $w=1.62e-07 $l=1.7e-07 $layer=LI1_cond $X=1.93 $Y=1.74
+ $X2=1.93 $Y2=1.91
r57 25 42 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=3.465 $Y=1.995
+ $X2=3.465 $Y2=2.255
r58 22 37 0.0901955 $w=2.6e-07 $l=1.38687e-07 $layer=LI1_cond $X=3.465 $Y=1.735
+ $X2=3.42 $Y2=1.617
r59 22 25 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=3.465 $Y=1.735
+ $X2=3.465 $Y2=1.995
r60 21 28 4.19673 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=1.585
+ $X2=2.52 $Y2=1.585
r61 21 38 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.685 $Y=1.585
+ $X2=3.22 $Y2=1.585
r62 19 34 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.48 $Y=1.995
+ $X2=2.48 $Y2=2.255
r63 16 31 3.83435 $w=3.07e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.48 $Y=1.825
+ $X2=2.52 $Y2=1.74
r64 16 19 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.48 $Y=1.825
+ $X2=2.48 $Y2=1.995
r65 15 26 0.420406 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=1.74
+ $X2=1.93 $Y2=1.74
r66 14 31 4.19673 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=1.74
+ $X2=2.52 $Y2=1.74
r67 14 15 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.355 $Y=1.74
+ $X2=2.015 $Y2=1.74
r68 10 27 0.420406 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=1.91
+ $X2=1.93 $Y2=1.91
r69 10 12 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=1.91
+ $X2=1.68 $Y2=1.91
r70 3 41 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=2.34
r71 3 37 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.65
r72 3 25 600 $w=1.7e-07 $l=5.73542e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.995
r73 2 33 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.485 $X2=2.52 $Y2=2.34
r74 2 30 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.485 $X2=2.52 $Y2=1.65
r75 2 19 600 $w=1.7e-07 $l=5.73542e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.485 $X2=2.52 $Y2=1.995
r76 1 12 600 $w=1.7e-07 $l=4.83477e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.485 $X2=1.68 $Y2=1.91
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%VPWR 1 7 9 12 13 14 24 25 31
r45 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 22 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 22 31 0.170725 $w=4.8e-07 $l=6e-07 $layer=MET1_cond $X=2.53 $Y=2.72 $X2=1.93
+ $Y2=2.72
r48 21 22 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 17 21 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 17 18 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 14 31 0.0256088 $w=4.8e-07 $l=9e-08 $layer=MET1_cond $X=1.84 $Y=2.72
+ $X2=1.93 $Y2=2.72
r52 14 18 0.458112 $w=4.8e-07 $l=1.61e-06 $layer=MET1_cond $X=1.84 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 12 21 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.855 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 12 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=2.72
+ $X2=2.94 $Y2=2.72
r55 11 24 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.025 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 11 13 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=2.72
+ $X2=2.94 $Y2=2.72
r57 5 13 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=2.635 $X2=2.94
+ $Y2=2.72
r58 5 7 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.94 $Y=2.635 $X2=2.94
+ $Y2=2.34
r59 4 9 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=2.075 $X2=2.94
+ $Y2=1.99
r60 4 7 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.94 $Y=2.075
+ $X2=2.94 $Y2=2.34
r61 1 9 600 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.485 $X2=2.94 $Y2=1.99
r62 1 7 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.485 $X2=2.94 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A222OI_1%VGND 1 2 7 9 11 18 29 32 35 42
r47 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r48 31 32 11.1368 $w=5.48e-07 $l=2.25e-07 $layer=LI1_cond $X=1.38 $Y=0.19
+ $X2=1.605 $Y2=0.19
r49 27 31 5.00178 $w=5.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.15 $Y=0.19
+ $X2=1.38 $Y2=0.19
r50 27 29 12.2241 $w=5.48e-07 $l=2.75e-07 $layer=LI1_cond $X=1.15 $Y=0.19
+ $X2=0.875 $Y2=0.19
r51 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r52 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r53 25 42 0.23617 $w=4.8e-07 $l=8.3e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.16
+ $Y2=0
r54 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r56 21 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r57 21 32 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.605
+ $Y2=0
r58 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r59 18 34 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.467
+ $Y2=0
r60 18 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=2.99
+ $Y2=0
r61 16 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r62 15 29 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=0.875
+ $Y2=0
r63 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r64 11 42 0.0910533 $w=4.8e-07 $l=3.2e-07 $layer=MET1_cond $X=1.84 $Y=0 $X2=2.16
+ $Y2=0
r65 11 22 0.0654446 $w=4.8e-07 $l=2.3e-07 $layer=MET1_cond $X=1.84 $Y=0 $X2=1.61
+ $Y2=0
r66 7 34 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.467 $Y2=0
r67 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.38
r68 2 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.38
r69 1 31 91 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_NDIFF $count=2 $X=0.905
+ $Y=0.235 $X2=1.38 $Y2=0.38
.ends


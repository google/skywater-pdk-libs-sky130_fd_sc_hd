* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
M1000 Y A KAPWR VPB phighvt w=1e+06u l=150000u
+  ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u
M1001 KAPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nshort w=420000u l=150000u
+  ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u
M1003 VGND A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 KAPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A KAPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 KAPWR A Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A KAPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__ebufn_1.spice.pex
* Created: Thu Aug 27 14:19:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EBUFN_1%A 3 7 9 10 17
r27 14 17 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.27 $Y=1.16 $X2=0.47
+ $Y2=1.16
r28 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.16 $X2=0.22
+ $Y2=1.53
r29 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r30 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r31 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.165
r32 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r33 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_1%TE_B 3 5 7 10 13 14 15 16
r49 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.075 $Y=1.16
+ $X2=1.075 $Y2=1.53
r50 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.16 $X2=1.075 $Y2=1.16
r51 14 20 120.654 $w=3.3e-07 $l=6.9e-07 $layer=POLY_cond $X=1.765 $Y=1.16
+ $X2=1.075 $Y2=1.16
r52 12 20 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.05 $Y=1.16
+ $X2=1.075 $Y2=1.16
r53 12 13 5.03009 $w=3.3e-07 $l=1.18e-07 $layer=POLY_cond $X=1.05 $Y=1.16
+ $X2=0.932 $Y2=1.16
r54 8 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.765 $Y2=1.16
r55 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.985
r56 5 13 37.0704 $w=1.5e-07 $l=1.85257e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.932 $Y2=1.16
r57 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=0.675
r58 1 13 37.0704 $w=1.5e-07 $l=1.84811e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.932 $Y2=1.16
r59 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_1%A_193_369# 1 2 7 9 12 15 17 20 28 31 34
c56 20 0 1.89939e-19 $X=2.37 $Y=1.16
r57 28 30 4.71941 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.52 $Y=0.76
+ $X2=1.52 $Y2=0.885
r58 21 34 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.37 $Y=1.16
+ $X2=2.58 $Y2=1.16
r59 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.16 $X2=2.37 $Y2=1.16
r60 18 31 2.41475 $w=2.5e-07 $l=1.98e-07 $layer=LI1_cond $X=1.805 $Y=1.2
+ $X2=1.607 $Y2=1.2
r61 18 20 26.0452 $w=2.48e-07 $l=5.65e-07 $layer=LI1_cond $X=1.805 $Y=1.2
+ $X2=2.37 $Y2=1.2
r62 16 31 4.02345 $w=3.35e-07 $l=1.25e-07 $layer=LI1_cond $X=1.607 $Y=1.325
+ $X2=1.607 $Y2=1.2
r63 16 17 13.8585 $w=3.93e-07 $l=4.75e-07 $layer=LI1_cond $X=1.607 $Y=1.325
+ $X2=1.607 $Y2=1.8
r64 15 31 4.02345 $w=3.35e-07 $l=1.52069e-07 $layer=LI1_cond $X=1.547 $Y=1.075
+ $X2=1.607 $Y2=1.2
r65 15 30 7.96233 $w=2.73e-07 $l=1.9e-07 $layer=LI1_cond $X=1.547 $Y=1.075
+ $X2=1.547 $Y2=0.885
r66 10 17 25.1574 $w=2.03e-07 $l=4.65e-07 $layer=LI1_cond $X=1.142 $Y=1.902
+ $X2=1.607 $Y2=1.902
r67 10 12 11.7504 $w=2.53e-07 $l=2.6e-07 $layer=LI1_cond $X=1.142 $Y=2.005
+ $X2=1.142 $Y2=2.265
r68 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=0.995
+ $X2=2.58 $Y2=1.16
r69 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.58 $Y=0.995 $X2=2.58
+ $Y2=0.56
r70 2 12 600 $w=1.7e-07 $l=4.82804e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.845 $X2=1.1 $Y2=2.265
r71 1 28 182 $w=1.7e-07 $l=5.99625e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.465 $X2=1.52 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_1%A_27_47# 1 2 9 12 16 20 23 24 25 27 28 29 31
+ 32 33 39 41 44 46
c111 44 0 1.89939e-19 $X=3 $Y=1.16
r112 44 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3 $Y=1.16 $X2=3
+ $Y2=1.325
r113 44 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3 $Y=1.16 $X2=3
+ $Y2=0.995
r114 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=1.16
+ $X2=3 $Y2=1.16
r115 41 43 12.882 $w=3.22e-07 $l=3.4e-07 $layer=LI1_cond $X=2.895 $Y=0.82
+ $X2=2.895 $Y2=1.16
r116 32 41 4.47834 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.705 $Y=0.82
+ $X2=2.895 $Y2=0.82
r117 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.705 $Y=0.82
+ $X2=2.025 $Y2=0.82
r118 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=0.735
+ $X2=2.025 $Y2=0.82
r119 30 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.94 $Y=0.465
+ $X2=1.94 $Y2=0.735
r120 28 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.855 $Y=0.36
+ $X2=1.94 $Y2=0.465
r121 28 29 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=0.36
+ $X2=1.185 $Y2=0.36
r122 26 29 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.1 $Y=0.465
+ $X2=1.185 $Y2=0.36
r123 26 27 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.1 $Y=0.465 $X2=1.1
+ $Y2=0.615
r124 25 36 5.7039 $w=2.08e-07 $l=1.08e-07 $layer=LI1_cond $X=0.74 $Y=0.72
+ $X2=0.632 $Y2=0.72
r125 24 27 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.015 $Y=0.72
+ $X2=1.1 $Y2=0.615
r126 24 25 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.015 $Y=0.72
+ $X2=0.74 $Y2=0.72
r127 23 39 0.884026 $w=2.15e-07 $l=1.1e-07 $layer=LI1_cond $X=0.632 $Y=1.785
+ $X2=0.632 $Y2=1.895
r128 22 36 0.601528 $w=2.15e-07 $l=1.05e-07 $layer=LI1_cond $X=0.632 $Y=0.825
+ $X2=0.632 $Y2=0.72
r129 22 23 51.4579 $w=2.13e-07 $l=9.6e-07 $layer=LI1_cond $X=0.632 $Y=0.825
+ $X2=0.632 $Y2=1.785
r130 18 39 21.844 $w=2.18e-07 $l=4.17e-07 $layer=LI1_cond $X=0.215 $Y=1.895
+ $X2=0.632 $Y2=1.895
r131 18 20 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.215 $Y=2.005
+ $X2=0.215 $Y2=2.22
r132 14 36 22.0234 $w=2.08e-07 $l=4.17e-07 $layer=LI1_cond $X=0.215 $Y=0.72
+ $X2=0.632 $Y2=0.72
r133 14 16 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.445
r134 12 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.94 $Y=1.985
+ $X2=2.94 $Y2=1.325
r135 9 46 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.94 $Y=0.56
+ $X2=2.94 $Y2=0.995
r136 2 20 600 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.22
r137 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_1%VPWR 1 2 9 13 15 17 22 32 33 36 39
r43 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 30 33 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 29 32 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r49 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 27 39 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.622 $Y2=2.72
r51 27 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r56 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 22 39 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.622 $Y2=2.72
r58 22 25 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.44 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r60 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r61 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 11 39 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.622 $Y=2.635
+ $X2=1.622 $Y2=2.72
r64 11 13 11.8402 $w=3.63e-07 $l=3.75e-07 $layer=LI1_cond $X=1.622 $Y=2.635
+ $X2=1.622 $Y2=2.26
r65 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.72
r66 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.36
r67 2 13 600 $w=1.7e-07 $l=8.35165e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.485 $X2=1.62 $Y2=2.26
r68 1 9 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_1%Z 1 2 7 9 11 13 14 15 16 33 47 49 55
r30 49 60 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=3.425 $Y=0.85
+ $X2=3.425 $Y2=0.825
r31 33 45 0.628866 $w=9.68e-07 $l=5e-08 $layer=LI1_cond $X=3.255 $Y=1.98
+ $X2=3.205 $Y2=1.98
r32 16 47 6.74114 $w=3.4e-07 $l=4.85e-07 $layer=LI1_cond $X=3.425 $Y=1.98
+ $X2=3.425 $Y2=1.495
r33 16 33 2.36288 $w=9.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.425 $Y=1.98
+ $X2=3.255 $Y2=1.98
r34 16 47 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=3.425 $Y=1.47
+ $X2=3.425 $Y2=1.495
r35 15 16 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=3.425 $Y=1.19
+ $X2=3.425 $Y2=1.47
r36 14 60 1.69879 $w=4.68e-07 $l=3e-08 $layer=LI1_cond $X=3.36 $Y=0.795 $X2=3.36
+ $Y2=0.825
r37 14 15 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=3.425 $Y=0.88
+ $X2=3.425 $Y2=1.19
r38 14 49 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=3.425 $Y=0.88
+ $X2=3.425 $Y2=0.85
r39 13 14 7.25282 $w=4.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.36 $Y=0.51
+ $X2=3.36 $Y2=0.795
r40 13 55 3.81727 $w=4.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.36 $Y=0.51
+ $X2=3.36 $Y2=0.36
r41 11 45 2.64124 $w=9.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.995 $Y=1.98
+ $X2=3.205 $Y2=1.98
r42 9 11 5.78557 $w=9.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.98
+ $X2=2.995 $Y2=1.98
r43 7 9 5.78557 $w=9.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.075 $Y=1.98
+ $X2=2.535 $Y2=1.98
r44 2 45 300 $w=1.7e-07 $l=4.14246e-07 $layer=licon1_PDIFF $count=2 $X=3.015
+ $Y=1.485 $X2=3.205 $Y2=1.815
r45 1 55 91 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=2 $X=3.015
+ $Y=0.235 $X2=3.29 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__EBUFN_1%VGND 1 2 9 11 13 28 29 32 36 40
r46 38 40 15.2662 $w=6.48e-07 $l=4.25e-07 $layer=LI1_cond $X=2.53 $Y=0.24
+ $X2=2.955 $Y2=0.24
r47 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r48 35 38 4.6003 $w=6.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.28 $Y=0.24 $X2=2.53
+ $Y2=0.24
r49 35 36 9.00983 $w=6.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.24
+ $X2=2.195 $Y2=0.24
r50 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 29 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r52 28 40 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.955
+ $Y2=0
r53 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r54 25 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r55 24 36 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.195
+ $Y2=0
r56 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r57 22 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r58 22 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r59 21 24 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r60 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 19 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r62 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r63 13 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r64 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r65 11 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r66 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r67 7 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r68 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r69 2 35 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.28 $Y2=0.38
r70 1 9 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


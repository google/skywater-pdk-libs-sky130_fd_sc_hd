* File: sky130_fd_sc_hd__nand3b_1.spice.pex
* Created: Thu Aug 27 14:29:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND3B_1%A_N 3 6 8 11 13
r30 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r31 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r33 8 12 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.51
+ $Y2=1.16
r34 6 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.6 $Y=1.695 $X2=0.6
+ $Y2=1.325
r35 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.6 $Y=0.675 $X2=0.6
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_1%C 3 6 8 11 13
r31 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.16
+ $X2=1.05 $Y2=1.325
r32 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.16
+ $X2=1.05 $Y2=0.995
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r34 8 12 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.15 $Y=1.16 $X2=1.05
+ $Y2=1.16
r35 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.085 $Y=1.985
+ $X2=1.085 $Y2=1.325
r36 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.085 $Y=0.56
+ $X2=1.085 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_1%B 3 6 8 11 13
r36 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.16
+ $X2=1.59 $Y2=1.325
r37 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.16
+ $X2=1.59 $Y2=0.995
r38 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.59
+ $Y=1.16 $X2=1.59 $Y2=1.16
r39 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.505 $Y=1.985
+ $X2=1.505 $Y2=1.325
r40 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.505 $Y=0.56
+ $X2=1.505 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_1%A_53_93# 1 2 9 12 15 16 20 21 27 31 34
r71 28 31 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.17 $Y=1.76
+ $X2=0.39 $Y2=1.76
r72 26 27 7.20646 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=0.39 $Y=0.635
+ $X2=0.51 $Y2=0.635
r73 23 26 6.67204 $w=3.78e-07 $l=2.2e-07 $layer=LI1_cond $X=0.17 $Y=0.635
+ $X2=0.39 $Y2=0.635
r74 21 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.16
+ $X2=2.13 $Y2=1.325
r75 21 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.16
+ $X2=2.13 $Y2=0.995
r76 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.16 $X2=2.13 $Y2=1.16
r77 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.13 $Y=0.825
+ $X2=2.13 $Y2=1.16
r78 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=0.74
+ $X2=2.13 $Y2=0.825
r79 16 27 100.144 $w=1.68e-07 $l=1.535e-06 $layer=LI1_cond $X=2.045 $Y=0.74
+ $X2=0.51 $Y2=0.74
r80 15 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=1.595
+ $X2=0.17 $Y2=1.76
r81 14 23 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.635
r82 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.595
r83 12 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.04 $Y=1.985
+ $X2=2.04 $Y2=1.325
r84 9 34 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.04 $Y=0.56 $X2=2.04
+ $Y2=0.995
r85 2 31 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.485 $X2=0.39 $Y2=1.76
r86 1 26 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.265
+ $Y=0.465 $X2=0.39 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_1%VPWR 1 2 9 15 18 19 21 22 23 33 34
r34 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r35 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r37 27 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r38 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r39 23 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 21 30 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.63 $Y=2.72 $X2=1.61
+ $Y2=2.72
r41 21 22 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.63 $Y=2.72
+ $X2=1.772 $Y2=2.72
r42 20 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 20 22 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.772 $Y2=2.72
r44 18 26 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.71 $Y=2.72 $X2=0.69
+ $Y2=2.72
r45 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.71 $Y=2.72
+ $X2=0.835 $Y2=2.72
r46 17 30 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=1.61 $Y2=2.72
r47 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=0.835 $Y2=2.72
r48 13 22 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.772 $Y=2.635
+ $X2=1.772 $Y2=2.72
r49 13 15 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=1.772 $Y=2.635
+ $X2=1.772 $Y2=2
r50 9 12 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.835 $Y=1.66
+ $X2=0.835 $Y2=2
r51 7 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=2.635
+ $X2=0.835 $Y2=2.72
r52 7 12 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.835 $Y=2.635
+ $X2=0.835 $Y2=2
r53 2 15 300 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=1.485 $X2=1.775 $Y2=2
r54 1 12 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=0.675
+ $Y=1.485 $X2=0.875 $Y2=2
r55 1 9 600 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.485 $X2=0.875 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_1%Y 1 2 3 10 12 14 16 22 23 24 25 26 27 36 39
r48 36 39 0.993485 $w=2.88e-07 $l=2.5e-08 $layer=LI1_cond $X=2.53 $Y=0.485
+ $X2=2.53 $Y2=0.51
r49 27 52 2.53406 $w=5.88e-07 $l=1.25e-07 $layer=LI1_cond $X=2.38 $Y=2.21
+ $X2=2.38 $Y2=2.335
r50 26 27 6.89266 $w=5.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.38 $Y=1.87
+ $X2=2.38 $Y2=2.21
r51 26 46 4.15587 $w=5.88e-07 $l=2.05e-07 $layer=LI1_cond $X=2.38 $Y=1.87
+ $X2=2.38 $Y2=1.665
r52 25 37 2.21278 $w=4.4e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.38 $Y=1.58
+ $X2=2.53 $Y2=1.495
r53 25 46 2.21278 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=1.58 $X2=2.38
+ $Y2=1.665
r54 25 37 0.993485 $w=2.88e-07 $l=2.5e-08 $layer=LI1_cond $X=2.53 $Y=1.47
+ $X2=2.53 $Y2=1.495
r55 24 25 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=2.53 $Y=1.19 $X2=2.53
+ $Y2=1.47
r56 23 24 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.53 $Y=0.85
+ $X2=2.53 $Y2=1.19
r57 22 36 3.06749 $w=2.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.53 $Y=0.37
+ $X2=2.53 $Y2=0.485
r58 22 23 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.53 $Y=0.54
+ $X2=2.53 $Y2=0.85
r59 22 39 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=2.53 $Y=0.54 $X2=2.53
+ $Y2=0.51
r60 16 22 3.86771 $w=2.3e-07 $l=1.45e-07 $layer=LI1_cond $X=2.385 $Y=0.37
+ $X2=2.53 $Y2=0.37
r61 16 18 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.385 $Y=0.37
+ $X2=2.25 $Y2=0.37
r62 15 21 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=1.58
+ $X2=1.295 $Y2=1.58
r63 14 25 4.90852 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.085 $Y=1.58
+ $X2=2.38 $Y2=1.58
r64 14 15 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.085 $Y=1.58
+ $X2=1.46 $Y2=1.58
r65 10 21 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=1.665
+ $X2=1.295 $Y2=1.58
r66 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.295 $Y=1.665
+ $X2=1.295 $Y2=2.34
r67 3 25 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.485 $X2=2.25 $Y2=1.655
r68 3 52 400 $w=1.7e-07 $l=9.15014e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.485 $X2=2.25 $Y2=2.335
r69 2 21 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.485 $X2=1.295 $Y2=1.66
r70 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.485 $X2=1.295 $Y2=2.34
r71 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.25 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3B_1%VGND 1 6 9 10 11 21 22
r31 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r32 19 22 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r33 18 21 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r34 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r35 15 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r36 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r37 11 15 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r38 9 14 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.69
+ $Y2=0
r39 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.875
+ $Y2=0
r40 8 18 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=1.15
+ $Y2=0
r41 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.875
+ $Y2=0
r42 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=0.085
+ $X2=0.875 $Y2=0
r43 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.875 $Y=0.085
+ $X2=0.875 $Y2=0.38
r44 1 6 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=0.675
+ $Y=0.465 $X2=0.875 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
M1000 a_212_413# a_27_413# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.218e+11p pd=1.42e+06u as=8.712e+11p ps=7.58e+06u
M1001 VPWR a_212_413# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1002 VGND B a_297_47# VNB nshort w=420000u l=150000u
+  ad=4.8845e+11p pd=5.18e+06u as=1.134e+11p ps=1.38e+06u
M1003 a_297_47# a_27_413# a_212_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1004 X a_212_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A_N a_27_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1006 VPWR B a_212_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_212_413# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1008 a_27_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1009 X a_212_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


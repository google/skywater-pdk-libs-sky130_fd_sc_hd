* File: sky130_fd_sc_hd__o31a_1.spice
* Created: Tue Sep  1 19:25:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o31a_1.pex.spice"
.subckt sky130_fd_sc_hd__o31a_1  VNB VPB A1 A2 A3 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_103_199#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.234 PD=1.04 PS=2.02 NRD=10.152 NRS=13.836 M=1 R=4.33333
+ SA=75000.3 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_253_47#_M1003_d N_A1_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75000.8 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_253_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_253_47#_M1007_d N_A3_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=4.608 NRS=4.608 M=1 R=4.33333
+ SA=75001.7 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_A_103_199#_M1009_d N_B1_M1009_g N_A_253_47#_M1007_d VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.10725 PD=1.92 PS=0.98 NRD=4.608 NRS=4.608 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_103_199#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.36 PD=1.39 PS=2.72 NRD=10.8153 NRS=14.7553 M=1 R=6.66667
+ SA=75000.3 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1005 A_253_297# N_A1_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.195 PD=1.27 PS=1.39 NRD=15.7403 NRS=10.8153 M=1 R=6.66667 SA=75000.8
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1004 A_337_297# N_A2_M1004_g A_253_297# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=15.7403 M=1 R=6.66667 SA=75001.2
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1000 N_A_103_199#_M1000_d N_A3_M1000_g A_337_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.2125 AS=0.165 PD=1.425 PS=1.33 NRD=28.565 NRS=21.6503 M=1 R=6.66667
+ SA=75001.7 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g N_A_103_199#_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.345 AS=0.2125 PD=2.69 PS=1.425 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__o31a_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a211oi_1.pex.spice
* Created: Tue Sep  1 18:51:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A211OI_1%A2 1 3 6 8 9 16
c27 8 0 1.7283e-19 $X=0.23 $Y=0.85
r28 13 16 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.35 $Y=1.16
+ $X2=0.62 $Y2=1.16
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.16 $X2=0.35 $Y2=1.16
r30 9 14 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=0.265 $Y=1.19 $X2=0.265
+ $Y2=1.16
r31 8 14 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.265 $Y=0.85
+ $X2=0.265 $Y2=1.16
r32 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.62 $Y=1.325
+ $X2=0.62 $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.62 $Y=1.325 $X2=0.62
+ $Y2=1.985
r34 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.62 $Y=0.995
+ $X2=0.62 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.62 $Y=0.995 $X2=0.62
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_1%A1 3 6 8 9 10 11 17 19
c36 17 0 1.7283e-19 $X=1.04 $Y=1.16
r37 21 30 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0.995
+ $X2=0.73 $Y2=1.16
r38 18 30 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.04 $Y=1.16 $X2=0.73
+ $Y2=1.16
r39 17 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.16
+ $X2=1.04 $Y2=1.325
r40 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.16
+ $X2=1.04 $Y2=0.995
r41 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.16 $X2=1.04 $Y2=1.16
r42 11 18 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.04 $Y2=1.16
r43 10 30 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.73
+ $Y2=1.16
r44 9 21 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=0.73 $Y=0.85
+ $X2=0.73 $Y2=0.995
r45 8 9 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.73 $Y=0.51 $X2=0.73
+ $Y2=0.85
r46 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.05 $Y=1.985
+ $X2=1.05 $Y2=1.325
r47 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.05 $Y=0.56 $X2=1.05
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_1%B1 3 6 8 9 10 11 17 18 19
c35 18 0 1.20783e-19 $X=1.52 $Y=1.16
r36 17 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.52 $Y2=1.325
r37 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.16
+ $X2=1.52 $Y2=0.995
r38 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r39 10 11 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.64 $Y=1.87
+ $X2=1.64 $Y2=2.21
r40 9 10 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.64 $Y=1.53 $X2=1.64
+ $Y2=1.87
r41 9 33 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.64 $Y=1.53
+ $X2=1.64 $Y2=1.325
r42 8 33 5.78494 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.59 $Y=1.19
+ $X2=1.59 $Y2=1.325
r43 8 18 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.59 $Y=1.19 $X2=1.59
+ $Y2=1.16
r44 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.48 $Y=1.985
+ $X2=1.48 $Y2=1.325
r45 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.56 $X2=1.48
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_1%C1 1 3 6 8 9 15
r30 12 15 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.94 $Y=1.16
+ $X2=2.15 $Y2=1.16
r31 8 9 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.085 $Y=1.16
+ $X2=2.085 $Y2=1.53
r32 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.16 $X2=2.15 $Y2=1.16
r33 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.94 $Y=1.325
+ $X2=1.94 $Y2=1.16
r34 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.94 $Y=1.325 $X2=1.94
+ $Y2=1.985
r35 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.94 $Y=0.995
+ $X2=1.94 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.94 $Y=0.995 $X2=1.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_1%A_56_297# 1 2 9 11 12 15
r16 13 15 7.49386 $w=1.83e-07 $l=1.25e-07 $layer=LI1_cond $X=1.262 $Y=1.725
+ $X2=1.262 $Y2=1.85
r17 11 13 6.82996 $w=2e-07 $l=1.38564e-07 $layer=LI1_cond $X=1.17 $Y=1.625
+ $X2=1.262 $Y2=1.725
r18 11 12 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=1.17 $Y=1.625
+ $X2=0.5 $Y2=1.625
r19 7 12 6.92652 $w=2e-07 $l=1.67705e-07 $layer=LI1_cond $X=0.375 $Y=1.725
+ $X2=0.5 $Y2=1.625
r20 7 9 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.375 $Y=1.725
+ $X2=0.375 $Y2=1.85
r21 2 15 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=1.125
+ $Y=1.485 $X2=1.265 $Y2=1.85
r22 1 9 300 $w=1.7e-07 $l=4.22907e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=1.485 $X2=0.405 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_1%VPWR 1 8 10 17 18 21
r30 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r32 15 18 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r33 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r34 14 17 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r35 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r36 12 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=0.835
+ $Y2=2.72
r37 12 14 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1 $Y=2.72 $X2=1.15
+ $Y2=2.72
r38 10 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r39 6 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=2.635
+ $X2=0.835 $Y2=2.72
r40 6 8 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.835 $Y=2.635
+ $X2=0.835 $Y2=2.02
r41 1 8 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=0.695
+ $Y=1.485 $X2=0.835 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_1%Y 1 2 3 12 14 15 18 20 22 23 24 25 36 39 55
r35 36 39 1.87607 $w=2.13e-07 $l=3.5e-08 $layer=LI1_cond $X=2.552 $Y=0.815
+ $X2=2.552 $Y2=0.85
r36 25 55 0.392742 $w=6.68e-07 $l=2.2e-08 $layer=LI1_cond $X=2.53 $Y=2.12
+ $X2=2.552 $Y2=2.12
r37 25 55 7.5304 $w=2.15e-07 $l=3.35e-07 $layer=LI1_cond $X=2.552 $Y=1.785
+ $X2=2.552 $Y2=2.12
r38 25 51 6.69447 $w=6.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.53 $Y=2.12
+ $X2=2.155 $Y2=2.12
r39 24 25 9.86223 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=2.552 $Y=1.53
+ $X2=2.552 $Y2=1.785
r40 23 24 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.552 $Y=1.19
+ $X2=2.552 $Y2=1.53
r41 22 36 1.28421 $w=1.88e-07 $l=2.2e-08 $layer=LI1_cond $X=2.53 $Y=0.72
+ $X2=2.552 $Y2=0.72
r42 22 23 16.8846 $w=2.13e-07 $l=3.15e-07 $layer=LI1_cond $X=2.552 $Y=0.875
+ $X2=2.552 $Y2=1.19
r43 22 39 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=2.552 $Y=0.875
+ $X2=2.552 $Y2=0.85
r44 20 51 1.51741 $w=6.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.12
+ $X2=2.155 $Y2=2.12
r45 16 22 21.1895 $w=1.88e-07 $l=3.63e-07 $layer=LI1_cond $X=2.167 $Y=0.72
+ $X2=2.53 $Y2=0.72
r46 16 18 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=2.167 $Y=0.625
+ $X2=2.167 $Y2=0.53
r47 14 16 6.5378 $w=1.88e-07 $l=1.12e-07 $layer=LI1_cond $X=2.055 $Y=0.72
+ $X2=2.167 $Y2=0.72
r48 14 15 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=2.055 $Y=0.72
+ $X2=1.365 $Y2=0.72
r49 10 15 6.81807 $w=1.9e-07 $l=1.33641e-07 $layer=LI1_cond $X=1.272 $Y=0.625
+ $X2=1.365 $Y2=0.72
r50 10 12 5.69533 $w=1.83e-07 $l=9.5e-08 $layer=LI1_cond $X=1.272 $Y=0.625
+ $X2=1.272 $Y2=0.53
r51 3 51 300 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.155 $Y2=1.87
r52 2 18 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.235 $X2=2.155 $Y2=0.53
r53 1 12 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.265 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_1%VGND 1 2 7 9 13 15 17 24 25 31
r38 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r39 25 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r40 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r41 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r42 22 24 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.53
+ $Y2=0
r43 21 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r44 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 18 28 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r46 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r47 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r48 17 20 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=0.69
+ $Y2=0
r49 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r50 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r52 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.36
r53 7 28 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.212 $Y2=0
r54 7 9 14.4055 $w=3.38e-07 $l=4.25e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.51
r55 2 13 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.71 $Y2=0.36
r56 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends


* File: sky130_fd_sc_hd__and3_4.pxi.spice
* Created: Tue Sep  1 18:57:38 2020
* 
x_PM_SKY130_FD_SC_HD__AND3_4%A N_A_M1006_g N_A_M1004_g A A A A A N_A_c_66_n
+ N_A_c_67_n N_A_c_68_n N_A_c_69_n PM_SKY130_FD_SC_HD__AND3_4%A
x_PM_SKY130_FD_SC_HD__AND3_4%B N_B_M1005_g N_B_M1009_g B B N_B_c_100_n
+ N_B_c_101_n PM_SKY130_FD_SC_HD__AND3_4%B
x_PM_SKY130_FD_SC_HD__AND3_4%C N_C_M1007_g N_C_M1013_g C N_C_c_134_n N_C_c_135_n
+ N_C_c_136_n PM_SKY130_FD_SC_HD__AND3_4%C
x_PM_SKY130_FD_SC_HD__AND3_4%A_94_47# N_A_94_47#_M1006_s N_A_94_47#_M1004_s
+ N_A_94_47#_M1009_d N_A_94_47#_c_174_n N_A_94_47#_M1000_g N_A_94_47#_M1001_g
+ N_A_94_47#_c_175_n N_A_94_47#_M1003_g N_A_94_47#_M1002_g N_A_94_47#_c_176_n
+ N_A_94_47#_M1010_g N_A_94_47#_M1008_g N_A_94_47#_c_177_n N_A_94_47#_M1011_g
+ N_A_94_47#_M1012_g N_A_94_47#_c_190_n N_A_94_47#_c_191_n N_A_94_47#_c_193_n
+ N_A_94_47#_c_196_n N_A_94_47#_c_244_p N_A_94_47#_c_214_n N_A_94_47#_c_216_n
+ N_A_94_47#_c_178_n N_A_94_47#_c_186_n N_A_94_47#_c_187_n N_A_94_47#_c_179_n
+ N_A_94_47#_c_222_n N_A_94_47#_c_209_n N_A_94_47#_c_180_n N_A_94_47#_c_181_n
+ PM_SKY130_FD_SC_HD__AND3_4%A_94_47#
x_PM_SKY130_FD_SC_HD__AND3_4%VPWR N_VPWR_M1004_d N_VPWR_M1013_d N_VPWR_M1002_s
+ N_VPWR_M1012_s N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n
+ N_VPWR_c_315_n VPWR N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n
+ N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_310_n
+ PM_SKY130_FD_SC_HD__AND3_4%VPWR
x_PM_SKY130_FD_SC_HD__AND3_4%X N_X_M1000_d N_X_M1010_d N_X_M1001_d N_X_M1008_d
+ N_X_c_400_n N_X_c_377_n N_X_c_380_n N_X_c_384_n N_X_c_420_p N_X_c_404_n
+ N_X_c_386_n N_X_c_375_n N_X_c_390_n N_X_c_392_n N_X_c_394_n X N_X_c_373_n X
+ PM_SKY130_FD_SC_HD__AND3_4%X
x_PM_SKY130_FD_SC_HD__AND3_4%VGND N_VGND_M1007_d N_VGND_M1003_s N_VGND_M1011_s
+ N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n VGND
+ N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n
+ N_VGND_c_444_n PM_SKY130_FD_SC_HD__AND3_4%VGND
cc_1 VNB N_A_c_66_n 0.0257419f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.16
cc_2 VNB N_A_c_67_n 0.00681569f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.16
cc_3 VNB N_A_c_68_n 0.0232356f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.995
cc_4 VNB N_A_c_69_n 0.0256738f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.34
cc_5 VNB B 0.00302691f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_B_c_100_n 0.0245622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_101_n 0.0163111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_C_c_134_n 0.0213314f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=2.125
cc_9 VNB N_C_c_135_n 0.00333403f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_10 VNB N_C_c_136_n 0.0171317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_94_47#_c_174_n 0.0169849f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.785
cc_12 VNB N_A_94_47#_c_175_n 0.0159983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_94_47#_c_176_n 0.0160024f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.53
cc_14 VNB N_A_94_47#_c_177_n 0.0184169f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.167
cc_15 VNB N_A_94_47#_c_178_n 0.00127837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_94_47#_c_179_n 0.0206169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_94_47#_c_180_n 0.00171227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_94_47#_c_181_n 0.0667411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_310_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_373_n 0.0108749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB X 0.0235754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_435_n 0.00498867f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_23 VNB N_VGND_c_436_n 3.16879e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_437_n 0.0115115f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.16
cc_25 VNB N_VGND_c_438_n 0.0107852f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.16
cc_26 VNB N_VGND_c_439_n 0.0517833f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.53
cc_27 VNB N_VGND_c_440_n 0.0151313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_441_n 0.0113516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_442_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_443_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_444_n 0.233861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_M1004_g 0.0240456f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=1.985
cc_33 VPB A 0.0554181f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_34 VPB N_A_c_66_n 0.00488865f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.16
cc_35 VPB N_A_c_67_n 0.00926757f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.16
cc_36 VPB N_A_c_69_n 0.00174909f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.34
cc_37 VPB N_B_M1009_g 0.020226f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=1.985
cc_38 VPB B 0.00291181f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_39 VPB N_B_c_100_n 0.00651756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_C_M1013_g 0.0201219f $X=-0.19 $Y=1.305 $X2=0.85 $Y2=1.985
cc_41 VPB N_C_c_134_n 0.00438033f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=2.125
cc_42 VPB N_C_c_135_n 0.0017826f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_43 VPB N_A_94_47#_M1001_g 0.0188029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_94_47#_M1002_g 0.018288f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.325
cc_45 VPB N_A_94_47#_M1008_g 0.0183103f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.167
cc_46 VPB N_A_94_47#_M1012_g 0.0210399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_94_47#_c_186_n 0.00127073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_94_47#_c_187_n 0.00920717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_94_47#_c_180_n 4.55278e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_94_47#_c_181_n 0.0124075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_311_n 5.98722e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_312_n 0.00431378f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.16
cc_53 VPB N_VPWR_c_313_n 3.16049e-19 $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.34
cc_54 VPB N_VPWR_c_314_n 0.0117752f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.87
cc_55 VPB N_VPWR_c_315_n 0.0236962f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_316_n 0.026081f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.167
cc_57 VPB N_VPWR_c_317_n 0.0151808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_318_n 0.0152595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_319_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_320_n 0.00617384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_321_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_322_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_310_n 0.0527447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_375_n 0.0124234f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.167
cc_65 VPB X 0.0114218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_B_M1009_g 0.0291441f $X=0.85 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_c_67_n B 0.0261614f $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_c_68_n B 0.00740956f $X=0.79 $Y=0.995 $X2=0 $Y2=0
cc_69 N_A_c_66_n N_B_c_100_n 0.0202499f $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_c_67_n N_B_c_100_n 3.29962e-19 $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_68_n N_B_c_101_n 0.0255029f $X=0.79 $Y=0.995 $X2=0 $Y2=0
cc_72 A N_A_94_47#_c_190_n 0.0429321f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_A_94_47#_c_191_n 0.017726f $X=0.85 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_c_67_n N_A_94_47#_c_191_n 0.0070886f $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_75 A N_A_94_47#_c_193_n 0.0138544f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_76 N_A_c_66_n N_A_94_47#_c_193_n 4.8941e-19 $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_67_n N_A_94_47#_c_193_n 0.0119615f $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_c_67_n N_A_94_47#_c_196_n 0.00255951f $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_c_68_n N_A_94_47#_c_196_n 0.0113389f $X=0.79 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_c_66_n N_A_94_47#_c_179_n 0.0025703f $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_c_67_n N_A_94_47#_c_179_n 0.0233015f $X=0.79 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_c_68_n N_A_94_47#_c_179_n 0.00832591f $X=0.79 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_M1004_g N_VPWR_c_311_n 0.0208021f $X=0.85 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1004_g N_VPWR_c_316_n 0.0046653f $X=0.85 $Y=1.985 $X2=0 $Y2=0
cc_85 A N_VPWR_c_316_n 0.00971455f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_VPWR_c_310_n 0.00921786f $X=0.85 $Y=1.985 $X2=0 $Y2=0
cc_87 A N_VPWR_c_310_n 0.00888181f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_88 N_A_c_68_n N_VGND_c_439_n 0.00379209f $X=0.79 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_c_68_n N_VGND_c_444_n 0.00693391f $X=0.79 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B_M1009_g N_C_M1013_g 0.0266737f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_91 B N_C_c_134_n 2.57509e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_92 N_B_c_100_n N_C_c_134_n 0.0377243f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_93 B N_C_c_135_n 0.026106f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_94 N_B_c_100_n N_C_c_135_n 0.00237503f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_95 B N_C_c_136_n 0.00102386f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_96 N_B_c_101_n N_C_c_136_n 0.0377243f $X=1.302 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B_M1009_g N_A_94_47#_c_191_n 0.0184853f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_98 B N_A_94_47#_c_191_n 0.0166254f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_99 N_B_c_100_n N_A_94_47#_c_191_n 0.00102608f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_100 B N_A_94_47#_c_196_n 0.0170032f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_101 N_B_c_100_n N_A_94_47#_c_196_n 6.64467e-19 $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B_c_101_n N_A_94_47#_c_196_n 0.0138739f $X=1.302 $Y=0.995 $X2=0 $Y2=0
cc_103 B N_A_94_47#_c_179_n 0.00328445f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_104 N_B_c_101_n N_A_94_47#_c_179_n 0.00153016f $X=1.302 $Y=0.995 $X2=0 $Y2=0
cc_105 B N_A_94_47#_c_209_n 0.00423161f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_106 N_B_c_101_n N_A_94_47#_c_209_n 0.00481831f $X=1.302 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B_M1009_g N_VPWR_c_311_n 0.0102669f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B_M1009_g N_VPWR_c_317_n 0.00486043f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_109 N_B_M1009_g N_VPWR_c_310_n 0.00825064f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_110 B A_185_47# 0.00404137f $X=1.065 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_111 N_B_c_101_n N_VGND_c_439_n 0.00381696f $X=1.302 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B_c_101_n N_VGND_c_444_n 0.00553654f $X=1.302 $Y=0.995 $X2=0 $Y2=0
cc_113 N_C_c_136_n N_A_94_47#_c_174_n 0.0183637f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_114 N_C_M1013_g N_A_94_47#_M1001_g 0.0204163f $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_115 N_C_c_135_n N_A_94_47#_c_196_n 3.68376e-19 $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C_M1013_g N_A_94_47#_c_214_n 0.0158815f $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_117 N_C_c_135_n N_A_94_47#_c_214_n 0.00910494f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C_c_134_n N_A_94_47#_c_216_n 0.00354699f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_119 N_C_c_135_n N_A_94_47#_c_216_n 0.00975994f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C_c_136_n N_A_94_47#_c_216_n 0.00927457f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_121 N_C_c_135_n N_A_94_47#_c_178_n 0.0018209f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_122 N_C_c_136_n N_A_94_47#_c_178_n 0.00398737f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_123 N_C_M1013_g N_A_94_47#_c_186_n 0.00498595f $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_124 N_C_c_134_n N_A_94_47#_c_222_n 4.90425e-19 $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_125 N_C_c_135_n N_A_94_47#_c_222_n 0.0109419f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_126 N_C_c_135_n N_A_94_47#_c_209_n 0.0120193f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_127 N_C_c_136_n N_A_94_47#_c_209_n 0.00938493f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_128 N_C_M1013_g N_A_94_47#_c_180_n 8.45385e-19 $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_129 N_C_c_134_n N_A_94_47#_c_180_n 0.00243438f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_130 N_C_c_135_n N_A_94_47#_c_180_n 0.025987f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_131 N_C_c_134_n N_A_94_47#_c_181_n 0.0124263f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_132 N_C_c_135_n N_A_94_47#_c_181_n 2.86813e-19 $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_133 N_C_M1013_g N_VPWR_c_311_n 6.18944e-19 $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_134 N_C_M1013_g N_VPWR_c_312_n 0.00171766f $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_135 N_C_M1013_g N_VPWR_c_317_n 0.00585385f $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_136 N_C_M1013_g N_VPWR_c_310_n 0.0107105f $X=1.825 $Y=1.985 $X2=0 $Y2=0
cc_137 N_C_c_136_n N_VGND_c_435_n 0.00746301f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_138 N_C_c_136_n N_VGND_c_439_n 0.0041129f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_139 N_C_c_136_n N_VGND_c_444_n 0.00585729f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_94_47#_c_191_n N_VPWR_M1004_d 0.0087476f $X=1.52 $Y=1.665 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_94_47#_c_214_n N_VPWR_M1013_d 0.00696425f $X=2.07 $Y=1.665 $X2=0
+ $Y2=0
cc_142 N_A_94_47#_c_186_n N_VPWR_M1013_d 0.00111849f $X=2.175 $Y=1.58 $X2=0
+ $Y2=0
cc_143 N_A_94_47#_c_191_n N_VPWR_c_311_n 0.0251938f $X=1.52 $Y=1.665 $X2=0 $Y2=0
cc_144 N_A_94_47#_M1001_g N_VPWR_c_312_n 0.00170185f $X=2.33 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_94_47#_c_214_n N_VPWR_c_312_n 0.0193839f $X=2.07 $Y=1.665 $X2=0 $Y2=0
cc_146 N_A_94_47#_M1001_g N_VPWR_c_313_n 6.10667e-19 $X=2.33 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_94_47#_M1002_g N_VPWR_c_313_n 0.00979109f $X=2.76 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_94_47#_M1008_g N_VPWR_c_313_n 0.00969908f $X=3.19 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_94_47#_M1012_g N_VPWR_c_313_n 5.94761e-19 $X=3.62 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_94_47#_M1008_g N_VPWR_c_315_n 5.94761e-19 $X=3.19 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_94_47#_M1012_g N_VPWR_c_315_n 0.0107575f $X=3.62 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_94_47#_c_190_n N_VPWR_c_316_n 0.012308f $X=0.635 $Y=1.96 $X2=0 $Y2=0
cc_153 N_A_94_47#_c_244_p N_VPWR_c_317_n 0.012099f $X=1.61 $Y=1.96 $X2=0 $Y2=0
cc_154 N_A_94_47#_M1001_g N_VPWR_c_318_n 0.00585385f $X=2.33 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_94_47#_M1002_g N_VPWR_c_318_n 0.00486043f $X=2.76 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A_94_47#_M1008_g N_VPWR_c_319_n 0.00486043f $X=3.19 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_94_47#_M1012_g N_VPWR_c_319_n 0.00486043f $X=3.62 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_94_47#_M1004_s N_VPWR_c_310_n 0.00683628f $X=0.47 $Y=1.485 $X2=0
+ $Y2=0
cc_159 N_A_94_47#_M1009_d N_VPWR_c_310_n 0.00570388f $X=1.47 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_94_47#_M1001_g N_VPWR_c_310_n 0.0106977f $X=2.33 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_94_47#_M1002_g N_VPWR_c_310_n 0.00822531f $X=2.76 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_94_47#_M1008_g N_VPWR_c_310_n 0.00822531f $X=3.19 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_94_47#_M1012_g N_VPWR_c_310_n 0.00822531f $X=3.62 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_94_47#_c_190_n N_VPWR_c_310_n 0.00685509f $X=0.635 $Y=1.96 $X2=0
+ $Y2=0
cc_165 N_A_94_47#_c_244_p N_VPWR_c_310_n 0.00685509f $X=1.61 $Y=1.96 $X2=0 $Y2=0
cc_166 N_A_94_47#_c_175_n N_X_c_377_n 0.011111f $X=2.76 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_94_47#_c_176_n N_X_c_377_n 0.0110478f $X=3.19 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_94_47#_c_181_n N_X_c_377_n 0.00231838f $X=3.62 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_94_47#_M1002_g N_X_c_380_n 0.016114f $X=2.76 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_94_47#_M1008_g N_X_c_380_n 0.0139045f $X=3.19 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_94_47#_c_187_n N_X_c_380_n 0.0417385f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_94_47#_c_181_n N_X_c_380_n 6.56764e-19 $X=3.62 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_94_47#_c_187_n N_X_c_384_n 0.0147839f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_94_47#_c_181_n N_X_c_384_n 7.2697e-19 $X=3.62 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_94_47#_c_177_n N_X_c_386_n 0.0160286f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_94_47#_c_187_n N_X_c_386_n 0.00590462f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_94_47#_M1012_g N_X_c_375_n 0.019007f $X=3.62 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_94_47#_c_187_n N_X_c_375_n 0.00595992f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_94_47#_c_187_n N_X_c_390_n 0.0546247f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_94_47#_c_181_n N_X_c_390_n 0.00234013f $X=3.62 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_94_47#_c_187_n N_X_c_392_n 0.0141519f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_94_47#_c_181_n N_X_c_392_n 0.00238051f $X=3.62 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_94_47#_c_187_n N_X_c_394_n 0.0147839f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_94_47#_c_181_n N_X_c_394_n 7.2697e-19 $X=3.62 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_94_47#_c_177_n X 0.0240627f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_94_47#_c_187_n X 0.0275568f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_94_47#_c_196_n A_185_47# 0.0089404f $X=1.535 $Y=0.47 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_94_47#_c_196_n A_294_47# 6.80594e-19 $X=1.535 $Y=0.47 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_94_47#_c_209_n A_294_47# 0.00503015f $X=1.63 $Y=0.47 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_94_47#_c_216_n N_VGND_M1007_d 0.00931057f $X=2.07 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_191 N_A_94_47#_c_178_n N_VGND_M1007_d 9.90294e-19 $X=2.175 $Y=1.02 $X2=-0.19
+ $Y2=-0.24
cc_192 N_A_94_47#_c_174_n N_VGND_c_435_n 0.00178881f $X=2.33 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_94_47#_c_216_n N_VGND_c_435_n 0.0232062f $X=2.07 $Y=0.71 $X2=0 $Y2=0
cc_194 N_A_94_47#_c_209_n N_VGND_c_435_n 0.00499547f $X=1.63 $Y=0.47 $X2=0 $Y2=0
cc_195 N_A_94_47#_c_174_n N_VGND_c_436_n 0.00107213f $X=2.33 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_94_47#_c_175_n N_VGND_c_436_n 0.00789008f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_94_47#_c_176_n N_VGND_c_436_n 0.00625485f $X=3.19 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_94_47#_c_177_n N_VGND_c_436_n 4.98572e-19 $X=3.62 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_94_47#_c_176_n N_VGND_c_438_n 4.98572e-19 $X=3.19 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_94_47#_c_177_n N_VGND_c_438_n 0.00731833f $X=3.62 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_94_47#_c_196_n N_VGND_c_439_n 0.0235175f $X=1.535 $Y=0.47 $X2=0 $Y2=0
cc_202 N_A_94_47#_c_216_n N_VGND_c_439_n 0.00272277f $X=2.07 $Y=0.71 $X2=0 $Y2=0
cc_203 N_A_94_47#_c_179_n N_VGND_c_439_n 0.0210562f $X=0.635 $Y=0.38 $X2=0 $Y2=0
cc_204 N_A_94_47#_c_209_n N_VGND_c_439_n 0.00612925f $X=1.63 $Y=0.47 $X2=0 $Y2=0
cc_205 N_A_94_47#_c_174_n N_VGND_c_440_n 0.00558147f $X=2.33 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_94_47#_c_175_n N_VGND_c_440_n 0.00351072f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_94_47#_c_216_n N_VGND_c_440_n 6.66898e-19 $X=2.07 $Y=0.71 $X2=0 $Y2=0
cc_208 N_A_94_47#_c_176_n N_VGND_c_441_n 0.00351072f $X=3.19 $Y=0.995 $X2=0
+ $Y2=0
cc_209 N_A_94_47#_c_177_n N_VGND_c_441_n 0.00351072f $X=3.62 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_94_47#_M1006_s N_VGND_c_444_n 0.0024621f $X=0.47 $Y=0.235 $X2=0 $Y2=0
cc_211 N_A_94_47#_c_174_n N_VGND_c_444_n 0.0101288f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_94_47#_c_175_n N_VGND_c_444_n 0.00411677f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_94_47#_c_176_n N_VGND_c_444_n 0.0040731f $X=3.19 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_94_47#_c_177_n N_VGND_c_444_n 0.0040731f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_94_47#_c_196_n N_VGND_c_444_n 0.0240682f $X=1.535 $Y=0.47 $X2=0 $Y2=0
cc_216 N_A_94_47#_c_216_n N_VGND_c_444_n 0.00754187f $X=2.07 $Y=0.71 $X2=0 $Y2=0
cc_217 N_A_94_47#_c_179_n N_VGND_c_444_n 0.0125723f $X=0.635 $Y=0.38 $X2=0 $Y2=0
cc_218 N_A_94_47#_c_209_n N_VGND_c_444_n 0.00645546f $X=1.63 $Y=0.47 $X2=0 $Y2=0
cc_219 N_VPWR_c_310_n N_X_M1001_d 0.00535672f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_c_310_n N_X_M1008_d 0.00535672f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_c_318_n N_X_c_400_n 0.0124538f $X=2.81 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_310_n N_X_c_400_n 0.00724021f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_M1002_s N_X_c_380_n 0.00340327f $X=2.835 $Y=1.485 $X2=0 $Y2=0
cc_224 N_VPWR_c_313_n N_X_c_380_n 0.0170296f $X=2.975 $Y=2.02 $X2=0 $Y2=0
cc_225 N_VPWR_c_319_n N_X_c_404_n 0.0124538f $X=3.67 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_c_310_n N_X_c_404_n 0.00724021f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_M1012_s N_X_c_375_n 0.00470097f $X=3.695 $Y=1.485 $X2=0 $Y2=0
cc_228 N_VPWR_c_315_n N_X_c_375_n 0.0239152f $X=3.835 $Y=2.02 $X2=0 $Y2=0
cc_229 N_VPWR_M1012_s X 8.60883e-19 $X=3.695 $Y=1.485 $X2=0 $Y2=0
cc_230 N_X_c_377_n N_VGND_M1003_s 0.00327388f $X=3.31 $Y=0.73 $X2=0 $Y2=0
cc_231 N_X_c_386_n N_VGND_M1011_s 0.0010969f $X=3.775 $Y=0.73 $X2=0 $Y2=0
cc_232 N_X_c_373_n N_VGND_M1011_s 0.00351052f $X=3.915 $Y=0.845 $X2=0 $Y2=0
cc_233 X N_VGND_M1011_s 6.85193e-19 $X=3.91 $Y=0.85 $X2=0 $Y2=0
cc_234 N_X_c_377_n N_VGND_c_436_n 0.0162283f $X=3.31 $Y=0.73 $X2=0 $Y2=0
cc_235 N_X_c_373_n N_VGND_c_437_n 0.00116793f $X=3.915 $Y=0.845 $X2=0 $Y2=0
cc_236 N_X_c_386_n N_VGND_c_438_n 0.00344107f $X=3.775 $Y=0.73 $X2=0 $Y2=0
cc_237 N_X_c_373_n N_VGND_c_438_n 0.0188167f $X=3.915 $Y=0.845 $X2=0 $Y2=0
cc_238 N_X_c_377_n N_VGND_c_440_n 0.00263122f $X=3.31 $Y=0.73 $X2=0 $Y2=0
cc_239 N_X_c_390_n N_VGND_c_440_n 0.00436709f $X=2.64 $Y=0.68 $X2=0 $Y2=0
cc_240 N_X_c_377_n N_VGND_c_441_n 0.00263122f $X=3.31 $Y=0.73 $X2=0 $Y2=0
cc_241 N_X_c_420_p N_VGND_c_441_n 0.0123333f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_242 N_X_c_386_n N_VGND_c_441_n 0.00263122f $X=3.775 $Y=0.73 $X2=0 $Y2=0
cc_243 N_X_M1000_d N_VGND_c_444_n 0.00434391f $X=2.405 $Y=0.235 $X2=0 $Y2=0
cc_244 N_X_M1010_d N_VGND_c_444_n 0.00251209f $X=3.265 $Y=0.235 $X2=0 $Y2=0
cc_245 N_X_c_377_n N_VGND_c_444_n 0.0101713f $X=3.31 $Y=0.73 $X2=0 $Y2=0
cc_246 N_X_c_420_p N_VGND_c_444_n 0.00721345f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_247 N_X_c_386_n N_VGND_c_444_n 0.00477848f $X=3.775 $Y=0.73 $X2=0 $Y2=0
cc_248 N_X_c_390_n N_VGND_c_444_n 0.00604783f $X=2.64 $Y=0.68 $X2=0 $Y2=0
cc_249 N_X_c_373_n N_VGND_c_444_n 0.00289812f $X=3.915 $Y=0.845 $X2=0 $Y2=0
cc_250 A_185_47# N_VGND_c_444_n 0.00338691f $X=0.925 $Y=0.235 $X2=0 $Y2=0
cc_251 A_294_47# N_VGND_c_444_n 0.00179095f $X=1.47 $Y=0.235 $X2=2.07 $Y2=1.665

* File: sky130_fd_sc_hd__fa_4.pex.spice
* Created: Thu Aug 27 14:21:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__FA_4%A_79_21# 1 2 7 9 12 14 16 19 21 23 26 28 30 33
+ 37 41 43 52 54 55 56 57 60 61 62 63 69 70 73 76 85 88 89
c256 88 0 5.62553e-20 $X=6.34 $Y=1.04
c257 76 0 1.85285e-19 $X=6.695 $Y=0.85
c258 70 0 1.9888e-19 $X=3.14 $Y=0.85
c259 60 0 1.83284e-19 $X=2.225 $Y=1.91
c260 54 0 1.81094e-19 $X=1.825 $Y=1.43
r261 88 91 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.34 $Y=1.04
+ $X2=6.34 $Y2=1.205
r262 88 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.34 $Y=1.04
+ $X2=6.34 $Y2=0.875
r263 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.34
+ $Y=1.04 $X2=6.34 $Y2=1.04
r264 82 83 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r265 77 89 13.8814 $w=3.12e-07 $l=3.99687e-07 $layer=LI1_cond $X=6.695 $Y=0.945
+ $X2=6.34 $Y2=1.04
r266 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.695 $Y=0.85
+ $X2=6.695 $Y2=0.85
r267 73 94 0.20132 $w=6.06e-07 $l=1e-08 $layer=LI1_cond $X=2.995 $Y=0.595
+ $X2=3.005 $Y2=0.595
r268 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.995 $Y=0.85
+ $X2=2.995 $Y2=0.85
r269 70 72 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.14 $Y=0.85
+ $X2=2.995 $Y2=0.85
r270 69 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.55 $Y=0.85
+ $X2=6.695 $Y2=0.85
r271 69 70 4.22029 $w=1.4e-07 $l=3.41e-06 $layer=MET1_cond $X=6.55 $Y=0.85
+ $X2=3.14 $Y2=0.85
r272 61 62 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.735 $Y=1.995
+ $X2=2.31 $Y2=1.995
r273 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.225 $Y=1.91
+ $X2=2.31 $Y2=1.995
r274 59 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.225 $Y=1.665
+ $X2=2.225 $Y2=1.91
r275 58 64 1.54022 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.945 $Y=1.58
+ $X2=1.842 $Y2=1.58
r276 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=1.58
+ $X2=2.225 $Y2=1.665
r277 57 58 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.14 $Y=1.58
+ $X2=1.945 $Y2=1.58
r278 55 73 19.6598 $w=6.06e-07 $l=6.93722e-07 $layer=LI1_cond $X=2.37 $Y=0.74
+ $X2=2.995 $Y2=0.595
r279 55 56 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.37 $Y=0.74
+ $X2=1.91 $Y2=0.74
r280 54 64 9.61743 $w=1.95e-07 $l=1.58272e-07 $layer=LI1_cond $X=1.825 $Y=1.43
+ $X2=1.842 $Y2=1.58
r281 53 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=1.245
+ $X2=1.825 $Y2=1.16
r282 53 54 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.825 $Y=1.245
+ $X2=1.825 $Y2=1.43
r283 52 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=1.075
+ $X2=1.825 $Y2=1.16
r284 51 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.825 $Y=0.825
+ $X2=1.91 $Y2=0.74
r285 51 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.825 $Y=0.825
+ $X2=1.825 $Y2=1.075
r286 50 85 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=1.45 $Y=1.16
+ $X2=1.73 $Y2=1.16
r287 50 83 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.45 $Y=1.16
+ $X2=1.31 $Y2=1.16
r288 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.16 $X2=1.45 $Y2=1.16
r289 46 82 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=0.77 $Y=1.16
+ $X2=0.89 $Y2=1.16
r290 46 79 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=0.77 $Y=1.16 $X2=0.47
+ $Y2=1.16
r291 45 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.77 $Y=1.16
+ $X2=1.45 $Y2=1.16
r292 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.16 $X2=0.77 $Y2=1.16
r293 43 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=1.16
+ $X2=1.825 $Y2=1.16
r294 43 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.74 $Y=1.16
+ $X2=1.45 $Y2=1.16
r295 41 91 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.28 $Y=2.165
+ $X2=6.28 $Y2=1.205
r296 37 90 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.28 $Y=0.445
+ $X2=6.28 $Y2=0.875
r297 31 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r298 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r299 28 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r300 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r301 24 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r302 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r303 21 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r304 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r305 17 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r306 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r307 14 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r308 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r309 10 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r310 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r311 7 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r312 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r313 2 61 300 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.855 $X2=2.94 $Y2=1.995
r314 1 94 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.235 $X2=3.005 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%A 1 3 7 11 15 19 23 27 31 38 39 41 42 43 44 45
+ 46 53 58 63 68 69 73 74
c268 69 0 3.76974e-20 $X=5.84 $Y=1.04
c269 53 0 1.2547e-19 $X=3.915 $Y=1.19
c270 44 0 3.10095e-19 $X=4.06 $Y=1.19
c271 43 0 1.21386e-19 $X=5.63 $Y=1.19
c272 42 0 3.35945e-19 $X=2.68 $Y=1.19
c273 39 0 1.39197e-19 $X=2.535 $Y=1.19
c274 23 0 7.10647e-20 $X=5.835 $Y=2.165
c275 11 0 1.9888e-19 $X=3.635 $Y=0.445
r276 73 75 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.72 $Y=1.16
+ $X2=7.72 $Y2=0.995
r277 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.72
+ $Y=1.16 $X2=7.72 $Y2=1.16
r278 68 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=1.04
+ $X2=5.84 $Y2=1.205
r279 68 70 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=1.04
+ $X2=5.84 $Y2=0.875
r280 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.04 $X2=5.84 $Y2=1.04
r281 63 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.195
+ $X2=3.695 $Y2=1.36
r282 63 65 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.195
+ $X2=3.695 $Y2=1.03
r283 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.195 $X2=3.695 $Y2=1.195
r284 59 74 23.2547 $w=2.78e-07 $l=5.65e-07 $layer=LI1_cond $X=7.155 $Y=1.135
+ $X2=7.72 $Y2=1.135
r285 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.155 $Y=1.19
+ $X2=7.155 $Y2=1.19
r286 55 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.775 $Y=1.19
+ $X2=5.775 $Y2=1.19
r287 53 64 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.915 $Y=1.195
+ $X2=3.695 $Y2=1.195
r288 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.915 $Y=1.19
+ $X2=3.915 $Y2=1.19
r289 46 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.92 $Y=1.19
+ $X2=5.775 $Y2=1.19
r290 45 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.01 $Y=1.19
+ $X2=7.155 $Y2=1.19
r291 45 46 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=7.01 $Y=1.19
+ $X2=5.92 $Y2=1.19
r292 44 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.06 $Y=1.19
+ $X2=3.915 $Y2=1.19
r293 43 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.63 $Y=1.19
+ $X2=5.775 $Y2=1.19
r294 43 44 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=5.63 $Y=1.19
+ $X2=4.06 $Y2=1.19
r295 42 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.68 $Y=1.19
+ $X2=2.535 $Y2=1.19
r296 41 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.77 $Y=1.19
+ $X2=3.915 $Y2=1.19
r297 41 42 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=3.77 $Y=1.19
+ $X2=2.68 $Y2=1.19
r298 39 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.535 $Y=1.19
+ $X2=2.535 $Y2=1.19
r299 38 39 8.02594 $w=2.78e-07 $l=1.95e-07 $layer=LI1_cond $X=2.34 $Y=1.135
+ $X2=2.535 $Y2=1.135
r300 35 38 6.40917 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.165 $Y=1.16
+ $X2=2.34 $Y2=1.16
r301 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.16 $X2=2.165 $Y2=1.16
r302 29 73 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.72 $Y=1.325
+ $X2=7.72 $Y2=1.16
r303 29 31 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=7.72 $Y=1.325
+ $X2=7.72 $Y2=2.17
r304 27 75 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.66 $Y=0.445
+ $X2=7.66 $Y2=0.995
r305 23 71 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=5.835 $Y=2.165
+ $X2=5.835 $Y2=1.205
r306 19 70 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.835 $Y=0.445
+ $X2=5.835 $Y2=0.875
r307 15 66 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.635 $Y=2.165
+ $X2=3.635 $Y2=1.36
r308 11 65 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=3.635 $Y=0.445
+ $X2=3.635 $Y2=1.03
r309 5 36 38.8629 $w=2.72e-07 $l=1.93959e-07 $layer=POLY_cond $X=2.23 $Y=0.995
+ $X2=2.167 $Y2=1.16
r310 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.23 $Y=0.995
+ $X2=2.23 $Y2=0.445
r311 1 36 38.8629 $w=2.72e-07 $l=1.83016e-07 $layer=POLY_cond $X=2.205 $Y=1.325
+ $X2=2.167 $Y2=1.16
r312 1 3 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=2.205 $Y=1.325
+ $X2=2.205 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%B 3 7 9 11 12 14 15 16 17 18 19 21 26 29 33 35
+ 36 38 39 40 41 50 51 54 59 60 61 63 65
c231 54 0 4.27861e-19 $X=2.645 $Y=1.53
c232 51 0 2.28652e-19 $X=7.615 $Y=1.53
c233 50 0 3.77214e-20 $X=7.615 $Y=1.53
c234 41 0 5.10808e-21 $X=5 $Y=1.53
c235 40 0 1.7744e-19 $X=7.47 $Y=1.53
c236 29 0 1.47587e-19 $X=7.18 $Y=0.445
c237 18 0 1.2547e-19 $X=4.13 $Y=1.695
r238 65 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.24 $Y=1.53
+ $X2=7.24 $Y2=1.695
r239 65 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.24 $Y=1.53
+ $X2=7.24 $Y2=1.365
r240 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.24
+ $Y=1.53 $X2=7.24 $Y2=1.53
r241 59 61 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.882 $Y=1.52
+ $X2=4.882 $Y2=1.355
r242 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.83
+ $Y=1.52 $X2=4.83 $Y2=1.52
r243 54 57 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.53
+ $X2=2.645 $Y2=1.695
r244 54 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.53
+ $X2=2.645 $Y2=1.365
r245 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.53 $X2=2.645 $Y2=1.53
r246 51 66 14.9023 $w=2.88e-07 $l=3.75e-07 $layer=LI1_cond $X=7.615 $Y=1.59
+ $X2=7.24 $Y2=1.59
r247 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.615 $Y=1.53
+ $X2=7.615 $Y2=1.53
r248 47 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.855 $Y=1.53
+ $X2=4.855 $Y2=1.53
r249 41 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5 $Y=1.53
+ $X2=4.855 $Y2=1.53
r250 40 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.47 $Y=1.53
+ $X2=7.615 $Y2=1.53
r251 40 41 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=7.47 $Y=1.53 $X2=5
+ $Y2=1.53
r252 39 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.14 $Y=1.53
+ $X2=2.995 $Y2=1.53
r253 38 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.71 $Y=1.53
+ $X2=4.855 $Y2=1.53
r254 38 39 1.94307 $w=1.4e-07 $l=1.57e-06 $layer=MET1_cond $X=4.71 $Y=1.53
+ $X2=3.14 $Y2=1.53
r255 36 55 16.4635 $w=2.43e-07 $l=3.5e-07 $layer=LI1_cond $X=2.995 $Y=1.567
+ $X2=2.645 $Y2=1.567
r256 36 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.995 $Y=1.53
+ $X2=2.995 $Y2=1.53
r257 33 68 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=7.18 $Y=2.17
+ $X2=7.18 $Y2=1.695
r258 29 67 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=7.18 $Y=0.445
+ $X2=7.18 $Y2=1.365
r259 26 63 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.995 $Y=2.165
+ $X2=4.995 $Y2=1.77
r260 22 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.995 $Y=0.88
+ $X2=4.995 $Y2=0.805
r261 22 61 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.995 $Y=0.88
+ $X2=4.995 $Y2=1.355
r262 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.995 $Y=0.73
+ $X2=4.995 $Y2=0.805
r263 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.995 $Y=0.73
+ $X2=4.995 $Y2=0.445
r264 17 63 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=4.882 $Y=1.695
+ $X2=4.882 $Y2=1.77
r265 17 59 25.9538 $w=3.75e-07 $l=1.75e-07 $layer=POLY_cond $X=4.882 $Y=1.695
+ $X2=4.882 $Y2=1.52
r266 17 18 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=4.695 $Y=1.695
+ $X2=4.13 $Y2=1.695
r267 15 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.92 $Y=0.805
+ $X2=4.995 $Y2=0.805
r268 15 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.92 $Y=0.805
+ $X2=4.13 $Y2=0.805
r269 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.055 $Y=1.77
+ $X2=4.13 $Y2=1.695
r270 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.055 $Y=1.77
+ $X2=4.055 $Y2=2.165
r271 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.055 $Y=0.73
+ $X2=4.13 $Y2=0.805
r272 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.055 $Y=0.73
+ $X2=4.055 $Y2=0.445
r273 7 56 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.705 $Y=0.445
+ $X2=2.705 $Y2=1.365
r274 3 57 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=2.65 $Y=2.17
+ $X2=2.65 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%CIN 3 7 11 14 20 24 26 27 29 30 31 33 34 35 37
+ 38 42 44 50 51 52 56 58 59
c228 50 0 2.2917e-19 $X=5.415 $Y=1.52
c229 44 0 1.55247e-19 $X=3.335 $Y=1.19
c230 42 0 1.79381e-19 $X=3.215 $Y=1.19
c231 34 0 7.10647e-20 $X=5.22 $Y=1.107
c232 31 0 1.25839e-19 $X=3.42 $Y=1.655
c233 29 0 2.73586e-19 $X=3.335 $Y=1.57
c234 20 0 1.8774e-19 $X=6.705 $Y=2.165
c235 3 0 1.39197e-19 $X=3.215 $Y=0.445
r236 59 64 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=6.72 $Y=1.52 $X2=6.72
+ $Y2=1.6
r237 58 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.76 $Y=1.52
+ $X2=6.76 $Y2=1.685
r238 58 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.76 $Y=1.52
+ $X2=6.76 $Y2=1.355
r239 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.76
+ $Y=1.52 $X2=6.76 $Y2=1.52
r240 52 64 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=6.72 $Y=1.87
+ $X2=6.72 $Y2=1.6
r241 50 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=1.52
+ $X2=5.415 $Y2=1.355
r242 49 51 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=1.56
+ $X2=5.58 $Y2=1.56
r243 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.415
+ $Y=1.52 $X2=5.415 $Y2=1.52
r244 46 49 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.305 $Y=1.56
+ $X2=5.415 $Y2=1.56
r245 41 44 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.215 $Y=1.19
+ $X2=3.335 $Y2=1.19
r246 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=1.19 $X2=3.215 $Y2=1.19
r247 38 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.595 $Y=1.6
+ $X2=6.72 $Y2=1.6
r248 38 51 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=6.595 $Y=1.6
+ $X2=5.58 $Y2=1.6
r249 37 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.305 $Y=1.435
+ $X2=5.305 $Y2=1.56
r250 36 37 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.305 $Y=1.25
+ $X2=5.305 $Y2=1.435
r251 34 36 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=5.22 $Y=1.107
+ $X2=5.305 $Y2=1.25
r252 34 35 35.5842 $w=2.83e-07 $l=8.8e-07 $layer=LI1_cond $X=5.22 $Y=1.107
+ $X2=4.34 $Y2=1.107
r253 32 35 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=4.255 $Y=1.25
+ $X2=4.34 $Y2=1.107
r254 32 33 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.255 $Y=1.25
+ $X2=4.255 $Y2=1.57
r255 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.17 $Y=1.655
+ $X2=4.255 $Y2=1.57
r256 30 31 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.17 $Y=1.655
+ $X2=3.42 $Y2=1.655
r257 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=1.57
+ $X2=3.42 $Y2=1.655
r258 28 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=1.275
+ $X2=3.335 $Y2=1.19
r259 28 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.335 $Y=1.275
+ $X2=3.335 $Y2=1.57
r260 27 56 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=5.42 $Y=0.88
+ $X2=5.42 $Y2=1.355
r261 26 27 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=5.417 $Y=0.73
+ $X2=5.417 $Y2=0.88
r262 24 60 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=6.82 $Y=0.445
+ $X2=6.82 $Y2=1.355
r263 20 61 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.705 $Y=2.165
+ $X2=6.705 $Y2=1.685
r264 12 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=1.685
+ $X2=5.415 $Y2=1.52
r265 12 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.415 $Y=1.685
+ $X2=5.415 $Y2=2.165
r266 11 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.415 $Y=0.445
+ $X2=5.415 $Y2=0.73
r267 5 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.355
+ $X2=3.215 $Y2=1.19
r268 5 7 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.215 $Y=1.355
+ $X2=3.215 $Y2=2.165
r269 1 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.025
+ $X2=3.215 $Y2=1.19
r270 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.215 $Y=1.025
+ $X2=3.215 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%A_1271_47# 1 2 7 9 12 16 18 20 21 23 26 28 30
+ 33 35 39 42 43 44 45 48 50 52 58 64 65 71 73 81
c178 65 0 1.7744e-19 $X=7.525 $Y=2.02
c179 64 0 5.62553e-20 $X=6.635 $Y=0.425
c180 48 0 3.77214e-20 $X=8.02 $Y=1.935
r181 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.695 $Y=1.16
+ $X2=9.115 $Y2=1.16
r182 77 78 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=8.615 $Y=1.16
+ $X2=8.695 $Y2=1.16
r183 69 71 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.02 $Y=1.555
+ $X2=8.14 $Y2=1.555
r184 62 64 3.71115 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=0.425
+ $X2=6.635 $Y2=0.425
r185 59 81 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=9.28 $Y=1.16
+ $X2=9.535 $Y2=1.16
r186 59 79 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.28 $Y=1.16
+ $X2=9.115 $Y2=1.16
r187 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.28
+ $Y=1.16 $X2=9.28 $Y2=1.16
r188 56 77 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.26 $Y=1.16
+ $X2=8.615 $Y2=1.16
r189 56 74 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=8.26 $Y=1.16
+ $X2=8.195 $Y2=1.16
r190 55 58 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.26 $Y=1.16
+ $X2=9.28 $Y2=1.16
r191 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.26
+ $Y=1.16 $X2=8.26 $Y2=1.16
r192 53 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.225 $Y=1.16
+ $X2=8.14 $Y2=1.16
r193 53 55 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=8.225 $Y=1.16
+ $X2=8.26 $Y2=1.16
r194 52 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.14 $Y=1.47
+ $X2=8.14 $Y2=1.555
r195 51 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.14 $Y=1.245
+ $X2=8.14 $Y2=1.16
r196 51 52 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.14 $Y=1.245
+ $X2=8.14 $Y2=1.47
r197 50 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.14 $Y=1.075
+ $X2=8.14 $Y2=1.16
r198 49 50 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.14 $Y=0.825
+ $X2=8.14 $Y2=1.075
r199 47 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=1.64
+ $X2=8.02 $Y2=1.555
r200 47 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.02 $Y=1.64
+ $X2=8.02 $Y2=1.935
r201 46 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.61 $Y=2.02
+ $X2=7.525 $Y2=2.02
r202 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.935 $Y=2.02
+ $X2=8.02 $Y2=1.935
r203 45 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.935 $Y=2.02
+ $X2=7.61 $Y2=2.02
r204 43 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.055 $Y=0.74
+ $X2=8.14 $Y2=0.825
r205 43 44 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=8.055 $Y=0.74
+ $X2=7.475 $Y2=0.74
r206 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.39 $Y=0.655
+ $X2=7.475 $Y2=0.74
r207 41 42 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.39 $Y=0.505
+ $X2=7.39 $Y2=0.655
r208 39 41 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.305 $Y=0.38
+ $X2=7.39 $Y2=0.505
r209 39 64 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.305 $Y=0.38
+ $X2=6.635 $Y2=0.38
r210 35 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.525 $Y=2.295
+ $X2=7.525 $Y2=2.02
r211 35 37 32.0311 $w=3.38e-07 $l=9.45e-07 $layer=LI1_cond $X=7.44 $Y=2.295
+ $X2=6.495 $Y2=2.295
r212 31 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.535 $Y=1.325
+ $X2=9.535 $Y2=1.16
r213 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.535 $Y=1.325
+ $X2=9.535 $Y2=1.985
r214 28 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.535 $Y=0.995
+ $X2=9.535 $Y2=1.16
r215 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.535 $Y=0.995
+ $X2=9.535 $Y2=0.56
r216 24 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=1.325
+ $X2=9.115 $Y2=1.16
r217 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.115 $Y=1.325
+ $X2=9.115 $Y2=1.985
r218 21 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=0.995
+ $X2=9.115 $Y2=1.16
r219 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.115 $Y=0.995
+ $X2=9.115 $Y2=0.56
r220 18 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.695 $Y=0.995
+ $X2=8.695 $Y2=1.16
r221 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.695 $Y=0.995
+ $X2=8.695 $Y2=0.56
r222 14 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.615 $Y=1.325
+ $X2=8.615 $Y2=1.16
r223 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.615 $Y=1.325
+ $X2=8.615 $Y2=1.985
r224 10 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=1.325
+ $X2=8.195 $Y2=1.16
r225 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.195 $Y=1.325
+ $X2=8.195 $Y2=1.985
r226 7 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=0.995
+ $X2=8.195 $Y2=1.16
r227 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.195 $Y=0.995
+ $X2=8.195 $Y2=0.56
r228 2 37 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=6.355
+ $Y=1.845 $X2=6.495 $Y2=2.3
r229 1 62 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.235 $X2=6.55 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54 58
+ 61 62 64 65 67 68 69 72 78 82 87 92 97 110 111 119 122 125 128 131 134
r165 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r166 128 129 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r167 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r168 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r169 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r170 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r171 108 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r172 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r173 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r174 105 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r175 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r176 102 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.145 $Y=2.72
+ $X2=7.98 $Y2=2.72
r177 102 104 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.145 $Y=2.72
+ $X2=8.51 $Y2=2.72
r178 101 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r179 101 129 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=5.75 $Y2=2.72
r180 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r181 98 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.79 $Y=2.72
+ $X2=5.625 $Y2=2.72
r182 98 100 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=5.79 $Y=2.72
+ $X2=7.59 $Y2=2.72
r183 97 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=2.72
+ $X2=7.98 $Y2=2.72
r184 97 100 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.815 $Y=2.72
+ $X2=7.59 $Y2=2.72
r185 96 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r186 96 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r187 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r188 93 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=4.785 $Y2=2.72
r189 93 95 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=5.29 $Y2=2.72
r190 92 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=2.72
+ $X2=5.625 $Y2=2.72
r191 92 95 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.46 $Y=2.72
+ $X2=5.29 $Y2=2.72
r192 91 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r193 91 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r194 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r195 88 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=2.72
+ $X2=3.845 $Y2=2.72
r196 88 90 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.01 $Y=2.72
+ $X2=4.37 $Y2=2.72
r197 87 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.785 $Y2=2.72
r198 87 90 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.62 $Y=2.72
+ $X2=4.37 $Y2=2.72
r199 86 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r200 86 120 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r201 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r202 83 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=1.98 $Y2=2.72
r203 83 85 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=3.45 $Y2=2.72
r204 82 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.68 $Y=2.72
+ $X2=3.845 $Y2=2.72
r205 82 85 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.68 $Y=2.72
+ $X2=3.45 $Y2=2.72
r206 81 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r207 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r208 78 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.98 $Y2=2.72
r209 78 80 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.61 $Y2=2.72
r210 77 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r211 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r212 74 76 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r213 72 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r214 69 134 27.1212 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=1.96
r215 69 74 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=2.72
+ $X2=0.345 $Y2=2.72
r216 69 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r217 67 107 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.66 $Y=2.72
+ $X2=9.43 $Y2=2.72
r218 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.72
+ $X2=9.745 $Y2=2.72
r219 66 110 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=9.83 $Y=2.72
+ $X2=9.89 $Y2=2.72
r220 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=2.72
+ $X2=9.745 $Y2=2.72
r221 64 104 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.74 $Y=2.72
+ $X2=8.51 $Y2=2.72
r222 64 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.74 $Y=2.72
+ $X2=8.825 $Y2=2.72
r223 63 107 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.91 $Y=2.72
+ $X2=9.43 $Y2=2.72
r224 63 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=2.72
+ $X2=8.825 $Y2=2.72
r225 61 76 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r226 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r227 60 80 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r228 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r229 56 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.745 $Y=2.635
+ $X2=9.745 $Y2=2.72
r230 56 58 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=9.745 $Y=2.635
+ $X2=9.745 $Y2=1.96
r231 52 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.825 $Y=2.635
+ $X2=8.825 $Y2=2.72
r232 52 54 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=8.825 $Y=2.635
+ $X2=8.825 $Y2=1.96
r233 48 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=2.635
+ $X2=7.98 $Y2=2.72
r234 48 50 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.98 $Y=2.635
+ $X2=7.98 $Y2=2.36
r235 44 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=2.635
+ $X2=5.625 $Y2=2.72
r236 44 46 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.625 $Y=2.635
+ $X2=5.625 $Y2=2.36
r237 40 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.635
+ $X2=4.785 $Y2=2.72
r238 40 42 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.785 $Y=2.635
+ $X2=4.785 $Y2=2
r239 36 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.72
r240 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.845 $Y=2.635
+ $X2=3.845 $Y2=2.36
r241 32 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.72
r242 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.36
r243 28 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r244 28 30 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=1.96
r245 9 58 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=9.61
+ $Y=1.485 $X2=9.745 $Y2=1.96
r246 8 54 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.69
+ $Y=1.485 $X2=8.825 $Y2=1.96
r247 7 50 600 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.855 $X2=7.98 $Y2=2.36
r248 6 46 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=5.49
+ $Y=1.845 $X2=5.625 $Y2=2.36
r249 5 42 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=4.66
+ $Y=1.845 $X2=4.785 $Y2=2
r250 4 38 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.845 $X2=3.845 $Y2=2.36
r251 3 34 600 $w=1.7e-07 $l=9.58514e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.98 $Y2=2.36
r252 2 30 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r253 1 134 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%COUT 1 2 3 4 14 17 19 20 21 22 24 29 40 42 43
+ 44 47
r77 44 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=2.3
r78 44 47 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=1.62
r79 42 43 9.41323 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=1.522 $Y=1.78
+ $X2=1.522 $Y2=1.95
r80 37 47 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.68 $Y=1.585
+ $X2=0.68 $Y2=1.62
r81 29 43 0.528139 $w=2.08e-07 $l=1e-08 $layer=LI1_cond $X=1.54 $Y=1.96 $X2=1.54
+ $Y2=1.95
r82 25 42 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.485 $Y=1.585
+ $X2=1.485 $Y2=1.78
r83 23 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=0.485
+ $X2=1.44 $Y2=0.4
r84 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.44 $Y=0.485
+ $X2=1.44 $Y2=0.735
r85 22 37 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.5
+ $X2=0.68 $Y2=1.5
r86 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.4 $Y=1.5
+ $X2=1.485 $Y2=1.585
r87 21 22 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.4 $Y=1.5
+ $X2=0.845 $Y2=1.5
r88 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.355 $Y=0.82
+ $X2=1.44 $Y2=0.735
r89 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=0.82
+ $X2=0.845 $Y2=0.82
r90 15 20 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.82
+ $X2=0.845 $Y2=0.82
r91 15 17 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.735
+ $X2=0.68 $Y2=0.4
r92 14 37 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.26 $Y=1.5 $X2=0.68
+ $Y2=1.5
r93 13 15 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.26 $Y=0.82
+ $X2=0.68 $Y2=0.82
r94 13 14 16.7927 $w=3.48e-07 $l=5.1e-07 $layer=LI1_cond $X=0.26 $Y=0.905
+ $X2=0.26 $Y2=1.415
r95 4 29 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r96 3 51 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.3
r97 3 47 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.62
r98 2 40 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r99 1 17 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%A_658_369# 1 2 7 10 11 12
c23 11 0 2.45299e-20 $X=3.51 $Y=2.02
r24 12 14 4.67234 $w=2.35e-07 $l=9e-08 $layer=LI1_cond $X=4.297 $Y=2.105
+ $X2=4.297 $Y2=2.195
r25 10 12 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=4.18 $Y=2.02
+ $X2=4.297 $Y2=2.105
r26 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.18 $Y=2.02
+ $X2=3.51 $Y2=2.02
r27 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.425 $Y=2.105
+ $X2=3.51 $Y2=2.02
r28 7 9 6.45882 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.425 $Y=2.105 $X2=3.425
+ $Y2=2.195
r29 2 14 600 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=1 $X=4.13
+ $Y=1.845 $X2=4.265 $Y2=2.195
r30 1 9 600 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.845 $X2=3.425 $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%A_1014_369# 1 2 9 11 12 15
c20 12 0 1.96224e-19 $X=5.29 $Y=2.02
r21 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.045 $Y=2.105
+ $X2=6.045 $Y2=2.275
r22 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.96 $Y=2.02
+ $X2=6.045 $Y2=2.105
r23 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.96 $Y=2.02
+ $X2=5.29 $Y2=2.02
r24 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.205 $Y=2.105
+ $X2=5.29 $Y2=2.02
r25 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.205 $Y=2.105
+ $X2=5.205 $Y2=2.275
r26 2 15 600 $w=1.7e-07 $l=4.929e-07 $layer=licon1_PDIFF $count=1 $X=5.91
+ $Y=1.845 $X2=6.045 $Y2=2.275
r27 1 9 600 $w=1.7e-07 $l=4.929e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=1.845 $X2=5.205 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%SUM 1 2 3 4 16 19 20 21 25 29 33 35 38 42 43 47
+ 48 51
c86 43 0 1.80183e-20 $X=8.445 $Y=1.795
c87 20 0 2.28938e-20 $X=8.57 $Y=1.5
r88 50 51 7.74029 $w=3.33e-07 $l=2.25e-07 $layer=LI1_cond $X=9.867 $Y=1.415
+ $X2=9.867 $Y2=1.19
r89 49 51 9.80437 $w=3.33e-07 $l=2.85e-07 $layer=LI1_cond $X=9.867 $Y=0.905
+ $X2=9.867 $Y2=1.19
r90 42 43 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.445 $Y=1.96
+ $X2=8.445 $Y2=1.795
r91 38 40 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.485 $Y=0.4
+ $X2=8.485 $Y2=0.485
r92 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.49 $Y=1.5
+ $X2=9.325 $Y2=1.5
r93 35 50 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=9.7 $Y=1.5
+ $X2=9.867 $Y2=1.415
r94 35 36 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.7 $Y=1.5 $X2=9.49
+ $Y2=1.5
r95 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.49 $Y=0.82
+ $X2=9.325 $Y2=0.82
r96 33 49 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=9.7 $Y=0.82
+ $X2=9.867 $Y2=0.905
r97 33 34 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.7 $Y=0.82 $X2=9.49
+ $Y2=0.82
r98 29 31 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.325 $Y=1.62
+ $X2=9.325 $Y2=2.3
r99 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=1.585
+ $X2=9.325 $Y2=1.5
r100 27 29 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=9.325 $Y=1.585
+ $X2=9.325 $Y2=1.62
r101 23 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=0.735
+ $X2=9.325 $Y2=0.82
r102 23 25 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.325 $Y=0.735
+ $X2=9.325 $Y2=0.4
r103 22 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.65 $Y=0.82
+ $X2=8.525 $Y2=0.82
r104 21 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.16 $Y=0.82
+ $X2=9.325 $Y2=0.82
r105 21 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.16 $Y=0.82
+ $X2=8.65 $Y2=0.82
r106 19 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.16 $Y=1.5
+ $X2=9.325 $Y2=1.5
r107 19 20 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.16 $Y=1.5 $X2=8.57
+ $Y2=1.5
r108 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.485 $Y=1.585
+ $X2=8.57 $Y2=1.5
r109 17 43 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.485 $Y=1.585
+ $X2=8.485 $Y2=1.795
r110 16 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=0.735
+ $X2=8.525 $Y2=0.82
r111 16 40 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=8.525 $Y=0.735
+ $X2=8.525 $Y2=0.485
r112 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.485 $X2=9.325 $Y2=2.3
r113 4 29 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.485 $X2=9.325 $Y2=1.62
r114 3 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.27
+ $Y=1.485 $X2=8.405 $Y2=1.96
r115 2 25 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=9.19
+ $Y=0.235 $X2=9.325 $Y2=0.4
r116 1 46 182 $w=1.7e-07 $l=6.02993e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.235 $X2=8.485 $Y2=0.74
r117 1 38 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.235 $X2=8.485 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54 58
+ 61 62 64 65 67 68 70 71 72 75 81 85 93 98 114 115 123 126 129 132 135
r183 132 133 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r184 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r185 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r186 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r187 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r188 112 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r189 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r190 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r191 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r192 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r193 106 133 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=5.75 $Y2=0
r194 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r195 103 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.79 $Y=0
+ $X2=5.625 $Y2=0
r196 103 105 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=5.79 $Y=0
+ $X2=7.59 $Y2=0
r197 102 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r198 102 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r199 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r200 99 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.95 $Y=0
+ $X2=4.785 $Y2=0
r201 99 101 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.95 $Y=0 $X2=5.29
+ $Y2=0
r202 98 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=0
+ $X2=5.625 $Y2=0
r203 98 101 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.46 $Y=0 $X2=5.29
+ $Y2=0
r204 97 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r205 97 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r206 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r207 94 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=0
+ $X2=3.845 $Y2=0
r208 94 96 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.01 $Y=0 $X2=4.37
+ $Y2=0
r209 93 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=0
+ $X2=4.785 $Y2=0
r210 93 96 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.62 $Y=0 $X2=4.37
+ $Y2=0
r211 92 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r212 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r213 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r214 89 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r215 88 91 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r216 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r217 86 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.02 $Y2=0
r218 86 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.53
+ $Y2=0
r219 85 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.68 $Y=0
+ $X2=3.845 $Y2=0
r220 85 91 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.68 $Y=0 $X2=3.45
+ $Y2=0
r221 84 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r222 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r223 81 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=2.02 $Y2=0
r224 81 83 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r225 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r226 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r227 77 79 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r228 75 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r229 72 135 13.9504 $w=3.13e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r230 72 77 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.172 $Y=0
+ $X2=0.345 $Y2=0
r231 72 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r232 70 111 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.66 $Y=0 $X2=9.43
+ $Y2=0
r233 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=0 $X2=9.745
+ $Y2=0
r234 69 114 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=9.83 $Y=0 $X2=9.89
+ $Y2=0
r235 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=0 $X2=9.745
+ $Y2=0
r236 67 108 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.82 $Y=0 $X2=8.51
+ $Y2=0
r237 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=0 $X2=8.905
+ $Y2=0
r238 66 111 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=8.99 $Y=0 $X2=9.43
+ $Y2=0
r239 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=0 $X2=8.905
+ $Y2=0
r240 64 105 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.705 $Y=0
+ $X2=7.59 $Y2=0
r241 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.705 $Y=0 $X2=7.87
+ $Y2=0
r242 63 108 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=8.035 $Y=0
+ $X2=8.51 $Y2=0
r243 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.035 $Y=0 $X2=7.87
+ $Y2=0
r244 61 79 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r245 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r246 60 83 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r247 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r248 56 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.745 $Y=0.085
+ $X2=9.745 $Y2=0
r249 56 58 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.745 $Y=0.085
+ $X2=9.745 $Y2=0.4
r250 52 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=0.085
+ $X2=8.905 $Y2=0
r251 52 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.905 $Y=0.085
+ $X2=8.905 $Y2=0.4
r252 48 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0
r253 48 50 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0.36
r254 44 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=0.085
+ $X2=5.625 $Y2=0
r255 44 46 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.625 $Y=0.085
+ $X2=5.625 $Y2=0.36
r256 40 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=0.085
+ $X2=4.785 $Y2=0
r257 40 42 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.785 $Y=0.085
+ $X2=4.785 $Y2=0.405
r258 36 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=0.085
+ $X2=3.845 $Y2=0
r259 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.845 $Y=0.085
+ $X2=3.845 $Y2=0.36
r260 32 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r261 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.38
r262 28 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r263 28 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.4
r264 9 58 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=9.61
+ $Y=0.235 $X2=9.745 $Y2=0.4
r265 8 54 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.77
+ $Y=0.235 $X2=8.905 $Y2=0.4
r266 7 50 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.735
+ $Y=0.235 $X2=7.87 $Y2=0.36
r267 6 46 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.49
+ $Y=0.235 $X2=5.625 $Y2=0.36
r268 5 42 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=4.66
+ $Y=0.235 $X2=4.785 $Y2=0.405
r269 4 38 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.235 $X2=3.845 $Y2=0.36
r270 3 34 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=2.02 $Y2=0.38
r271 2 30 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r272 1 135 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%A_658_47# 1 2 9 11 12 15
r35 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.265 $Y=0.615
+ $X2=4.265 $Y2=0.445
r36 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.18 $Y=0.7
+ $X2=4.265 $Y2=0.615
r37 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.18 $Y=0.7 $X2=3.51
+ $Y2=0.7
r38 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.425 $Y=0.615
+ $X2=3.51 $Y2=0.7
r39 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.425 $Y=0.615
+ $X2=3.425 $Y2=0.445
r40 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=4.13
+ $Y=0.235 $X2=4.265 $Y2=0.445
r41 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.235 $X2=3.425 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__FA_4%A_1014_47# 1 2 9 11 12 15
c32 12 0 1.49223e-19 $X=5.29 $Y=0.7
r33 13 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.045 $Y=0.615
+ $X2=6.045 $Y2=0.445
r34 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.96 $Y=0.7
+ $X2=6.045 $Y2=0.615
r35 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.96 $Y=0.7 $X2=5.29
+ $Y2=0.7
r36 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.205 $Y=0.615
+ $X2=5.29 $Y2=0.7
r37 7 9 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.205 $Y=0.615
+ $X2=5.205 $Y2=0.445
r38 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.235 $X2=6.045 $Y2=0.445
r39 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.07
+ $Y=0.235 $X2=5.205 $Y2=0.445
.ends


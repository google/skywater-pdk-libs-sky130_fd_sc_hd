* NGSPICE file created from sky130_fd_sc_hd__dlrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=1.8528e+12p ps=1.785e+07u
M1001 a_561_413# a_27_47# a_465_369# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=1.936e+11p ps=1.94e+06u
M1002 a_711_307# a_561_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1003 Q a_711_307# VGND VNB nshort w=650000u l=150000u
+  ad=1.885e+11p pd=1.88e+06u as=1.076e+12p ps=1.165e+07u
M1004 Q_N a_1316_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1005 VGND D a_299_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1006 a_659_47# a_27_47# a_561_413# VNB nshort w=360000u l=150000u
+  ad=1.32e+11p pd=1.49e+06u as=1.008e+11p ps=1.28e+06u
M1007 a_942_47# a_561_413# a_711_307# VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=1.69e+11p ps=1.82e+06u
M1008 VPWR RESET_B a_711_307# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_1316_47# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_465_47# a_299_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.554e+11p pd=1.62e+06u as=0p ps=0u
M1011 VPWR a_711_307# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 VPWR GATE a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1013 VPWR a_711_307# a_645_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1014 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1015 a_465_369# a_299_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND RESET_B a_942_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_1316_47# Q_N VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1018 a_561_413# a_193_47# a_465_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_711_307# a_659_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR D a_299_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1021 VGND a_711_307# a_1316_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1022 Q_N a_1316_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_711_307# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND GATE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1025 VPWR a_711_307# a_1316_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1026 a_645_413# a_193_47# a_561_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q a_711_307# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


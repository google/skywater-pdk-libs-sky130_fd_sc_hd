# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__einvn_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.765000 1.755000 1.955000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.650000 1.725000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.275600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.160000 0.255000 1.755000 0.595000 ;
        RECT 1.160000 0.595000 1.330000 2.125000 ;
        RECT 1.160000 2.125000 1.755000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.255000 0.360000 0.655000 ;
      RECT 0.085000  0.655000 0.990000 0.825000 ;
      RECT 0.085000  1.895000 0.990000 2.065000 ;
      RECT 0.085000  2.065000 0.400000 2.465000 ;
      RECT 0.530000  0.085000 0.990000 0.485000 ;
      RECT 0.570000  2.235000 0.990000 2.635000 ;
      RECT 0.820000  0.825000 0.990000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_0
END LIBRARY

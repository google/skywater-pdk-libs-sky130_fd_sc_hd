* File: sky130_fd_sc_hd__nor3b_1.pex.spice
* Created: Thu Aug 27 14:32:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR3B_1%A_91_199# 1 2 9 12 14 17 20 21 22 26 28 31
r63 28 29 15.549 $w=2.55e-07 $l=3.25e-07 $layer=LI1_cond $X=2.265 $Y=0.655
+ $X2=2.59 $Y2=0.655
r64 25 29 3.11056 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.59 $Y=0.825
+ $X2=2.59 $Y2=0.655
r65 25 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.59 $Y=0.825
+ $X2=2.59 $Y2=1.785
r66 22 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.885 $Y=1.87
+ $X2=2.265 $Y2=1.87
r67 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=1.87
+ $X2=2.59 $Y2=1.785
r68 21 24 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.505 $Y=1.87
+ $X2=2.265 $Y2=1.87
r69 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.8 $Y=1.785
+ $X2=0.885 $Y2=1.87
r70 19 20 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.8 $Y=1.245 $X2=0.8
+ $Y2=1.785
r71 17 32 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.16
+ $X2=0.63 $Y2=1.325
r72 17 31 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.16
+ $X2=0.63 $Y2=0.995
r73 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r74 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.715 $Y=1.16
+ $X2=0.8 $Y2=1.245
r75 14 16 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.715 $Y=1.16
+ $X2=0.59 $Y2=1.16
r76 12 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=1.325
r77 9 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.73 $Y=0.56 $X2=0.73
+ $Y2=0.995
r78 2 24 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.65 $X2=2.265 $Y2=1.87
r79 1 28 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=2.13
+ $Y=0.465 $X2=2.265 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_1%B 1 3 6 8 11
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.16 $X2=1.15 $Y2=1.16
r38 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.325
+ $X2=1.15 $Y2=1.16
r39 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.15 $Y=1.325 $X2=1.15
+ $Y2=1.985
r40 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=0.995
+ $X2=1.15 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.15 $Y=0.995 $X2=1.15
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_1%A 3 6 8 11 13
r34 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=1.63 $Y2=1.325
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=1.63 $Y2=0.995
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.16 $X2=1.63 $Y2=1.16
r37 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.57 $Y=1.985
+ $X2=1.57 $Y2=1.325
r38 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.57 $Y=0.56 $X2=1.57
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_1%C_N 3 6 8 11 13
r30 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.16
+ $X2=2.11 $Y2=1.325
r31 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.16
+ $X2=2.11 $Y2=0.995
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.16 $X2=2.11 $Y2=1.16
r33 6 14 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.055 $Y=1.86
+ $X2=2.055 $Y2=1.325
r34 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.055 $Y=0.675
+ $X2=2.055 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_1%Y 1 2 3 10 14 18 22 23
r31 27 35 0.650043 $w=4.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.315 $Y=1.675
+ $X2=0.315 $Y2=1.65
r32 23 27 5.17174 $w=4.6e-07 $l=1.95e-07 $layer=LI1_cond $X=0.315 $Y=1.87
+ $X2=0.315 $Y2=1.675
r33 22 35 3.1202 $w=4.58e-07 $l=1.2e-07 $layer=LI1_cond $X=0.315 $Y=1.53
+ $X2=0.315 $Y2=1.65
r34 21 22 26.7323 $w=2.78e-07 $l=6.2e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.445
r35 20 21 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.345 $Y2=0.825
r36 18 20 8.05053 $w=5.18e-07 $l=3.5e-07 $layer=LI1_cond $X=0.345 $Y=0.39
+ $X2=0.345 $Y2=0.74
r37 12 14 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.36 $Y=0.655
+ $X2=1.36 $Y2=0.495
r38 11 20 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.74
+ $X2=0.345 $Y2=0.74
r39 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.275 $Y=0.74
+ $X2=1.36 $Y2=0.655
r40 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.275 $Y=0.74
+ $X2=0.605 $Y2=0.74
r41 3 35 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.335
+ $Y=1.485 $X2=0.46 $Y2=1.65
r42 2 14 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.235 $X2=1.36 $Y2=0.495
r43 1 18 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.315
+ $Y=0.235 $X2=0.44 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_1%VPWR 1 6 9 10 11 21 22
r27 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r28 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r29 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 14 18 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r31 11 19 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r32 11 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r33 9 18 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.615 $Y=2.72 $X2=1.61
+ $Y2=2.72
r34 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=2.72
+ $X2=1.78 $Y2=2.72
r35 8 21 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.945 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=2.72
+ $X2=1.78 $Y2=2.72
r37 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=2.635 $X2=1.78
+ $Y2=2.72
r38 4 6 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.78 $Y=2.635
+ $X2=1.78 $Y2=2.21
r39 1 6 600 $w=1.7e-07 $l=7.8962e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.485 $X2=1.78 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__NOR3B_1%VGND 1 2 9 13 16 17 19 20 21 31 32
r38 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r39 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r40 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r41 25 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r42 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r43 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r44 19 28 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.61
+ $Y2=0
r45 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r46 18 31 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.53
+ $Y2=0
r47 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r48 16 24 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.69
+ $Y2=0
r49 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.94
+ $Y2=0
r50 15 28 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=1.61
+ $Y2=0
r51 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=0.94
+ $Y2=0
r52 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r53 11 13 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.39
r54 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=0.085 $X2=0.94
+ $Y2=0
r55 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.94 $Y=0.085
+ $X2=0.94 $Y2=0.39
r56 2 13 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.645
+ $Y=0.235 $X2=1.78 $Y2=0.39
r57 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.805
+ $Y=0.235 $X2=0.94 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__clkbuf_8.pex.spice
* Created: Tue Sep  1 19:00:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKBUF_8%A 3 5 7 10 12 14 15 16 24
c39 15 0 1.46759e-19 $X=0.23 $Y=0.85
r40 23 24 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.155
+ $X2=0.905 $Y2=1.155
r41 20 23 21.5061 $w=5.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.155
+ $X2=0.475 $Y2=1.155
r42 16 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r43 15 16 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=0.242 $Y=0.85
+ $X2=0.242 $Y2=1.16
r44 12 24 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.155
r45 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.985
r46 8 24 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=1.155
r47 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=0.445
r48 5 23 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.155
r49 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.985
r50 1 23 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=1.155
r51 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_8%A_110_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 49 53 57 61 63 65 69 73 77 84 87
r146 84 85 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.245
+ $Y=1.16 $X2=3.245 $Y2=1.16
r147 81 84 78.3661 $w=2.48e-07 $l=1.7e-06 $layer=LI1_cond $X=1.545 $Y=1.2
+ $X2=3.245 $Y2=1.2
r148 81 82 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.545
+ $Y=1.16 $X2=1.545 $Y2=1.16
r149 79 87 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=1.2
+ $X2=0.695 $Y2=1.2
r150 79 81 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=0.82 $Y=1.2
+ $X2=1.545 $Y2=1.2
r151 75 87 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.695 $Y2=1.2
r152 75 77 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.695 $Y2=1.69
r153 71 87 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.075
+ $X2=0.695 $Y2=1.2
r154 71 73 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=0.695 $Y=1.075
+ $X2=0.695 $Y2=0.445
r155 67 69 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.345 $Y=1.325
+ $X2=4.345 $Y2=1.985
r156 63 67 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=4.345 $Y=1.137
+ $X2=4.345 $Y2=1.325
r157 63 65 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.345 $Y=0.95
+ $X2=4.345 $Y2=0.445
r158 59 61 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.915 $Y=1.325
+ $X2=3.915 $Y2=1.985
r159 55 63 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=4.345 $Y2=1.137
r160 55 59 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=3.915 $Y2=1.325
r161 55 57 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.915 $Y=0.95
+ $X2=3.915 $Y2=0.445
r162 51 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.485 $Y=1.325
+ $X2=3.485 $Y2=1.985
r163 47 55 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.915 $Y2=1.137
r164 47 51 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.485 $Y2=1.325
r165 47 85 35.5938 $w=3.75e-07 $l=2.4e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.245 $Y2=1.137
r166 47 49 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.485 $Y=0.95
+ $X2=3.485 $Y2=0.445
r167 43 45 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.055 $Y=1.325
+ $X2=3.055 $Y2=1.985
r168 39 85 28.1785 $w=3.75e-07 $l=1.9e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.245 $Y2=1.137
r169 39 43 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.055 $Y2=1.325
r170 39 41 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.055 $Y=0.95
+ $X2=3.055 $Y2=0.445
r171 35 37 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.625 $Y=1.325
+ $X2=2.625 $Y2=1.985
r172 31 39 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=3.055 $Y2=1.137
r173 31 35 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=2.625 $Y2=1.325
r174 31 33 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.625 $Y=0.95
+ $X2=2.625 $Y2=0.445
r175 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.195 $Y=1.325
+ $X2=2.195 $Y2=1.985
r176 23 31 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.625 $Y2=1.137
r177 23 27 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.195 $Y2=1.325
r178 23 25 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.195 $Y=0.95
+ $X2=2.195 $Y2=0.445
r179 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=1.325
+ $X2=1.765 $Y2=1.985
r180 15 23 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=1.765 $Y=1.137
+ $X2=2.195 $Y2=1.137
r181 15 19 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=1.765 $Y=1.137
+ $X2=1.765 $Y2=1.325
r182 15 82 32.6277 $w=3.75e-07 $l=2.2e-07 $layer=POLY_cond $X=1.765 $Y=1.137
+ $X2=1.545 $Y2=1.137
r183 15 17 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.765 $Y=0.95
+ $X2=1.765 $Y2=0.445
r184 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.325
+ $X2=1.335 $Y2=1.985
r185 7 82 31.1446 $w=3.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.335 $Y=1.137
+ $X2=1.545 $Y2=1.137
r186 7 11 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=1.335 $Y=1.137
+ $X2=1.335 $Y2=1.325
r187 7 9 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.335 $Y=0.95
+ $X2=1.335 $Y2=0.445
r188 2 77 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.69
r189 1 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_8%VPWR 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 55 57 76 77 83
c78 6 0 4.2343e-20 $X=4.42 $Y=1.485
c79 5 0 1.26035e-19 $X=3.56 $Y=1.485
r80 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r81 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r82 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r83 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r84 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r85 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r86 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r87 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r88 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 65 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r90 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r91 62 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=2.72 $X2=1.12
+ $Y2=2.72
r92 62 64 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 61 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 58 80 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=0.195 $Y2=2.72
r96 58 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=2.72 $X2=0.69
+ $Y2=2.72
r97 57 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=1.12
+ $Y2=2.72
r98 57 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=2.72 $X2=0.69
+ $Y2=2.72
r99 55 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r100 55 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r101 53 73 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.43 $Y=2.72 $X2=4.37
+ $Y2=2.72
r102 53 54 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.43 $Y=2.72
+ $X2=4.577 $Y2=2.72
r103 52 76 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.725 $Y=2.72
+ $X2=4.83 $Y2=2.72
r104 52 54 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=4.725 $Y=2.72
+ $X2=4.577 $Y2=2.72
r105 50 70 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=2.72
+ $X2=3.45 $Y2=2.72
r106 50 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=2.72 $X2=3.7
+ $Y2=2.72
r107 49 73 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r108 49 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=2.72 $X2=3.7
+ $Y2=2.72
r109 47 67 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=2.72
+ $X2=2.53 $Y2=2.72
r110 47 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=2.72
+ $X2=2.84 $Y2=2.72
r111 46 70 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.97 $Y=2.72
+ $X2=3.45 $Y2=2.72
r112 46 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=2.72
+ $X2=2.84 $Y2=2.72
r113 44 64 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.98 $Y2=2.72
r115 43 67 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=2.72
+ $X2=2.53 $Y2=2.72
r116 43 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=2.72
+ $X2=1.98 $Y2=2.72
r117 39 54 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.577 $Y=2.635
+ $X2=4.577 $Y2=2.72
r118 39 41 16.2123 $w=2.93e-07 $l=4.15e-07 $layer=LI1_cond $X=4.577 $Y=2.635
+ $X2=4.577 $Y2=2.22
r119 35 51 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=2.635
+ $X2=3.7 $Y2=2.72
r120 35 37 18.3948 $w=2.58e-07 $l=4.15e-07 $layer=LI1_cond $X=3.7 $Y=2.635
+ $X2=3.7 $Y2=2.22
r121 31 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=2.635
+ $X2=2.84 $Y2=2.72
r122 31 33 18.3948 $w=2.58e-07 $l=4.15e-07 $layer=LI1_cond $X=2.84 $Y=2.635
+ $X2=2.84 $Y2=2.22
r123 27 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.72
r124 27 29 18.3948 $w=2.58e-07 $l=4.15e-07 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.22
r125 23 83 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r126 23 25 41.8869 $w=2.58e-07 $l=9.45e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=1.69
r127 19 80 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.195 $Y2=2.72
r128 19 21 36.9172 $w=2.93e-07 $l=9.45e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=1.69
r129 6 41 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.485 $X2=4.56 $Y2=2.22
r130 5 37 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.485 $X2=3.7 $Y2=2.22
r131 4 33 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.485 $X2=2.84 $Y2=2.22
r132 3 29 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.485 $X2=1.98 $Y2=2.22
r133 2 25 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=1.69
r134 1 21 300 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.69
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_8%X 1 2 3 4 5 6 7 8 27 31 32 33 37 41 43 47
+ 51 53 57 62 63 65 66 68 69 70 71
c117 69 0 1.68378e-19 $X=4.37 $Y=0.85
r118 71 86 2.23356 $w=6.15e-07 $l=1.2e-07 $layer=LI1_cond $X=4.245 $Y=1.615
+ $X2=4.245 $Y2=1.495
r119 71 86 0.314433 $w=9.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.245 $Y=1.47
+ $X2=4.245 $Y2=1.495
r120 70 71 3.52165 $w=9.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.245 $Y=1.19
+ $X2=4.245 $Y2=1.47
r121 69 85 1.61223 $w=6.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.82
+ $X2=4.245 $Y2=0.905
r122 69 70 3.39588 $w=9.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.245 $Y=0.92
+ $X2=4.245 $Y2=1.19
r123 69 85 0.18866 $w=9.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.245 $Y=0.92
+ $X2=4.245 $Y2=0.905
r124 55 69 1.61223 $w=6.15e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.245 $Y2=0.82
r125 55 57 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.445
r126 54 68 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=1.615
+ $X2=3.27 $Y2=1.615
r127 53 71 4.87019 $w=2.4e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=1.615
+ $X2=4.245 $Y2=1.615
r128 53 54 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=1.615
+ $X2=3.4 $Y2=1.615
r129 52 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=0.82 $X2=3.27
+ $Y2=0.82
r130 51 69 6.19726 $w=1.7e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=0.82
+ $X2=4.245 $Y2=0.82
r131 51 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=0.82
+ $X2=3.4 $Y2=0.82
r132 45 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.82
r133 45 47 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.445
r134 44 65 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=1.615
+ $X2=2.41 $Y2=1.615
r135 43 68 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=3.27 $Y2=1.615
r136 43 44 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=2.54 $Y2=1.615
r137 42 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=0.82
+ $X2=2.41 $Y2=0.82
r138 41 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=0.82
+ $X2=3.27 $Y2=0.82
r139 41 42 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=0.82 $X2=2.54
+ $Y2=0.82
r140 35 63 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.82
r141 35 37 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.445
r142 34 62 3.55196 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=1.55 $Y2=1.615
r143 33 65 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=1.615
+ $X2=2.41 $Y2=1.615
r144 33 34 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=1.615
+ $X2=1.68 $Y2=1.615
r145 31 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=0.82
+ $X2=2.41 $Y2=0.82
r146 31 32 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=0.82 $X2=1.68
+ $Y2=0.82
r147 25 32 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.68 $Y2=0.82
r148 25 27 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.55 $Y2=0.445
r149 8 71 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.485 $X2=4.13 $Y2=1.69
r150 7 68 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=1.485 $X2=3.27 $Y2=1.69
r151 6 65 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.485 $X2=2.41 $Y2=1.69
r152 5 62 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.485 $X2=1.55 $Y2=1.69
r153 4 57 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.445
r154 3 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.445
r155 2 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.445
r156 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_8%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 55 57 76 77 83
c84 57 0 1.46759e-19 $X=0.99 $Y=0
r85 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r86 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r87 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r88 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r89 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r90 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r91 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r92 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r93 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r94 65 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r95 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r96 62 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.12
+ $Y2=0
r97 62 64 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.61
+ $Y2=0
r98 61 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r99 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r100 58 80 3.93884 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r101 58 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.69
+ $Y2=0
r102 57 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.12
+ $Y2=0
r103 57 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.69
+ $Y2=0
r104 55 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r105 55 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r106 53 73 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.37
+ $Y2=0
r107 53 54 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.58
+ $Y2=0
r108 52 76 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.83
+ $Y2=0
r109 52 54 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.58
+ $Y2=0
r110 50 70 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.45
+ $Y2=0
r111 50 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.7
+ $Y2=0
r112 49 73 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.37
+ $Y2=0
r113 49 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.7
+ $Y2=0
r114 47 67 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.53
+ $Y2=0
r115 47 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.84
+ $Y2=0
r116 46 70 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=3.45
+ $Y2=0
r117 46 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.84
+ $Y2=0
r118 44 64 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.61
+ $Y2=0
r119 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.98
+ $Y2=0
r120 43 67 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.53
+ $Y2=0
r121 43 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.98
+ $Y2=0
r122 39 54 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r123 39 41 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.4
r124 35 51 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r125 35 37 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.4
r126 31 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r127 31 33 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.4
r128 27 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r129 27 29 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.4
r130 23 83 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r131 23 25 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.445
r132 19 80 3.17127 $w=2.45e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.195 $Y2=0
r133 19 21 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.267 $Y2=0.38
r134 6 41 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.235 $X2=4.565 $Y2=0.4
r135 5 37 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.4
r136 4 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.4
r137 3 29 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.4
r138 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.445
r139 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__a21oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_113_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.45e+11p pd=5.09e+06u as=2.95e+11p ps=2.59e+06u
M1001 VGND A2 a_199_47# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=3.66e+06u as=1.9175e+11p ps=1.89e+06u
M1002 a_113_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1003 Y B1 VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1004 VPWR A1 a_113_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_199_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


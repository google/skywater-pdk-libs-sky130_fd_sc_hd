# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlygate4sd3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.775000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.255000 3.595000 0.825000 ;
        RECT 3.210000 1.495000 3.595000 2.465000 ;
        RECT 3.315000 0.825000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.655000  0.085000 0.925000 0.545000 ;
        RECT 2.715000  0.085000 3.040000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.655000 2.175000 0.925000 2.635000 ;
        RECT 2.715000 2.175000 3.040000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.200000 0.255000 0.485000 0.715000 ;
      RECT 0.200000 0.715000 1.155000 0.885000 ;
      RECT 0.200000 1.785000 1.155000 2.005000 ;
      RECT 0.200000 2.005000 0.485000 2.465000 ;
      RECT 0.945000 0.885000 1.155000 1.785000 ;
      RECT 1.325000 0.255000 1.725000 1.055000 ;
      RECT 1.325000 1.055000 2.420000 1.615000 ;
      RECT 1.325000 1.615000 1.725000 2.465000 ;
      RECT 1.915000 0.255000 2.195000 0.715000 ;
      RECT 1.915000 0.715000 3.040000 0.885000 ;
      RECT 1.915000 1.785000 3.040000 2.005000 ;
      RECT 1.915000 2.005000 2.195000 2.465000 ;
      RECT 2.590000 0.885000 3.040000 0.995000 ;
      RECT 2.590000 0.995000 3.145000 1.325000 ;
      RECT 2.590000 1.325000 3.040000 1.785000 ;
  END
END sky130_fd_sc_hd__dlygate4sd3_1

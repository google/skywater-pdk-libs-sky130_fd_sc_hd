* File: sky130_fd_sc_hd__o21ai_0.pex.spice
* Created: Thu Aug 27 14:35:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21AI_0%A1 1 3 4 6 10 15 17 20 21
c36 10 0 1.75383e-19 $X=0.5 $Y=0.805
r37 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.25
+ $Y=1.04 $X2=0.25 $Y2=1.04
r38 17 21 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.25 $Y=1.53 $X2=0.25
+ $Y2=1.04
r39 13 20 121.085 $w=2.7e-07 $l=5.45e-07 $layer=POLY_cond $X=0.25 $Y=1.585
+ $X2=0.25 $Y2=1.04
r40 13 15 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.25 $Y=1.66
+ $X2=0.525 $Y2=1.66
r41 8 20 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.25 $Y=0.88 $X2=0.25
+ $Y2=1.04
r42 8 10 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.25 $Y=0.805 $X2=0.5
+ $Y2=0.805
r43 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.525 $Y=1.735
+ $X2=0.525 $Y2=1.66
r44 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.525 $Y=1.735
+ $X2=0.525 $Y2=2.165
r45 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.5 $Y=0.73 $X2=0.5
+ $Y2=0.805
r46 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=0.73 $X2=0.5
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_0%A2 3 7 11 14 15
c43 14 0 8.8227e-20 $X=0.84 $Y=1.21
c44 11 0 2.87357e-20 $X=0.69 $Y=1.19
c45 3 0 9.73357e-20 $X=0.915 $Y=2.165
r46 14 17 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.855 $Y=1.21
+ $X2=0.855 $Y2=1.375
r47 14 16 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.855 $Y=1.21
+ $X2=0.855 $Y2=1.045
r48 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.84
+ $Y=1.21 $X2=0.84 $Y2=1.21
r49 11 15 7.20277 $w=2.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=1.22
+ $X2=0.84 $Y2=1.22
r50 7 16 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.93 $Y=0.445 $X2=0.93
+ $Y2=1.045
r51 3 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.915 $Y=2.165
+ $X2=0.915 $Y2=1.375
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_0%B1 3 7 9 15
c28 15 0 1.66457e-20 $X=1.6 $Y=1.52
c29 9 0 9.73357e-20 $X=1.61 $Y=1.53
c30 7 0 1.209e-20 $X=1.36 $Y=0.445
r31 13 15 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.36 $Y=1.52 $X2=1.6
+ $Y2=1.52
r32 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.345 $Y=1.52
+ $X2=1.36 $Y2=1.52
r33 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6 $Y=1.52
+ $X2=1.6 $Y2=1.52
r34 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.355
+ $X2=1.36 $Y2=1.52
r35 5 7 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.36 $Y=1.355 $X2=1.36
+ $Y2=0.445
r36 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.685
+ $X2=1.345 $Y2=1.52
r37 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.345 $Y=1.685
+ $X2=1.345 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_0%VPWR 1 2 7 9 11 13 15 17 27
r25 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r26 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r27 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r28 18 23 4.66755 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=2.72
+ $X2=0.237 $Y2=2.72
r29 18 20 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.475 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 17 26 4.04813 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.655 $Y2=2.72
r31 17 20 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.47 $Y=2.72 $X2=1.15
+ $Y2=2.72
r32 15 21 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r33 15 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r34 11 26 3.1291 $w=2.55e-07 $l=1.1025e-07 $layer=LI1_cond $X=1.597 $Y=2.635
+ $X2=1.655 $Y2=2.72
r35 11 13 27.7942 $w=2.53e-07 $l=6.15e-07 $layer=LI1_cond $X=1.597 $Y=2.635
+ $X2=1.597 $Y2=2.02
r36 7 23 3.09863 $w=3.3e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.31 $Y=2.635
+ $X2=0.237 $Y2=2.72
r37 7 9 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=0.31 $Y=2.635 $X2=0.31
+ $Y2=1.99
r38 2 13 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=1.42
+ $Y=1.845 $X2=1.56 $Y2=2.02
r39 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=1.845 $X2=0.31 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_0%Y 1 2 9 11 14 15 20 23
c37 9 0 8.8227e-20 $X=1.597 $Y=0.955
r38 20 23 7.56828 $w=3.33e-07 $l=2.2e-07 $layer=LI1_cond $X=1.132 $Y=2.21
+ $X2=1.132 $Y2=1.99
r39 15 23 10.6644 $w=3.33e-07 $l=3.1e-07 $layer=LI1_cond $X=1.132 $Y=1.68
+ $X2=1.132 $Y2=1.99
r40 14 15 8.63814 $w=3.33e-07 $l=1.7e-07 $layer=LI1_cond $X=1.155 $Y=1.51
+ $X2=1.155 $Y2=1.68
r41 9 16 21.9861 $w=1.68e-07 $l=3.37e-07 $layer=LI1_cond $X=1.597 $Y=1.04
+ $X2=1.26 $Y2=1.04
r42 9 11 20.6227 $w=2.83e-07 $l=5.1e-07 $layer=LI1_cond $X=1.597 $Y=0.955
+ $X2=1.597 $Y2=0.445
r43 7 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=1.125
+ $X2=1.26 $Y2=1.04
r44 7 14 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.26 $Y=1.125
+ $X2=1.26 $Y2=1.51
r45 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.99
+ $Y=1.845 $X2=1.13 $Y2=1.99
r46 1 11 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.575 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_0%A_32_47# 1 2 9 11 12 15
r25 13 15 8.33682 $w=2.33e-07 $l=1.7e-07 $layer=LI1_cond $X=1.167 $Y=0.615
+ $X2=1.167 $Y2=0.445
r26 11 13 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=1.05 $Y=0.7
+ $X2=1.167 $Y2=0.615
r27 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.05 $Y=0.7 $X2=0.38
+ $Y2=0.7
r28 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.25 $Y=0.615
+ $X2=0.38 $Y2=0.7
r29 7 9 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.25 $Y=0.615 $X2=0.25
+ $Y2=0.445
r30 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.145 $Y2=0.445
r31 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_0%VGND 1 6 8 10 17 18 21
c29 18 0 1.75383e-19 $X=1.61 $Y=0
r30 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r31 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r32 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r33 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.715
+ $Y2=0
r34 15 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.61
+ $Y2=0
r35 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.715
+ $Y2=0
r36 10 12 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.23
+ $Y2=0
r37 8 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r38 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r39 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r40 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.36
r41 1 6 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.36
.ends


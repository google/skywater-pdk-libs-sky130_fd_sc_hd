* File: sky130_fd_sc_hd__o21ai_0.spice.SKY130_FD_SC_HD__O21AI_0.pxi
* Created: Thu Aug 27 14:35:31 2020
* 
x_PM_SKY130_FD_SC_HD__O21AI_0%A1 N_A1_c_41_n N_A1_M1005_g N_A1_c_45_n
+ N_A1_M1001_g N_A1_c_42_n N_A1_c_46_n A1 N_A1_c_43_n N_A1_c_44_n
+ PM_SKY130_FD_SC_HD__O21AI_0%A1
x_PM_SKY130_FD_SC_HD__O21AI_0%A2 N_A2_M1003_g N_A2_M1004_g A2 N_A2_c_78_n
+ N_A2_c_79_n PM_SKY130_FD_SC_HD__O21AI_0%A2
x_PM_SKY130_FD_SC_HD__O21AI_0%B1 N_B1_M1000_g N_B1_M1002_g B1 N_B1_c_124_n
+ PM_SKY130_FD_SC_HD__O21AI_0%B1
x_PM_SKY130_FD_SC_HD__O21AI_0%VPWR N_VPWR_M1001_s N_VPWR_M1000_d N_VPWR_c_149_n
+ N_VPWR_c_150_n N_VPWR_c_151_n N_VPWR_c_152_n VPWR N_VPWR_c_153_n
+ N_VPWR_c_148_n PM_SKY130_FD_SC_HD__O21AI_0%VPWR
x_PM_SKY130_FD_SC_HD__O21AI_0%Y N_Y_M1002_d N_Y_M1003_d N_Y_c_174_n N_Y_c_175_n
+ N_Y_c_176_n N_Y_c_178_n Y N_Y_c_180_n PM_SKY130_FD_SC_HD__O21AI_0%Y
x_PM_SKY130_FD_SC_HD__O21AI_0%A_32_47# N_A_32_47#_M1005_s N_A_32_47#_M1004_d
+ N_A_32_47#_c_211_n N_A_32_47#_c_212_n N_A_32_47#_c_213_n N_A_32_47#_c_230_p
+ PM_SKY130_FD_SC_HD__O21AI_0%A_32_47#
x_PM_SKY130_FD_SC_HD__O21AI_0%VGND N_VGND_M1005_d N_VGND_c_236_n VGND
+ N_VGND_c_237_n N_VGND_c_238_n N_VGND_c_239_n N_VGND_c_240_n
+ PM_SKY130_FD_SC_HD__O21AI_0%VGND
cc_1 VNB N_A1_c_41_n 0.017348f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.73
cc_2 VNB N_A1_c_42_n 0.0323624f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.805
cc_3 VNB N_A1_c_43_n 0.0315837f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.04
cc_4 VNB N_A1_c_44_n 0.0175838f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.04
cc_5 VNB N_A2_M1004_g 0.0327073f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=0.805
cc_6 VNB N_A2_c_78_n 0.0201472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A2_c_79_n 0.00379687f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.66
cc_8 VNB N_B1_M1002_g 0.0530437f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=0.805
cc_9 VNB N_VPWR_c_148_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_Y_c_174_n 0.0145493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_175_n 0.0306185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_Y_c_176_n 0.00139074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_32_47#_c_211_n 0.012774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_32_47#_c_212_n 0.0111597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_32_47#_c_213_n 0.00468366f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.66
cc_16 VNB N_VGND_c_236_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=2.165
cc_17 VNB N_VGND_c_237_n 0.0154802f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=0.805
cc_18 VNB N_VGND_c_238_n 0.0262158f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_19 VNB N_VGND_c_239_n 0.125064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_240_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.04
cc_21 VPB N_A1_c_45_n 0.0206581f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.735
cc_22 VPB N_A1_c_46_n 0.0338372f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.66
cc_23 VPB N_A1_c_43_n 0.0192887f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.04
cc_24 VPB N_A1_c_44_n 0.0147077f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.04
cc_25 VPB N_A2_M1003_g 0.03431f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=0.445
cc_26 VPB A2 0.0112066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A2_c_78_n 0.0101189f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A2_c_79_n 7.20874e-19 $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.66
cc_29 VPB N_B1_M1000_g 0.0254883f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=0.445
cc_30 VPB N_B1_M1002_g 0.00372857f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=0.805
cc_31 VPB B1 0.0043162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_B1_c_124_n 0.0568805f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.66
cc_33 VPB N_VPWR_c_149_n 0.0119347f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=0.805
cc_34 VPB N_VPWR_c_150_n 0.030433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_151_n 0.010745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_152_n 0.02835f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.585
cc_37 VPB N_VPWR_c_153_n 0.0271923f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_38 VPB N_VPWR_c_148_n 0.0457041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_176_n 0.00158118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_Y_c_178_n 0.00701444f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.66
cc_41 N_A1_c_46_n N_A2_M1003_g 0.0527348f $X=0.525 $Y=1.66 $X2=0 $Y2=0
cc_42 N_A1_c_43_n N_A2_M1003_g 0.00236039f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_43 N_A1_c_41_n N_A2_M1004_g 0.0212891f $X=0.5 $Y=0.73 $X2=0 $Y2=0
cc_44 N_A1_c_43_n N_A2_M1004_g 0.00154274f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_45 N_A1_c_44_n N_A2_M1004_g 0.00179655f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_46 N_A1_c_46_n A2 0.00104575f $X=0.525 $Y=1.66 $X2=0 $Y2=0
cc_47 N_A1_c_43_n A2 5.17965e-19 $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_48 N_A1_c_44_n A2 0.0200336f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_49 N_A1_c_43_n N_A2_c_78_n 0.0125056f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_50 N_A1_c_44_n N_A2_c_78_n 0.00199379f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_51 N_A1_c_43_n N_A2_c_79_n 8.5058e-19 $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_52 N_A1_c_44_n N_A2_c_79_n 0.0186676f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_53 N_A1_c_45_n N_VPWR_c_150_n 0.0183211f $X=0.525 $Y=1.735 $X2=0 $Y2=0
cc_54 N_A1_c_46_n N_VPWR_c_150_n 0.00961874f $X=0.525 $Y=1.66 $X2=0 $Y2=0
cc_55 N_A1_c_44_n N_VPWR_c_150_n 0.020316f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_56 N_A1_c_45_n N_VPWR_c_153_n 0.00486043f $X=0.525 $Y=1.735 $X2=0 $Y2=0
cc_57 N_A1_c_45_n N_VPWR_c_148_n 0.00822386f $X=0.525 $Y=1.735 $X2=0 $Y2=0
cc_58 N_A1_c_46_n N_Y_c_178_n 0.00138735f $X=0.525 $Y=1.66 $X2=0 $Y2=0
cc_59 N_A1_c_45_n N_Y_c_180_n 0.00138735f $X=0.525 $Y=1.735 $X2=0 $Y2=0
cc_60 N_A1_c_41_n N_A_32_47#_c_212_n 0.00779725f $X=0.5 $Y=0.73 $X2=0 $Y2=0
cc_61 N_A1_c_42_n N_A_32_47#_c_212_n 0.00858629f $X=0.5 $Y=0.805 $X2=0 $Y2=0
cc_62 N_A1_c_44_n N_A_32_47#_c_212_n 0.00267933f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_63 N_A1_c_42_n N_A_32_47#_c_213_n 0.0130813f $X=0.5 $Y=0.805 $X2=0 $Y2=0
cc_64 N_A1_c_44_n N_A_32_47#_c_213_n 0.0214759f $X=0.25 $Y=1.04 $X2=0 $Y2=0
cc_65 N_A1_c_41_n N_VGND_c_236_n 0.00867088f $X=0.5 $Y=0.73 $X2=0 $Y2=0
cc_66 N_A1_c_41_n N_VGND_c_237_n 0.00351072f $X=0.5 $Y=0.73 $X2=0 $Y2=0
cc_67 N_A1_c_42_n N_VGND_c_237_n 8.86695e-19 $X=0.5 $Y=0.805 $X2=0 $Y2=0
cc_68 N_A1_c_41_n N_VGND_c_239_n 0.00510895f $X=0.5 $Y=0.73 $X2=0 $Y2=0
cc_69 N_A2_M1004_g N_B1_M1002_g 0.039044f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A2_c_79_n N_B1_M1002_g 2.51827e-19 $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A2_M1003_g N_B1_c_124_n 0.0271657f $X=0.915 $Y=2.165 $X2=0 $Y2=0
cc_72 N_A2_c_78_n N_B1_c_124_n 9.21608e-19 $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A2_M1003_g N_VPWR_c_150_n 0.00298263f $X=0.915 $Y=2.165 $X2=0 $Y2=0
cc_74 N_A2_M1003_g N_VPWR_c_153_n 0.0054895f $X=0.915 $Y=2.165 $X2=0 $Y2=0
cc_75 N_A2_M1003_g N_VPWR_c_148_n 0.00988587f $X=0.915 $Y=2.165 $X2=0 $Y2=0
cc_76 N_A2_M1004_g N_Y_c_174_n 0.00383318f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A2_c_79_n N_Y_c_174_n 0.00194545f $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A2_M1003_g N_Y_c_176_n 0.00104671f $X=0.915 $Y=2.165 $X2=0 $Y2=0
cc_79 A2 N_Y_c_176_n 0.00690341f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A2_c_78_n N_Y_c_176_n 9.92215e-19 $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A2_c_79_n N_Y_c_176_n 0.0164027f $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A2_M1003_g N_Y_c_178_n 0.00444285f $X=0.915 $Y=2.165 $X2=0 $Y2=0
cc_83 A2 N_Y_c_178_n 0.00943104f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_84 N_A2_c_78_n N_Y_c_178_n 4.25964e-19 $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A2_c_79_n N_Y_c_178_n 0.00311069f $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A2_M1003_g N_Y_c_180_n 0.0152308f $X=0.915 $Y=2.165 $X2=0 $Y2=0
cc_87 N_A2_M1004_g N_A_32_47#_c_212_n 0.0119679f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A2_c_78_n N_A_32_47#_c_212_n 0.00329224f $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A2_c_79_n N_A_32_47#_c_212_n 0.0183711f $X=0.84 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A2_M1004_g N_VGND_c_236_n 0.00757764f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A2_M1004_g N_VGND_c_238_n 0.00351072f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A2_M1004_g N_VGND_c_239_n 0.00414308f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_93 N_B1_M1000_g N_VPWR_c_152_n 0.00450113f $X=1.345 $Y=2.165 $X2=0 $Y2=0
cc_94 B1 N_VPWR_c_152_n 0.0172962f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_95 N_B1_c_124_n N_VPWR_c_152_n 0.00350097f $X=1.6 $Y=1.52 $X2=0 $Y2=0
cc_96 N_B1_M1000_g N_VPWR_c_153_n 0.00541359f $X=1.345 $Y=2.165 $X2=0 $Y2=0
cc_97 N_B1_M1000_g N_VPWR_c_148_n 0.0105306f $X=1.345 $Y=2.165 $X2=0 $Y2=0
cc_98 N_B1_M1002_g N_Y_c_174_n 0.017654f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_99 B1 N_Y_c_174_n 0.0128134f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_100 N_B1_c_124_n N_Y_c_174_n 0.00453252f $X=1.6 $Y=1.52 $X2=0 $Y2=0
cc_101 N_B1_M1002_g N_Y_c_175_n 0.0106162f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_102 N_B1_M1002_g N_Y_c_176_n 0.0115309f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_103 B1 N_Y_c_176_n 0.0231565f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_104 N_B1_c_124_n N_Y_c_176_n 0.00437126f $X=1.6 $Y=1.52 $X2=0 $Y2=0
cc_105 N_B1_c_124_n N_Y_c_178_n 0.00784516f $X=1.6 $Y=1.52 $X2=0 $Y2=0
cc_106 N_B1_M1000_g N_Y_c_180_n 0.0162104f $X=1.345 $Y=2.165 $X2=0 $Y2=0
cc_107 B1 N_Y_c_180_n 2.7028e-19 $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_108 N_B1_M1002_g N_A_32_47#_c_212_n 0.00131663f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_109 N_B1_M1002_g N_VGND_c_236_n 0.00121802f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_110 N_B1_M1002_g N_VGND_c_238_n 0.00585385f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_111 N_B1_M1002_g N_VGND_c_239_n 0.0118661f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_112 N_VPWR_c_148_n A_120_369# 0.0102589f $X=1.61 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_113 N_VPWR_c_148_n N_Y_M1003_d 0.00223231f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_114 N_VPWR_c_150_n N_Y_c_180_n 0.020299f $X=0.31 $Y=1.99 $X2=0 $Y2=0
cc_115 N_VPWR_c_153_n N_Y_c_180_n 0.0192662f $X=1.47 $Y=2.72 $X2=0 $Y2=0
cc_116 N_VPWR_c_148_n N_Y_c_180_n 0.0124371f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_117 N_Y_c_174_n N_A_32_47#_c_212_n 0.00906817f $X=1.597 $Y=0.955 $X2=0 $Y2=0
cc_118 N_Y_c_175_n N_A_32_47#_c_212_n 0.0125455f $X=1.575 $Y=0.445 $X2=0 $Y2=0
cc_119 N_Y_c_175_n N_VGND_c_238_n 0.0161202f $X=1.575 $Y=0.445 $X2=0 $Y2=0
cc_120 N_Y_M1002_d N_VGND_c_239_n 0.00288166f $X=1.435 $Y=0.235 $X2=0 $Y2=0
cc_121 N_Y_c_175_n N_VGND_c_239_n 0.0107647f $X=1.575 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_32_47#_c_212_n N_VGND_M1005_d 0.00169105f $X=1.05 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_32_47#_c_212_n N_VGND_c_236_n 0.0159085f $X=1.05 $Y=0.7 $X2=0 $Y2=0
cc_124 N_A_32_47#_c_211_n N_VGND_c_237_n 0.0150357f $X=0.285 $Y=0.445 $X2=0
+ $Y2=0
cc_125 N_A_32_47#_c_212_n N_VGND_c_237_n 0.0025909f $X=1.05 $Y=0.7 $X2=0 $Y2=0
cc_126 N_A_32_47#_c_212_n N_VGND_c_238_n 0.0025909f $X=1.05 $Y=0.7 $X2=0 $Y2=0
cc_127 N_A_32_47#_c_230_p N_VGND_c_238_n 0.0119167f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_128 N_A_32_47#_M1005_s N_VGND_c_239_n 0.00229482f $X=0.16 $Y=0.235 $X2=0
+ $Y2=0
cc_129 N_A_32_47#_M1004_d N_VGND_c_239_n 0.00239355f $X=1.005 $Y=0.235 $X2=0
+ $Y2=0
cc_130 N_A_32_47#_c_211_n N_VGND_c_239_n 0.00973428f $X=0.285 $Y=0.445 $X2=0
+ $Y2=0
cc_131 N_A_32_47#_c_212_n N_VGND_c_239_n 0.0100658f $X=1.05 $Y=0.7 $X2=0 $Y2=0
cc_132 N_A_32_47#_c_230_p N_VGND_c_239_n 0.00879104f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__ha_4.spice.pex
* Created: Thu Aug 27 14:22:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__HA_4%A_79_21# 1 2 3 10 12 15 17 19 22 24 26 29 31 33
+ 36 38 44 47 50 52 53 55 59 61 62 64 65 67 69
c140 55 0 9.8674e-20 $X=2.88 $Y=0.73
c141 47 0 1.06093e-19 $X=2.225 $Y=1.16
c142 29 0 9.33312e-20 $X=1.31 $Y=1.985
c143 22 0 1.29575e-19 $X=0.89 $Y=1.985
c144 3 0 1.59207e-19 $X=4.03 $Y=1.485
r145 70 73 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.665 $Y=1.85
+ $X2=2.855 $Y2=1.85
r146 65 67 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.7 $Y=2.29
+ $X2=4.165 $Y2=2.29
r147 64 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=2.205
+ $X2=3.7 $Y2=2.29
r148 63 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.615 $Y=1.935
+ $X2=3.615 $Y2=2.205
r149 62 73 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=1.85
+ $X2=2.855 $Y2=1.85
r150 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.53 $Y=1.85
+ $X2=3.615 $Y2=1.935
r151 61 62 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.53 $Y=1.85
+ $X2=2.94 $Y2=1.85
r152 57 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=1.935
+ $X2=2.855 $Y2=1.85
r153 57 59 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.855 $Y=1.935
+ $X2=2.855 $Y2=2.19
r154 53 55 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.75 $Y=0.73
+ $X2=2.88 $Y2=0.73
r155 52 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=1.765
+ $X2=2.665 $Y2=1.85
r156 51 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=1.245
+ $X2=2.665 $Y2=1.16
r157 51 52 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.665 $Y=1.245
+ $X2=2.665 $Y2=1.765
r158 50 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=1.075
+ $X2=2.665 $Y2=1.16
r159 49 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.665 $Y=0.815
+ $X2=2.75 $Y2=0.73
r160 49 50 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.665 $Y=0.815
+ $X2=2.665 $Y2=1.075
r161 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.225
+ $Y=1.16 $X2=2.225 $Y2=1.16
r162 44 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=1.16
+ $X2=2.665 $Y2=1.16
r163 44 46 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.58 $Y=1.16
+ $X2=2.225 $Y2=1.16
r164 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r165 41 42 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r166 39 41 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r167 38 47 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.805 $Y=1.16
+ $X2=2.225 $Y2=1.16
r168 38 43 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=1.16
+ $X2=1.73 $Y2=1.16
r169 34 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r170 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r171 31 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r172 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r173 27 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r174 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r175 24 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r176 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r177 20 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r178 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r179 17 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r180 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r181 13 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r182 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r183 10 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r184 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r185 3 67 600 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.485 $X2=4.165 $Y2=2.29
r186 2 73 600 $w=1.7e-07 $l=4.272e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.485 $X2=2.855 $Y2=1.85
r187 2 59 600 $w=1.7e-07 $l=7.69545e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.485 $X2=2.855 $Y2=2.19
r188 1 55 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%A_514_199# 1 2 3 12 14 16 19 21 23 24 26 29 31
+ 33 36 38 40 43 45 47 50 54 57 58 60 61 62 65 67 69 75 78 79 81 82 84 86 89 92
+ 93 94 100 107
c220 107 0 1.47169e-19 $X=8.73 $Y=1.16
c221 93 0 1.51157e-19 $X=6.76 $Y=1.94
c222 54 0 1.06093e-19 $X=3.005 $Y=1.16
r223 106 107 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.31 $Y=1.16
+ $X2=8.73 $Y2=1.16
r224 102 104 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=7.47 $Y=1.16
+ $X2=7.89 $Y2=1.16
r225 99 100 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.065 $Y=1.16
+ $X2=3.09 $Y2=1.16
r226 95 97 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.645 $Y=1.16
+ $X2=2.67 $Y2=1.16
r227 90 106 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=8.06 $Y=1.16
+ $X2=8.31 $Y2=1.16
r228 90 104 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=8.06 $Y=1.16
+ $X2=7.89 $Y2=1.16
r229 89 90 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.06
+ $Y=1.16 $X2=8.06 $Y2=1.16
r230 87 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=1.16
+ $X2=7.31 $Y2=1.16
r231 87 89 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.395 $Y=1.16
+ $X2=8.06 $Y2=1.16
r232 85 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=1.245
+ $X2=7.31 $Y2=1.16
r233 85 86 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.31 $Y=1.245
+ $X2=7.31 $Y2=1.855
r234 84 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=1.075
+ $X2=7.31 $Y2=1.16
r235 83 84 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.31 $Y=0.815
+ $X2=7.31 $Y2=1.075
r236 81 83 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.225 $Y=0.73
+ $X2=7.31 $Y2=0.815
r237 81 82 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.225 $Y=0.73
+ $X2=6.875 $Y2=0.73
r238 80 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=1.94
+ $X2=6.76 $Y2=1.94
r239 79 86 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.225 $Y=1.94
+ $X2=7.31 $Y2=1.855
r240 79 80 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.225 $Y=1.94
+ $X2=6.845 $Y2=1.94
r241 78 82 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.79 $Y=0.645
+ $X2=6.875 $Y2=0.73
r242 77 78 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.79 $Y=0.465
+ $X2=6.79 $Y2=0.645
r243 73 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=2.025
+ $X2=6.76 $Y2=1.94
r244 73 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.76 $Y=2.025
+ $X2=6.76 $Y2=2.19
r245 69 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.705 $Y=0.38
+ $X2=6.79 $Y2=0.465
r246 69 71 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.705 $Y=0.38
+ $X2=6.34 $Y2=0.38
r247 68 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=1.94
+ $X2=5.92 $Y2=1.94
r248 67 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=1.94
+ $X2=6.76 $Y2=1.94
r249 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.675 $Y=1.94
+ $X2=6.005 $Y2=1.94
r250 63 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.025
+ $X2=5.92 $Y2=1.94
r251 63 65 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.92 $Y=2.025
+ $X2=5.92 $Y2=2.19
r252 61 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=1.94
+ $X2=5.92 $Y2=1.94
r253 61 62 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=5.835 $Y=1.94
+ $X2=4.04 $Y2=1.94
r254 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.955 $Y=1.855
+ $X2=4.04 $Y2=1.94
r255 59 60 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.955 $Y=1.595
+ $X2=3.955 $Y2=1.855
r256 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.87 $Y=1.51
+ $X2=3.955 $Y2=1.595
r257 57 58 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.87 $Y=1.51
+ $X2=3.09 $Y2=1.51
r258 55 99 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.005 $Y=1.16
+ $X2=3.065 $Y2=1.16
r259 55 97 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=3.005 $Y=1.16
+ $X2=2.67 $Y2=1.16
r260 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.005
+ $Y=1.16 $X2=3.005 $Y2=1.16
r261 52 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.005 $Y=1.425
+ $X2=3.09 $Y2=1.51
r262 52 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.005 $Y=1.425
+ $X2=3.005 $Y2=1.16
r263 48 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.73 $Y=1.325
+ $X2=8.73 $Y2=1.16
r264 48 50 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.73 $Y=1.325
+ $X2=8.73 $Y2=1.985
r265 45 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.73 $Y=0.995
+ $X2=8.73 $Y2=1.16
r266 45 47 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.73 $Y=0.995
+ $X2=8.73 $Y2=0.56
r267 41 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.31 $Y=1.325
+ $X2=8.31 $Y2=1.16
r268 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.31 $Y=1.325
+ $X2=8.31 $Y2=1.985
r269 38 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.31 $Y=0.995
+ $X2=8.31 $Y2=1.16
r270 38 40 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.31 $Y=0.995
+ $X2=8.31 $Y2=0.56
r271 34 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.89 $Y=1.325
+ $X2=7.89 $Y2=1.16
r272 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.89 $Y=1.325
+ $X2=7.89 $Y2=1.985
r273 31 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.89 $Y=0.995
+ $X2=7.89 $Y2=1.16
r274 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.89 $Y=0.995
+ $X2=7.89 $Y2=0.56
r275 27 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.47 $Y=1.325
+ $X2=7.47 $Y2=1.16
r276 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.47 $Y=1.325
+ $X2=7.47 $Y2=1.985
r277 24 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.47 $Y=0.995
+ $X2=7.47 $Y2=1.16
r278 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.47 $Y=0.995
+ $X2=7.47 $Y2=0.56
r279 21 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=1.16
r280 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=0.56
r281 17 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.325
+ $X2=3.065 $Y2=1.16
r282 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.065 $Y=1.325
+ $X2=3.065 $Y2=1.985
r283 14 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=1.16
r284 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=0.56
r285 10 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.325
+ $X2=2.645 $Y2=1.16
r286 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.645 $Y=1.325
+ $X2=2.645 $Y2=1.985
r287 3 75 600 $w=1.7e-07 $l=7.69545e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.485 $X2=6.76 $Y2=2.19
r288 2 65 600 $w=1.7e-07 $l=7.69545e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.485 $X2=5.92 $Y2=2.19
r289 1 71 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.205
+ $Y=0.235 $X2=6.34 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%A 1 3 6 10 12 14 17 19 21 22 24 27 29 32 35 36
+ 37 40 41 44 45 46 57 58 60
c156 58 0 1.47169e-19 $X=6.97 $Y=1.16
c157 57 0 3.40373e-19 $X=6.97 $Y=1.16
c158 46 0 1.38713e-19 $X=6.665 $Y=1.53
c159 35 0 1.59207e-19 $X=4.295 $Y=1.505
c160 1 0 9.8674e-20 $X=3.51 $Y=0.995
r161 59 67 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=1.325
+ $X2=6.695 $Y2=1.16
r162 58 67 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.97 $Y=1.16
+ $X2=6.695 $Y2=1.16
r163 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.97
+ $Y=1.16 $X2=6.97 $Y2=1.16
r164 46 60 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.695 $Y=1.59
+ $X2=6.695 $Y2=1.505
r165 46 60 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=6.695 $Y=1.475
+ $X2=6.695 $Y2=1.505
r166 46 59 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.695 $Y=1.475
+ $X2=6.695 $Y2=1.325
r167 45 67 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=6.665 $Y=1.16
+ $X2=6.695 $Y2=1.16
r168 43 46 33.5235 $w=2.78e-07 $l=7.85e-07 $layer=LI1_cond $X=5.795 $Y=1.59
+ $X2=6.58 $Y2=1.59
r169 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.795 $Y=1.59
+ $X2=5.71 $Y2=1.59
r170 41 55 8.36806 $w=2.88e-07 $l=5e-08 $layer=POLY_cond $X=5.71 $Y=1.16
+ $X2=5.76 $Y2=1.16
r171 41 53 61.9236 $w=2.88e-07 $l=3.7e-07 $layer=POLY_cond $X=5.71 $Y=1.16
+ $X2=5.34 $Y2=1.16
r172 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.71
+ $Y=1.16 $X2=5.71 $Y2=1.16
r173 38 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=1.505
+ $X2=5.71 $Y2=1.59
r174 38 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.71 $Y=1.505
+ $X2=5.71 $Y2=1.16
r175 36 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=1.59
+ $X2=5.71 $Y2=1.59
r176 36 37 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=5.625 $Y=1.59
+ $X2=4.38 $Y2=1.59
r177 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.295 $Y=1.505
+ $X2=4.38 $Y2=1.59
r178 34 35 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.295 $Y=1.245
+ $X2=4.295 $Y2=1.505
r179 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.51
+ $Y=1.16 $X2=3.51 $Y2=1.16
r180 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.21 $Y=1.16
+ $X2=4.295 $Y2=1.245
r181 29 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.21 $Y=1.16 $X2=3.51
+ $Y2=1.16
r182 25 57 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=1.325
+ $X2=6.97 $Y2=1.16
r183 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.97 $Y=1.325
+ $X2=6.97 $Y2=1.985
r184 22 57 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=1.16
r185 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=0.56
r186 19 55 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.76 $Y=0.995
+ $X2=5.76 $Y2=1.16
r187 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.76 $Y=0.995
+ $X2=5.76 $Y2=0.56
r188 15 41 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.71 $Y=1.325
+ $X2=5.71 $Y2=1.16
r189 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.71 $Y=1.325
+ $X2=5.71 $Y2=1.985
r190 12 53 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.34 $Y=0.995
+ $X2=5.34 $Y2=1.16
r191 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.34 $Y=0.995
+ $X2=5.34 $Y2=0.56
r192 8 53 40.1667 $w=2.88e-07 $l=3.11769e-07 $layer=POLY_cond $X=5.1 $Y=1.325
+ $X2=5.34 $Y2=1.16
r193 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.1 $Y=1.325 $X2=5.1
+ $Y2=1.985
r194 4 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=1.325
+ $X2=3.51 $Y2=1.16
r195 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.51 $Y=1.325
+ $X2=3.51 $Y2=1.985
r196 1 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.16
r197 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 33 35 39
+ 40 42 44 45 56 58 60
c128 60 0 3.71106e-19 $X=6.205 $Y=0.85
c129 56 0 1.38713e-19 $X=6.55 $Y=1.16
r130 58 60 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.2 $Y=0.825
+ $X2=6.2 $Y2=0.85
r131 54 56 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=6.23 $Y=1.16
+ $X2=6.55 $Y2=1.16
r132 51 54 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.13 $Y=1.16 $X2=6.23
+ $Y2=1.16
r133 45 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.23
+ $Y=1.16 $X2=6.23 $Y2=1.16
r134 44 58 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.2 $Y=0.74 $X2=6.2
+ $Y2=0.825
r135 44 45 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.2 $Y=0.88 $X2=6.2
+ $Y2=1.16
r136 44 60 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=6.2 $Y=0.88 $X2=6.2
+ $Y2=0.85
r137 42 43 21.1633 $w=1.96e-07 $l=3.4e-07 $layer=LI1_cond $X=5.41 $Y=0.74
+ $X2=5.41 $Y2=1.08
r138 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.16 $X2=4.635 $Y2=1.16
r139 36 42 1.57051 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.535 $Y=0.74
+ $X2=5.41 $Y2=0.74
r140 35 44 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.085 $Y=0.74
+ $X2=6.2 $Y2=0.74
r141 35 36 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.085 $Y=0.74
+ $X2=5.535 $Y2=0.74
r142 34 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.72 $Y=1.08
+ $X2=4.635 $Y2=1.08
r143 33 43 1.57051 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.285 $Y=1.08
+ $X2=5.41 $Y2=1.08
r144 33 34 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.285 $Y=1.08
+ $X2=4.72 $Y2=1.08
r145 30 32 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.955 $Y=1.16
+ $X2=4.375 $Y2=1.16
r146 29 40 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=4.45 $Y=1.16
+ $X2=4.635 $Y2=1.16
r147 29 32 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.45 $Y=1.16
+ $X2=4.375 $Y2=1.16
r148 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=1.325
+ $X2=6.55 $Y2=1.16
r149 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.55 $Y=1.325
+ $X2=6.55 $Y2=1.985
r150 22 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=0.995
+ $X2=6.55 $Y2=1.16
r151 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.55 $Y=0.995
+ $X2=6.55 $Y2=0.56
r152 18 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=1.325
+ $X2=6.13 $Y2=1.16
r153 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.13 $Y=1.325
+ $X2=6.13 $Y2=1.985
r154 15 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=1.16
r155 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=0.56
r156 11 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.325
+ $X2=4.375 $Y2=1.16
r157 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.375 $Y=1.325
+ $X2=4.375 $Y2=1.985
r158 8 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=0.995
+ $X2=4.375 $Y2=1.16
r159 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.375 $Y=0.995
+ $X2=4.375 $Y2=0.56
r160 4 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=1.325
+ $X2=3.955 $Y2=1.16
r161 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.955 $Y=1.325
+ $X2=3.955 $Y2=1.985
r162 1 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=0.995
+ $X2=3.955 $Y2=1.16
r163 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.955 $Y=0.995
+ $X2=3.955 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 42 48 52 54 58
+ 60 64 68 70 72 77 78 80 81 82 88 96 100 105 114 117 120 123 126 130
r145 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r146 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r147 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r148 121 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r149 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r150 118 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r151 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r152 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r153 109 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r154 109 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r155 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r156 106 126 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=8.225 $Y=2.72
+ $X2=8.08 $Y2=2.72
r157 106 108 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.225 $Y=2.72
+ $X2=8.51 $Y2=2.72
r158 105 129 3.67103 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=9.027 $Y2=2.72
r159 105 108 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=8.51 $Y2=2.72
r160 104 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r161 104 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r162 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r163 101 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.385 $Y=2.72
+ $X2=7.22 $Y2=2.72
r164 101 103 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.385 $Y=2.72
+ $X2=7.59 $Y2=2.72
r165 100 126 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.935 $Y=2.72
+ $X2=8.08 $Y2=2.72
r166 100 103 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=2.72
+ $X2=7.59 $Y2=2.72
r167 99 118 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=5.29 $Y2=2.72
r168 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r169 96 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.24 $Y=2.72
+ $X2=5.405 $Y2=2.72
r170 96 98 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=5.24 $Y=2.72
+ $X2=3.45 $Y2=2.72
r171 95 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r172 95 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r173 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r174 92 114 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.365 $Y=2.72
+ $X2=2.11 $Y2=2.72
r175 92 94 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.365 $Y=2.72
+ $X2=2.99 $Y2=2.72
r176 91 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r177 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r178 88 114 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=2.11 $Y2=2.72
r179 88 90 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r180 87 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r181 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r182 84 111 3.66972 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r183 84 86 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 82 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r185 82 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r186 80 94 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.19 $Y=2.72 $X2=2.99
+ $Y2=2.72
r187 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=2.72
+ $X2=3.275 $Y2=2.72
r188 79 98 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.36 $Y=2.72 $X2=3.45
+ $Y2=2.72
r189 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=2.72
+ $X2=3.275 $Y2=2.72
r190 77 86 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r191 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r192 76 90 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r193 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r194 72 75 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=8.96 $Y=1.66
+ $X2=8.96 $Y2=2.34
r195 70 129 3.24416 $w=2.1e-07 $l=1.13666e-07 $layer=LI1_cond $X=8.96 $Y=2.635
+ $X2=9.027 $Y2=2.72
r196 70 75 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=8.96 $Y=2.635
+ $X2=8.96 $Y2=2.34
r197 66 126 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.08 $Y=2.635
+ $X2=8.08 $Y2=2.72
r198 66 68 28.4137 $w=2.88e-07 $l=7.15e-07 $layer=LI1_cond $X=8.08 $Y=2.635
+ $X2=8.08 $Y2=1.92
r199 62 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.635
+ $X2=7.22 $Y2=2.72
r200 62 64 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=7.22 $Y=2.635
+ $X2=7.22 $Y2=2.29
r201 61 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.34 $Y2=2.72
r202 60 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=2.72
+ $X2=7.22 $Y2=2.72
r203 60 61 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.055 $Y=2.72
+ $X2=6.505 $Y2=2.72
r204 56 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.34 $Y=2.635
+ $X2=6.34 $Y2=2.72
r205 56 58 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.34 $Y=2.635
+ $X2=6.34 $Y2=2.29
r206 55 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=2.72
+ $X2=5.405 $Y2=2.72
r207 54 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=2.72
+ $X2=6.34 $Y2=2.72
r208 54 55 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.175 $Y=2.72
+ $X2=5.57 $Y2=2.72
r209 50 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=2.635
+ $X2=5.405 $Y2=2.72
r210 50 52 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=5.405 $Y=2.635
+ $X2=5.405 $Y2=2.29
r211 46 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=2.635
+ $X2=3.275 $Y2=2.72
r212 46 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.275 $Y=2.635
+ $X2=3.275 $Y2=2.27
r213 42 45 15.9477 $w=5.08e-07 $l=6.8e-07 $layer=LI1_cond $X=2.11 $Y=1.66
+ $X2=2.11 $Y2=2.34
r214 40 114 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=2.635
+ $X2=2.11 $Y2=2.72
r215 40 45 6.91849 $w=5.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.11 $Y=2.635
+ $X2=2.11 $Y2=2.34
r216 36 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.1 $Y=1.68 $X2=1.1
+ $Y2=2.36
r217 34 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r218 34 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2.36
r219 30 33 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=1.66
+ $X2=0.24 $Y2=2.34
r220 28 111 3.24547 $w=2.1e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.172 $Y2=2.72
r221 28 33 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.34
r222 9 75 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.805
+ $Y=1.485 $X2=8.94 $Y2=2.34
r223 9 72 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.805
+ $Y=1.485 $X2=8.94 $Y2=1.66
r224 8 68 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=7.965
+ $Y=1.485 $X2=8.1 $Y2=1.92
r225 7 64 600 $w=1.7e-07 $l=8.882e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=1.485 $X2=7.22 $Y2=2.29
r226 6 58 600 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=2.29
r227 5 52 600 $w=1.7e-07 $l=9.12784e-07 $layer=licon1_PDIFF $count=1 $X=5.175
+ $Y=1.485 $X2=5.405 $Y2=2.29
r228 4 48 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.485 $X2=3.275 $Y2=2.27
r229 3 45 200 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=3 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.34
r230 3 42 200 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=3 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.66
r231 2 39 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.36
r232 2 36 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.68
r233 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r234 1 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%SUM 1 2 3 4 13 17 20 25 27 28 30 31 32 33 34 35
+ 36 37 46
c49 34 0 1.29575e-19 $X=0.695 $Y=1.19
c50 28 0 2.02904e-19 $X=1.452 $Y=1.2
r51 37 62 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.68 $Y=2.21 $X2=0.68
+ $Y2=2.33
r52 36 37 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=2.21
r53 36 56 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.68 $Y=1.87
+ $X2=0.68 $Y2=1.65
r54 35 56 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.68 $Y=1.53 $X2=0.68
+ $Y2=1.65
r55 35 52 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.68 $Y=1.53
+ $X2=0.68 $Y2=1.335
r56 34 44 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=0.68 $Y=1.2 $X2=0.68
+ $Y2=1.065
r57 34 52 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=0.68 $Y=1.2 $X2=0.68
+ $Y2=1.335
r58 33 44 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=0.85
+ $X2=0.68 $Y2=1.065
r59 32 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.68 $Y=0.51
+ $X2=0.68 $Y2=0.85
r60 32 46 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.68 $Y=0.51
+ $X2=0.68 $Y2=0.4
r61 30 31 4.88132 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.65
+ $X2=1.52 $Y2=1.565
r62 23 30 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.52 $Y=1.73 $X2=1.52
+ $Y2=1.65
r63 23 25 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=1.52 $Y=1.73 $X2=1.52
+ $Y2=2.33
r64 21 28 6.71073 $w=1.95e-07 $l=1.35e-07 $layer=LI1_cond $X=1.452 $Y=1.335
+ $X2=1.452 $Y2=1.2
r65 21 31 13.0816 $w=1.93e-07 $l=2.3e-07 $layer=LI1_cond $X=1.452 $Y=1.335
+ $X2=1.452 $Y2=1.565
r66 20 28 6.71073 $w=1.95e-07 $l=1.35e-07 $layer=LI1_cond $X=1.452 $Y=1.065
+ $X2=1.452 $Y2=1.2
r67 20 27 13.6503 $w=1.93e-07 $l=2.4e-07 $layer=LI1_cond $X=1.452 $Y=1.065
+ $X2=1.452 $Y2=0.825
r68 15 27 7.67512 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0.66
+ $X2=1.52 $Y2=0.825
r69 15 17 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.52 $Y=0.66
+ $X2=1.52 $Y2=0.4
r70 14 34 2.07418 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.2
+ $X2=0.68 $Y2=1.2
r71 13 28 0.201498 $w=2.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.355 $Y=1.2
+ $X2=1.452 $Y2=1.2
r72 13 14 21.7684 $w=2.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.2
+ $X2=0.845 $Y2=1.2
r73 4 30 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.65
r74 4 25 400 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.33
r75 3 62 400 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.33
r76 3 56 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.65
r77 2 17 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.4
r78 1 46 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%COUT 1 2 3 4 15 19 21 22 23 24 25 26 27 28 29
+ 30
r52 29 30 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=8.545 $Y=1.87
+ $X2=8.545 $Y2=2.21
r53 29 52 6.58539 $w=2.78e-07 $l=1.6e-07 $layer=LI1_cond $X=8.545 $Y=1.87
+ $X2=8.545 $Y2=1.71
r54 28 45 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=1.5 $X2=8.545
+ $Y2=1.415
r55 28 49 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=1.5 $X2=8.545
+ $Y2=1.585
r56 28 52 4.52745 $w=2.78e-07 $l=1.1e-07 $layer=LI1_cond $X=8.545 $Y=1.6
+ $X2=8.545 $Y2=1.71
r57 28 49 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=8.545 $Y=1.6
+ $X2=8.545 $Y2=1.585
r58 27 45 9.2607 $w=2.78e-07 $l=2.25e-07 $layer=LI1_cond $X=8.545 $Y=1.19
+ $X2=8.545 $Y2=1.415
r59 26 39 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=0.82 $X2=8.545
+ $Y2=0.735
r60 26 44 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=0.82 $X2=8.545
+ $Y2=0.905
r61 26 27 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=8.545 $Y=0.92
+ $X2=8.545 $Y2=1.19
r62 26 44 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=8.545 $Y=0.92
+ $X2=8.545 $Y2=0.905
r63 25 39 9.2607 $w=2.78e-07 $l=2.25e-07 $layer=LI1_cond $X=8.545 $Y=0.51
+ $X2=8.545 $Y2=0.735
r64 23 26 3.18746 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.405 $Y=0.82
+ $X2=8.545 $Y2=0.82
r65 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.405 $Y=0.82
+ $X2=7.845 $Y2=0.82
r66 21 28 3.18746 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.405 $Y=1.5
+ $X2=8.545 $Y2=1.5
r67 21 22 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.405 $Y=1.5
+ $X2=7.765 $Y2=1.5
r68 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.68 $Y=1.585
+ $X2=7.765 $Y2=1.5
r69 17 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.68 $Y=1.585
+ $X2=7.68 $Y2=1.71
r70 13 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.72 $Y=0.735
+ $X2=7.845 $Y2=0.82
r71 13 15 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.72 $Y=0.735
+ $X2=7.72 $Y2=0.57
r72 4 52 300 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=2 $X=8.385
+ $Y=1.485 $X2=8.52 $Y2=1.71
r73 3 19 300 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=2 $X=7.545
+ $Y=1.485 $X2=7.68 $Y2=1.71
r74 2 25 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=8.385
+ $Y=0.235 $X2=8.52 $Y2=0.57
r75 1 15 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=7.545
+ $Y=0.235 $X2=7.68 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50 54
+ 56 60 62 64 67 68 70 71 73 74 76 77 78 84 98 102 111 114 117 121
r151 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r152 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r153 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r154 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r155 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r156 106 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r157 106 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r158 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r159 103 117 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.225 $Y=0
+ $X2=8.12 $Y2=0
r160 103 105 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.225 $Y=0
+ $X2=8.51 $Y2=0
r161 102 120 3.67103 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=8.855 $Y=0
+ $X2=9.027 $Y2=0
r162 102 105 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.855 $Y=0
+ $X2=8.51 $Y2=0
r163 101 115 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=7.13 $Y2=0
r164 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r165 98 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=0
+ $X2=7.22 $Y2=0
r166 98 100 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=7.055 $Y=0
+ $X2=5.75 $Y2=0
r167 97 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r168 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r169 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r170 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r171 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r172 91 112 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.07 $Y2=0
r173 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r174 88 111 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.095 $Y=0
+ $X2=1.975 $Y2=0
r175 88 90 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=2.095 $Y=0
+ $X2=3.45 $Y2=0
r176 87 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r177 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r178 84 111 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.975 $Y2=0
r179 84 86 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r180 83 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r181 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r182 80 108 3.66972 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r183 80 82 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r184 78 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r185 78 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r186 76 96 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.29
+ $Y2=0
r187 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.55
+ $Y2=0
r188 75 100 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.715 $Y=0
+ $X2=5.75 $Y2=0
r189 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.55
+ $Y2=0
r190 73 93 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.37
+ $Y2=0
r191 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.585
+ $Y2=0
r192 72 96 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=5.29
+ $Y2=0
r193 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.585
+ $Y2=0
r194 70 90 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.45 $Y2=0
r195 70 71 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.732 $Y2=0
r196 69 93 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r197 69 71 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=3.732
+ $Y2=0
r198 67 82 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r199 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r200 66 86 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r201 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r202 62 120 3.24416 $w=2.1e-07 $l=1.13666e-07 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=9.027 $Y2=0
r203 62 64 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0.38
r204 58 117 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.12 $Y=0.085
+ $X2=8.12 $Y2=0
r205 58 60 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=8.12 $Y=0.085
+ $X2=8.12 $Y2=0.4
r206 57 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.385 $Y=0
+ $X2=7.22 $Y2=0
r207 56 117 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.015 $Y=0
+ $X2=8.12 $Y2=0
r208 56 57 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=8.015 $Y=0
+ $X2=7.385 $Y2=0
r209 52 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=0.085
+ $X2=7.22 $Y2=0
r210 52 54 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.22 $Y=0.085
+ $X2=7.22 $Y2=0.38
r211 48 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0
r212 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0.38
r213 44 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=0.085
+ $X2=4.585 $Y2=0
r214 44 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.585 $Y=0.085
+ $X2=4.585 $Y2=0.38
r215 40 71 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.732 $Y=0.085
+ $X2=3.732 $Y2=0
r216 40 42 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=3.732 $Y=0.085
+ $X2=3.732 $Y2=0.38
r217 36 111 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0
r218 36 38 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0.38
r219 32 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r220 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r221 28 108 3.24547 $w=2.1e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.172 $Y2=0
r222 28 30 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r223 9 64 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=8.805
+ $Y=0.235 $X2=8.94 $Y2=0.38
r224 8 60 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.965
+ $Y=0.235 $X2=8.1 $Y2=0.4
r225 7 54 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=7.045
+ $Y=0.235 $X2=7.22 $Y2=0.38
r226 6 50 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.235 $X2=5.55 $Y2=0.38
r227 5 46 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.235 $X2=4.585 $Y2=0.38
r228 4 42 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.73 $Y2=0.38
r229 3 38 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r230 2 34 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r231 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__HA_4%A_467_47# 1 2 3 4 13 21 22 25 27 29 31
r52 31 32 15.8243 $w=2.39e-07 $l=3.1e-07 $layer=LI1_cond $X=5.055 $Y=0.42
+ $X2=5.055 $Y2=0.73
r53 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=0.73
+ $X2=4.165 $Y2=0.73
r54 27 32 2.73298 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.92 $Y=0.73
+ $X2=5.055 $Y2=0.73
r55 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.92 $Y=0.73
+ $X2=4.25 $Y2=0.73
r56 23 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.645
+ $X2=4.165 $Y2=0.73
r57 23 25 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.165 $Y=0.645
+ $X2=4.165 $Y2=0.51
r58 21 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=0.73
+ $X2=4.165 $Y2=0.73
r59 21 22 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.08 $Y=0.73
+ $X2=3.385 $Y2=0.73
r60 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.3 $Y=0.645
+ $X2=3.385 $Y2=0.73
r61 18 20 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.3 $Y=0.645
+ $X2=3.3 $Y2=0.51
r62 17 20 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.3 $Y=0.475 $X2=3.3
+ $Y2=0.51
r63 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.215 $Y=0.39
+ $X2=3.3 $Y2=0.475
r64 13 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.215 $Y=0.39
+ $X2=2.46 $Y2=0.39
r65 4 31 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.98
+ $Y=0.235 $X2=5.105 $Y2=0.42
r66 3 25 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.235 $X2=4.165 $Y2=0.51
r67 2 20 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.51
r68 1 15 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.39
.ends


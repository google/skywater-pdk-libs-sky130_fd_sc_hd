* File: sky130_fd_sc_hd__o21ai_1.pex.spice
* Created: Thu Aug 27 14:35:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21AI_1%A1 3 6 8 11 12 13
r25 11 14 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.16
+ $X2=0.367 $Y2=1.325
r26 11 13 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.367 $Y=1.16
+ $X2=0.367 $Y2=0.995
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.325
+ $Y=1.16 $X2=0.325 $Y2=1.16
r28 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.235 $Y=1.16 $X2=0.325
+ $Y2=1.16
r29 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r30 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_1%A2 3 7 8 9 10 11 17 18 19
r42 21 29 3.83364 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.687 $Y=1.325
+ $X2=0.687 $Y2=1.16
r43 17 20 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.16
+ $X2=0.895 $Y2=1.325
r44 17 19 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.16
+ $X2=0.895 $Y2=0.995
r45 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r46 10 11 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=0.687 $Y=1.87
+ $X2=0.687 $Y2=2.21
r47 9 10 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=0.687 $Y=1.53
+ $X2=0.687 $Y2=1.87
r48 9 21 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=0.687 $Y=1.53
+ $X2=0.687 $Y2=1.325
r49 8 18 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.89 $Y2=1.16
r50 8 29 0.27938 $w=3.28e-07 $l=8e-09 $layer=LI1_cond $X=0.695 $Y=1.16 $X2=0.687
+ $Y2=1.16
r51 7 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.95 $Y=0.56 $X2=0.95
+ $Y2=0.995
r52 3 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.83 $Y=1.985
+ $X2=0.83 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_1%B1 3 7 9 14
r31 11 14 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.37 $Y=1.46 $X2=1.6
+ $Y2=1.46
r32 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6 $Y=1.46
+ $X2=1.6 $Y2=1.46
r33 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.625
+ $X2=1.37 $Y2=1.46
r34 5 7 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.37 $Y=1.625 $X2=1.37
+ $Y2=2.135
r35 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.295
+ $X2=1.37 $Y2=1.46
r36 1 3 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.37 $Y=1.295
+ $X2=1.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_1%VPWR 1 2 7 9 13 15 17 19 29
r27 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r28 23 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r29 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 20 25 4.70099 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=2.72
+ $X2=0.205 $Y2=2.72
r31 20 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r32 19 28 4.08769 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.495 $Y=2.72
+ $X2=1.667 $Y2=2.72
r33 19 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.495 $Y=2.72
+ $X2=1.15 $Y2=2.72
r34 17 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r36 13 28 3.08953 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.622 $Y=2.635
+ $X2=1.667 $Y2=2.72
r37 13 15 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=1.622 $Y=2.635
+ $X2=1.622 $Y2=2
r38 9 12 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=0.25 $Y=1.66 $X2=0.25
+ $Y2=2.34
r39 7 25 2.98112 $w=3.2e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.25 $Y=2.635
+ $X2=0.205 $Y2=2.72
r40 7 12 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.25 $Y=2.635
+ $X2=0.25 $Y2=2.34
r41 2 15 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.785 $X2=1.58 $Y2=2
r42 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r43 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_1%Y 1 2 9 10 13 15 16 28
r34 16 24 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.13 $Y=2.21
+ $X2=1.13 $Y2=2
r35 15 28 10.3022 $w=4.98e-07 $l=2.8e-07 $layer=LI1_cond $X=1.14 $Y=1.785
+ $X2=1.14 $Y2=1.505
r36 15 24 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.13 $Y=1.87
+ $X2=1.13 $Y2=2
r37 11 13 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.58 $Y=0.955 $X2=1.58
+ $Y2=0.555
r38 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=1.04
+ $X2=1.58 $Y2=0.955
r39 9 10 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.495 $Y=1.04
+ $X2=1.315 $Y2=1.04
r40 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=1.125
+ $X2=1.315 $Y2=1.04
r41 7 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.23 $Y=1.125
+ $X2=1.23 $Y2=1.505
r42 2 24 300 $w=1.7e-07 $l=6.17333e-07 $layer=licon1_PDIFF $count=2 $X=0.905
+ $Y=1.485 $X2=1.13 $Y2=2
r43 1 13 182 $w=1.7e-07 $l=3.81576e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_1%A_27_47# 1 2 9 11 12 15
r23 13 15 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.19 $Y=0.615
+ $X2=1.19 $Y2=0.475
r24 11 13 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.075 $Y=0.7
+ $X2=1.19 $Y2=0.615
r25 11 12 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.075 $Y=0.7
+ $X2=0.38 $Y2=0.7
r26 7 12 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.235 $Y=0.615
+ $X2=0.38 $Y2=0.7
r27 7 9 7.35179 $w=2.88e-07 $l=1.85e-07 $layer=LI1_cond $X=0.235 $Y=0.615
+ $X2=0.235 $Y2=0.43
r28 2 15 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=1.025 $Y=0.235
+ $X2=1.16 $Y2=0.475
r29 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_1%VGND 1 6 8 10 17 18 21
r28 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r29 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r30 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r31 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r32 15 17 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.61
+ $Y2=0
r33 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r34 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.23
+ $Y2=0
r35 8 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r36 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r37 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r38 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.36
r39 1 6 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.74 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__o32a_4.pex.spice
* Created: Thu Aug 27 14:41:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O32A_4%A1 5 9 13 17 19 20 24 27
c41 20 0 1.52846e-19 $X=0.695 $Y=1.19
r42 26 27 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.89
+ $Y2=1.16
r43 24 26 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=0.465 $Y=1.16 $X2=0.47
+ $Y2=1.16
r44 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.465
+ $Y=1.16 $X2=0.465 $Y2=1.16
r45 20 25 12.7545 $w=1.98e-07 $l=2.3e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.465 $Y2=1.175
r46 19 25 12.7545 $w=1.98e-07 $l=2.3e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.465 $Y2=1.175
r47 15 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.16
r48 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r49 11 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=1.16
r50 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r51 7 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r52 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295 $X2=0.47
+ $Y2=1.985
r53 3 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r54 3 5 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%A2 3 7 11 15 17 18 26
c41 26 0 1.52846e-19 $X=1.73 $Y=1.16
c42 18 0 1.89941e-19 $X=1.615 $Y=1.19
c43 15 0 1.63215e-19 $X=1.73 $Y=1.985
r44 24 26 43.3239 $w=2.7e-07 $l=1.95e-07 $layer=POLY_cond $X=1.535 $Y=1.16
+ $X2=1.73 $Y2=1.16
r45 21 24 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.535 $Y2=1.16
r46 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.535
+ $Y=1.16 $X2=1.535 $Y2=1.16
r47 17 18 21.0727 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.535 $Y2=1.175
r48 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.16
r49 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r50 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=1.16
r51 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r52 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.16
r53 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295 $X2=1.31
+ $Y2=1.985
r54 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=1.16
r55 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%A3 3 7 11 15 17 23 26
c45 26 0 1.89941e-19 $X=3.09 $Y=1.16
r46 25 26 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.67 $Y=1.16 $X2=3.09
+ $Y2=1.16
r47 24 25 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=2.59 $Y=1.16 $X2=2.67
+ $Y2=1.16
r48 22 24 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.59 $Y2=1.16
r49 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r50 19 22 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.17 $Y=1.16 $X2=2.26
+ $Y2=1.16
r51 17 23 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=1.175
+ $X2=2.26 $Y2=1.175
r52 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.16
r53 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.985
r54 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.16
r55 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.985
r56 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.59 $Y=1.025
+ $X2=2.59 $Y2=1.16
r57 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.59 $Y=1.025
+ $X2=2.59 $Y2=0.56
r58 1 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.17 $Y=1.025
+ $X2=2.17 $Y2=1.16
r59 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.17 $Y=1.025
+ $X2=2.17 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%B1 3 7 11 15 17 23 24
r57 22 24 85.5369 $w=2.7e-07 $l=3.85e-07 $layer=POLY_cond $X=4.065 $Y=1.16
+ $X2=4.45 $Y2=1.16
r58 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.065
+ $Y=1.16 $X2=4.065 $Y2=1.16
r59 19 22 7.77608 $w=2.7e-07 $l=3.5e-08 $layer=POLY_cond $X=4.03 $Y=1.16
+ $X2=4.065 $Y2=1.16
r60 17 23 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=3.955 $Y=1.175 $X2=4.065
+ $Y2=1.175
r61 13 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.45 $Y=1.295
+ $X2=4.45 $Y2=1.16
r62 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.45 $Y=1.295
+ $X2=4.45 $Y2=1.985
r63 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.45 $Y=1.025
+ $X2=4.45 $Y2=1.16
r64 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.45 $Y=1.025
+ $X2=4.45 $Y2=0.56
r65 5 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.03 $Y=1.295
+ $X2=4.03 $Y2=1.16
r66 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.03 $Y=1.295 $X2=4.03
+ $Y2=1.985
r67 1 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.03 $Y=1.025
+ $X2=4.03 $Y2=1.16
r68 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.03 $Y=1.025
+ $X2=4.03 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%B2 3 7 11 15 18 19 20 21 25
c51 25 0 1.77246e-19 $X=5.095 $Y=1.16
r52 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.095
+ $Y=1.16 $X2=5.095 $Y2=1.16
r53 21 25 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=4.875 $Y=1.175
+ $X2=5.095 $Y2=1.175
r54 19 24 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=5.245 $Y=1.16
+ $X2=5.095 $Y2=1.16
r55 19 20 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.245 $Y=1.16
+ $X2=5.32 $Y2=1.16
r56 17 24 33.3261 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=4.945 $Y=1.16
+ $X2=5.095 $Y2=1.16
r57 17 18 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.945 $Y=1.16
+ $X2=4.87 $Y2=1.16
r58 13 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.32 $Y=1.295
+ $X2=5.32 $Y2=1.16
r59 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.32 $Y=1.295
+ $X2=5.32 $Y2=1.985
r60 9 20 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.32 $Y=1.025
+ $X2=5.32 $Y2=1.16
r61 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.32 $Y=1.025
+ $X2=5.32 $Y2=0.56
r62 5 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.87 $Y=1.295
+ $X2=4.87 $Y2=1.16
r63 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.87 $Y=1.295 $X2=4.87
+ $Y2=1.985
r64 1 18 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.87 $Y=1.025
+ $X2=4.87 $Y2=1.16
r65 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.87 $Y=1.025
+ $X2=4.87 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%A_549_297# 1 2 3 4 5 18 22 26 30 34 38 42 46
+ 50 52 53 55 56 57 61 62 66 67 70 72 73 74 75 78 81 88 95
c174 88 0 1.77246e-19 $X=6.185 $Y=1.16
c175 50 0 1.81415e-19 $X=2.88 $Y=1.865
r176 92 93 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.68 $Y=1.16 $X2=7.1
+ $Y2=1.16
r177 91 92 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.26 $Y=1.16
+ $X2=6.68 $Y2=1.16
r178 88 91 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.185 $Y=1.16
+ $X2=6.26 $Y2=1.16
r179 86 88 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=6.055 $Y=1.16
+ $X2=6.185 $Y2=1.16
r180 85 87 4.81805 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=6.055 $Y=1.17
+ $X2=6.135 $Y2=1.17
r181 85 86 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.055
+ $Y=1.16 $X2=6.055 $Y2=1.16
r182 79 95 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=7.31 $Y=1.16
+ $X2=7.52 $Y2=1.16
r183 79 93 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=7.31 $Y=1.16
+ $X2=7.1 $Y2=1.16
r184 78 87 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=7.31 $Y=1.16
+ $X2=6.135 $Y2=1.16
r185 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.31
+ $Y=1.16 $X2=7.31 $Y2=1.16
r186 74 85 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=6.04 $Y=1.17
+ $X2=6.055 $Y2=1.17
r187 74 75 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=6.04 $Y=1.17
+ $X2=5.775 $Y2=1.17
r188 73 75 7.00737 $w=1.9e-07 $l=1.6895e-07 $layer=LI1_cond $X=5.647 $Y=1.075
+ $X2=5.775 $Y2=1.17
r189 72 83 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.647 $Y=0.805
+ $X2=5.647 $Y2=0.72
r190 72 73 12.2023 $w=2.53e-07 $l=2.7e-07 $layer=LI1_cond $X=5.647 $Y=0.805
+ $X2=5.647 $Y2=1.075
r191 68 70 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.11 $Y=1.615
+ $X2=5.11 $Y2=1.95
r192 66 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.025 $Y=1.53
+ $X2=5.11 $Y2=1.615
r193 66 67 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.025 $Y=1.53
+ $X2=4.62 $Y2=1.53
r194 63 81 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.62 $Y=0.72
+ $X2=4.51 $Y2=0.72
r195 63 65 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=4.62 $Y=0.72 $X2=4.66
+ $Y2=0.72
r196 62 83 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=5.52 $Y=0.72
+ $X2=5.647 $Y2=0.72
r197 62 65 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.52 $Y=0.72
+ $X2=4.66 $Y2=0.72
r198 61 67 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.51 $Y=1.445
+ $X2=4.62 $Y2=1.53
r199 60 81 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=0.805
+ $X2=4.51 $Y2=0.72
r200 60 61 33.5256 $w=2.18e-07 $l=6.4e-07 $layer=LI1_cond $X=4.51 $Y=0.805
+ $X2=4.51 $Y2=1.445
r201 57 59 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.645 $Y=0.72
+ $X2=3.82 $Y2=0.72
r202 56 81 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.4 $Y=0.72 $X2=4.51
+ $Y2=0.72
r203 56 59 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.4 $Y=0.72
+ $X2=3.82 $Y2=0.72
r204 54 57 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.55 $Y=0.805
+ $X2=3.645 $Y2=0.72
r205 54 55 17.512 $w=1.88e-07 $l=3e-07 $layer=LI1_cond $X=3.55 $Y=0.805 $X2=3.55
+ $Y2=1.105
r206 52 55 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.455 $Y=1.19
+ $X2=3.55 $Y2=1.105
r207 52 53 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.455 $Y=1.19
+ $X2=2.965 $Y2=1.19
r208 48 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.88 $Y=1.275
+ $X2=2.965 $Y2=1.19
r209 48 50 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.88 $Y=1.275
+ $X2=2.88 $Y2=1.865
r210 44 95 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.52 $Y=1.295
+ $X2=7.52 $Y2=1.16
r211 44 46 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.52 $Y=1.295
+ $X2=7.52 $Y2=1.985
r212 40 95 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.52 $Y=1.025
+ $X2=7.52 $Y2=1.16
r213 40 42 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.52 $Y=1.025
+ $X2=7.52 $Y2=0.56
r214 36 93 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.1 $Y=1.295
+ $X2=7.1 $Y2=1.16
r215 36 38 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.1 $Y=1.295
+ $X2=7.1 $Y2=1.985
r216 32 93 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.1 $Y=1.025
+ $X2=7.1 $Y2=1.16
r217 32 34 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.1 $Y=1.025
+ $X2=7.1 $Y2=0.56
r218 28 92 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.68 $Y=1.295
+ $X2=6.68 $Y2=1.16
r219 28 30 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.68 $Y=1.295
+ $X2=6.68 $Y2=1.985
r220 24 92 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.68 $Y=1.025
+ $X2=6.68 $Y2=1.16
r221 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.68 $Y=1.025
+ $X2=6.68 $Y2=0.56
r222 20 91 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.26 $Y=1.295
+ $X2=6.26 $Y2=1.16
r223 20 22 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.26 $Y=1.295
+ $X2=6.26 $Y2=1.985
r224 16 91 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.26 $Y=1.025
+ $X2=6.26 $Y2=1.16
r225 16 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.26 $Y=1.025
+ $X2=6.26 $Y2=0.56
r226 5 70 600 $w=1.7e-07 $l=5.41249e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.485 $X2=5.11 $Y2=1.95
r227 4 50 600 $w=1.7e-07 $l=4.4238e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.865
r228 3 83 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.53 $Y2=0.72
r229 2 65 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.235 $X2=4.66 $Y2=0.72
r230 1 59 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.235 $X2=3.82 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%A_27_297# 1 2 3 10 12 14 16 17 18 22
c48 16 0 1.63215e-19 $X=1.1 $Y=1.665
r49 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=1.94 $Y2=2
r50 19 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.38
+ $X2=1.1 $Y2=2.38
r51 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.775 $Y=2.38
+ $X2=1.94 $Y2=2.295
r52 18 19 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=2.38
+ $X2=1.265 $Y2=2.38
r53 17 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.295 $X2=1.1
+ $Y2=2.38
r54 16 27 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.1 $Y=1.665 $X2=1.1
+ $Y2=1.555
r55 16 17 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=1.1 $Y=1.665 $X2=1.1
+ $Y2=2.295
r56 15 25 4.39066 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=0.425 $Y=1.555
+ $X2=0.255 $Y2=1.555
r57 14 27 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.555
+ $X2=1.1 $Y2=1.555
r58 14 15 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=0.935 $Y=1.555
+ $X2=0.425 $Y2=1.555
r59 10 25 2.84101 $w=3.4e-07 $l=1.1e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.555
r60 10 12 22.8794 $w=3.38e-07 $l=6.75e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.34
r61 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r62 2 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r63 2 27 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.66
r64 1 25 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r65 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 46 47 48 50 72 73 76
r106 76 77 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r107 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r108 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r109 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r110 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r111 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r112 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r113 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r114 61 64 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 60 63 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=5.75 $Y2=2.72
r116 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r117 58 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r118 58 77 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 57 58 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r120 55 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.68 $Y2=2.72
r121 55 57 205.182 $w=1.68e-07 $l=3.145e-06 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=3.91 $Y2=2.72
r122 50 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.68 $Y2=2.72
r123 50 52 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 48 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 48 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 46 69 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.645 $Y=2.72
+ $X2=7.59 $Y2=2.72
r127 46 47 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.645 $Y=2.72
+ $X2=7.772 $Y2=2.72
r128 45 72 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.9 $Y=2.72 $X2=8.05
+ $Y2=2.72
r129 45 47 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.9 $Y=2.72
+ $X2=7.772 $Y2=2.72
r130 43 66 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=6.67 $Y2=2.72
r131 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=6.89 $Y2=2.72
r132 42 69 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.975 $Y=2.72
+ $X2=7.59 $Y2=2.72
r133 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=2.72
+ $X2=6.89 $Y2=2.72
r134 40 63 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.965 $Y=2.72
+ $X2=5.75 $Y2=2.72
r135 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=2.72
+ $X2=6.05 $Y2=2.72
r136 39 66 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.135 $Y=2.72
+ $X2=6.67 $Y2=2.72
r137 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.135 $Y=2.72
+ $X2=6.05 $Y2=2.72
r138 37 57 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=3.91 $Y2=2.72
r139 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.24 $Y2=2.72
r140 36 60 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.325 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.325 $Y=2.72
+ $X2=4.24 $Y2=2.72
r142 32 47 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.772 $Y=2.635
+ $X2=7.772 $Y2=2.72
r143 32 34 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=7.772 $Y=2.635
+ $X2=7.772 $Y2=2
r144 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=2.635
+ $X2=6.89 $Y2=2.72
r145 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.89 $Y=2.635
+ $X2=6.89 $Y2=2
r146 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.05 $Y=2.635
+ $X2=6.05 $Y2=2.72
r147 24 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.05 $Y=2.635
+ $X2=6.05 $Y2=2
r148 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=2.635
+ $X2=4.24 $Y2=2.72
r149 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.24 $Y=2.635
+ $X2=4.24 $Y2=2.29
r150 16 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r151 16 18 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2
r152 5 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=7.595
+ $Y=1.485 $X2=7.73 $Y2=2
r153 4 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.755
+ $Y=1.485 $X2=6.89 $Y2=2
r154 3 26 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=5.925
+ $Y=1.485 $X2=6.05 $Y2=2
r155 2 22 600 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.485 $X2=4.24 $Y2=2.29
r156 1 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%A_277_297# 1 2 3 12 14 15 16 17 18 20 22
r52 20 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.295 $X2=3.3
+ $Y2=2.38
r53 20 22 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.3 $Y=2.295
+ $X2=3.3 $Y2=1.66
r54 19 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=2.38
+ $X2=2.46 $Y2=2.38
r55 18 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=2.38
+ $X2=3.3 $Y2=2.38
r56 18 19 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.135 $Y=2.38
+ $X2=2.625 $Y2=2.38
r57 17 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.295 $X2=2.46
+ $Y2=2.38
r58 16 25 2.99472 $w=3.3e-07 $l=1.23e-07 $layer=LI1_cond $X=2.46 $Y=1.69
+ $X2=2.46 $Y2=1.567
r59 16 17 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=2.46 $Y=1.69
+ $X2=2.46 $Y2=2.295
r60 14 25 4.01731 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=1.567
+ $X2=2.46 $Y2=1.567
r61 14 15 32.4566 $w=2.43e-07 $l=6.9e-07 $layer=LI1_cond $X=2.295 $Y=1.567
+ $X2=1.605 $Y2=1.567
r62 10 15 7.11011 $w=2.45e-07 $l=1.5995e-07 $layer=LI1_cond $X=1.52 $Y=1.69
+ $X2=1.605 $Y2=1.567
r63 10 12 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.52 $Y=1.69
+ $X2=1.52 $Y2=1.865
r64 3 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=2.34
r65 3 22 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=1.66
r66 2 27 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=2.34
r67 2 25 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=1.66
r68 1 12 600 $w=1.7e-07 $l=4.4238e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.865
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%A_739_297# 1 2 3 12 16 18 23 24 25 26 28 30
r66 26 32 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.53 $Y=2.285 $X2=5.53
+ $Y2=2.375
r67 26 28 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=5.53 $Y=2.285
+ $X2=5.53 $Y2=1.66
r68 24 32 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=2.375
+ $X2=5.53 $Y2=2.375
r69 24 25 33.2727 $w=1.78e-07 $l=5.4e-07 $layer=LI1_cond $X=5.365 $Y=2.375
+ $X2=4.825 $Y2=2.375
r70 21 25 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.66 $Y=2.285
+ $X2=4.825 $Y2=2.375
r71 21 23 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.66 $Y=2.285
+ $X2=4.66 $Y2=2
r72 20 23 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.66 $Y=1.955
+ $X2=4.66 $Y2=2
r73 19 30 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=1.87
+ $X2=3.82 $Y2=1.87
r74 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.495 $Y=1.87
+ $X2=4.66 $Y2=1.955
r75 18 19 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.495 $Y=1.87
+ $X2=3.985 $Y2=1.87
r76 14 30 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=1.955
+ $X2=3.82 $Y2=1.87
r77 14 16 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.82 $Y=1.955
+ $X2=3.82 $Y2=2.34
r78 10 30 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=1.785
+ $X2=3.82 $Y2=1.87
r79 10 12 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.82 $Y=1.785
+ $X2=3.82 $Y2=1.66
r80 3 32 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.485 $X2=5.53 $Y2=2.34
r81 3 28 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.485 $X2=5.53 $Y2=1.66
r82 2 23 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.525
+ $Y=1.485 $X2=4.66 $Y2=2
r83 1 16 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.695
+ $Y=1.485 $X2=3.82 $Y2=2.34
r84 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=3.695
+ $Y=1.485 $X2=3.82 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%X 1 2 3 4 15 17 19 21 22 23 27 31 35 36 37
r69 44 55 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.89 $Y=1.58
+ $X2=7.31 $Y2=1.58
r70 37 44 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=8.05 $Y=1.58
+ $X2=7.89 $Y2=1.58
r71 37 44 0.610244 $w=4.88e-07 $l=2.5e-08 $layer=LI1_cond $X=7.89 $Y=1.47
+ $X2=7.89 $Y2=1.495
r72 36 37 6.83473 $w=4.88e-07 $l=2.8e-07 $layer=LI1_cond $X=7.89 $Y=1.19
+ $X2=7.89 $Y2=1.47
r73 35 43 9.33971 $w=1.88e-07 $l=1.6e-07 $layer=LI1_cond $X=8.05 $Y=0.81
+ $X2=7.89 $Y2=0.81
r74 35 36 6.59064 $w=4.88e-07 $l=2.7e-07 $layer=LI1_cond $X=7.89 $Y=0.92
+ $X2=7.89 $Y2=1.19
r75 35 43 0.366146 $w=4.88e-07 $l=1.5e-08 $layer=LI1_cond $X=7.89 $Y=0.92
+ $X2=7.89 $Y2=0.905
r76 31 55 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.31 $Y=2.34
+ $X2=7.31 $Y2=1.665
r77 25 43 33.8565 $w=1.88e-07 $l=5.8e-07 $layer=LI1_cond $X=7.31 $Y=0.81
+ $X2=7.89 $Y2=0.81
r78 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.31 $Y=0.715
+ $X2=7.31 $Y2=0.38
r79 24 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.635 $Y=1.58
+ $X2=6.47 $Y2=1.58
r80 23 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=1.58
+ $X2=7.31 $Y2=1.58
r81 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.145 $Y=1.58
+ $X2=6.635 $Y2=1.58
r82 21 25 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=0.81
+ $X2=7.31 $Y2=0.81
r83 21 22 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=7.145 $Y=0.81
+ $X2=6.635 $Y2=0.81
r84 17 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=1.665 $X2=6.47
+ $Y2=1.58
r85 17 19 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.47 $Y=1.665
+ $X2=6.47 $Y2=2.34
r86 13 22 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=6.47 $Y=0.715
+ $X2=6.635 $Y2=0.81
r87 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.47 $Y=0.715
+ $X2=6.47 $Y2=0.38
r88 4 55 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.175
+ $Y=1.485 $X2=7.31 $Y2=1.66
r89 4 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.175
+ $Y=1.485 $X2=7.31 $Y2=2.34
r90 3 34 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.335
+ $Y=1.485 $X2=6.47 $Y2=1.66
r91 3 19 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.335
+ $Y=1.485 $X2=6.47 $Y2=2.34
r92 2 27 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.175
+ $Y=0.235 $X2=7.31 $Y2=0.38
r93 1 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.335
+ $Y=0.235 $X2=6.47 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%A_27_47# 1 2 3 4 5 6 21 23 24 32 33 37
r64 35 37 45.9481 $w=2.08e-07 $l=8.7e-07 $layer=LI1_cond $X=4.24 $Y=0.36
+ $X2=5.11 $Y2=0.36
r65 33 35 67.3377 $w=2.08e-07 $l=1.275e-06 $layer=LI1_cond $X=2.965 $Y=0.36
+ $X2=4.24 $Y2=0.36
r66 30 32 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.84 $Y=0.635
+ $X2=2.84 $Y2=0.505
r67 29 33 6.88375 $w=2.1e-07 $l=1.69558e-07 $layer=LI1_cond $X=2.84 $Y=0.465
+ $X2=2.965 $Y2=0.36
r68 29 32 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=2.84 $Y=0.465 $X2=2.84
+ $Y2=0.505
r69 26 28 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=1.1 $Y=0.76 $X2=1.96
+ $Y2=0.76
r70 24 26 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=0.345 $Y=0.76
+ $X2=1.1 $Y2=0.76
r71 23 30 6.81649 $w=2.5e-07 $l=1.76777e-07 $layer=LI1_cond $X=2.715 $Y=0.76
+ $X2=2.84 $Y2=0.635
r72 23 28 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=2.715 $Y=0.76
+ $X2=1.96 $Y2=0.76
r73 19 24 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.76
r74 19 21 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.505
r75 6 37 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.945
+ $Y=0.235 $X2=5.11 $Y2=0.38
r76 5 35 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.105
+ $Y=0.235 $X2=4.24 $Y2=0.38
r77 4 32 182 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.505
r78 3 28 182 $w=1.7e-07 $l=5.57136e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.96 $Y2=0.72
r79 2 26 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.72
r80 1 21 182 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_4%VGND 1 2 3 4 5 6 21 25 29 32 33 35 36 38 39
+ 40 47 48 68 69 73 82
r91 80 82 6.56995 $w=5.48e-07 $l=1.5e-08 $layer=LI1_cond $X=2.53 $Y=0.19
+ $X2=2.545 $Y2=0.19
r92 80 81 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r93 78 80 3.26203 $w=5.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.38 $Y=0.19
+ $X2=2.53 $Y2=0.19
r94 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r95 72 75 0.217469 $w=5.48e-07 $l=1e-08 $layer=LI1_cond $X=0.68 $Y=0.19 $X2=0.69
+ $Y2=0.19
r96 72 73 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.19
+ $X2=0.515 $Y2=0.19
r97 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r98 66 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r99 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r100 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r101 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r102 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r103 60 81 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=2.53 $Y2=0
r104 59 82 209.096 $w=1.68e-07 $l=3.205e-06 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=2.545 $Y2=0
r105 59 60 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r106 56 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r107 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r108 53 55 11.9608 $w=5.48e-07 $l=5.5e-07 $layer=LI1_cond $X=1.52 $Y=0.19
+ $X2=2.07 $Y2=0.19
r109 51 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r110 51 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r111 50 53 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.19
+ $X2=1.52 $Y2=0.19
r112 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r113 48 75 8.15508 $w=5.48e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0.19
+ $X2=0.69 $Y2=0.19
r114 48 50 1.84848 $w=5.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=0.19
+ $X2=1.15 $Y2=0.19
r115 47 78 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=2.27 $Y=0.19
+ $X2=2.38 $Y2=0.19
r116 47 55 4.34938 $w=5.48e-07 $l=2e-07 $layer=LI1_cond $X=2.27 $Y=0.19 $X2=2.07
+ $Y2=0.19
r117 44 73 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r118 40 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 40 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 38 65 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.645 $Y=0 $X2=7.59
+ $Y2=0
r121 38 39 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.645 $Y=0
+ $X2=7.772 $Y2=0
r122 37 68 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.9 $Y=0 $X2=8.05
+ $Y2=0
r123 37 39 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.9 $Y=0 $X2=7.772
+ $Y2=0
r124 35 62 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.805 $Y=0
+ $X2=6.67 $Y2=0
r125 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=0 $X2=6.89
+ $Y2=0
r126 34 65 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.975 $Y=0 $X2=7.59
+ $Y2=0
r127 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=0 $X2=6.89
+ $Y2=0
r128 32 59 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=5.75 $Y2=0
r129 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=0 $X2=6.05
+ $Y2=0
r130 31 62 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.135 $Y=0
+ $X2=6.67 $Y2=0
r131 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.135 $Y=0 $X2=6.05
+ $Y2=0
r132 27 39 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.772 $Y=0.085
+ $X2=7.772 $Y2=0
r133 27 29 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=7.772 $Y=0.085
+ $X2=7.772 $Y2=0.38
r134 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=0.085
+ $X2=6.89 $Y2=0
r135 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.89 $Y=0.085
+ $X2=6.89 $Y2=0.38
r136 19 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.05 $Y=0.085
+ $X2=6.05 $Y2=0
r137 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.05 $Y=0.085
+ $X2=6.05 $Y2=0.38
r138 6 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.595
+ $Y=0.235 $X2=7.73 $Y2=0.38
r139 5 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.755
+ $Y=0.235 $X2=6.89 $Y2=0.38
r140 4 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.925
+ $Y=0.235 $X2=6.05 $Y2=0.38
r141 3 78 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.38
r142 2 53 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r143 1 72 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


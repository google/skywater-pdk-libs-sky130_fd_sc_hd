* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
M1000 VPWR A a_573_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.05225e+11p pd=5.16e+06u as=2.7e+11p ps=2.54e+06u
M1001 a_573_297# B a_477_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1002 VGND C_N a_27_410# VNB nshort w=420000u l=150000u
+  ad=6.743e+11p pd=7.02e+06u as=1.092e+11p ps=1.36e+06u
M1003 Y a_205_93# VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=0p ps=0u
M1004 a_477_297# a_27_410# a_393_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 VGND a_27_410# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_393_297# a_205_93# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.559e+11p ps=2.52e+06u
M1008 a_205_93# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1009 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C_N a_27_410# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 a_205_93# D_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.085e+11p pd=1.36e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__a311oi_1.spice.SKY130_FD_SC_HD__A311OI_1.pxi
* Created: Thu Aug 27 14:04:14 2020
* 
x_PM_SKY130_FD_SC_HD__A311OI_1%A3 N_A3_M1009_g N_A3_M1006_g A3 N_A3_c_53_n
+ N_A3_c_54_n N_A3_c_57_n PM_SKY130_FD_SC_HD__A311OI_1%A3
x_PM_SKY130_FD_SC_HD__A311OI_1%A2 N_A2_M1002_g N_A2_M1000_g A2 A2 A2 N_A2_c_78_n
+ N_A2_c_79_n N_A2_c_80_n PM_SKY130_FD_SC_HD__A311OI_1%A2
x_PM_SKY130_FD_SC_HD__A311OI_1%A1 N_A1_M1005_g N_A1_M1008_g N_A1_c_117_n
+ N_A1_c_118_n N_A1_c_119_n A1 N_A1_c_120_n N_A1_c_132_n
+ PM_SKY130_FD_SC_HD__A311OI_1%A1
x_PM_SKY130_FD_SC_HD__A311OI_1%B1 N_B1_M1004_g N_B1_M1001_g N_B1_c_159_n
+ N_B1_c_160_n N_B1_c_175_p B1 N_B1_c_161_n PM_SKY130_FD_SC_HD__A311OI_1%B1
x_PM_SKY130_FD_SC_HD__A311OI_1%C1 N_C1_M1007_g N_C1_c_203_n N_C1_M1003_g C1
+ N_C1_c_205_n PM_SKY130_FD_SC_HD__A311OI_1%C1
x_PM_SKY130_FD_SC_HD__A311OI_1%VPWR N_VPWR_M1006_s N_VPWR_M1000_d N_VPWR_c_232_n
+ N_VPWR_c_233_n N_VPWR_c_234_n VPWR N_VPWR_c_235_n N_VPWR_c_236_n
+ N_VPWR_c_231_n N_VPWR_c_238_n PM_SKY130_FD_SC_HD__A311OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A311OI_1%A_109_297# N_A_109_297#_M1006_d
+ N_A_109_297#_M1008_d N_A_109_297#_c_287_n N_A_109_297#_c_272_n
+ N_A_109_297#_c_274_n N_A_109_297#_c_276_n N_A_109_297#_c_281_n
+ PM_SKY130_FD_SC_HD__A311OI_1%A_109_297#
x_PM_SKY130_FD_SC_HD__A311OI_1%Y N_Y_M1005_d N_Y_M1003_d N_Y_M1007_d N_Y_c_302_n
+ N_Y_c_306_n N_Y_c_304_n N_Y_c_298_n N_Y_c_319_n N_Y_c_300_n Y Y Y N_Y_c_301_n
+ PM_SKY130_FD_SC_HD__A311OI_1%Y
x_PM_SKY130_FD_SC_HD__A311OI_1%VGND N_VGND_M1009_s N_VGND_M1001_d N_VGND_c_344_n
+ N_VGND_c_345_n N_VGND_c_346_n VGND N_VGND_c_347_n N_VGND_c_348_n
+ N_VGND_c_349_n N_VGND_c_350_n PM_SKY130_FD_SC_HD__A311OI_1%VGND
cc_1 VNB A3 0.015257f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_2 VNB N_A3_c_53_n 0.0367666f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_3 VNB N_A3_c_54_n 0.0209915f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=0.995
cc_4 VNB A2 0.00222805f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_5 VNB N_A2_c_78_n 0.0191065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A2_c_79_n 0.00419979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A2_c_80_n 0.0165744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_c_117_n 0.00101987f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_9 VNB N_A1_c_118_n 0.00197434f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.41
cc_10 VNB N_A1_c_119_n 0.0229329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_120_n 0.0166833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_159_n 0.00280001f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_13 VNB N_B1_c_160_n 0.0206793f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_14 VNB N_B1_c_161_n 0.0178452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_C1_c_203_n 0.0222526f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_16 VNB C1 0.0142618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_C1_c_205_n 0.0349829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_231_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_298_n 0.00289819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_344_n 0.0103361f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_21 VNB N_VGND_c_345_n 0.0250316f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_22 VNB N_VGND_c_346_n 0.00561423f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.41
cc_23 VNB N_VGND_c_347_n 0.038076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_348_n 0.0306352f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_349_n 0.199386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_350_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB A3 0.00101659f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_28 VPB N_A3_c_53_n 0.0188217f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_29 VPB N_A3_c_57_n 0.0185091f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.41
cc_30 VPB N_A2_M1000_g 0.0190678f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_31 VPB N_A2_c_78_n 0.0040131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A2_c_79_n 0.00188913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A1_M1008_g 0.0199041f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_34 VPB N_A1_c_118_n 5.43096e-19 $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.41
cc_35 VPB N_A1_c_119_n 0.00414814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_B1_M1004_g 0.0187617f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_37 VPB N_B1_c_159_n 0.00292545f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_38 VPB N_B1_c_160_n 0.0046629f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_39 VPB N_C1_M1007_g 0.026191f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_40 VPB C1 0.00386774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_C1_c_205_n 0.00973546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_232_n 0.0102077f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_43 VPB N_VPWR_c_233_n 0.0411758f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_44 VPB N_VPWR_c_234_n 0.00231034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_235_n 0.0130631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_236_n 0.0591683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_231_n 0.0630723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_238_n 0.00368061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_Y_c_298_n 0.0010993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_Y_c_300_n 0.00687849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_Y_c_301_n 0.024518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_A3_c_53_n N_A2_M1000_g 0.0269575f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_53 A3 A2 0.00141892f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A3_c_54_n A2 0.00488584f $X=0.325 $Y=0.995 $X2=0 $Y2=0
cc_55 A3 N_A2_c_78_n 2.55747e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A3_c_53_n N_A2_c_78_n 0.0208026f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_57 A3 N_A2_c_79_n 0.0254894f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A3_c_53_n N_A2_c_79_n 0.00254955f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A3_c_54_n N_A2_c_80_n 0.0341897f $X=0.325 $Y=0.995 $X2=0 $Y2=0
cc_60 A3 N_VPWR_c_233_n 0.0243447f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_61 N_A3_c_53_n N_VPWR_c_233_n 0.00762665f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A3_c_57_n N_VPWR_c_233_n 0.0177289f $X=0.325 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A3_c_57_n N_VPWR_c_234_n 0.00100292f $X=0.325 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A3_c_57_n N_VPWR_c_235_n 0.0046653f $X=0.325 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A3_c_57_n N_VPWR_c_231_n 0.00800869f $X=0.325 $Y=1.41 $X2=0 $Y2=0
cc_66 A3 N_VGND_c_345_n 0.0255459f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A3_c_53_n N_VGND_c_345_n 0.00199688f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A3_c_54_n N_VGND_c_345_n 0.0128284f $X=0.325 $Y=0.995 $X2=0 $Y2=0
cc_69 N_A3_c_54_n N_VGND_c_347_n 0.0046653f $X=0.325 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A3_c_54_n N_VGND_c_349_n 0.00800869f $X=0.325 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A2_M1000_g N_A1_M1008_g 0.0406951f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_72 A2 N_A1_c_117_n 0.00457181f $X=0.615 $Y=0.425 $X2=0 $Y2=0
cc_73 N_A2_c_80_n N_A1_c_117_n 0.00146497f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A2_c_78_n N_A1_c_118_n 0.00103325f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A2_c_79_n N_A1_c_118_n 0.0262171f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A2_c_78_n N_A1_c_119_n 0.021383f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A2_c_79_n N_A1_c_119_n 3.77889e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A2_c_80_n N_A1_c_120_n 0.0395129f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A2_c_79_n N_A1_c_132_n 0.00141937f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A2_c_80_n N_A1_c_132_n 0.00816697f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A2_M1000_g N_VPWR_c_233_n 0.00152112f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A2_M1000_g N_VPWR_c_234_n 0.0129816f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A2_M1000_g N_VPWR_c_235_n 0.0046653f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A2_M1000_g N_VPWR_c_231_n 0.00800869f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A2_M1000_g N_A_109_297#_c_272_n 0.0128027f $X=0.895 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A2_c_79_n N_A_109_297#_c_272_n 0.0107666f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A2_c_78_n N_A_109_297#_c_274_n 3.08478e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A2_c_79_n N_A_109_297#_c_274_n 0.0107917f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A2_M1000_g N_A_109_297#_c_276_n 4.56265e-19 $X=0.895 $Y=1.985 $X2=0
+ $Y2=0
cc_90 N_A2_c_80_n N_VGND_c_345_n 0.00134278f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_91 A2 N_VGND_c_347_n 0.0117108f $X=0.615 $Y=0.425 $X2=0 $Y2=0
cc_92 N_A2_c_80_n N_VGND_c_347_n 0.00577871f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_93 A2 N_VGND_c_349_n 0.00739224f $X=0.615 $Y=0.425 $X2=0 $Y2=0
cc_94 N_A2_c_80_n N_VGND_c_349_n 0.0107215f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_95 A2 A_109_47# 0.00645918f $X=0.615 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_96 N_A1_M1008_g N_B1_M1004_g 0.0325694f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A1_M1008_g N_B1_c_159_n 0.00327232f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A1_c_118_n N_B1_c_159_n 0.0183536f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A1_c_119_n N_B1_c_159_n 0.00197545f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A1_c_118_n N_B1_c_160_n 3.8342e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A1_c_119_n N_B1_c_160_n 0.0204221f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A1_c_117_n N_B1_c_161_n 0.00109306f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A1_c_120_n N_B1_c_161_n 0.0217298f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A1_M1008_g N_VPWR_c_234_n 0.0037129f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A1_M1008_g N_VPWR_c_236_n 0.00544647f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A1_M1008_g N_VPWR_c_231_n 0.0098157f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A1_M1008_g N_A_109_297#_c_272_n 0.0135099f $X=1.325 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A1_c_118_n N_A_109_297#_c_272_n 0.0112204f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A1_c_119_n N_A_109_297#_c_272_n 0.00297344f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A1_M1008_g N_A_109_297#_c_276_n 0.00872609f $X=1.325 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A1_M1008_g N_A_109_297#_c_281_n 0.00225073f $X=1.325 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A1_c_120_n N_Y_c_302_n 0.00286888f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A1_c_132_n N_Y_c_302_n 0.0292673f $X=1.28 $Y=0.462 $X2=0 $Y2=0
cc_114 N_A1_c_117_n N_Y_c_304_n 0.0130236f $X=1.28 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A1_c_120_n N_Y_c_304_n 0.0014156f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A1_c_120_n N_VGND_c_347_n 0.00412562f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A1_c_132_n N_VGND_c_347_n 0.0216209f $X=1.28 $Y=0.462 $X2=0 $Y2=0
cc_118 N_A1_c_120_n N_VGND_c_349_n 0.00683533f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A1_c_132_n N_VGND_c_349_n 0.0145539f $X=1.28 $Y=0.462 $X2=0 $Y2=0
cc_120 N_A1_c_132_n A_194_47# 0.00864838f $X=1.28 $Y=0.462 $X2=-0.19 $Y2=-0.24
cc_121 N_B1_M1004_g N_C1_M1007_g 0.0438928f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_c_159_n N_C1_M1007_g 4.24083e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_123 N_B1_c_175_p N_C1_M1007_g 0.00400645f $X=2.09 $Y=2.005 $X2=0 $Y2=0
cc_124 B1 N_C1_M1007_g 0.0079764f $X=2.005 $Y=2.125 $X2=0 $Y2=0
cc_125 N_B1_c_161_n N_C1_c_203_n 0.0181419f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B1_c_159_n N_C1_c_205_n 3.08917e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B1_c_160_n N_C1_c_205_n 0.0170382f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_128 N_B1_M1004_g N_VPWR_c_236_n 0.00436487f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_129 N_B1_c_175_p N_VPWR_c_236_n 0.00288512f $X=2.09 $Y=2.005 $X2=0 $Y2=0
cc_130 B1 N_VPWR_c_236_n 0.00988361f $X=2.005 $Y=2.125 $X2=0 $Y2=0
cc_131 N_B1_M1004_g N_VPWR_c_231_n 0.00645608f $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_132 N_B1_c_175_p N_VPWR_c_231_n 0.00567281f $X=2.09 $Y=2.005 $X2=0 $Y2=0
cc_133 B1 N_VPWR_c_231_n 0.00984044f $X=2.005 $Y=2.125 $X2=0 $Y2=0
cc_134 N_B1_M1004_g N_A_109_297#_c_272_n 6.7616e-19 $X=1.805 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_B1_M1004_g N_A_109_297#_c_276_n 0.00183861f $X=1.805 $Y=1.985 $X2=0
+ $Y2=0
cc_136 B1 N_A_109_297#_c_276_n 0.00669549f $X=2.005 $Y=2.125 $X2=0 $Y2=0
cc_137 N_B1_c_175_p A_376_297# 0.00688394f $X=2.09 $Y=2.005 $X2=-0.19 $Y2=-0.24
cc_138 B1 A_376_297# 0.0078927f $X=2.005 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_139 N_B1_c_159_n N_Y_c_306_n 0.0145195f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_140 N_B1_c_160_n N_Y_c_306_n 0.00143037f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B1_c_161_n N_Y_c_306_n 0.0119923f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_M1004_g N_Y_c_298_n 4.95428e-19 $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B1_c_159_n N_Y_c_298_n 0.0367252f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B1_c_160_n N_Y_c_298_n 0.00201257f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_145 N_B1_c_161_n N_Y_c_298_n 0.00349461f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B1_M1004_g N_Y_c_300_n 5.91463e-19 $X=1.805 $Y=1.985 $X2=0 $Y2=0
cc_147 N_B1_c_175_p N_Y_c_300_n 0.00487848f $X=2.09 $Y=2.005 $X2=0 $Y2=0
cc_148 N_B1_c_161_n N_VGND_c_346_n 0.00325394f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_149 N_B1_c_161_n N_VGND_c_347_n 0.00427293f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B1_c_161_n N_VGND_c_349_n 0.00600587f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C1_M1007_g N_VPWR_c_236_n 0.00578905f $X=2.3 $Y=1.985 $X2=0 $Y2=0
cc_152 N_C1_M1007_g N_VPWR_c_231_n 0.0121667f $X=2.3 $Y=1.985 $X2=0 $Y2=0
cc_153 N_C1_M1007_g N_Y_c_298_n 0.00866449f $X=2.3 $Y=1.985 $X2=0 $Y2=0
cc_154 N_C1_c_203_n N_Y_c_298_n 0.00836622f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_155 C1 N_Y_c_298_n 0.0229763f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_156 N_C1_c_205_n N_Y_c_298_n 0.00834954f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_157 N_C1_c_203_n N_Y_c_319_n 0.0131003f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_158 C1 N_Y_c_319_n 0.0147377f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_159 N_C1_c_205_n N_Y_c_319_n 0.00141409f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_160 N_C1_M1007_g N_Y_c_300_n 0.0140795f $X=2.3 $Y=1.985 $X2=0 $Y2=0
cc_161 C1 N_Y_c_300_n 0.0151587f $X=2.455 $Y=1.105 $X2=0 $Y2=0
cc_162 N_C1_c_205_n N_Y_c_300_n 0.00307234f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_163 N_C1_c_203_n N_VGND_c_346_n 0.00319864f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_164 N_C1_c_203_n N_VGND_c_348_n 0.00428022f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_165 N_C1_c_203_n N_VGND_c_349_n 0.00724932f $X=2.325 $Y=0.995 $X2=0 $Y2=0
cc_166 N_VPWR_c_231_n N_A_109_297#_M1006_d 0.00607087f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_167 N_VPWR_c_231_n N_A_109_297#_M1008_d 0.00325684f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_235_n N_A_109_297#_c_287_n 0.00565015f $X=0.94 $Y=2.72 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_231_n N_A_109_297#_c_287_n 0.0058949f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_170 N_VPWR_M1000_d N_A_109_297#_c_272_n 0.00809843f $X=0.97 $Y=1.485 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_234_n N_A_109_297#_c_272_n 0.0156725f $X=1.105 $Y=2.08 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_236_n N_A_109_297#_c_281_n 0.0105131f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_231_n N_A_109_297#_c_281_n 0.0112095f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_231_n A_376_297# 0.00323933f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_175 N_VPWR_c_231_n N_Y_M1007_d 0.00348903f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_176 N_VPWR_c_236_n N_Y_c_301_n 0.00868346f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_177 N_VPWR_c_231_n N_Y_c_301_n 0.00851907f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_178 A_376_297# N_Y_c_298_n 2.68705e-19 $X=1.88 $Y=1.485 $X2=0 $Y2=0
cc_179 A_376_297# N_Y_c_300_n 0.00232693f $X=1.88 $Y=1.485 $X2=0 $Y2=0
cc_180 N_Y_c_306_n N_VGND_M1001_d 0.00626473f $X=2.105 $Y=0.74 $X2=0 $Y2=0
cc_181 N_Y_c_298_n N_VGND_M1001_d 9.6607e-19 $X=2.19 $Y=1.495 $X2=0 $Y2=0
cc_182 N_Y_c_319_n N_VGND_M1001_d 0.00116047f $X=2.527 $Y=0.655 $X2=0 $Y2=0
cc_183 N_Y_c_306_n N_VGND_c_346_n 0.0177002f $X=2.105 $Y=0.74 $X2=0 $Y2=0
cc_184 N_Y_c_302_n N_VGND_c_347_n 0.011459f $X=1.62 $Y=0.42 $X2=0 $Y2=0
cc_185 N_Y_c_306_n N_VGND_c_347_n 0.00279912f $X=2.105 $Y=0.74 $X2=0 $Y2=0
cc_186 N_Y_c_319_n N_VGND_c_348_n 0.00254024f $X=2.527 $Y=0.655 $X2=0 $Y2=0
cc_187 Y N_VGND_c_348_n 0.0117315f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_188 N_Y_M1005_d N_VGND_c_349_n 0.00774885f $X=1.4 $Y=0.235 $X2=0 $Y2=0
cc_189 N_Y_M1003_d N_VGND_c_349_n 0.00248504f $X=2.4 $Y=0.235 $X2=0 $Y2=0
cc_190 N_Y_c_302_n N_VGND_c_349_n 0.00644035f $X=1.62 $Y=0.42 $X2=0 $Y2=0
cc_191 N_Y_c_306_n N_VGND_c_349_n 0.00618703f $X=2.105 $Y=0.74 $X2=0 $Y2=0
cc_192 N_Y_c_319_n N_VGND_c_349_n 0.0039971f $X=2.527 $Y=0.655 $X2=0 $Y2=0
cc_193 Y N_VGND_c_349_n 0.00900857f $X=2.465 $Y=0.425 $X2=0 $Y2=0
cc_194 N_VGND_c_349_n A_109_47# 0.00505731f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_195 N_VGND_c_349_n A_194_47# 0.0022523f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__fahcin_1.spice
* Created: Tue Sep  1 19:09:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__fahcin_1.pex.spice"
.subckt sky130_fd_sc_hd__fahcin_1  VNB VPB A B CIN VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_67_199#_M1007_g N_A_27_47#_M1007_s VNB NSHORT L=0.15
+ W=0.64 AD=0.104434 AS=0.1696 PD=0.967442 PS=1.81 NRD=4.68 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1018 N_A_67_199#_M1018_d N_A_M1018_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.323715 AS=0.106066 PD=1.65775 PS=0.982558 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_434_49#_M1005_d N_B_M1005_g N_A_67_199#_M1018_d VNB NSHORT L=0.15
+ W=0.64 AD=0.088 AS=0.318735 PD=0.915 PS=1.63225 NRD=0 NRS=67.02 M=1 R=4.26667
+ SA=75001.8 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1026 N_A_27_47#_M1026_d N_A_489_21#_M1026_g N_A_434_49#_M1005_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.199825 AS=0.088 PD=1.91 PS=0.915 NRD=9.372 NRS=0 M=1
+ R=4.26667 SA=75002.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1028 N_A_721_47#_M1028_d N_A_489_21#_M1028_g N_A_67_199#_M1028_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.165675 AS=0.168125 PD=1.165 PS=1.83 NRD=44.988 NRS=1.872
+ M=1 R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 N_A_27_47#_M1012_d N_B_M1012_g N_A_721_47#_M1028_d VNB NSHORT L=0.15
+ W=0.64 AD=0.162825 AS=0.165675 PD=1.8 PS=1.165 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_B_M1015_g N_A_489_21#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.117353 AS=0.165325 PD=1.01783 PS=1.82 NRD=0.912 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1024 N_A_1142_49#_M1024_d N_A_489_21#_M1024_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1664 AS=0.115547 PD=1.8 PS=1.00217 NRD=0 NRS=14.052 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1031 N_COUT_M1031_d N_A_434_49#_M1031_g N_A_1251_49#_M1031_s VNB NSHORT L=0.15
+ W=0.64 AD=0.088 AS=0.192 PD=0.915 PS=1.88 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_A_1142_49#_M1014_d N_A_721_47#_M1014_g N_COUT_M1031_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1792 AS=0.088 PD=1.84 PS=0.915 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_1647_49#_M1029_d N_A_721_47#_M1029_g N_A_1565_49#_M1029_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0928 AS=0.1664 PD=0.93 PS=1.8 NRD=2.808 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1019 N_A_1636_315#_M1019_d N_A_434_49#_M1019_g N_A_1647_49#_M1029_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.4768 AS=0.0928 PD=2.77 PS=0.93 NRD=14.052 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A_1636_315#_M1001_g N_A_1565_49#_M1001_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.104434 AS=0.1728 PD=0.967442 PS=1.82 NRD=2.808 NRS=0.936
+ M=1 R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1022 N_A_1636_315#_M1022_d N_CIN_M1022_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.106066 PD=1.82 PS=0.982558 NRD=0 NRS=5.532 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_CIN_M1008_g N_A_1251_49#_M1008_s VNB NSHORT L=0.15
+ W=0.64 AD=0.104434 AS=0.1664 PD=0.967442 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1025 N_SUM_M1025_d N_A_1647_49#_M1025_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.65 AD=0.18525 AS=0.106066 PD=1.87 PS=0.982558 NRD=3.684 NRS=9.228 M=1
+ R=4.33333 SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_VPWR_M1013_d N_A_67_199#_M1013_g N_A_27_47#_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.265 PD=1.35 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1010 N_A_67_199#_M1010_d N_A_M1010_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.31175 AS=0.175 PD=2.88 PS=1.35 NRD=34.4553 NRS=14.7553 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1027 N_A_434_49#_M1027_d N_B_M1027_g N_A_27_47#_M1027_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1155 AS=0.2629 PD=1.115 PS=2.64 NRD=0 NRS=18.7544 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_A_67_199#_M1003_d N_A_489_21#_M1003_g N_A_434_49#_M1027_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2184 AS=0.1155 PD=2.2 PS=1.115 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 N_A_721_47#_M1020_d N_A_489_21#_M1020_g N_A_27_47#_M1020_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.152262 AS=0.3398 PD=1.3 PS=2.77 NRD=0 NRS=9.3772 M=1 R=5.6
+ SA=75000.3 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1011 N_A_67_199#_M1011_d N_B_M1011_g N_A_721_47#_M1020_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2814 AS=0.152262 PD=2.35 PS=1.3 NRD=0 NRS=14.0658 M=1 R=5.6
+ SA=75000.7 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_489_21#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.18 AS=0.26 PD=1.36 PS=2.52 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1006 N_A_1142_49#_M1006_d N_A_489_21#_M1006_g N_VPWR_M1004_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.41587 AS=0.18 PD=1.94565 PS=1.36 NRD=50.2153 NRS=0 M=1
+ R=6.66667 SA=75000.7 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1030 N_COUT_M1030_d N_A_434_49#_M1030_g N_A_1142_49#_M1006_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1134 AS=0.34933 PD=1.11 PS=1.63435 NRD=0 NRS=59.7895 M=1
+ R=5.6 SA=75001.6 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1009 N_A_1251_49#_M1009_d N_A_721_47#_M1009_g N_COUT_M1030_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.7033 AS=0.1134 PD=3.36 PS=1.11 NRD=59.7895 NRS=0 M=1 R=5.6
+ SA=75002.1 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1000 N_A_1647_49#_M1000_d N_A_721_47#_M1000_g N_A_1636_315#_M1000_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1134 AS=0.2184 PD=1.11 PS=2.2 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1023 N_A_1565_49#_M1023_d N_A_434_49#_M1023_g N_A_1647_49#_M1000_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.410139 AS=0.1134 PD=1.80783 PS=1.11 NRD=164.16 NRS=0 M=1
+ R=5.6 SA=75000.6 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_1636_315#_M1002_g N_A_1565_49#_M1023_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.488261 PD=1.27 PS=2.15217 NRD=0 NRS=0.9653 M=1
+ R=6.66667 SA=75001.5 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1016 N_A_1636_315#_M1016_d N_CIN_M1016_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.135 PD=2.53 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1021_d N_CIN_M1021_g N_A_1251_49#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_SUM_M1017_d N_A_1647_49#_M1017_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.135 PD=2.57 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.544 P=28.81
pX33_noxref noxref_20 B B PROBETYPE=1
c_209 VPB 0 1.75206e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__fahcin_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__clkinv_8.spice.SKY130_FD_SC_HD__CLKINV_8.pxi
* Created: Thu Aug 27 14:12:50 2020
* 
x_PM_SKY130_FD_SC_HD__CLKINV_8%A N_A_c_100_n N_A_M1000_g N_A_c_101_n N_A_M1003_g
+ N_A_c_102_n N_A_M1004_g N_A_M1001_g N_A_c_103_n N_A_M1006_g N_A_M1002_g
+ N_A_c_104_n N_A_M1007_g N_A_M1005_g N_A_c_105_n N_A_M1010_g N_A_M1008_g
+ N_A_c_106_n N_A_M1012_g N_A_M1009_g N_A_c_107_n N_A_M1013_g N_A_M1011_g
+ N_A_c_108_n N_A_M1014_g N_A_M1016_g N_A_c_109_n N_A_M1015_g N_A_M1017_g
+ N_A_c_110_n N_A_M1018_g N_A_c_111_n N_A_M1019_g A A A A A A A A A N_A_c_149_p
+ N_A_c_99_n PM_SKY130_FD_SC_HD__CLKINV_8%A
x_PM_SKY130_FD_SC_HD__CLKINV_8%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1006_s
+ N_VPWR_M1010_s N_VPWR_M1013_s N_VPWR_M1015_s N_VPWR_M1019_s N_VPWR_c_260_n
+ N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_265_n
+ N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n
+ N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n VPWR
+ N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_259_n N_VPWR_c_279_n
+ N_VPWR_c_280_n N_VPWR_c_281_n PM_SKY130_FD_SC_HD__CLKINV_8%VPWR
x_PM_SKY130_FD_SC_HD__CLKINV_8%Y N_Y_M1001_d N_Y_M1005_d N_Y_M1009_d N_Y_M1016_d
+ N_Y_M1000_d N_Y_M1004_d N_Y_M1007_d N_Y_M1012_d N_Y_M1014_d N_Y_M1018_d
+ N_Y_c_352_n N_Y_c_353_n N_Y_c_354_n N_Y_c_366_n N_Y_c_367_n N_Y_c_463_n
+ N_Y_c_368_n N_Y_c_467_n N_Y_c_355_n N_Y_c_369_n N_Y_c_356_n N_Y_c_471_n
+ N_Y_c_357_n N_Y_c_370_n N_Y_c_358_n N_Y_c_475_n N_Y_c_359_n N_Y_c_371_n
+ N_Y_c_360_n N_Y_c_479_n N_Y_c_361_n N_Y_c_372_n N_Y_c_362_n N_Y_c_483_n
+ N_Y_c_373_n N_Y_c_374_n N_Y_c_434_n N_Y_c_375_n N_Y_c_438_n N_Y_c_376_n
+ N_Y_c_442_n N_Y_c_377_n N_Y_c_446_n Y Y Y N_Y_c_364_n N_Y_c_379_n
+ PM_SKY130_FD_SC_HD__CLKINV_8%Y
x_PM_SKY130_FD_SC_HD__CLKINV_8%VGND N_VGND_M1001_s N_VGND_M1002_s N_VGND_M1008_s
+ N_VGND_M1011_s N_VGND_M1017_s N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n
+ N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n
+ N_VGND_c_531_n VGND N_VGND_c_532_n N_VGND_c_533_n N_VGND_c_534_n
+ N_VGND_c_535_n N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n N_VGND_c_539_n
+ VGND PM_SKY130_FD_SC_HD__CLKINV_8%VGND
cc_1 VNB N_A_M1001_g 0.0222492f $X=-0.19 $Y=-0.24 $X2=1.415 $Y2=0.445
cc_2 VNB N_A_M1002_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=1.845 $Y2=0.445
cc_3 VNB N_A_M1005_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=2.275 $Y2=0.445
cc_4 VNB N_A_M1008_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.445
cc_5 VNB N_A_M1009_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=3.135 $Y2=0.445
cc_6 VNB N_A_M1011_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=0.445
cc_7 VNB N_A_M1016_g 0.0173004f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.445
cc_8 VNB N_A_M1017_g 0.0222492f $X=-0.19 $Y=-0.24 $X2=4.425 $Y2=0.445
cc_9 VNB N_A_c_99_n 0.342075f $X=-0.19 $Y=-0.24 $X2=5.095 $Y2=1.097
cc_10 VNB N_VPWR_c_259_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_352_n 0.0204208f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.445
cc_12 VNB N_Y_c_353_n 0.0150647f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=0.445
cc_13 VNB N_Y_c_354_n 0.00997812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_355_n 6.75361e-19 $X=-0.19 $Y=-0.24 $X2=3.835 $Y2=1.385
cc_15 VNB N_Y_c_356_n 0.0035731f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.445
cc_16 VNB N_Y_c_357_n 6.52615e-19 $X=-0.19 $Y=-0.24 $X2=4.425 $Y2=0.445
cc_17 VNB N_Y_c_358_n 0.0035731f $X=-0.19 $Y=-0.24 $X2=4.675 $Y2=1.985
cc_18 VNB N_Y_c_359_n 6.52615e-19 $X=-0.19 $Y=-0.24 $X2=2.45 $Y2=1.105
cc_19 VNB N_Y_c_360_n 0.0035731f $X=-0.19 $Y=-0.24 $X2=4.29 $Y2=1.105
cc_20 VNB N_Y_c_361_n 6.75361e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_362_n 0.00820216f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.097
cc_22 VNB Y 0.0225434f $X=-0.19 $Y=-0.24 $X2=3.565 $Y2=1.097
cc_23 VNB N_Y_c_364_n 0.0113484f $X=-0.19 $Y=-0.24 $X2=4.7 $Y2=1.16
cc_24 VNB N_VGND_c_523_n 0.0141137f $X=-0.19 $Y=-0.24 $X2=1.845 $Y2=0.445
cc_25 VNB N_VGND_c_524_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=2.155 $Y2=1.985
cc_26 VNB N_VGND_c_525_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=2.275 $Y2=0.445
cc_27 VNB N_VGND_c_526_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=1.985
cc_28 VNB N_VGND_c_527_n 0.0141137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_528_n 0.011666f $X=-0.19 $Y=-0.24 $X2=2.995 $Y2=1.985
cc_30 VNB N_VGND_c_529_n 0.00436502f $X=-0.19 $Y=-0.24 $X2=3.135 $Y2=0.81
cc_31 VNB N_VGND_c_530_n 0.011666f $X=-0.19 $Y=-0.24 $X2=3.135 $Y2=0.445
cc_32 VNB N_VGND_c_531_n 0.00510476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_532_n 0.0314546f $X=-0.19 $Y=-0.24 $X2=3.415 $Y2=1.985
cc_34 VNB N_VGND_c_533_n 0.011666f $X=-0.19 $Y=-0.24 $X2=3.835 $Y2=1.385
cc_35 VNB N_VGND_c_534_n 0.011666f $X=-0.19 $Y=-0.24 $X2=3.995 $Y2=0.445
cc_36 VNB N_VGND_c_535_n 0.0370325f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_37 VNB N_VGND_c_536_n 0.332673f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_38 VNB N_VGND_c_537_n 0.00510476f $X=-0.19 $Y=-0.24 $X2=2.91 $Y2=1.105
cc_39 VNB N_VGND_c_538_n 0.00436502f $X=-0.19 $Y=-0.24 $X2=4.29 $Y2=1.105
cc_40 VNB N_VGND_c_539_n 0.00436502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VPB N_A_c_100_n 0.0186165f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.385
cc_42 VPB N_A_c_101_n 0.0152912f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.385
cc_43 VPB N_A_c_102_n 0.0153104f $X=-0.19 $Y=1.305 $X2=1.315 $Y2=1.385
cc_44 VPB N_A_c_103_n 0.0152623f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=1.385
cc_45 VPB N_A_c_104_n 0.0152623f $X=-0.19 $Y=1.305 $X2=2.155 $Y2=1.385
cc_46 VPB N_A_c_105_n 0.0152623f $X=-0.19 $Y=1.305 $X2=2.575 $Y2=1.385
cc_47 VPB N_A_c_106_n 0.0152623f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.385
cc_48 VPB N_A_c_107_n 0.0152623f $X=-0.19 $Y=1.305 $X2=3.415 $Y2=1.385
cc_49 VPB N_A_c_108_n 0.0152623f $X=-0.19 $Y=1.305 $X2=3.835 $Y2=1.385
cc_50 VPB N_A_c_109_n 0.0152623f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.385
cc_51 VPB N_A_c_110_n 0.0152408f $X=-0.19 $Y=1.305 $X2=4.675 $Y2=1.385
cc_52 VPB N_A_c_111_n 0.0186132f $X=-0.19 $Y=1.305 $X2=5.095 $Y2=1.385
cc_53 VPB N_A_c_99_n 0.0693682f $X=-0.19 $Y=1.305 $X2=5.095 $Y2=1.097
cc_54 VPB N_VPWR_c_260_n 0.0114824f $X=-0.19 $Y=1.305 $X2=2.155 $Y2=1.985
cc_55 VPB N_VPWR_c_261_n 0.0046049f $X=-0.19 $Y=1.305 $X2=2.275 $Y2=0.81
cc_56 VPB N_VPWR_c_262_n 0.00395987f $X=-0.19 $Y=1.305 $X2=2.575 $Y2=1.385
cc_57 VPB N_VPWR_c_263_n 0.00397229f $X=-0.19 $Y=1.305 $X2=2.705 $Y2=0.445
cc_58 VPB N_VPWR_c_264_n 0.00389651f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.985
cc_59 VPB N_VPWR_c_265_n 0.00395746f $X=-0.19 $Y=1.305 $X2=3.135 $Y2=0.445
cc_60 VPB N_VPWR_c_266_n 0.0166258f $X=-0.19 $Y=1.305 $X2=3.415 $Y2=1.385
cc_61 VPB N_VPWR_c_267_n 0.00392376f $X=-0.19 $Y=1.305 $X2=3.565 $Y2=0.445
cc_62 VPB N_VPWR_c_268_n 0.00457723f $X=-0.19 $Y=1.305 $X2=3.835 $Y2=1.985
cc_63 VPB N_VPWR_c_269_n 0.0161792f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=0.445
cc_64 VPB N_VPWR_c_270_n 0.00497514f $X=-0.19 $Y=1.305 $X2=3.995 $Y2=0.445
cc_65 VPB N_VPWR_c_271_n 0.0164599f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.385
cc_66 VPB N_VPWR_c_272_n 0.00468662f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.985
cc_67 VPB N_VPWR_c_273_n 0.0163451f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.985
cc_68 VPB N_VPWR_c_274_n 0.00487897f $X=-0.19 $Y=1.305 $X2=4.425 $Y2=0.81
cc_69 VPB N_VPWR_c_275_n 0.0162816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_276_n 0.0161407f $X=-0.19 $Y=1.305 $X2=4.29 $Y2=1.105
cc_71 VPB N_VPWR_c_277_n 0.0196454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_259_n 0.063808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_279_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_74 VPB N_VPWR_c_280_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.415 $Y2=1.097
cc_75 VPB N_VPWR_c_281_n 0.00487897f $X=-0.19 $Y=1.305 $X2=2.155 $Y2=1.097
cc_76 VPB N_Y_c_352_n 0.00728169f $X=-0.19 $Y=1.305 $X2=2.705 $Y2=0.445
cc_77 VPB N_Y_c_366_n 0.00171067f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.385
cc_78 VPB N_Y_c_367_n 0.00789722f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.985
cc_79 VPB N_Y_c_368_n 0.00241699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_Y_c_369_n 0.00243386f $X=-0.19 $Y=1.305 $X2=3.835 $Y2=1.985
cc_81 VPB N_Y_c_370_n 0.00225932f $X=-0.19 $Y=1.305 $X2=4.675 $Y2=1.385
cc_82 VPB N_Y_c_371_n 0.00238793f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.105
cc_83 VPB N_Y_c_372_n 0.00230525f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.097
cc_84 VPB N_Y_c_373_n 0.00194324f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=1.097
cc_85 VPB N_Y_c_374_n 0.00194324f $X=-0.19 $Y=1.305 $X2=1.845 $Y2=1.097
cc_86 VPB N_Y_c_375_n 0.00203715f $X=-0.19 $Y=1.305 $X2=2.275 $Y2=1.097
cc_87 VPB N_Y_c_376_n 0.00199019f $X=-0.19 $Y=1.305 $X2=2.705 $Y2=1.097
cc_88 VPB N_Y_c_377_n 0.0020841f $X=-0.19 $Y=1.305 $X2=3.135 $Y2=1.097
cc_89 VPB Y 0.00839106f $X=-0.19 $Y=1.305 $X2=3.565 $Y2=1.097
cc_90 VPB N_Y_c_379_n 0.0106811f $X=-0.19 $Y=1.305 $X2=5.095 $Y2=1.097
cc_91 N_A_c_100_n N_VPWR_c_261_n 0.00342588f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_92 N_A_c_101_n N_VPWR_c_262_n 0.00157835f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_93 N_A_c_102_n N_VPWR_c_262_n 0.00159968f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_94 N_A_c_103_n N_VPWR_c_263_n 0.00159118f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_95 N_A_c_104_n N_VPWR_c_263_n 0.00160491f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_96 N_A_c_105_n N_VPWR_c_264_n 0.00155476f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_97 N_A_c_106_n N_VPWR_c_264_n 0.00156899f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A_c_107_n N_VPWR_c_265_n 0.00159548f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A_c_108_n N_VPWR_c_265_n 0.0015877f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_100 N_A_c_108_n N_VPWR_c_266_n 0.00585385f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_101 N_A_c_109_n N_VPWR_c_266_n 0.00585385f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_102 N_A_c_109_n N_VPWR_c_267_n 0.00156401f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_103 N_A_c_110_n N_VPWR_c_267_n 0.00158601f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_104 N_A_c_111_n N_VPWR_c_268_n 0.00340482f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_105 N_A_c_102_n N_VPWR_c_269_n 0.00585385f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_106 N_A_c_103_n N_VPWR_c_269_n 0.00585385f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_107 N_A_c_104_n N_VPWR_c_271_n 0.00585385f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_108 N_A_c_105_n N_VPWR_c_271_n 0.00585385f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_109 N_A_c_106_n N_VPWR_c_273_n 0.00585385f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_110 N_A_c_107_n N_VPWR_c_273_n 0.00585385f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A_c_100_n N_VPWR_c_275_n 0.00583607f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_112 N_A_c_101_n N_VPWR_c_275_n 0.00585385f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_113 N_A_c_110_n N_VPWR_c_276_n 0.00585385f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_114 N_A_c_111_n N_VPWR_c_276_n 0.00585385f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_115 N_A_c_100_n N_VPWR_c_259_n 0.0114285f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_116 N_A_c_101_n N_VPWR_c_259_n 0.0105259f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_117 N_A_c_102_n N_VPWR_c_259_n 0.0105133f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_118 N_A_c_103_n N_VPWR_c_259_n 0.0105001f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_119 N_A_c_104_n N_VPWR_c_259_n 0.0105001f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_120 N_A_c_105_n N_VPWR_c_259_n 0.0105252f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_121 N_A_c_106_n N_VPWR_c_259_n 0.0105126f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_122 N_A_c_107_n N_VPWR_c_259_n 0.0105001f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_123 N_A_c_108_n N_VPWR_c_259_n 0.0105126f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_124 N_A_c_109_n N_VPWR_c_259_n 0.0105252f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A_c_110_n N_VPWR_c_259_n 0.0105001f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A_c_111_n N_VPWR_c_259_n 0.0118261f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_127 N_A_c_149_p N_Y_c_352_n 0.0202172f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_c_99_n N_Y_c_352_n 0.0216629f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_129 N_A_M1001_g N_Y_c_353_n 0.0090634f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A_c_149_p N_Y_c_353_n 0.0755218f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_99_n N_Y_c_353_n 0.0388808f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_132 N_A_c_100_n N_Y_c_366_n 0.017106f $X=0.47 $Y=1.385 $X2=0 $Y2=0
cc_133 N_A_c_149_p N_Y_c_366_n 0.00773305f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_101_n N_Y_c_368_n 0.0149361f $X=0.89 $Y=1.385 $X2=0 $Y2=0
cc_135 N_A_c_102_n N_Y_c_368_n 0.0149803f $X=1.315 $Y=1.385 $X2=0 $Y2=0
cc_136 N_A_c_149_p N_Y_c_368_n 0.0430258f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_99_n N_Y_c_368_n 0.0026718f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_138 N_A_M1001_g N_Y_c_355_n 0.00101119f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_M1002_g N_Y_c_355_n 5.8681e-19 $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A_c_103_n N_Y_c_369_n 0.0149489f $X=1.735 $Y=1.385 $X2=0 $Y2=0
cc_141 N_A_c_104_n N_Y_c_369_n 0.0149489f $X=2.155 $Y=1.385 $X2=0 $Y2=0
cc_142 N_A_c_149_p N_Y_c_369_n 0.0430259f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_c_99_n N_Y_c_369_n 0.00265179f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_144 N_A_M1002_g N_Y_c_356_n 0.0076909f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_M1005_g N_Y_c_356_n 0.0076909f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_c_149_p N_Y_c_356_n 0.0468048f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_99_n N_Y_c_356_n 0.014197f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_Y_c_357_n 5.8681e-19 $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_M1008_g N_Y_c_357_n 5.8681e-19 $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_c_105_n N_Y_c_370_n 0.0149489f $X=2.575 $Y=1.385 $X2=0 $Y2=0
cc_151 N_A_c_106_n N_Y_c_370_n 0.0149489f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_152 N_A_c_149_p N_Y_c_370_n 0.0419202f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_c_99_n N_Y_c_370_n 0.00265179f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_154 N_A_M1008_g N_Y_c_358_n 0.0076909f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A_M1009_g N_Y_c_358_n 0.0076909f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A_c_149_p N_Y_c_358_n 0.0468048f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_c_99_n N_Y_c_358_n 0.0141423f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_158 N_A_M1009_g N_Y_c_359_n 5.8681e-19 $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_M1011_g N_Y_c_359_n 5.8681e-19 $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_c_107_n N_Y_c_371_n 0.0149489f $X=3.415 $Y=1.385 $X2=0 $Y2=0
cc_161 N_A_c_108_n N_Y_c_371_n 0.0149489f $X=3.835 $Y=1.385 $X2=0 $Y2=0
cc_162 N_A_c_149_p N_Y_c_371_n 0.0426573f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_c_99_n N_Y_c_371_n 0.00265179f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_164 N_A_M1011_g N_Y_c_360_n 0.0076909f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_M1016_g N_Y_c_360_n 0.0076909f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_c_149_p N_Y_c_360_n 0.0468048f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_c_99_n N_Y_c_360_n 0.014197f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_168 N_A_M1016_g N_Y_c_361_n 5.8681e-19 $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_M1017_g N_Y_c_361_n 0.00101119f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_170 N_A_c_109_n N_Y_c_372_n 0.0149489f $X=4.255 $Y=1.385 $X2=0 $Y2=0
cc_171 N_A_c_110_n N_Y_c_372_n 0.0149047f $X=4.675 $Y=1.385 $X2=0 $Y2=0
cc_172 N_A_c_149_p N_Y_c_372_n 0.0496601f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_99_n N_Y_c_372_n 0.00263839f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_174 N_A_M1017_g N_Y_c_362_n 0.0090634f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A_c_149_p N_Y_c_362_n 0.0391432f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_c_99_n N_Y_c_362_n 0.0310808f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_177 N_A_c_149_p N_Y_c_373_n 0.0198915f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_99_n N_Y_c_373_n 0.00262698f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_179 N_A_c_149_p N_Y_c_374_n 0.0198915f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_c_99_n N_Y_c_374_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_181 N_A_c_149_p N_Y_c_434_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_c_99_n N_Y_c_434_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_183 N_A_c_149_p N_Y_c_375_n 0.0207204f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_c_99_n N_Y_c_375_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_185 N_A_c_149_p N_Y_c_438_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_99_n N_Y_c_438_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_187 N_A_c_149_p N_Y_c_376_n 0.020306f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_c_99_n N_Y_c_376_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_189 N_A_c_149_p N_Y_c_442_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_c_99_n N_Y_c_442_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_191 N_A_c_149_p N_Y_c_377_n 0.0211349f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_c_99_n N_Y_c_377_n 0.00274773f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_193 N_A_c_149_p N_Y_c_446_n 0.0147099f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_c_99_n N_Y_c_446_n 0.00596888f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_195 N_A_c_149_p Y 0.0134731f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_c_99_n Y 0.0260425f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_197 N_A_c_99_n N_Y_c_364_n 0.00106081f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_198 N_A_c_111_n N_Y_c_379_n 0.0182383f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_199 N_A_c_99_n N_Y_c_379_n 0.00286303f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_200 N_A_M1001_g N_VGND_c_523_n 0.00831231f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_201 N_A_M1002_g N_VGND_c_523_n 5.62611e-19 $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A_c_99_n N_VGND_c_523_n 0.00163226f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_203 N_A_M1001_g N_VGND_c_524_n 5.62611e-19 $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_204 N_A_M1002_g N_VGND_c_524_n 0.00724882f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A_M1005_g N_VGND_c_524_n 0.00724882f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A_M1008_g N_VGND_c_524_n 5.62611e-19 $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A_c_99_n N_VGND_c_524_n 5.80335e-19 $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_208 N_A_M1005_g N_VGND_c_525_n 5.62611e-19 $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_209 N_A_M1008_g N_VGND_c_525_n 0.00724882f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_210 N_A_M1009_g N_VGND_c_525_n 0.00724882f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_211 N_A_M1011_g N_VGND_c_525_n 5.62611e-19 $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_212 N_A_c_99_n N_VGND_c_525_n 5.80335e-19 $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_213 N_A_M1009_g N_VGND_c_526_n 5.62611e-19 $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A_M1011_g N_VGND_c_526_n 0.00724882f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A_M1016_g N_VGND_c_526_n 0.00724882f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A_M1017_g N_VGND_c_526_n 5.62611e-19 $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A_c_99_n N_VGND_c_526_n 5.80335e-19 $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_218 N_A_M1016_g N_VGND_c_527_n 5.62611e-19 $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A_M1017_g N_VGND_c_527_n 0.00831231f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_c_99_n N_VGND_c_527_n 0.0016306f $X=5.095 $Y=1.097 $X2=0 $Y2=0
cc_221 N_A_M1009_g N_VGND_c_528_n 0.00360664f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_M1011_g N_VGND_c_528_n 0.00360664f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A_M1016_g N_VGND_c_530_n 0.00360664f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_224 N_A_M1017_g N_VGND_c_530_n 0.00360664f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_M1001_g N_VGND_c_533_n 0.00360664f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_226 N_A_M1002_g N_VGND_c_533_n 0.00360664f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_227 N_A_M1005_g N_VGND_c_534_n 0.00360664f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_228 N_A_M1008_g N_VGND_c_534_n 0.00360664f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_M1001_g N_VGND_c_536_n 0.00428048f $X=1.415 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A_M1002_g N_VGND_c_536_n 0.00428048f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_231 N_A_M1005_g N_VGND_c_536_n 0.00428048f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_232 N_A_M1008_g N_VGND_c_536_n 0.00428048f $X=2.705 $Y=0.445 $X2=0 $Y2=0
cc_233 N_A_M1009_g N_VGND_c_536_n 0.00428048f $X=3.135 $Y=0.445 $X2=0 $Y2=0
cc_234 N_A_M1011_g N_VGND_c_536_n 0.00428048f $X=3.565 $Y=0.445 $X2=0 $Y2=0
cc_235 N_A_M1016_g N_VGND_c_536_n 0.00428048f $X=3.995 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A_M1017_g N_VGND_c_536_n 0.00428048f $X=4.425 $Y=0.445 $X2=0 $Y2=0
cc_237 N_VPWR_c_259_n N_Y_M1000_d 0.00329227f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_238 N_VPWR_c_259_n N_Y_M1004_d 0.00329227f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_239 N_VPWR_c_259_n N_Y_M1007_d 0.00294567f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_240 N_VPWR_c_259_n N_Y_M1012_d 0.00311897f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_241 N_VPWR_c_259_n N_Y_M1014_d 0.00277237f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_242 N_VPWR_c_259_n N_Y_M1018_d 0.00329227f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_243 N_VPWR_M1000_s N_Y_c_366_n 5.5277e-19 $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_244 N_VPWR_c_261_n N_Y_c_366_n 0.00427553f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_245 N_VPWR_M1000_s N_Y_c_367_n 0.00229093f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_246 N_VPWR_c_261_n N_Y_c_367_n 0.0134341f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_247 N_VPWR_c_275_n N_Y_c_463_n 0.0116691f $X=0.975 $Y=2.72 $X2=0 $Y2=0
cc_248 N_VPWR_c_259_n N_Y_c_463_n 0.00903178f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_249 N_VPWR_M1003_s N_Y_c_368_n 0.00171146f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_250 N_VPWR_c_262_n N_Y_c_368_n 0.0130987f $X=1.105 $Y=1.965 $X2=0 $Y2=0
cc_251 N_VPWR_c_269_n N_Y_c_467_n 0.0116691f $X=1.815 $Y=2.72 $X2=0 $Y2=0
cc_252 N_VPWR_c_259_n N_Y_c_467_n 0.00903178f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_253 N_VPWR_M1006_s N_Y_c_369_n 0.00165831f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_254 N_VPWR_c_263_n N_Y_c_369_n 0.0126919f $X=1.945 $Y=1.965 $X2=0 $Y2=0
cc_255 N_VPWR_c_271_n N_Y_c_471_n 0.0119709f $X=2.665 $Y=2.72 $X2=0 $Y2=0
cc_256 N_VPWR_c_259_n N_Y_c_471_n 0.00941127f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_257 N_VPWR_M1010_s N_Y_c_370_n 0.00165831f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_258 N_VPWR_c_264_n N_Y_c_370_n 0.0126919f $X=2.785 $Y=1.965 $X2=0 $Y2=0
cc_259 N_VPWR_c_273_n N_Y_c_475_n 0.01182f $X=3.495 $Y=2.72 $X2=0 $Y2=0
cc_260 N_VPWR_c_259_n N_Y_c_475_n 0.00922153f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_261 N_VPWR_M1013_s N_Y_c_371_n 0.00165831f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_262 N_VPWR_c_265_n N_Y_c_371_n 0.0126919f $X=3.625 $Y=1.965 $X2=0 $Y2=0
cc_263 N_VPWR_c_266_n N_Y_c_479_n 0.0121219f $X=4.345 $Y=2.72 $X2=0 $Y2=0
cc_264 N_VPWR_c_259_n N_Y_c_479_n 0.00960102f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_265 N_VPWR_M1015_s N_Y_c_372_n 0.00165831f $X=4.33 $Y=1.485 $X2=0 $Y2=0
cc_266 N_VPWR_c_267_n N_Y_c_372_n 0.0126919f $X=4.465 $Y=1.965 $X2=0 $Y2=0
cc_267 N_VPWR_c_276_n N_Y_c_483_n 0.0116691f $X=5.175 $Y=2.72 $X2=0 $Y2=0
cc_268 N_VPWR_c_259_n N_Y_c_483_n 0.00903178f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_M1019_s N_Y_c_379_n 0.00278493f $X=5.17 $Y=1.485 $X2=0 $Y2=0
cc_270 N_VPWR_c_268_n N_Y_c_379_n 0.0164344f $X=5.305 $Y=1.965 $X2=0 $Y2=0
cc_271 N_Y_c_353_n N_VGND_c_523_n 0.0232314f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_272 N_Y_c_356_n N_VGND_c_524_n 0.020457f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_273 N_Y_c_358_n N_VGND_c_525_n 0.020457f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_274 N_Y_c_360_n N_VGND_c_526_n 0.020457f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_275 N_Y_c_362_n N_VGND_c_527_n 0.0232314f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_276 N_Y_c_358_n N_VGND_c_528_n 0.00249722f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_277 N_Y_c_359_n N_VGND_c_528_n 0.0106278f $X=3.35 $Y=0.445 $X2=0 $Y2=0
cc_278 N_Y_c_360_n N_VGND_c_528_n 0.00249722f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_279 N_Y_c_360_n N_VGND_c_530_n 0.00249722f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_280 N_Y_c_361_n N_VGND_c_530_n 0.0106278f $X=4.21 $Y=0.445 $X2=0 $Y2=0
cc_281 N_Y_c_362_n N_VGND_c_530_n 0.00249722f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_282 N_Y_c_353_n N_VGND_c_532_n 0.0121037f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_283 N_Y_c_354_n N_VGND_c_532_n 0.0030627f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_284 N_Y_c_353_n N_VGND_c_533_n 0.00249722f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_285 N_Y_c_355_n N_VGND_c_533_n 0.0106278f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_286 N_Y_c_356_n N_VGND_c_533_n 0.00249722f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_287 N_Y_c_356_n N_VGND_c_534_n 0.00249722f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_288 N_Y_c_357_n N_VGND_c_534_n 0.0106278f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_289 N_Y_c_358_n N_VGND_c_534_n 0.00249722f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_290 N_Y_c_362_n N_VGND_c_535_n 0.00588215f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_291 N_Y_c_364_n N_VGND_c_535_n 0.0048643f $X=5.305 $Y=0.865 $X2=0 $Y2=0
cc_292 N_Y_M1001_d N_VGND_c_536_n 0.00264766f $X=1.49 $Y=0.235 $X2=0 $Y2=0
cc_293 N_Y_M1005_d N_VGND_c_536_n 0.00264766f $X=2.35 $Y=0.235 $X2=0 $Y2=0
cc_294 N_Y_M1009_d N_VGND_c_536_n 0.00264766f $X=3.21 $Y=0.235 $X2=0 $Y2=0
cc_295 N_Y_M1016_d N_VGND_c_536_n 0.00264766f $X=4.07 $Y=0.235 $X2=0 $Y2=0
cc_296 N_Y_c_353_n N_VGND_c_536_n 0.0256198f $X=1.535 $Y=0.78 $X2=0 $Y2=0
cc_297 N_Y_c_354_n N_VGND_c_536_n 0.00489372f $X=0.285 $Y=0.78 $X2=0 $Y2=0
cc_298 N_Y_c_355_n N_VGND_c_536_n 0.00712214f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_299 N_Y_c_356_n N_VGND_c_536_n 0.00929518f $X=2.395 $Y=0.78 $X2=0 $Y2=0
cc_300 N_Y_c_357_n N_VGND_c_536_n 0.00712214f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_301 N_Y_c_358_n N_VGND_c_536_n 0.00929518f $X=3.255 $Y=0.78 $X2=0 $Y2=0
cc_302 N_Y_c_359_n N_VGND_c_536_n 0.00712214f $X=3.35 $Y=0.445 $X2=0 $Y2=0
cc_303 N_Y_c_360_n N_VGND_c_536_n 0.00929518f $X=4.115 $Y=0.78 $X2=0 $Y2=0
cc_304 N_Y_c_361_n N_VGND_c_536_n 0.00712214f $X=4.21 $Y=0.445 $X2=0 $Y2=0
cc_305 N_Y_c_362_n N_VGND_c_536_n 0.0152079f $X=5.17 $Y=0.78 $X2=0 $Y2=0
cc_306 N_Y_c_364_n N_VGND_c_536_n 0.00777238f $X=5.305 $Y=0.865 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__a32o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_93_21# A1 a_346_47# VNB nshort w=650000u l=150000u
+  ad=2.86e+11p pd=2.18e+06u as=2.925e+11p ps=2.2e+06u
M1001 a_250_297# B2 a_93_21# VPB phighvt w=1e+06u l=150000u
+  ad=9.65e+11p pd=7.93e+06u as=2.8e+11p ps=2.56e+06u
M1002 a_584_47# B1 a_93_21# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=0p ps=0u
M1003 VGND B2 a_584_47# VNB nshort w=650000u l=150000u
+  ad=5.07e+11p pd=4.16e+06u as=0p ps=0u
M1004 VPWR a_93_21# X VPB phighvt w=1e+06u l=150000u
+  ad=9.35e+11p pd=5.87e+06u as=3.3e+11p ps=2.66e+06u
M1005 VGND a_93_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.145e+11p ps=1.96e+06u
M1006 a_93_21# B1 a_250_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A2 a_250_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_256_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=1.95e+11p pd=1.9e+06u as=0p ps=0u
M1009 a_346_47# A2 a_256_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_250_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_250_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__a32oi_4.pex.spice
* Created: Tue Sep  1 18:56:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A32OI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 34 50 51
c79 22 0 1.16491e-19 $X=1.73 $Y=0.995
r80 49 50 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.73 $Y2=1.16
r81 47 49 2.23839 $w=3.23e-07 $l=1.5e-08 $layer=POLY_cond $X=1.295 $Y=1.16
+ $X2=1.31 $Y2=1.16
r82 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.295
+ $Y=1.16 $X2=1.295 $Y2=1.16
r83 45 47 60.4365 $w=3.23e-07 $l=4.05e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.295 $Y2=1.16
r84 44 45 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.89 $Y2=1.16
r85 42 44 29.0991 $w=3.23e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r86 34 48 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.615 $Y=1.19
+ $X2=1.295 $Y2=1.19
r87 33 48 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=1.295 $Y2=1.19
r88 32 33 23.0489 $w=2.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.19
+ $X2=1.155 $Y2=1.19
r89 32 57 18.2888 $w=2.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.695 $Y=1.19
+ $X2=0.33 $Y2=1.19
r90 30 31 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=0.22 $Y=1.53
+ $X2=0.22 $Y2=1.87
r91 30 51 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=0.22 $Y=1.53
+ $X2=0.22 $Y2=1.305
r92 29 51 3.48622 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=0.22 $Y=1.19
+ $X2=0.22 $Y2=1.305
r93 29 57 3.33465 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.22 $Y=1.19 $X2=0.33
+ $Y2=1.19
r94 29 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r95 25 50 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r96 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r97 22 50 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r98 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r99 18 49 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r100 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r101 15 49 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r102 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r103 11 45 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r104 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r105 8 45 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r106 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r107 4 44 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r108 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r109 1 44 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r110 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 43
r78 41 43 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.35 $Y=1.16 $X2=3.41
+ $Y2=1.16
r79 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.16 $X2=3.35 $Y2=1.16
r80 39 41 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.35 $Y2=1.16
r81 37 39 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.99 $Y2=1.16
r82 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.16 $X2=2.67 $Y2=1.16
r83 35 37 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.57 $Y=1.16 $X2=2.67
+ $Y2=1.16
r84 33 35 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r85 30 42 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.455 $Y=1.16
+ $X2=3.35 $Y2=1.16
r86 29 42 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=3.35 $Y2=1.16
r87 29 38 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=2.67 $Y2=1.16
r88 25 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r89 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r90 22 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r92 18 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r93 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r94 15 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r95 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r96 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r97 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r98 8 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r99 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r100 4 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r101 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r102 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%A1 3 7 9 11 14 16 18 19 21 24 26 28 29 30 31
+ 32 49
c66 32 0 1.83742e-19 $X=5.315 $Y=1.19
c67 3 0 1.23524e-19 $X=3.85 $Y=1.985
r68 47 49 30.0377 $w=3.45e-07 $l=2.15e-07 $layer=POLY_cond $X=5.3 $Y=1.17
+ $X2=5.515 $Y2=1.17
r69 45 47 15.3681 $w=3.45e-07 $l=1.1e-07 $layer=POLY_cond $X=5.19 $Y=1.17
+ $X2=5.3 $Y2=1.17
r70 44 45 58.6783 $w=3.45e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.17
+ $X2=5.19 $Y2=1.17
r71 43 44 11.1768 $w=3.45e-07 $l=8e-08 $layer=POLY_cond $X=4.69 $Y=1.17 $X2=4.77
+ $Y2=1.17
r72 42 43 47.5014 $w=3.45e-07 $l=3.4e-07 $layer=POLY_cond $X=4.35 $Y=1.17
+ $X2=4.69 $Y2=1.17
r73 41 42 11.1768 $w=3.45e-07 $l=8e-08 $layer=POLY_cond $X=4.27 $Y=1.17 $X2=4.35
+ $Y2=1.17
r74 39 41 46.1043 $w=3.45e-07 $l=3.3e-07 $layer=POLY_cond $X=3.94 $Y=1.17
+ $X2=4.27 $Y2=1.17
r75 37 39 12.5739 $w=3.45e-07 $l=9e-08 $layer=POLY_cond $X=3.85 $Y=1.17 $X2=3.94
+ $Y2=1.17
r76 32 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.3
+ $Y=1.16 $X2=5.3 $Y2=1.16
r77 31 32 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=4.855 $Y=1.18
+ $X2=5.3 $Y2=1.18
r78 30 31 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=4.395 $Y=1.18
+ $X2=4.855 $Y2=1.18
r79 29 30 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=3.935 $Y=1.18
+ $X2=4.395 $Y2=1.18
r80 29 39 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.94
+ $Y=1.16 $X2=3.94 $Y2=1.16
r81 26 49 13.2725 $w=3.45e-07 $l=9.5e-08 $layer=POLY_cond $X=5.61 $Y=1.17
+ $X2=5.515 $Y2=1.17
r82 26 28 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.61 $Y=1.01 $X2=5.61
+ $Y2=0.56
r83 22 49 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.515 $Y=1.345
+ $X2=5.515 $Y2=1.17
r84 22 24 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.515 $Y=1.345
+ $X2=5.515 $Y2=1.985
r85 19 45 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.17
r86 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r87 16 44 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.17
r88 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r89 12 43 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.69 $Y=1.345
+ $X2=4.69 $Y2=1.17
r90 12 14 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.69 $Y=1.345
+ $X2=4.69 $Y2=1.985
r91 9 42 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.17
r92 9 11 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
r93 5 41 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.27 $Y=1.345
+ $X2=4.27 $Y2=1.17
r94 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.27 $Y=1.345 $X2=4.27
+ $Y2=1.985
r95 1 37 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.85 $Y=1.345
+ $X2=3.85 $Y2=1.17
r96 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.85 $Y=1.345 $X2=3.85
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32
c63 22 0 1.83742e-19 $X=7.43 $Y=1.01
r64 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.28
+ $Y=1.16 $X2=7.28 $Y2=1.16
r65 42 44 37.7217 $w=3.45e-07 $l=2.7e-07 $layer=POLY_cond $X=7.01 $Y=1.17
+ $X2=7.28 $Y2=1.17
r66 41 42 58.6783 $w=3.45e-07 $l=4.2e-07 $layer=POLY_cond $X=6.59 $Y=1.17
+ $X2=7.01 $Y2=1.17
r67 39 41 46.1043 $w=3.45e-07 $l=3.3e-07 $layer=POLY_cond $X=6.26 $Y=1.17
+ $X2=6.59 $Y2=1.17
r68 37 39 12.5739 $w=3.45e-07 $l=9e-08 $layer=POLY_cond $X=6.17 $Y=1.17 $X2=6.26
+ $Y2=1.17
r69 32 45 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=7.575 $Y=1.187
+ $X2=7.28 $Y2=1.187
r70 31 45 8.45125 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=1.187
+ $X2=7.28 $Y2=1.187
r71 30 31 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=6.655 $Y=1.187
+ $X2=7.115 $Y2=1.187
r72 29 30 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=6.195 $Y=1.187
+ $X2=6.655 $Y2=1.187
r73 29 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.26
+ $Y=1.16 $X2=6.26 $Y2=1.16
r74 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.43 $Y=1.345
+ $X2=7.43 $Y2=1.985
r75 22 25 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.43 $Y=1.17
+ $X2=7.43 $Y2=1.345
r76 22 44 20.9565 $w=3.45e-07 $l=1.5e-07 $layer=POLY_cond $X=7.43 $Y=1.17
+ $X2=7.28 $Y2=1.17
r77 22 24 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.43 $Y=1.01 $X2=7.43
+ $Y2=0.56
r78 18 42 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.01 $Y=1.345
+ $X2=7.01 $Y2=1.17
r79 18 20 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.01 $Y=1.345
+ $X2=7.01 $Y2=1.985
r80 15 42 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.01 $Y=0.995
+ $X2=7.01 $Y2=1.17
r81 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.01 $Y=0.995
+ $X2=7.01 $Y2=0.56
r82 11 41 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.59 $Y=1.345
+ $X2=6.59 $Y2=1.17
r83 11 13 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.59 $Y=1.345
+ $X2=6.59 $Y2=1.985
r84 8 41 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.59 $Y=0.995
+ $X2=6.59 $Y2=1.17
r85 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.59 $Y=0.995
+ $X2=6.59 $Y2=0.56
r86 4 37 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.17 $Y=1.345
+ $X2=6.17 $Y2=1.17
r87 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.17 $Y=1.345 $X2=6.17
+ $Y2=1.985
r88 1 37 22.2839 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.17 $Y=0.995
+ $X2=6.17 $Y2=1.17
r89 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.17 $Y=0.995 $X2=6.17
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 45 49 57
r70 45 47 28.3529 $w=3.23e-07 $l=1.9e-07 $layer=POLY_cond $X=9.63 $Y=1.16
+ $X2=9.82 $Y2=1.16
r71 44 45 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=9.21 $Y=1.16
+ $X2=9.63 $Y2=1.16
r72 43 44 62.6749 $w=3.23e-07 $l=4.2e-07 $layer=POLY_cond $X=8.79 $Y=1.16
+ $X2=9.21 $Y2=1.16
r73 41 43 49.2446 $w=3.23e-07 $l=3.3e-07 $layer=POLY_cond $X=8.46 $Y=1.16
+ $X2=8.79 $Y2=1.16
r74 39 41 13.4303 $w=3.23e-07 $l=9e-08 $layer=POLY_cond $X=8.37 $Y=1.16 $X2=8.46
+ $Y2=1.16
r75 33 57 3.64116 $w=1.8e-07 $l=1.02e-07 $layer=LI1_cond $X=9.895 $Y=1.177
+ $X2=9.895 $Y2=1.075
r76 33 49 3.21279 $w=2.05e-07 $l=9e-08 $layer=LI1_cond $X=9.895 $Y=1.177
+ $X2=9.805 $Y2=1.177
r77 33 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.82
+ $Y=1.16 $X2=9.82 $Y2=1.16
r78 32 57 13.8636 $w=1.78e-07 $l=2.25e-07 $layer=LI1_cond $X=9.895 $Y=0.85
+ $X2=9.895 $Y2=1.075
r79 31 49 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=9.435 $Y=1.177
+ $X2=9.805 $Y2=1.177
r80 30 31 24.8869 $w=2.03e-07 $l=4.6e-07 $layer=LI1_cond $X=8.975 $Y=1.177
+ $X2=9.435 $Y2=1.177
r81 29 30 27.8625 $w=2.03e-07 $l=5.15e-07 $layer=LI1_cond $X=8.46 $Y=1.177
+ $X2=8.975 $Y2=1.177
r82 29 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.46
+ $Y=1.16 $X2=8.46 $Y2=1.16
r83 25 45 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=1.325
+ $X2=9.63 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.63 $Y=1.325
+ $X2=9.63 $Y2=1.985
r85 22 45 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=0.995
+ $X2=9.63 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.63 $Y=0.995
+ $X2=9.63 $Y2=0.56
r87 18 44 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.21 $Y=1.325
+ $X2=9.21 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.21 $Y=1.325
+ $X2=9.21 $Y2=1.985
r89 15 44 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.21 $Y=0.995
+ $X2=9.21 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.21 $Y=0.995
+ $X2=9.21 $Y2=0.56
r91 11 43 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.79 $Y=1.325
+ $X2=8.79 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.79 $Y=1.325
+ $X2=8.79 $Y2=1.985
r93 8 43 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.79 $Y=0.995
+ $X2=8.79 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.79 $Y=0.995
+ $X2=8.79 $Y2=0.56
r95 4 39 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.37 $Y=1.325
+ $X2=8.37 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.37 $Y=1.325 $X2=8.37
+ $Y2=1.985
r97 1 39 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.37 $Y=0.995
+ $X2=8.37 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.37 $Y=0.995 $X2=8.37
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%A_27_297# 1 2 3 4 5 6 7 8 9 10 11 34 45 46
+ 47 50 52 56 58 62 64 68 70 74 76 80 84 85 86 87 88
r105 78 80 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.84 $Y=1.745
+ $X2=9.84 $Y2=1.96
r106 77 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.085 $Y=1.66 $X2=9
+ $Y2=1.66
r107 76 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.755 $Y=1.66
+ $X2=9.84 $Y2=1.745
r108 76 77 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.755 $Y=1.66
+ $X2=9.085 $Y2=1.66
r109 72 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9 $Y=1.745 $X2=9
+ $Y2=1.66
r110 72 74 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9 $Y=1.745 $X2=9
+ $Y2=1.96
r111 71 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=1.66
+ $X2=7.64 $Y2=1.66
r112 70 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.915 $Y=1.66 $X2=9
+ $Y2=1.66
r113 70 71 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=8.915 $Y=1.66
+ $X2=7.725 $Y2=1.66
r114 66 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.64 $Y=1.745
+ $X2=7.64 $Y2=1.66
r115 66 68 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.64 $Y=1.745
+ $X2=7.64 $Y2=1.96
r116 65 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.885 $Y=1.66
+ $X2=6.8 $Y2=1.66
r117 64 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=1.66
+ $X2=7.64 $Y2=1.66
r118 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.555 $Y=1.66
+ $X2=6.885 $Y2=1.66
r119 60 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=1.745 $X2=6.8
+ $Y2=1.66
r120 60 62 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.8 $Y=1.745
+ $X2=6.8 $Y2=1.96
r121 59 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.81 $Y=1.66
+ $X2=5.725 $Y2=1.66
r122 58 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=1.66
+ $X2=6.8 $Y2=1.66
r123 58 59 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.715 $Y=1.66
+ $X2=5.81 $Y2=1.66
r124 54 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.725 $Y=1.745
+ $X2=5.725 $Y2=1.66
r125 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.725 $Y=1.745
+ $X2=5.725 $Y2=1.96
r126 53 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=1.66
+ $X2=4.48 $Y2=1.66
r127 52 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=1.66
+ $X2=5.725 $Y2=1.66
r128 52 53 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=5.64 $Y=1.66
+ $X2=4.565 $Y2=1.66
r129 48 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=1.745
+ $X2=4.48 $Y2=1.66
r130 48 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.48 $Y=1.745
+ $X2=4.48 $Y2=1.96
r131 46 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.395 $Y=1.66
+ $X2=4.48 $Y2=1.66
r132 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.395 $Y=1.66
+ $X2=3.705 $Y2=1.66
r133 45 83 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.255
+ $X2=3.62 $Y2=2.34
r134 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.62 $Y=1.745
+ $X2=3.705 $Y2=1.66
r135 44 45 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.62 $Y=1.745
+ $X2=3.62 $Y2=2.255
r136 41 43 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.94 $Y=2.34
+ $X2=2.78 $Y2=2.34
r137 39 41 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=2.34
+ $X2=1.94 $Y2=2.34
r138 36 39 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.26 $Y=2.34
+ $X2=1.1 $Y2=2.34
r139 34 83 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.34
+ $X2=3.62 $Y2=2.34
r140 34 43 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.535 $Y=2.34
+ $X2=2.78 $Y2=2.34
r141 11 80 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=9.705
+ $Y=1.485 $X2=9.84 $Y2=1.96
r142 10 74 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.865
+ $Y=1.485 $X2=9 $Y2=1.96
r143 9 68 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.505
+ $Y=1.485 $X2=7.64 $Y2=1.96
r144 8 62 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.665
+ $Y=1.485 $X2=6.8 $Y2=1.96
r145 7 56 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.59
+ $Y=1.485 $X2=5.725 $Y2=1.96
r146 6 50 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.48 $Y2=1.96
r147 5 83 600 $w=1.7e-07 $l=8.39792e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2.26
r148 4 43 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2.34
r149 3 41 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.34
r150 2 39 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r151 1 36 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%Y 1 2 3 4 5 6 7 8 27 31 33 41 43 48 50 54 55
+ 56 57 66 70 72
c103 54 0 1.23524e-19 $X=3.2 $Y=1.66
c104 33 0 1.16491e-19 $X=2.28 $Y=0.805
r105 70 74 1.32974 $w=3.88e-07 $l=4.5e-08 $layer=LI1_cond $X=2.17 $Y=1.53
+ $X2=2.17 $Y2=1.575
r106 63 66 0.147749 $w=3.88e-07 $l=5e-09 $layer=LI1_cond $X=2.17 $Y=1.185
+ $X2=2.17 $Y2=1.19
r107 57 76 4.56684 $w=5.48e-07 $l=2.1e-07 $layer=LI1_cond $X=2.25 $Y=1.87
+ $X2=2.25 $Y2=1.66
r108 56 76 1.41355 $w=5.48e-07 $l=6.5e-08 $layer=LI1_cond $X=2.25 $Y=1.595
+ $X2=2.25 $Y2=1.66
r109 56 74 1.46339 $w=5.48e-07 $l=2e-08 $layer=LI1_cond $X=2.25 $Y=1.595
+ $X2=2.25 $Y2=1.575
r110 56 70 0.590996 $w=3.88e-07 $l=2e-08 $layer=LI1_cond $X=2.17 $Y=1.51
+ $X2=2.17 $Y2=1.53
r111 55 63 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=2.17 $Y=1.145
+ $X2=2.17 $Y2=1.185
r112 55 72 8.31213 $w=3.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.17 $Y=1.145
+ $X2=2.17 $Y2=0.99
r113 55 56 8.27395 $w=3.88e-07 $l=2.8e-07 $layer=LI1_cond $X=2.17 $Y=1.23
+ $X2=2.17 $Y2=1.51
r114 55 66 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=2.17 $Y=1.23 $X2=2.17
+ $Y2=1.19
r115 44 76 7.75927 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.525 $Y=1.66
+ $X2=2.25 $Y2=1.66
r116 43 54 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=1.66
+ $X2=3.2 $Y2=1.66
r117 43 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.035 $Y=1.66
+ $X2=2.525 $Y2=1.66
r118 39 41 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.56 $Y=0.72
+ $X2=5.4 $Y2=0.72
r119 37 39 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.2 $Y=0.72
+ $X2=4.56 $Y2=0.72
r120 35 52 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=0.72
+ $X2=2.28 $Y2=0.72
r121 35 37 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.365 $Y=0.72
+ $X2=3.2 $Y2=0.72
r122 33 52 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.805
+ $X2=2.28 $Y2=0.72
r123 33 72 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.28 $Y=0.805
+ $X2=2.28 $Y2=0.99
r124 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.66
+ $X2=1.52 $Y2=1.66
r125 31 76 7.75927 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=1.975 $Y=1.66
+ $X2=2.25 $Y2=1.66
r126 31 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.975 $Y=1.66
+ $X2=1.685 $Y2=1.66
r127 28 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.66
+ $X2=0.68 $Y2=1.66
r128 27 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.66
+ $X2=1.52 $Y2=1.66
r129 27 28 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.66
+ $X2=0.845 $Y2=1.66
r130 8 54 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.66
r131 7 76 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.66
r132 6 50 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r133 5 48 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r134 4 41 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.72
r135 3 39 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.72
r136 2 37 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.72
r137 1 52 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%VPWR 1 2 3 4 5 6 21 23 27 31 33 37 41 45 47
+ 48 49 51 60 65 72 73 76 79 84 87 90
r125 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r126 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r127 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r128 80 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r129 79 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r130 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r131 77 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r132 76 77 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r133 73 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r134 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r135 70 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.585 $Y=2.72
+ $X2=9.42 $Y2=2.72
r136 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.585 $Y=2.72
+ $X2=9.89 $Y2=2.72
r137 69 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r138 69 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r139 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r140 66 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.745 $Y=2.72
+ $X2=8.58 $Y2=2.72
r141 66 68 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.745 $Y=2.72
+ $X2=8.97 $Y2=2.72
r142 65 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=2.72
+ $X2=9.42 $Y2=2.72
r143 65 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.255 $Y=2.72
+ $X2=8.97 $Y2=2.72
r144 64 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r145 64 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.13 $Y2=2.72
r146 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r147 61 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.385 $Y=2.72
+ $X2=7.22 $Y2=2.72
r148 61 63 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.385 $Y=2.72
+ $X2=8.05 $Y2=2.72
r149 60 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.415 $Y=2.72
+ $X2=8.58 $Y2=2.72
r150 60 63 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.415 $Y=2.72
+ $X2=8.05 $Y2=2.72
r151 59 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r152 59 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.29 $Y2=2.72
r153 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r154 56 79 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.44 $Y=2.72
+ $X2=5.105 $Y2=2.72
r155 56 58 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.44 $Y=2.72
+ $X2=6.21 $Y2=2.72
r156 51 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=4.06 $Y2=2.72
r157 51 53 239.107 $w=1.68e-07 $l=3.665e-06 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=0.23 $Y2=2.72
r158 49 77 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.91 $Y2=2.72
r159 49 53 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r160 47 58 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.215 $Y=2.72
+ $X2=6.21 $Y2=2.72
r161 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.215 $Y=2.72
+ $X2=6.38 $Y2=2.72
r162 43 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.42 $Y=2.635
+ $X2=9.42 $Y2=2.72
r163 43 45 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=9.42 $Y=2.635
+ $X2=9.42 $Y2=2
r164 39 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.58 $Y=2.635
+ $X2=8.58 $Y2=2.72
r165 39 41 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=8.58 $Y=2.635
+ $X2=8.58 $Y2=2
r166 35 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.635
+ $X2=7.22 $Y2=2.72
r167 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.22 $Y=2.635
+ $X2=7.22 $Y2=2.34
r168 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=6.38 $Y2=2.72
r169 33 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=2.72
+ $X2=7.22 $Y2=2.72
r170 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.055 $Y=2.72
+ $X2=6.545 $Y2=2.72
r171 29 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=2.635
+ $X2=6.38 $Y2=2.72
r172 29 31 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.38 $Y=2.635
+ $X2=6.38 $Y2=2
r173 25 79 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=2.635
+ $X2=5.105 $Y2=2.72
r174 25 27 11.336 $w=6.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.105 $Y=2.635
+ $X2=5.105 $Y2=2
r175 24 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.06 $Y2=2.72
r176 23 79 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.77 $Y=2.72
+ $X2=5.105 $Y2=2.72
r177 23 24 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.77 $Y=2.72
+ $X2=4.225 $Y2=2.72
r178 19 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=2.635
+ $X2=4.06 $Y2=2.72
r179 19 21 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.06 $Y=2.635
+ $X2=4.06 $Y2=2
r180 6 45 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.285
+ $Y=1.485 $X2=9.42 $Y2=2
r181 5 41 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.445
+ $Y=1.485 $X2=8.58 $Y2=2
r182 4 37 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.085
+ $Y=1.485 $X2=7.22 $Y2=2.34
r183 3 31 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.245
+ $Y=1.485 $X2=6.38 $Y2=2
r184 2 27 150 $w=1.7e-07 $l=7.2655e-07 $layer=licon1_PDIFF $count=4 $X=4.765
+ $Y=1.485 $X2=5.275 $Y2=2
r185 1 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.485 $X2=4.06 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 28 34 36
r51 32 34 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.78 $Y=0.38
+ $X2=3.62 $Y2=0.38
r52 30 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.38
+ $X2=1.94 $Y2=0.38
r53 30 32 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.025 $Y=0.38
+ $X2=2.78 $Y2=0.38
r54 28 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.465
+ $X2=1.94 $Y2=0.38
r55 28 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.94 $Y=0.465
+ $X2=1.94 $Y2=0.635
r56 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.72 $X2=1.1
+ $Y2=0.72
r57 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.855 $Y=0.72
+ $X2=1.94 $Y2=0.635
r58 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.855 $Y=0.72
+ $X2=1.185 $Y2=0.72
r59 22 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.635 $X2=1.1
+ $Y2=0.72
r60 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.1 $Y=0.635
+ $X2=1.1 $Y2=0.42
r61 20 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.72 $X2=1.1
+ $Y2=0.72
r62 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.72
+ $X2=0.345 $Y2=0.72
r63 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r64 16 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.42
r65 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.38
r66 4 32 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.38
r67 3 38 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.46
r68 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.42
r69 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%VGND 1 2 3 4 5 18 22 24 28 32 34 36 38 40 45
+ 50 55 61 64 67 70 74
r132 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r133 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r134 67 68 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r135 65 68 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=8.05
+ $Y2=0
r136 64 65 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r137 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r138 59 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=9.89
+ $Y2=0
r139 59 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=8.97
+ $Y2=0
r140 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r141 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.165 $Y=0 $X2=9
+ $Y2=0
r142 56 58 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.165 $Y=0
+ $X2=9.43 $Y2=0
r143 55 73 4.88166 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=9.685 $Y=0
+ $X2=9.902 $Y2=0
r144 55 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.685 $Y=0
+ $X2=9.43 $Y2=0
r145 54 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.97
+ $Y2=0
r146 54 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.05
+ $Y2=0
r147 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r148 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.325 $Y=0 $X2=8.16
+ $Y2=0
r149 51 53 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.51 $Y2=0
r150 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.835 $Y=0 $X2=9
+ $Y2=0
r151 50 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.835 $Y=0
+ $X2=8.51 $Y2=0
r152 49 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r153 49 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r154 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r155 46 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r156 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r157 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.52
+ $Y2=0
r158 45 48 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.15 $Y2=0
r159 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r160 40 42 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r161 38 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r162 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r163 34 73 2.96949 $w=3.4e-07 $l=1.05924e-07 $layer=LI1_cond $X=9.855 $Y=0.085
+ $X2=9.902 $Y2=0
r164 34 36 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=9.855 $Y=0.085
+ $X2=9.855 $Y2=0.38
r165 30 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9 $Y=0.085 $X2=9
+ $Y2=0
r166 30 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9 $Y=0.085 $X2=9
+ $Y2=0.38
r167 26 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.16 $Y=0.085
+ $X2=8.16 $Y2=0
r168 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.16 $Y=0.085
+ $X2=8.16 $Y2=0.38
r169 25 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0 $X2=1.52
+ $Y2=0
r170 24 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=8.16
+ $Y2=0
r171 24 25 411.668 $w=1.68e-07 $l=6.31e-06 $layer=LI1_cond $X=7.995 $Y=0
+ $X2=1.685 $Y2=0
r172 20 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0
r173 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.52 $Y=0.085
+ $X2=1.52 $Y2=0.38
r174 16 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r175 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r176 5 36 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=9.705
+ $Y=0.235 $X2=9.85 $Y2=0.38
r177 4 32 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.865
+ $Y=0.235 $X2=9 $Y2=0.38
r178 3 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=8.035
+ $Y=0.235 $X2=8.16 $Y2=0.38
r179 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.38
r180 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%A_803_47# 1 2 3 4 5 26
r29 24 26 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.8 $Y=0.38 $X2=7.64
+ $Y2=0.38
r30 22 24 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.82 $Y=0.38 $X2=6.8
+ $Y2=0.38
r31 20 22 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.98 $Y=0.38
+ $X2=5.82 $Y2=0.38
r32 17 20 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.14 $Y=0.38
+ $X2=4.98 $Y2=0.38
r33 5 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.505
+ $Y=0.235 $X2=7.64 $Y2=0.38
r34 4 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.665
+ $Y=0.235 $X2=6.8 $Y2=0.38
r35 3 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.38
r36 2 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.38
r37 1 17 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A32OI_4%A_1249_47# 1 2 3 4 13 21 23 27 29
r39 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.42 $Y=0.635
+ $X2=9.42 $Y2=0.42
r40 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=0.72
+ $X2=8.58 $Y2=0.72
r41 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.335 $Y=0.72
+ $X2=9.42 $Y2=0.635
r42 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.335 $Y=0.72
+ $X2=8.665 $Y2=0.72
r43 19 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.58 $Y=0.635
+ $X2=8.58 $Y2=0.72
r44 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.58 $Y=0.635
+ $X2=8.58 $Y2=0.42
r45 15 18 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.38 $Y=0.72
+ $X2=7.22 $Y2=0.72
r46 13 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.495 $Y=0.72
+ $X2=8.58 $Y2=0.72
r47 13 18 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=8.495 $Y=0.72
+ $X2=7.22 $Y2=0.72
r48 4 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.285
+ $Y=0.235 $X2=9.42 $Y2=0.42
r49 3 21 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.445
+ $Y=0.235 $X2=8.58 $Y2=0.42
r50 2 18 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=7.085
+ $Y=0.235 $X2=7.22 $Y2=0.72
r51 1 15 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=6.245
+ $Y=0.235 $X2=6.38 $Y2=0.72
.ends


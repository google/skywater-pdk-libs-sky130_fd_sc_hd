* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_1.spice.SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1.pxi
* Created: Thu Aug 27 14:23:21 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%A_75_212# N_A_75_212#_M1001_d
+ N_A_75_212#_M1002_d N_A_75_212#_M1003_g N_A_75_212#_M1000_g N_A_75_212#_c_40_n
+ N_A_75_212#_c_35_n N_A_75_212#_c_63_p N_A_75_212#_c_41_n N_A_75_212#_c_65_p
+ N_A_75_212#_c_98_p N_A_75_212#_c_57_p N_A_75_212#_c_36_n N_A_75_212#_c_37_n
+ N_A_75_212#_c_38_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%A_75_212#
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%A N_A_c_107_n N_A_M1001_g N_A_M1002_g
+ N_A_c_108_n N_A_c_111_n N_A_c_112_n A
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%X N_X_M1003_s N_X_M1000_s N_X_c_139_n
+ N_X_c_142_n N_X_c_140_n X X X PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%X
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%KAPWR N_KAPWR_M1000_d N_KAPWR_c_167_n
+ N_KAPWR_c_168_n KAPWR N_KAPWR_c_176_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%VGND N_VGND_M1003_d N_VGND_c_194_n
+ VGND N_VGND_c_196_n N_VGND_c_197_n N_VGND_c_198_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%VPWR VPWR N_VPWR_c_222_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_1%VPWR
cc_1 VNB N_A_75_212#_M1003_g 0.0289893f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_2 VNB N_A_75_212#_c_35_n 0.00771329f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=0.72
cc_3 VNB N_A_75_212#_c_36_n 0.00163395f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.225
cc_4 VNB N_A_75_212#_c_37_n 0.0191693f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.225
cc_5 VNB N_A_75_212#_c_38_n 0.0021693f $X=-0.19 $Y=-0.24 $X2=0.567 $Y2=1.06
cc_6 VNB N_A_c_107_n 0.0179813f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=0.235
cc_7 VNB N_A_c_108_n 0.048966f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.06
cc_8 VNB A 0.0163436f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.39
cc_9 VNB N_X_c_139_n 0.00847523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_X_c_140_n 0.0254822f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.09
cc_11 VNB X 0.0145716f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.09
cc_12 VNB N_VGND_c_194_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB VGND 0.10585f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_14 VNB N_VGND_c_196_n 0.0153759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_197_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.39
cc_16 VNB N_VGND_c_198_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.62
cc_17 VNB VPWR 0.0609879f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=0.235
cc_18 VPB N_A_75_212#_M1000_g 0.0291084f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.09
cc_19 VPB N_A_75_212#_c_40_n 0.00135348f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.535
cc_20 VPB N_A_75_212#_c_41_n 0.0120187f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.62
cc_21 VPB N_A_75_212#_c_36_n 6.91362e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.225
cc_22 VPB N_A_75_212#_c_37_n 0.00918419f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.225
cc_23 VPB N_A_c_108_n 0.00829456f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.06
cc_24 VPB N_A_c_111_n 0.0136585f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.495
cc_25 VPB N_A_c_112_n 0.0275872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB A 0.00627368f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.39
cc_27 VPB N_X_c_142_n 0.0110375f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.39
cc_28 VPB N_X_c_140_n 0.0119115f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.09
cc_29 VPB X 0.0250115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_KAPWR_c_167_n 0.0107845f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.495
cc_31 VPB N_KAPWR_c_168_n 0.00876329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB VPWR 0.0420658f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=0.235
cc_33 VPB N_VPWR_c_222_n 0.0408481f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.495
cc_34 N_A_75_212#_M1003_g N_A_c_107_n 0.0209393f $X=0.47 $Y=0.495 $X2=-0.19
+ $Y2=-0.24
cc_35 N_A_75_212#_c_35_n N_A_c_107_n 0.015302f $X=1.035 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_36 N_A_75_212#_c_38_n N_A_c_107_n 0.00318324f $X=0.567 $Y=1.06 $X2=-0.19
+ $Y2=-0.24
cc_37 N_A_75_212#_M1003_g N_A_c_108_n 0.003841f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_38 N_A_75_212#_c_35_n N_A_c_108_n 0.00234783f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_39 N_A_75_212#_c_41_n N_A_c_108_n 0.00154723f $X=1.035 $Y=1.62 $X2=0 $Y2=0
cc_40 N_A_75_212#_c_37_n N_A_c_108_n 0.0193066f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_41 N_A_75_212#_c_38_n N_A_c_108_n 0.00324151f $X=0.567 $Y=1.06 $X2=0 $Y2=0
cc_42 N_A_75_212#_M1000_g N_A_c_111_n 0.00368068f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_43 N_A_75_212#_c_36_n N_A_c_111_n 0.00324151f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_44 N_A_75_212#_M1000_g N_A_c_112_n 0.0173618f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_45 N_A_75_212#_c_40_n N_A_c_112_n 7.5643e-19 $X=0.625 $Y=1.535 $X2=0 $Y2=0
cc_46 N_A_75_212#_c_41_n N_A_c_112_n 0.0161707f $X=1.035 $Y=1.62 $X2=0 $Y2=0
cc_47 N_A_75_212#_c_57_p N_A_c_112_n 0.00140798f $X=1.12 $Y=1.96 $X2=0 $Y2=0
cc_48 N_A_75_212#_c_35_n A 0.0207534f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_49 N_A_75_212#_c_41_n A 0.0208772f $X=1.035 $Y=1.62 $X2=0 $Y2=0
cc_50 N_A_75_212#_c_37_n A 2.94551e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_51 N_A_75_212#_c_38_n A 0.0224427f $X=0.567 $Y=1.06 $X2=0 $Y2=0
cc_52 N_A_75_212#_M1003_g N_X_c_139_n 0.00222896f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_53 N_A_75_212#_c_63_p N_X_c_139_n 0.00484499f $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_54 N_A_75_212#_M1000_g N_X_c_142_n 0.00373896f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_55 N_A_75_212#_c_65_p N_X_c_142_n 0.0108006f $X=0.71 $Y=1.62 $X2=0 $Y2=0
cc_56 N_A_75_212#_M1003_g N_X_c_140_n 0.00632981f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_57 N_A_75_212#_M1000_g N_X_c_140_n 0.00357773f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_58 N_A_75_212#_c_40_n N_X_c_140_n 0.0070136f $X=0.625 $Y=1.535 $X2=0 $Y2=0
cc_59 N_A_75_212#_c_63_p N_X_c_140_n 0.00240564f $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_60 N_A_75_212#_c_65_p N_X_c_140_n 0.00132477f $X=0.71 $Y=1.62 $X2=0 $Y2=0
cc_61 N_A_75_212#_c_36_n N_X_c_140_n 0.0245251f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_62 N_A_75_212#_c_37_n N_X_c_140_n 0.00753248f $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_63 N_A_75_212#_c_38_n N_X_c_140_n 0.0123683f $X=0.567 $Y=1.06 $X2=0 $Y2=0
cc_64 N_A_75_212#_c_41_n N_KAPWR_M1000_d 6.82533e-19 $X=1.035 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_75_212#_c_65_p N_KAPWR_M1000_d 0.00114523f $X=0.71 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_75_212#_M1002_d N_KAPWR_c_167_n 0.00258808f $X=0.985 $Y=1.695 $X2=0
+ $Y2=0
cc_67 N_A_75_212#_c_41_n N_KAPWR_c_167_n 0.00624624f $X=1.035 $Y=1.62 $X2=0
+ $Y2=0
cc_68 N_A_75_212#_c_65_p N_KAPWR_c_167_n 8.55177e-19 $X=0.71 $Y=1.62 $X2=0 $Y2=0
cc_69 N_A_75_212#_c_57_p N_KAPWR_c_167_n 0.0214905f $X=1.12 $Y=1.96 $X2=0 $Y2=0
cc_70 N_A_75_212#_M1000_g N_KAPWR_c_168_n 0.00629033f $X=0.47 $Y=2.09 $X2=0
+ $Y2=0
cc_71 N_A_75_212#_M1000_g N_KAPWR_c_176_n 0.00582352f $X=0.47 $Y=2.09 $X2=0
+ $Y2=0
cc_72 N_A_75_212#_c_41_n N_KAPWR_c_176_n 0.00649838f $X=1.035 $Y=1.62 $X2=0
+ $Y2=0
cc_73 N_A_75_212#_c_65_p N_KAPWR_c_176_n 0.00943796f $X=0.71 $Y=1.62 $X2=0 $Y2=0
cc_74 N_A_75_212#_c_57_p N_KAPWR_c_176_n 0.0234331f $X=1.12 $Y=1.96 $X2=0 $Y2=0
cc_75 N_A_75_212#_c_36_n N_KAPWR_c_176_n 4.70471e-19 $X=0.51 $Y=1.225 $X2=0
+ $Y2=0
cc_76 N_A_75_212#_c_37_n N_KAPWR_c_176_n 3.03855e-19 $X=0.51 $Y=1.225 $X2=0
+ $Y2=0
cc_77 N_A_75_212#_c_35_n N_VGND_M1003_d 6.85198e-19 $X=1.035 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_75_212#_c_63_p N_VGND_M1003_d 0.00114971f $X=0.71 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_75_212#_M1003_g N_VGND_c_194_n 0.00801602f $X=0.47 $Y=0.495 $X2=0
+ $Y2=0
cc_80 N_A_75_212#_c_35_n N_VGND_c_194_n 0.00647139f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_81 N_A_75_212#_c_63_p N_VGND_c_194_n 0.00945604f $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_82 N_A_75_212#_c_36_n N_VGND_c_194_n 3.89729e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_83 N_A_75_212#_c_37_n N_VGND_c_194_n 2.51407e-19 $X=0.51 $Y=1.225 $X2=0 $Y2=0
cc_84 N_A_75_212#_M1001_d VGND 0.00369894f $X=0.985 $Y=0.235 $X2=0 $Y2=0
cc_85 N_A_75_212#_M1003_g VGND 0.00957284f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_86 N_A_75_212#_c_35_n VGND 0.0050992f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_87 N_A_75_212#_c_63_p VGND 8.54935e-19 $X=0.71 $Y=0.72 $X2=0 $Y2=0
cc_88 N_A_75_212#_c_98_p VGND 0.00643448f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_75_212#_M1003_g N_VGND_c_196_n 0.00505556f $X=0.47 $Y=0.495 $X2=0
+ $Y2=0
cc_90 N_A_75_212#_c_35_n N_VGND_c_197_n 0.00260015f $X=1.035 $Y=0.72 $X2=0 $Y2=0
cc_91 N_A_75_212#_c_98_p N_VGND_c_197_n 0.01143f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_75_212#_M1002_d VPWR 0.00143721f $X=0.985 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_93 N_A_75_212#_M1000_g VPWR 0.00612094f $X=0.47 $Y=2.09 $X2=-0.19 $Y2=-0.24
cc_94 N_A_75_212#_c_57_p VPWR 0.00155926f $X=1.12 $Y=1.96 $X2=-0.19 $Y2=-0.24
cc_95 N_A_75_212#_M1000_g N_VPWR_c_222_n 0.0055654f $X=0.47 $Y=2.09 $X2=0 $Y2=0
cc_96 N_A_75_212#_c_57_p N_VPWR_c_222_n 0.0116048f $X=1.12 $Y=1.96 $X2=0 $Y2=0
cc_97 N_A_c_112_n N_KAPWR_c_167_n 0.00242504f $X=0.925 $Y=1.62 $X2=0 $Y2=0
cc_98 N_A_c_112_n N_KAPWR_c_176_n 0.00588034f $X=0.925 $Y=1.62 $X2=0 $Y2=0
cc_99 N_A_c_107_n N_VGND_c_194_n 0.00787353f $X=0.91 $Y=0.83 $X2=0 $Y2=0
cc_100 N_A_c_107_n VGND 0.00526324f $X=0.91 $Y=0.83 $X2=0 $Y2=0
cc_101 N_A_c_107_n N_VGND_c_197_n 0.00367706f $X=0.91 $Y=0.83 $X2=0 $Y2=0
cc_102 N_A_c_112_n VPWR 0.00612094f $X=0.925 $Y=1.62 $X2=-0.19 $Y2=-0.24
cc_103 N_A_c_112_n N_VPWR_c_222_n 0.0055654f $X=0.925 $Y=1.62 $X2=0 $Y2=0
cc_104 X N_KAPWR_c_167_n 4.3931e-19 $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_105 N_X_M1000_s N_KAPWR_c_168_n 0.00168005f $X=0.135 $Y=1.695 $X2=0 $Y2=0
cc_106 X N_KAPWR_c_168_n 0.0285517f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_107 X N_KAPWR_c_176_n 0.0247379f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_108 N_X_M1003_s VGND 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_109 X VGND 0.00990988f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_110 X N_VGND_c_196_n 0.0178762f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_111 N_X_M1000_s VPWR 0.00123164f $X=0.135 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_112 X VPWR 0.0024874f $X=0.145 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_113 X N_VPWR_c_222_n 0.0183559f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_114 N_KAPWR_M1000_d VPWR 0.0011753f $X=0.545 $Y=1.695 $X2=-0.19 $Y2=1.305
cc_115 N_KAPWR_c_168_n VPWR 0.127537f $X=0.55 $Y=2.21 $X2=-0.19 $Y2=1.305
cc_116 N_KAPWR_c_176_n VPWR 0.00292242f $X=0.69 $Y=1.96 $X2=-0.19 $Y2=1.305
cc_117 N_KAPWR_c_167_n N_VPWR_c_222_n 0.00159238f $X=0.695 $Y=2.21 $X2=0 $Y2=0
cc_118 N_KAPWR_c_168_n N_VPWR_c_222_n 0.00135211f $X=0.55 $Y=2.21 $X2=0 $Y2=0
cc_119 N_KAPWR_c_176_n N_VPWR_c_222_n 0.0187938f $X=0.69 $Y=1.96 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__or3_1.spice
* Created: Thu Aug 27 14:43:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or3_1.spice.pex"
.subckt sky130_fd_sc_hd__or3_1  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_C_M1004_g N_A_29_53#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_A_29_53#_M1000_d N_B_M1000_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_29_53#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0567 PD=0.777196 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_29_53#_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.123773 PD=1.86 PS=1.2028 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 A_111_297# N_C_M1003_g N_A_29_53#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 A_183_297# N_B_M1001_g A_111_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.0693
+ AS=0.0441 PD=0.75 PS=0.63 NRD=51.5943 NRS=23.443 M=1 R=2.8 SA=75000.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_183_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0876972 AS=0.0693 PD=0.792676 PS=0.75 NRD=72.1217 NRS=51.5943 M=1 R=2.8
+ SA=75001 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_29_53#_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.208803 PD=2.56 PS=1.88732 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
c_55 VPB 0 2.26204e-19 $X=0.14 $Y=2.635
*
.include "sky130_fd_sc_hd__or3_1.spice.SKY130_FD_SC_HD__OR3_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a21o_4.pxi.spice
* Created: Thu Aug 27 14:01:08 2020
* 
x_PM_SKY130_FD_SC_HD__A21O_4%A_84_21# N_A_84_21#_M1007_d N_A_84_21#_M1006_d
+ N_A_84_21#_M1017_s N_A_84_21#_c_82_n N_A_84_21#_M1001_g N_A_84_21#_M1002_g
+ N_A_84_21#_c_83_n N_A_84_21#_M1003_g N_A_84_21#_M1004_g N_A_84_21#_c_84_n
+ N_A_84_21#_M1005_g N_A_84_21#_M1011_g N_A_84_21#_c_85_n N_A_84_21#_M1014_g
+ N_A_84_21#_M1015_g N_A_84_21#_c_86_n N_A_84_21#_c_87_n N_A_84_21#_c_88_n
+ N_A_84_21#_c_98_p N_A_84_21#_c_150_p N_A_84_21#_c_186_p N_A_84_21#_c_89_n
+ N_A_84_21#_c_102_p N_A_84_21#_c_120_p PM_SKY130_FD_SC_HD__A21O_4%A_84_21#
x_PM_SKY130_FD_SC_HD__A21O_4%B1 N_B1_c_207_n N_B1_M1007_g N_B1_M1017_g
+ N_B1_c_208_n N_B1_M1010_g N_B1_M1019_g B1 N_B1_c_210_n
+ PM_SKY130_FD_SC_HD__A21O_4%B1
x_PM_SKY130_FD_SC_HD__A21O_4%A2 N_A2_M1012_g N_A2_M1009_g N_A2_M1016_g
+ N_A2_M1013_g N_A2_c_256_n N_A2_c_271_n N_A2_c_303_p N_A2_c_257_n N_A2_c_258_n
+ N_A2_c_259_n N_A2_c_260_n A2 N_A2_c_262_n N_A2_c_263_n N_A2_c_306_p
+ PM_SKY130_FD_SC_HD__A21O_4%A2
x_PM_SKY130_FD_SC_HD__A21O_4%A1 N_A1_c_341_n N_A1_M1006_g N_A1_M1000_g
+ N_A1_c_342_n N_A1_M1008_g N_A1_M1018_g A1 N_A1_c_344_n
+ PM_SKY130_FD_SC_HD__A21O_4%A1
x_PM_SKY130_FD_SC_HD__A21O_4%VPWR N_VPWR_M1002_s N_VPWR_M1004_s N_VPWR_M1015_s
+ N_VPWR_M1012_d N_VPWR_M1018_s N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n
+ N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_394_n
+ N_VPWR_c_395_n N_VPWR_c_396_n VPWR N_VPWR_c_397_n N_VPWR_c_398_n
+ N_VPWR_c_399_n N_VPWR_c_386_n N_VPWR_c_401_n N_VPWR_c_402_n
+ PM_SKY130_FD_SC_HD__A21O_4%VPWR
x_PM_SKY130_FD_SC_HD__A21O_4%X N_X_M1001_s N_X_M1005_s N_X_M1002_d N_X_M1011_d
+ N_X_c_508_n N_X_c_485_n N_X_c_486_n N_X_c_492_n N_X_c_496_n N_X_c_499_n X X
+ PM_SKY130_FD_SC_HD__A21O_4%X
x_PM_SKY130_FD_SC_HD__A21O_4%A_483_297# N_A_483_297#_M1017_d
+ N_A_483_297#_M1019_d N_A_483_297#_M1000_d N_A_483_297#_M1013_s
+ N_A_483_297#_c_536_n N_A_483_297#_c_531_n N_A_483_297#_c_570_n
+ N_A_483_297#_c_528_n N_A_483_297#_c_546_n N_A_483_297#_c_578_n
+ N_A_483_297#_c_550_n N_A_483_297#_c_529_n N_A_483_297#_c_557_n
+ N_A_483_297#_c_530_n PM_SKY130_FD_SC_HD__A21O_4%A_483_297#
x_PM_SKY130_FD_SC_HD__A21O_4%VGND N_VGND_M1001_d N_VGND_M1003_d N_VGND_M1014_d
+ N_VGND_M1010_s N_VGND_M1016_s N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n
+ N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n VGND
+ N_VGND_c_596_n N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n N_VGND_c_600_n
+ N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n PM_SKY130_FD_SC_HD__A21O_4%VGND
cc_1 VNB N_A_84_21#_c_82_n 0.0186908f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_2 VNB N_A_84_21#_c_83_n 0.0159846f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.995
cc_3 VNB N_A_84_21#_c_84_n 0.016003f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=0.995
cc_4 VNB N_A_84_21#_c_85_n 0.0193863f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=0.995
cc_5 VNB N_A_84_21#_c_86_n 0.00355803f $X=-0.19 $Y=-0.24 $X2=2.035 $Y2=1.16
cc_6 VNB N_A_84_21#_c_87_n 0.0783442f $X=-0.19 $Y=-0.24 $X2=1.84 $Y2=1.16
cc_7 VNB N_A_84_21#_c_88_n 0.00241867f $X=-0.19 $Y=-0.24 $X2=2.12 $Y2=0.995
cc_8 VNB N_A_84_21#_c_89_n 0.00192548f $X=-0.19 $Y=-0.24 $X2=2.96 $Y2=1.62
cc_9 VNB N_B1_c_207_n 0.0190753f $X=-0.19 $Y=-0.24 $X2=2.825 $Y2=0.235
cc_10 VNB N_B1_c_208_n 0.0165854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB B1 0.00312281f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_12 VNB N_B1_c_210_n 0.0438235f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_13 VNB N_A2_c_256_n 5.48114e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A2_c_257_n 0.0185455f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_15 VNB N_A2_c_258_n 0.00539737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_259_n 0.0152561f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=1.985
cc_17 VNB N_A2_c_260_n 0.027153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB A2 4.06108e-19 $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=0.56
cc_19 VNB N_A2_c_262_n 0.0161936f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.985
cc_20 VNB N_A2_c_263_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=2.035 $Y2=1.16
cc_21 VNB N_A1_c_341_n 0.0158558f $X=-0.19 $Y=-0.24 $X2=2.825 $Y2=0.235
cc_22 VNB N_A1_c_342_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB A1 0.00239074f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_24 VNB N_A1_c_344_n 0.0303857f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_25 VNB N_VPWR_c_386_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0191138f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=0.56
cc_27 VNB N_VGND_c_589_n 0.0108424f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_590_n 0.0119149f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.56
cc_29 VNB N_VGND_c_591_n 3.21528e-19 $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_30 VNB N_VGND_c_592_n 0.00215534f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=0.56
cc_31 VNB N_VGND_c_593_n 0.0329246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_594_n 0.0381373f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=0.56
cc_33 VNB N_VGND_c_595_n 0.00538573f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.325
cc_34 VNB N_VGND_c_596_n 0.0122657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_597_n 0.0136763f $X=-0.19 $Y=-0.24 $X2=2.12 $Y2=0.995
cc_36 VNB N_VGND_c_598_n 0.0115308f $X=-0.19 $Y=-0.24 $X2=2.96 $Y2=0.727
cc_37 VNB N_VGND_c_599_n 0.283827f $X=-0.19 $Y=-0.24 $X2=2.96 $Y2=0.76
cc_38 VNB N_VGND_c_600_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_39 VNB N_VGND_c_601_n 0.0161586f $X=-0.19 $Y=-0.24 $X2=1.785 $Y2=1.16
cc_40 VNB N_VGND_c_602_n 0.0184583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_603_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_A_84_21#_M1002_g 0.0215831f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_43 VPB N_A_84_21#_M1004_g 0.0185175f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_44 VPB N_A_84_21#_M1011_g 0.0185471f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=1.985
cc_45 VPB N_A_84_21#_M1015_g 0.0232145f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.985
cc_46 VPB N_A_84_21#_c_86_n 0.003676f $X=-0.19 $Y=1.305 $X2=2.035 $Y2=1.16
cc_47 VPB N_A_84_21#_c_87_n 0.0162427f $X=-0.19 $Y=1.305 $X2=1.84 $Y2=1.16
cc_48 VPB N_A_84_21#_c_89_n 0.00226264f $X=-0.19 $Y=1.305 $X2=2.96 $Y2=1.62
cc_49 VPB N_B1_M1017_g 0.0229722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_B1_M1019_g 0.018768f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_51 VPB B1 0.00372025f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_52 VPB N_B1_c_210_n 0.0103668f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_53 VPB N_A2_M1012_g 0.0179332f $X=-0.19 $Y=1.305 $X2=2.825 $Y2=1.485
cc_54 VPB N_A2_M1013_g 0.0221236f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_55 VPB N_A2_c_256_n 0.00167838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A2_c_257_n 0.00459096f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_57 VPB N_A2_c_260_n 0.00554505f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB A2 0.00690885f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=0.56
cc_59 VPB N_A1_M1000_g 0.0185163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A1_M1018_g 0.0185229f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_61 VPB N_A1_c_344_n 0.00412554f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_62 VPB N_VPWR_c_387_n 0.0109777f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_388_n 0.024292f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=0.56
cc_64 VPB N_VPWR_c_389_n 3.22457e-19 $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_65 VPB N_VPWR_c_390_n 0.0148075f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=0.56
cc_66 VPB N_VPWR_c_391_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.785 $Y2=0.56
cc_67 VPB N_VPWR_c_392_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=1.785 $Y2=1.985
cc_68 VPB N_VPWR_c_393_n 0.0352434f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.16
cc_69 VPB N_VPWR_c_394_n 0.00436029f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.16
cc_70 VPB N_VPWR_c_395_n 0.0111466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_396_n 0.00436029f $X=-0.19 $Y=1.305 $X2=1.84 $Y2=1.16
cc_72 VPB N_VPWR_c_397_n 0.0137965f $X=-0.19 $Y=1.305 $X2=2.12 $Y2=0.785
cc_73 VPB N_VPWR_c_398_n 0.0169549f $X=-0.19 $Y=1.305 $X2=2.96 $Y2=0.42
cc_74 VPB N_VPWR_c_399_n 0.0202711f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_75 VPB N_VPWR_c_386_n 0.0579736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_401_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_402_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB X 0.00946967f $X=-0.19 $Y=1.305 $X2=1.785 $Y2=0.56
cc_79 VPB N_A_483_297#_c_528_n 0.00330706f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_80 VPB N_A_483_297#_c_529_n 0.0223004f $X=-0.19 $Y=1.305 $X2=1.16 $Y2=1.16
cc_81 VPB N_A_483_297#_c_530_n 0.0219742f $X=-0.19 $Y=1.305 $X2=1.84 $Y2=1.16
cc_82 N_A_84_21#_c_88_n N_B1_c_207_n 0.0034583f $X=2.12 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_84_21#_c_98_p N_B1_c_207_n 0.0152609f $X=2.875 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_84_21#_c_89_n N_B1_c_207_n 0.00141942f $X=2.96 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_84_21#_c_89_n N_B1_M1017_g 0.0010989f $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_86 N_A_84_21#_c_89_n N_B1_c_208_n 0.00260329f $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_87 N_A_84_21#_c_102_p N_B1_c_208_n 0.0146368f $X=4.085 $Y=0.755 $X2=0 $Y2=0
cc_88 N_A_84_21#_c_89_n N_B1_M1019_g 0.0017889f $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_89 N_A_84_21#_M1015_g B1 0.00444188f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_84_21#_c_86_n B1 0.0268894f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_84_21#_c_87_n B1 8.0369e-19 $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_84_21#_c_98_p B1 0.0187508f $X=2.875 $Y=0.7 $X2=0 $Y2=0
cc_93 N_A_84_21#_c_89_n B1 0.0369083f $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_94 N_A_84_21#_c_86_n N_B1_c_210_n 0.00124369f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_84_21#_c_87_n N_B1_c_210_n 0.00624819f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_84_21#_c_98_p N_B1_c_210_n 0.00400852f $X=2.875 $Y=0.7 $X2=0 $Y2=0
cc_97 N_A_84_21#_c_89_n N_B1_c_210_n 0.0189867f $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_98 N_A_84_21#_c_89_n N_A2_c_256_n 0.00447131f $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_99 N_A_84_21#_c_102_p N_A2_c_271_n 0.00267108f $X=4.085 $Y=0.755 $X2=0 $Y2=0
cc_100 N_A_84_21#_c_89_n N_A2_c_257_n 4.5982e-19 $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_101 N_A_84_21#_c_102_p N_A2_c_257_n 0.00231315f $X=4.085 $Y=0.755 $X2=0 $Y2=0
cc_102 N_A_84_21#_c_89_n N_A2_c_258_n 0.0111268f $X=2.96 $Y=1.62 $X2=0 $Y2=0
cc_103 N_A_84_21#_c_102_p N_A2_c_258_n 0.0246715f $X=4.085 $Y=0.755 $X2=0 $Y2=0
cc_104 N_A_84_21#_c_102_p N_A2_c_262_n 0.0115203f $X=4.085 $Y=0.755 $X2=0 $Y2=0
cc_105 N_A_84_21#_c_120_p N_A2_c_263_n 0.00126506f $X=4.22 $Y=0.57 $X2=0 $Y2=0
cc_106 N_A_84_21#_c_102_p N_A1_c_341_n 0.0104547f $X=4.085 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_84_21#_c_120_p N_A1_c_342_n 0.0084371f $X=4.22 $Y=0.57 $X2=0 $Y2=0
cc_108 N_A_84_21#_c_102_p A1 0.00666638f $X=4.085 $Y=0.755 $X2=0 $Y2=0
cc_109 N_A_84_21#_c_120_p A1 0.0170411f $X=4.22 $Y=0.57 $X2=0 $Y2=0
cc_110 N_A_84_21#_c_120_p N_A1_c_344_n 0.0021041f $X=4.22 $Y=0.57 $X2=0 $Y2=0
cc_111 N_A_84_21#_M1002_g N_VPWR_c_388_n 0.0128801f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_A_84_21#_M1004_g N_VPWR_c_388_n 0.00131858f $X=0.925 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_84_21#_M1002_g N_VPWR_c_389_n 0.00131858f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_84_21#_M1004_g N_VPWR_c_389_n 0.0118176f $X=0.925 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_84_21#_M1011_g N_VPWR_c_389_n 0.0123474f $X=1.355 $Y=1.985 $X2=0
+ $Y2=0
cc_116 N_A_84_21#_M1015_g N_VPWR_c_389_n 0.00130238f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_84_21#_M1015_g N_VPWR_c_390_n 0.00311066f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_84_21#_c_86_n N_VPWR_c_390_n 0.0201913f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_84_21#_c_87_n N_VPWR_c_390_n 0.00135746f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_84_21#_M1002_g N_VPWR_c_397_n 0.00486043f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_84_21#_M1004_g N_VPWR_c_397_n 0.00486043f $X=0.925 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_84_21#_M1011_g N_VPWR_c_398_n 0.00486043f $X=1.355 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_84_21#_M1015_g N_VPWR_c_398_n 0.00557236f $X=1.785 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_84_21#_M1017_s N_VPWR_c_386_n 0.00216833f $X=2.825 $Y=1.485 $X2=0
+ $Y2=0
cc_125 N_A_84_21#_M1002_g N_VPWR_c_386_n 0.00830219f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_84_21#_M1004_g N_VPWR_c_386_n 0.00830219f $X=0.925 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_84_21#_M1011_g N_VPWR_c_386_n 0.00830219f $X=1.355 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_84_21#_M1015_g N_VPWR_c_386_n 0.011152f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_84_21#_c_82_n N_X_c_485_n 0.00884112f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_84_21#_c_83_n N_X_c_486_n 0.00972932f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_84_21#_c_84_n N_X_c_486_n 0.00972932f $X=1.355 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_84_21#_c_85_n N_X_c_486_n 0.00326174f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_84_21#_c_86_n N_X_c_486_n 0.0491543f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_84_21#_c_87_n N_X_c_486_n 0.00796547f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_84_21#_c_150_p N_X_c_486_n 0.00946301f $X=2.205 $Y=0.7 $X2=0 $Y2=0
cc_136 N_A_84_21#_M1004_g N_X_c_492_n 0.0127906f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_84_21#_M1011_g N_X_c_492_n 0.0127906f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_84_21#_c_86_n N_X_c_492_n 0.0299054f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_84_21#_c_87_n N_X_c_492_n 0.00210827f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_84_21#_M1015_g N_X_c_496_n 0.00227919f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_84_21#_c_86_n N_X_c_496_n 0.0127464f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_84_21#_c_87_n N_X_c_496_n 0.00220118f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_84_21#_M1015_g N_X_c_499_n 0.00513391f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_84_21#_c_82_n X 0.00755382f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_84_21#_M1002_g X 0.0220744f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_84_21#_c_83_n X 0.00470017f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_84_21#_M1004_g X 0.00589715f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_84_21#_c_86_n X 0.0269326f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_84_21#_c_87_n X 0.0216299f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_84_21#_M1017_s N_A_483_297#_c_531_n 0.00312348f $X=2.825 $Y=1.485
+ $X2=0 $Y2=0
cc_151 N_A_84_21#_c_89_n N_A_483_297#_c_531_n 0.0118865f $X=2.96 $Y=1.62 $X2=0
+ $Y2=0
cc_152 N_A_84_21#_c_89_n N_A_483_297#_c_528_n 0.00231527f $X=2.96 $Y=1.62 $X2=0
+ $Y2=0
cc_153 N_A_84_21#_c_102_p N_A_483_297#_c_528_n 0.00440519f $X=4.085 $Y=0.755
+ $X2=0 $Y2=0
cc_154 N_A_84_21#_c_88_n N_VGND_M1014_d 0.00322373f $X=2.12 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_98_p N_VGND_M1014_d 0.016382f $X=2.875 $Y=0.7 $X2=0 $Y2=0
cc_156 N_A_84_21#_c_150_p N_VGND_M1014_d 0.00525789f $X=2.205 $Y=0.7 $X2=0 $Y2=0
cc_157 N_A_84_21#_c_102_p N_VGND_M1010_s 0.00540394f $X=4.085 $Y=0.755 $X2=0
+ $Y2=0
cc_158 N_A_84_21#_c_82_n N_VGND_c_590_n 0.00873208f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_84_21#_c_83_n N_VGND_c_590_n 0.00104439f $X=0.925 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_84_21#_c_82_n N_VGND_c_591_n 0.00104385f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A_84_21#_c_83_n N_VGND_c_591_n 0.00765006f $X=0.925 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_84_21#_c_84_n N_VGND_c_591_n 0.00802115f $X=1.355 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_84_21#_c_85_n N_VGND_c_591_n 0.00109177f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_84_21#_c_102_p N_VGND_c_592_n 0.0133243f $X=4.085 $Y=0.755 $X2=0
+ $Y2=0
cc_165 N_A_84_21#_c_120_p N_VGND_c_592_n 0.00138436f $X=4.22 $Y=0.57 $X2=0 $Y2=0
cc_166 N_A_84_21#_c_102_p N_VGND_c_594_n 0.00696372f $X=4.085 $Y=0.755 $X2=0
+ $Y2=0
cc_167 N_A_84_21#_c_120_p N_VGND_c_594_n 0.00778691f $X=4.22 $Y=0.57 $X2=0 $Y2=0
cc_168 N_A_84_21#_c_82_n N_VGND_c_596_n 0.00350947f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_84_21#_c_83_n N_VGND_c_596_n 0.00351072f $X=0.925 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_84_21#_c_98_p N_VGND_c_597_n 0.00289974f $X=2.875 $Y=0.7 $X2=0 $Y2=0
cc_171 N_A_84_21#_c_186_p N_VGND_c_597_n 0.0113958f $X=2.96 $Y=0.42 $X2=0 $Y2=0
cc_172 N_A_84_21#_c_102_p N_VGND_c_597_n 0.00278663f $X=4.085 $Y=0.755 $X2=0
+ $Y2=0
cc_173 N_A_84_21#_M1007_d N_VGND_c_599_n 0.00250439f $X=2.825 $Y=0.235 $X2=0
+ $Y2=0
cc_174 N_A_84_21#_M1006_d N_VGND_c_599_n 0.00237222f $X=4.085 $Y=0.235 $X2=0
+ $Y2=0
cc_175 N_A_84_21#_c_82_n N_VGND_c_599_n 0.00411477f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_84_21#_c_83_n N_VGND_c_599_n 0.00411677f $X=0.925 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_84_21#_c_84_n N_VGND_c_599_n 0.00411677f $X=1.355 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_84_21#_c_85_n N_VGND_c_599_n 0.0112602f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_84_21#_c_98_p N_VGND_c_599_n 0.00692106f $X=2.875 $Y=0.7 $X2=0 $Y2=0
cc_180 N_A_84_21#_c_150_p N_VGND_c_599_n 8.9526e-19 $X=2.205 $Y=0.7 $X2=0 $Y2=0
cc_181 N_A_84_21#_c_186_p N_VGND_c_599_n 0.00646998f $X=2.96 $Y=0.42 $X2=0 $Y2=0
cc_182 N_A_84_21#_c_102_p N_VGND_c_599_n 0.0189434f $X=4.085 $Y=0.755 $X2=0
+ $Y2=0
cc_183 N_A_84_21#_c_120_p N_VGND_c_599_n 0.00961573f $X=4.22 $Y=0.57 $X2=0 $Y2=0
cc_184 N_A_84_21#_c_84_n N_VGND_c_601_n 0.00351072f $X=1.355 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_84_21#_c_85_n N_VGND_c_601_n 0.00558173f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_84_21#_c_85_n N_VGND_c_602_n 0.00729481f $X=1.785 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_84_21#_c_86_n N_VGND_c_602_n 0.00413883f $X=2.035 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_84_21#_c_87_n N_VGND_c_602_n 0.0011228f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_84_21#_c_98_p N_VGND_c_602_n 0.0317731f $X=2.875 $Y=0.7 $X2=0 $Y2=0
cc_190 N_A_84_21#_c_150_p N_VGND_c_602_n 0.0141996f $X=2.205 $Y=0.7 $X2=0 $Y2=0
cc_191 N_A_84_21#_c_102_p A_901_47# 0.00393556f $X=4.085 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_192 N_B1_M1019_g N_A2_M1012_g 0.0252159f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B1_c_210_n N_A2_c_256_n 5.41061e-19 $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B1_c_210_n N_A2_c_257_n 0.0221136f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_195 N_B1_c_210_n N_A2_c_258_n 0.00236109f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B1_c_208_n N_A2_c_262_n 0.0234488f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B1_M1017_g N_VPWR_c_390_n 0.00817358f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_198 B1 N_VPWR_c_390_n 5.93496e-19 $X=2.465 $Y=1.105 $X2=0 $Y2=0
cc_199 N_B1_M1019_g N_VPWR_c_391_n 0.00127615f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B1_M1017_g N_VPWR_c_393_n 0.00357877f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_201 N_B1_M1019_g N_VPWR_c_393_n 0.00357877f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B1_M1017_g N_VPWR_c_386_n 0.00664112f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B1_M1019_g N_VPWR_c_386_n 0.0052923f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_204 B1 N_A_483_297#_M1017_d 0.00366179f $X=2.465 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_205 B1 N_A_483_297#_c_536_n 0.0142739f $X=2.465 $Y=1.105 $X2=0 $Y2=0
cc_206 N_B1_c_210_n N_A_483_297#_c_536_n 6.82729e-19 $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_207 N_B1_M1017_g N_A_483_297#_c_531_n 0.0132518f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B1_M1019_g N_A_483_297#_c_531_n 0.013667f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B1_M1019_g N_A_483_297#_c_528_n 5.1213e-19 $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B1_c_208_n N_VGND_c_592_n 0.00165199f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B1_c_207_n N_VGND_c_597_n 0.00393283f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_c_208_n N_VGND_c_597_n 0.00430182f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_c_207_n N_VGND_c_599_n 0.00445457f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B1_c_208_n N_VGND_c_599_n 0.00577464f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B1_c_207_n N_VGND_c_602_n 0.00719299f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_208_n N_VGND_c_602_n 5.25906e-19 $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A2_c_262_n N_A1_c_341_n 0.0514295f $X=3.59 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_218 N_A2_M1012_g N_A1_M1000_g 0.0444243f $X=3.59 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A2_c_271_n N_A1_M1000_g 0.0114028f $X=4.685 $Y=1.595 $X2=0 $Y2=0
cc_220 N_A2_c_263_n N_A1_c_342_n 0.0340027f $X=4.91 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A2_M1013_g N_A1_M1018_g 0.0340027f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A2_c_271_n N_A1_M1018_g 0.0107085f $X=4.685 $Y=1.595 $X2=0 $Y2=0
cc_223 N_A2_c_271_n A1 0.025618f $X=4.685 $Y=1.595 $X2=0 $Y2=0
cc_224 N_A2_c_257_n A1 2.48288e-19 $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A2_c_258_n A1 0.0220504f $X=3.732 $Y=1.142 $X2=0 $Y2=0
cc_226 N_A2_c_259_n A1 0.0192998f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A2_c_260_n A1 0.00172154f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A2_c_256_n N_A1_c_344_n 0.00519415f $X=3.732 $Y=1.51 $X2=0 $Y2=0
cc_229 N_A2_c_271_n N_A1_c_344_n 0.00204885f $X=4.685 $Y=1.595 $X2=0 $Y2=0
cc_230 N_A2_c_257_n N_A1_c_344_n 0.0214987f $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A2_c_258_n N_A1_c_344_n 0.00180338f $X=3.732 $Y=1.142 $X2=0 $Y2=0
cc_232 N_A2_c_259_n N_A1_c_344_n 0.00114509f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A2_c_260_n N_A1_c_344_n 0.0340027f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_234 A2 N_A1_c_344_n 0.00483939f $X=4.765 $Y=1.445 $X2=0 $Y2=0
cc_235 N_A2_c_256_n N_VPWR_M1012_d 2.7057e-19 $X=3.732 $Y=1.51 $X2=0 $Y2=0
cc_236 N_A2_c_271_n N_VPWR_M1012_d 0.00181035f $X=4.685 $Y=1.595 $X2=0 $Y2=0
cc_237 N_A2_c_303_p N_VPWR_M1012_d 0.00105919f $X=3.82 $Y=1.595 $X2=0 $Y2=0
cc_238 N_A2_c_271_n N_VPWR_M1018_s 0.00595502f $X=4.685 $Y=1.595 $X2=0 $Y2=0
cc_239 A2 N_VPWR_M1018_s 2.9363e-19 $X=4.765 $Y=1.445 $X2=0 $Y2=0
cc_240 N_A2_c_306_p N_VPWR_M1018_s 3.4902e-19 $X=4.81 $Y=1.51 $X2=0 $Y2=0
cc_241 N_A2_M1012_g N_VPWR_c_391_n 0.00766759f $X=3.59 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A2_M1013_g N_VPWR_c_392_n 0.0106555f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A2_M1012_g N_VPWR_c_393_n 0.0034676f $X=3.59 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A2_M1013_g N_VPWR_c_399_n 0.0034676f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A2_M1012_g N_VPWR_c_386_n 0.00414378f $X=3.59 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A2_M1013_g N_VPWR_c_386_n 0.00525631f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A2_c_271_n N_A_483_297#_M1000_d 0.00332991f $X=4.685 $Y=1.595 $X2=0
+ $Y2=0
cc_248 N_A2_M1012_g N_A_483_297#_c_528_n 4.66965e-19 $X=3.59 $Y=1.985 $X2=0
+ $Y2=0
cc_249 N_A2_c_256_n N_A_483_297#_c_528_n 0.00350263f $X=3.732 $Y=1.51 $X2=0
+ $Y2=0
cc_250 N_A2_c_257_n N_A_483_297#_c_528_n 2.22737e-19 $X=3.59 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A2_c_258_n N_A_483_297#_c_528_n 0.00336061f $X=3.732 $Y=1.142 $X2=0
+ $Y2=0
cc_252 N_A2_M1012_g N_A_483_297#_c_546_n 0.0114928f $X=3.59 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A2_c_271_n N_A_483_297#_c_546_n 0.0143096f $X=4.685 $Y=1.595 $X2=0
+ $Y2=0
cc_254 N_A2_c_303_p N_A_483_297#_c_546_n 0.00902688f $X=3.82 $Y=1.595 $X2=0
+ $Y2=0
cc_255 N_A2_c_258_n N_A_483_297#_c_546_n 0.00403743f $X=3.732 $Y=1.142 $X2=0
+ $Y2=0
cc_256 N_A2_M1013_g N_A_483_297#_c_550_n 0.0134471f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A2_c_271_n N_A_483_297#_c_550_n 0.0190307f $X=4.685 $Y=1.595 $X2=0
+ $Y2=0
cc_258 N_A2_c_259_n N_A_483_297#_c_550_n 0.00200278f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A2_c_260_n N_A_483_297#_c_550_n 0.00149675f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A2_c_306_p N_A_483_297#_c_550_n 0.01344f $X=4.81 $Y=1.51 $X2=0 $Y2=0
cc_261 N_A2_M1013_g N_A_483_297#_c_529_n 0.00760973f $X=4.85 $Y=1.985 $X2=0
+ $Y2=0
cc_262 A2 N_A_483_297#_c_529_n 0.00292345f $X=4.765 $Y=1.445 $X2=0 $Y2=0
cc_263 N_A2_c_271_n N_A_483_297#_c_557_n 0.0125884f $X=4.685 $Y=1.595 $X2=0
+ $Y2=0
cc_264 N_A2_M1013_g N_A_483_297#_c_530_n 0.0127573f $X=4.85 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A2_c_259_n N_A_483_297#_c_530_n 0.00240172f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A2_c_260_n N_A_483_297#_c_530_n 2.75449e-19 $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A2_c_262_n N_VGND_c_592_n 0.00902354f $X=3.59 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A2_c_259_n N_VGND_c_593_n 0.0110232f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A2_c_260_n N_VGND_c_593_n 0.00235636f $X=4.91 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A2_c_263_n N_VGND_c_593_n 0.0047742f $X=4.91 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A2_c_262_n N_VGND_c_594_n 0.00343403f $X=3.59 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A2_c_263_n N_VGND_c_594_n 0.00585385f $X=4.91 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A2_c_262_n N_VGND_c_599_n 0.00397751f $X=3.59 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A2_c_263_n N_VGND_c_599_n 0.0116645f $X=4.91 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A1_M1000_g N_VPWR_c_391_n 0.00649906f $X=4.01 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A1_M1018_g N_VPWR_c_391_n 5.02907e-19 $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A1_M1000_g N_VPWR_c_392_n 5.02907e-19 $X=4.01 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A1_M1018_g N_VPWR_c_392_n 0.00649906f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A1_M1000_g N_VPWR_c_395_n 0.0034676f $X=4.01 $Y=1.985 $X2=0 $Y2=0
cc_280 N_A1_M1018_g N_VPWR_c_395_n 0.0034676f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A1_M1000_g N_VPWR_c_386_n 0.0040715f $X=4.01 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A1_M1018_g N_VPWR_c_386_n 0.0040715f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A1_M1000_g N_A_483_297#_c_546_n 0.00972199f $X=4.01 $Y=1.985 $X2=0
+ $Y2=0
cc_284 N_A1_M1018_g N_A_483_297#_c_550_n 0.00972199f $X=4.43 $Y=1.985 $X2=0
+ $Y2=0
cc_285 N_A1_c_341_n N_VGND_c_592_n 0.00206539f $X=4.01 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A1_c_341_n N_VGND_c_594_n 0.00430182f $X=4.01 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A1_c_342_n N_VGND_c_594_n 0.00573486f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A1_c_341_n N_VGND_c_599_n 0.00588392f $X=4.01 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A1_c_342_n N_VGND_c_599_n 0.010515f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_290 N_VPWR_c_386_n N_X_M1002_d 0.00651522f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_291 N_VPWR_c_386_n N_X_M1011_d 0.00469738f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_397_n N_X_c_508_n 0.00401379f $X=0.975 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_386_n N_X_c_508_n 0.00537716f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_M1004_s N_X_c_492_n 0.00368607f $X=1 $Y=1.485 $X2=0 $Y2=0
cc_295 N_VPWR_c_389_n N_X_c_492_n 0.0163515f $X=1.14 $Y=2.02 $X2=0 $Y2=0
cc_296 N_VPWR_c_398_n N_X_c_499_n 0.00529151f $X=1.915 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_c_386_n N_X_c_499_n 0.00783756f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_M1002_s X 0.0158247f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_299 N_VPWR_c_388_n X 0.0206836f $X=0.28 $Y=2.02 $X2=0 $Y2=0
cc_300 N_VPWR_c_386_n N_A_483_297#_M1017_d 0.0034899f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_301 N_VPWR_c_386_n N_A_483_297#_M1019_d 0.0023981f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_386_n N_A_483_297#_M1000_d 0.00258673f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_386_n N_A_483_297#_M1013_s 0.00374487f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_390_n N_A_483_297#_c_536_n 0.0312213f $X=2 $Y=1.68 $X2=0 $Y2=0
cc_305 N_VPWR_c_393_n N_A_483_297#_c_531_n 0.0473604f $X=3.635 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_386_n N_A_483_297#_c_531_n 0.0301315f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_390_n N_A_483_297#_c_570_n 0.00983759f $X=2 $Y=1.68 $X2=0 $Y2=0
cc_308 N_VPWR_c_393_n N_A_483_297#_c_570_n 0.0117106f $X=3.635 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_386_n N_A_483_297#_c_570_n 0.006547f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_310 N_VPWR_M1012_d N_A_483_297#_c_546_n 0.00353749f $X=3.665 $Y=1.485 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_391_n N_A_483_297#_c_546_n 0.0112304f $X=3.8 $Y=2.36 $X2=0 $Y2=0
cc_312 N_VPWR_c_393_n N_A_483_297#_c_546_n 0.00209524f $X=3.635 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_395_n N_A_483_297#_c_546_n 0.00209524f $X=4.475 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_386_n N_A_483_297#_c_546_n 0.00948897f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_395_n N_A_483_297#_c_578_n 0.0113154f $X=4.475 $Y=2.72 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_386_n N_A_483_297#_c_578_n 0.00645298f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_317 N_VPWR_M1018_s N_A_483_297#_c_550_n 0.00357106f $X=4.505 $Y=1.485 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_392_n N_A_483_297#_c_550_n 0.0112304f $X=4.64 $Y=2.36 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_395_n N_A_483_297#_c_550_n 0.00209524f $X=4.475 $Y=2.72 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_399_n N_A_483_297#_c_550_n 0.00288338f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_386_n N_A_483_297#_c_550_n 0.0109806f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_392_n N_A_483_297#_c_530_n 0.00751063f $X=4.64 $Y=2.36 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_399_n N_A_483_297#_c_530_n 0.015862f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_c_386_n N_A_483_297#_c_530_n 0.0121599f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_325 N_X_c_485_n N_VGND_M1001_d 0.0108744f $X=0.63 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_326 X N_VGND_M1001_d 0.00480177f $X=0.145 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_327 N_X_c_486_n N_VGND_M1003_d 0.00338318f $X=1.57 $Y=0.7 $X2=0 $Y2=0
cc_328 N_X_c_485_n N_VGND_c_590_n 0.0200973f $X=0.63 $Y=0.7 $X2=0 $Y2=0
cc_329 N_X_c_486_n N_VGND_c_591_n 0.0159085f $X=1.57 $Y=0.7 $X2=0 $Y2=0
cc_330 N_X_c_485_n N_VGND_c_596_n 0.00298323f $X=0.63 $Y=0.7 $X2=0 $Y2=0
cc_331 N_X_c_486_n N_VGND_c_596_n 0.00569019f $X=1.57 $Y=0.7 $X2=0 $Y2=0
cc_332 N_X_M1001_s N_VGND_c_599_n 0.00318884f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_333 N_X_M1005_s N_VGND_c_599_n 0.00318969f $X=1.43 $Y=0.235 $X2=0 $Y2=0
cc_334 N_X_c_485_n N_VGND_c_599_n 0.00658802f $X=0.63 $Y=0.7 $X2=0 $Y2=0
cc_335 N_X_c_486_n N_VGND_c_599_n 0.0224517f $X=1.57 $Y=0.7 $X2=0 $Y2=0
cc_336 N_X_c_486_n N_VGND_c_601_n 0.00676299f $X=1.57 $Y=0.7 $X2=0 $Y2=0
cc_337 N_A_483_297#_c_529_n N_VGND_c_593_n 0.00456504f $X=5.195 $Y=1.63 $X2=0
+ $Y2=0
cc_338 N_VGND_c_599_n A_901_47# 0.00280308f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24
cc_339 N_VGND_c_599_n A_741_47# 0.0115413f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o31a_1.spice.SKY130_FD_SC_HD__O31A_1.pxi
* Created: Thu Aug 27 14:39:50 2020
* 
x_PM_SKY130_FD_SC_HD__O31A_1%A_103_199# N_A_103_199#_M1009_d
+ N_A_103_199#_M1000_d N_A_103_199#_c_56_n N_A_103_199#_M1001_g
+ N_A_103_199#_M1002_g N_A_103_199#_c_57_n N_A_103_199#_c_58_n
+ N_A_103_199#_c_64_n N_A_103_199#_c_65_n N_A_103_199#_c_71_p
+ N_A_103_199#_c_82_p N_A_103_199#_c_72_p N_A_103_199#_c_86_p
+ N_A_103_199#_c_87_p N_A_103_199#_c_66_n N_A_103_199#_c_59_n
+ N_A_103_199#_c_60_n PM_SKY130_FD_SC_HD__O31A_1%A_103_199#
x_PM_SKY130_FD_SC_HD__O31A_1%A1 N_A1_M1003_g N_A1_M1005_g A1 N_A1_c_139_n
+ N_A1_c_140_n PM_SKY130_FD_SC_HD__O31A_1%A1
x_PM_SKY130_FD_SC_HD__O31A_1%A2 N_A2_c_171_n N_A2_M1006_g N_A2_M1004_g A2 A2 A2
+ N_A2_c_173_n PM_SKY130_FD_SC_HD__O31A_1%A2
x_PM_SKY130_FD_SC_HD__O31A_1%A3 N_A3_c_207_n N_A3_M1007_g N_A3_M1000_g A3
+ N_A3_c_209_n PM_SKY130_FD_SC_HD__O31A_1%A3
x_PM_SKY130_FD_SC_HD__O31A_1%B1 N_B1_M1009_g N_B1_M1008_g B1 N_B1_c_243_n
+ N_B1_c_244_n PM_SKY130_FD_SC_HD__O31A_1%B1
x_PM_SKY130_FD_SC_HD__O31A_1%X N_X_M1001_s N_X_M1002_s X X X X X X X N_X_c_276_n
+ X PM_SKY130_FD_SC_HD__O31A_1%X
x_PM_SKY130_FD_SC_HD__O31A_1%VPWR N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_c_292_n
+ N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n VPWR
+ N_VPWR_c_297_n N_VPWR_c_291_n PM_SKY130_FD_SC_HD__O31A_1%VPWR
x_PM_SKY130_FD_SC_HD__O31A_1%VGND N_VGND_M1001_d N_VGND_M1006_d N_VGND_c_337_n
+ N_VGND_c_338_n N_VGND_c_339_n VGND N_VGND_c_340_n N_VGND_c_341_n
+ N_VGND_c_342_n N_VGND_c_343_n PM_SKY130_FD_SC_HD__O31A_1%VGND
x_PM_SKY130_FD_SC_HD__O31A_1%A_253_47# N_A_253_47#_M1003_d N_A_253_47#_M1007_d
+ N_A_253_47#_c_397_n N_A_253_47#_c_384_n N_A_253_47#_c_385_n
+ N_A_253_47#_c_392_n PM_SKY130_FD_SC_HD__O31A_1%A_253_47#
cc_1 VNB N_A_103_199#_c_56_n 0.020295f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.995
cc_2 VNB N_A_103_199#_c_57_n 4.46663e-19 $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_3 VNB N_A_103_199#_c_58_n 0.0252531f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_4 VNB N_A_103_199#_c_59_n 0.0231706f $X=-0.19 $Y=-0.24 $X2=3.05 $Y2=1.495
cc_5 VNB N_A_103_199#_c_60_n 0.0275245f $X=-0.19 $Y=-0.24 $X2=2.81 $Y2=0.36
cc_6 VNB A1 0.00751177f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.56
cc_7 VNB N_A1_c_139_n 0.0190063f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.985
cc_8 VNB N_A1_c_140_n 0.017251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A2_c_171_n 0.0167675f $X=-0.19 $Y=-0.24 $X2=2.645 $Y2=0.235
cc_10 VNB A2 8.31138e-19 $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.56
cc_11 VNB N_A2_c_173_n 0.0222913f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_12 VNB N_A3_c_207_n 0.0171433f $X=-0.19 $Y=-0.24 $X2=2.645 $Y2=0.235
cc_13 VNB A3 0.00290055f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.56
cc_14 VNB N_A3_c_209_n 0.0203366f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.985
cc_15 VNB B1 0.00582402f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.56
cc_16 VNB N_B1_c_243_n 0.0264604f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.985
cc_17 VNB N_B1_c_244_n 0.0203297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0258296f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=2.38
cc_19 VNB N_X_c_276_n 0.0252463f $X=-0.19 $Y=-0.24 $X2=2.45 $Y2=1.66
cc_20 VNB N_VPWR_c_291_n 0.136896f $X=-0.19 $Y=-0.24 $X2=2.89 $Y2=0.36
cc_21 VNB N_VGND_c_337_n 5.61383e-19 $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.56
cc_22 VNB N_VGND_c_338_n 0.0191719f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.985
cc_23 VNB N_VGND_c_339_n 0.00617014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_340_n 0.0117788f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=1.53
cc_25 VNB N_VGND_c_341_n 0.0300713f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=2.295
cc_26 VNB N_VGND_c_342_n 0.182563f $X=-0.19 $Y=-0.24 $X2=2.965 $Y2=1.58
cc_27 VNB N_VGND_c_343_n 0.00598854f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=1.58
cc_28 VPB N_A_103_199#_M1002_g 0.0233522f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.985
cc_29 VPB N_A_103_199#_c_57_n 0.00245953f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_30 VPB N_A_103_199#_c_58_n 0.00548087f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_31 VPB N_A_103_199#_c_64_n 0.00599705f $X=-0.19 $Y=1.305 $X2=1.185 $Y2=1.53
cc_32 VPB N_A_103_199#_c_65_n 3.66229e-19 $X=-0.19 $Y=1.305 $X2=0.735 $Y2=1.53
cc_33 VPB N_A_103_199#_c_66_n 0.00801084f $X=-0.19 $Y=1.305 $X2=2.965 $Y2=1.58
cc_34 VPB N_A_103_199#_c_59_n 0.00935436f $X=-0.19 $Y=1.305 $X2=3.05 $Y2=1.495
cc_35 VPB N_A1_M1005_g 0.019844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A1_c_139_n 0.00406143f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.985
cc_37 VPB N_A2_M1004_g 0.0179385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB A2 0.00164103f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=0.56
cc_39 VPB A2 0.00256075f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=0.56
cc_40 VPB N_A2_c_173_n 0.00525592f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_41 VPB N_A3_M1000_g 0.0194949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB A3 0.00315937f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=0.56
cc_43 VPB N_A3_c_209_n 0.00566534f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.985
cc_44 VPB N_B1_M1008_g 0.0240351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB B1 0.0012295f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=0.56
cc_46 VPB N_B1_c_243_n 0.00531816f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.985
cc_47 VPB X 0.0245048f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=2.38
cc_48 VPB X 0.0282657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_292_n 0.00271285f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=0.56
cc_50 VPB N_VPWR_c_293_n 0.0115529f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.985
cc_51 VPB N_VPWR_c_294_n 0.0310364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_295_n 0.0192513f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_53 VPB N_VPWR_c_296_n 0.0048162f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_54 VPB N_VPWR_c_297_n 0.0426085f $X=-0.19 $Y=1.305 $X2=1.355 $Y2=2.38
cc_55 VPB N_VPWR_c_291_n 0.0441664f $X=-0.19 $Y=1.305 $X2=2.89 $Y2=0.36
cc_56 N_A_103_199#_M1002_g N_A1_M1005_g 0.0170252f $X=0.65 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A_103_199#_c_57_n N_A1_M1005_g 0.00201299f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_103_199#_c_64_n N_A1_M1005_g 0.0109966f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_59 N_A_103_199#_c_71_p N_A1_M1005_g 0.0147648f $X=1.27 $Y=2.295 $X2=0 $Y2=0
cc_60 N_A_103_199#_c_72_p N_A1_M1005_g 0.00500312f $X=1.355 $Y=2.38 $X2=0 $Y2=0
cc_61 N_A_103_199#_c_57_n A1 0.0214385f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_103_199#_c_58_n A1 0.00173297f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_103_199#_c_64_n A1 0.029767f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_64 N_A_103_199#_c_57_n N_A1_c_139_n 5.86485e-19 $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_103_199#_c_58_n N_A1_c_139_n 0.0203302f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_103_199#_c_64_n N_A1_c_139_n 0.00285216f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_67 N_A_103_199#_c_56_n N_A1_c_140_n 0.00783657f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_68 N_A_103_199#_c_64_n N_A2_M1004_g 6.63228e-19 $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_69 N_A_103_199#_c_71_p N_A2_M1004_g 0.00499689f $X=1.27 $Y=2.295 $X2=0 $Y2=0
cc_70 N_A_103_199#_c_82_p N_A2_M1004_g 0.00984966f $X=2.365 $Y=2.38 $X2=0 $Y2=0
cc_71 N_A_103_199#_c_64_n A2 0.00921084f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_72 N_A_103_199#_c_82_p A2 0.0106994f $X=2.365 $Y=2.38 $X2=0 $Y2=0
cc_73 N_A_103_199#_c_82_p N_A3_M1000_g 0.010625f $X=2.365 $Y=2.38 $X2=0 $Y2=0
cc_74 N_A_103_199#_c_86_p N_A3_M1000_g 7.54408e-19 $X=2.49 $Y=1.665 $X2=0 $Y2=0
cc_75 N_A_103_199#_c_87_p N_A3_M1000_g 0.00559579f $X=2.49 $Y=2.295 $X2=0 $Y2=0
cc_76 N_A_103_199#_c_82_p A3 0.0131377f $X=2.365 $Y=2.38 $X2=0 $Y2=0
cc_77 N_A_103_199#_c_82_p N_B1_M1008_g 0.00206775f $X=2.365 $Y=2.38 $X2=0 $Y2=0
cc_78 N_A_103_199#_c_86_p N_B1_M1008_g 7.32094e-19 $X=2.49 $Y=1.665 $X2=0 $Y2=0
cc_79 N_A_103_199#_c_87_p N_B1_M1008_g 0.0151299f $X=2.49 $Y=2.295 $X2=0 $Y2=0
cc_80 N_A_103_199#_c_66_n N_B1_M1008_g 0.0127303f $X=2.965 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_103_199#_c_86_p B1 0.0160964f $X=2.49 $Y=1.665 $X2=0 $Y2=0
cc_82 N_A_103_199#_c_66_n B1 0.0111826f $X=2.965 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A_103_199#_c_59_n B1 0.0265524f $X=3.05 $Y=1.495 $X2=0 $Y2=0
cc_84 N_A_103_199#_c_60_n B1 0.00990947f $X=2.81 $Y=0.36 $X2=0 $Y2=0
cc_85 N_A_103_199#_c_86_p N_B1_c_243_n 0.00381184f $X=2.49 $Y=1.665 $X2=0 $Y2=0
cc_86 N_A_103_199#_c_59_n N_B1_c_243_n 0.00748071f $X=3.05 $Y=1.495 $X2=0 $Y2=0
cc_87 N_A_103_199#_c_60_n N_B1_c_243_n 0.0023839f $X=2.81 $Y=0.36 $X2=0 $Y2=0
cc_88 N_A_103_199#_c_59_n N_B1_c_244_n 0.00406668f $X=3.05 $Y=1.495 $X2=0 $Y2=0
cc_89 N_A_103_199#_c_56_n X 0.0043528f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_103_199#_M1002_g X 0.00830335f $X=0.65 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_103_199#_c_57_n X 0.0342139f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_103_199#_c_58_n X 0.00765123f $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_103_199#_c_65_n X 0.00866322f $X=0.735 $Y=1.53 $X2=0 $Y2=0
cc_94 N_A_103_199#_c_58_n N_X_c_276_n 2.50771e-19 $X=0.65 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_103_199#_c_64_n N_VPWR_M1002_d 0.00434929f $X=1.185 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_103_199#_c_66_n N_VPWR_M1008_d 0.00797371f $X=2.965 $Y=1.58 $X2=0
+ $Y2=0
cc_97 N_A_103_199#_M1002_g N_VPWR_c_292_n 0.0148895f $X=0.65 $Y=1.985 $X2=0
+ $Y2=0
cc_98 N_A_103_199#_c_64_n N_VPWR_c_292_n 0.0188752f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_99 N_A_103_199#_c_65_n N_VPWR_c_292_n 0.00197512f $X=0.735 $Y=1.53 $X2=0
+ $Y2=0
cc_100 N_A_103_199#_c_71_p N_VPWR_c_292_n 0.0375609f $X=1.27 $Y=2.295 $X2=0
+ $Y2=0
cc_101 N_A_103_199#_c_72_p N_VPWR_c_292_n 0.0139612f $X=1.355 $Y=2.38 $X2=0
+ $Y2=0
cc_102 N_A_103_199#_c_66_n N_VPWR_c_294_n 0.0280603f $X=2.965 $Y=1.58 $X2=0
+ $Y2=0
cc_103 N_A_103_199#_M1002_g N_VPWR_c_295_n 0.00486043f $X=0.65 $Y=1.985 $X2=0
+ $Y2=0
cc_104 N_A_103_199#_c_82_p N_VPWR_c_297_n 0.0725033f $X=2.365 $Y=2.38 $X2=0
+ $Y2=0
cc_105 N_A_103_199#_c_72_p N_VPWR_c_297_n 0.00979741f $X=1.355 $Y=2.38 $X2=0
+ $Y2=0
cc_106 N_A_103_199#_M1000_d N_VPWR_c_291_n 0.00341579f $X=2.165 $Y=1.485 $X2=0
+ $Y2=0
cc_107 N_A_103_199#_M1002_g N_VPWR_c_291_n 0.00940435f $X=0.65 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_103_199#_c_82_p N_VPWR_c_291_n 0.0456869f $X=2.365 $Y=2.38 $X2=0
+ $Y2=0
cc_109 N_A_103_199#_c_72_p N_VPWR_c_291_n 0.00618115f $X=1.355 $Y=2.38 $X2=0
+ $Y2=0
cc_110 N_A_103_199#_c_64_n A_253_297# 0.00113639f $X=1.185 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_103_199#_c_71_p A_253_297# 0.00624788f $X=1.27 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_103_199#_c_82_p A_253_297# 0.00580081f $X=2.365 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_103_199#_c_72_p A_253_297# 3.22723e-19 $X=1.355 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_103_199#_c_82_p A_337_297# 0.00938948f $X=2.365 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_103_199#_c_56_n N_VGND_c_337_n 0.013122f $X=0.65 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_103_199#_c_57_n N_VGND_c_337_n 0.00277103f $X=0.65 $Y=1.16 $X2=0
+ $Y2=0
cc_117 N_A_103_199#_c_58_n N_VGND_c_337_n 0.00106074f $X=0.65 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_A_103_199#_c_64_n N_VGND_c_337_n 0.00469622f $X=1.185 $Y=1.53 $X2=0
+ $Y2=0
cc_119 N_A_103_199#_c_56_n N_VGND_c_338_n 0.0046653f $X=0.65 $Y=0.995 $X2=0
+ $Y2=0
cc_120 N_A_103_199#_c_60_n N_VGND_c_341_n 0.0323743f $X=2.81 $Y=0.36 $X2=0 $Y2=0
cc_121 N_A_103_199#_M1009_d N_VGND_c_342_n 0.00250309f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_122 N_A_103_199#_c_56_n N_VGND_c_342_n 0.00909722f $X=0.65 $Y=0.995 $X2=0
+ $Y2=0
cc_123 N_A_103_199#_c_60_n N_VGND_c_342_n 0.0187375f $X=2.81 $Y=0.36 $X2=0 $Y2=0
cc_124 N_A_103_199#_c_86_p N_A_253_47#_c_384_n 7.86906e-19 $X=2.49 $Y=1.665
+ $X2=0 $Y2=0
cc_125 N_A_103_199#_c_64_n N_A_253_47#_c_385_n 0.00130321f $X=1.185 $Y=1.53
+ $X2=0 $Y2=0
cc_126 N_A1_c_140_n N_A2_c_171_n 0.0235606f $X=1.13 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_127 N_A1_M1005_g N_A2_M1004_g 0.0602645f $X=1.19 $Y=1.985 $X2=0 $Y2=0
cc_128 A1 A2 0.0206392f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_129 N_A1_c_139_n A2 6.78235e-19 $X=1.13 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A1_M1005_g A2 0.00280499f $X=1.19 $Y=1.985 $X2=0 $Y2=0
cc_131 A1 N_A2_c_173_n 0.00159548f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A1_c_139_n N_A2_c_173_n 0.020542f $X=1.13 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A1_M1005_g N_VPWR_c_292_n 0.00510722f $X=1.19 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A1_M1005_g N_VPWR_c_297_n 0.00463936f $X=1.19 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A1_M1005_g N_VPWR_c_291_n 0.00809909f $X=1.19 $Y=1.985 $X2=0 $Y2=0
cc_136 A1 N_VGND_c_337_n 0.017196f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A1_c_139_n N_VGND_c_337_n 7.77033e-19 $X=1.13 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A1_c_140_n N_VGND_c_337_n 0.0108291f $X=1.13 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_c_140_n N_VGND_c_340_n 0.0046653f $X=1.13 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_c_140_n N_VGND_c_342_n 0.00799591f $X=1.13 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A1_c_140_n N_VGND_c_343_n 5.59196e-19 $X=1.13 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A2_c_171_n N_A3_c_207_n 0.0218007f $X=1.61 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_143 N_A2_M1004_g N_A3_M1000_g 0.0477842f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_144 A2 N_A3_M1000_g 9.18397e-19 $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_145 N_A2_M1004_g A3 0.00263562f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_146 A2 A3 0.0550984f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A2_c_173_n A3 0.00185237f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_148 A2 N_A3_c_209_n 3.8169e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A2_c_173_n N_A3_c_209_n 0.0203414f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_M1004_g N_VPWR_c_297_n 0.00357877f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A2_M1004_g N_VPWR_c_291_n 0.00546655f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A2_c_171_n N_VGND_c_337_n 6.91082e-19 $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A2_c_171_n N_VGND_c_340_n 0.00342417f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A2_c_171_n N_VGND_c_342_n 0.00405449f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A2_c_171_n N_VGND_c_343_n 0.00707893f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_c_171_n N_A_253_47#_c_384_n 0.0104349f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_157 A2 N_A_253_47#_c_384_n 0.0149998f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A2_c_173_n N_A_253_47#_c_384_n 4.76779e-19 $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A3_M1000_g N_B1_M1008_g 0.0231588f $X=2.09 $Y=1.985 $X2=0 $Y2=0
cc_160 A3 N_B1_M1008_g 0.00281575f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_161 A3 B1 0.0218001f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A3_c_209_n B1 0.00207544f $X=2.09 $Y=1.16 $X2=0 $Y2=0
cc_163 A3 N_B1_c_243_n 3.51722e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A3_c_209_n N_B1_c_243_n 0.0203288f $X=2.09 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A3_c_207_n N_B1_c_244_n 0.0188926f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A3_M1000_g N_VPWR_c_297_n 0.00357877f $X=2.09 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A3_M1000_g N_VPWR_c_291_n 0.00581352f $X=2.09 $Y=1.985 $X2=0 $Y2=0
cc_168 A3 A_337_297# 0.0062622f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_169 N_A3_c_207_n N_VGND_c_341_n 0.00256813f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A3_c_207_n N_VGND_c_342_n 0.00335748f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A3_c_207_n N_VGND_c_343_n 0.0101098f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A3_c_207_n N_A_253_47#_c_384_n 0.0103396f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_173 A3 N_A_253_47#_c_384_n 0.016853f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A3_c_209_n N_A_253_47#_c_384_n 0.00138218f $X=2.09 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A3_c_207_n N_A_253_47#_c_392_n 0.00462294f $X=2.09 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B1_M1008_g N_VPWR_c_294_n 0.0169743f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B1_M1008_g N_VPWR_c_297_n 0.00547432f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_178 N_B1_M1008_g N_VPWR_c_291_n 0.0111648f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_179 N_B1_c_244_n N_VGND_c_341_n 0.00585385f $X=2.587 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B1_c_244_n N_VGND_c_342_n 0.0119977f $X=2.587 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B1_c_244_n N_VGND_c_343_n 0.00119839f $X=2.587 $Y=0.995 $X2=0 $Y2=0
cc_182 B1 N_A_253_47#_c_384_n 0.0054881f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_183 N_B1_c_243_n N_A_253_47#_c_384_n 8.18609e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_184 X N_VPWR_c_295_n 0.0307205f $X=0.23 $Y=1.87 $X2=0 $Y2=0
cc_185 N_X_M1002_s N_VPWR_c_291_n 0.00469152f $X=0.215 $Y=1.485 $X2=0 $Y2=0
cc_186 X N_VPWR_c_291_n 0.0168582f $X=0.23 $Y=1.87 $X2=0 $Y2=0
cc_187 N_X_c_276_n N_VGND_c_338_n 0.0288089f $X=0.36 $Y=0.36 $X2=0 $Y2=0
cc_188 N_X_M1001_s N_VGND_c_342_n 0.00469537f $X=0.215 $Y=0.235 $X2=0 $Y2=0
cc_189 N_X_c_276_n N_VGND_c_342_n 0.0167626f $X=0.36 $Y=0.36 $X2=0 $Y2=0
cc_190 N_VPWR_c_291_n A_253_297# 0.00216824f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_191 N_VPWR_c_291_n A_337_297# 0.00265018f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_192 N_VGND_c_342_n N_A_253_47#_M1003_d 0.00412745f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_193 N_VGND_c_342_n N_A_253_47#_M1007_d 0.00370961f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_340_n N_A_253_47#_c_397_n 0.0112554f $X=1.655 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_342_n N_A_253_47#_c_397_n 0.00644035f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_M1006_d N_A_253_47#_c_384_n 0.00943141f $X=1.685 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_VGND_c_340_n N_A_253_47#_c_384_n 0.00233324f $X=1.655 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_341_n N_A_253_47#_c_384_n 0.00230733f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_342_n N_A_253_47#_c_384_n 0.0102298f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_c_343_n N_A_253_47#_c_384_n 0.022823f $X=2.07 $Y=0 $X2=0 $Y2=0
cc_201 N_VGND_c_341_n N_A_253_47#_c_392_n 0.0146061f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_342_n N_A_253_47#_c_392_n 0.00874048f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_c_343_n N_A_253_47#_c_392_n 0.0176937f $X=2.07 $Y=0 $X2=0 $Y2=0

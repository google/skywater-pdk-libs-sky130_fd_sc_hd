* File: sky130_fd_sc_hd__a211oi_1.spice
* Created: Thu Aug 27 13:59:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a211oi_1.pex.spice"
.subckt sky130_fd_sc_hd__a211oi_1  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 A_139_47# N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.2665 PD=0.93 PS=2.12 NRD=15.684 NRS=26.76 M=1 R=4.33333 SA=75000.3
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g A_139_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75000.8 SB=75001.1
+ A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.091 PD=0.96 PS=0.93 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_C1_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.10075 PD=1.83 PS=0.96 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_56_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1000 N_A_56_297#_M1000_d N_A1_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 A_311_297# N_B1_M1005_g N_A_56_297#_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.155 AS=0.14 PD=1.31 PS=1.28 NRD=19.6803 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1006_d N_C1_M1006_g A_311_297# VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.155 PD=2.53 PS=1.31 NRD=0 NRS=19.6803 M=1 R=6.66667 SA=75001.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
c_44 VPB 0 1.20783e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a211oi_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o2111ai_2.spice.SKY130_FD_SC_HD__O2111AI_2.pxi
* Created: Thu Aug 27 14:34:13 2020
* 
x_PM_SKY130_FD_SC_HD__O2111AI_2%D1 N_D1_c_93_n N_D1_M1006_g N_D1_M1005_g
+ N_D1_c_94_n N_D1_M1007_g N_D1_M1017_g N_D1_c_95_n N_D1_c_96_n D1
+ PM_SKY130_FD_SC_HD__O2111AI_2%D1
x_PM_SKY130_FD_SC_HD__O2111AI_2%C1 N_C1_M1004_g N_C1_M1000_g N_C1_M1016_g
+ N_C1_M1012_g N_C1_c_141_n N_C1_c_142_n N_C1_c_143_n C1 C1
+ PM_SKY130_FD_SC_HD__O2111AI_2%C1
x_PM_SKY130_FD_SC_HD__O2111AI_2%B1 N_B1_M1002_g N_B1_M1014_g N_B1_M1013_g
+ N_B1_M1019_g N_B1_c_191_n N_B1_c_192_n N_B1_c_193_n N_B1_c_194_n B1 B1
+ PM_SKY130_FD_SC_HD__O2111AI_2%B1
x_PM_SKY130_FD_SC_HD__O2111AI_2%A2 N_A2_M1009_g N_A2_M1003_g N_A2_M1018_g
+ N_A2_M1011_g N_A2_c_246_n N_A2_c_247_n N_A2_c_248_n A2 A2 A2
+ PM_SKY130_FD_SC_HD__O2111AI_2%A2
x_PM_SKY130_FD_SC_HD__O2111AI_2%A1 N_A1_M1010_g N_A1_M1001_g N_A1_M1015_g
+ N_A1_M1008_g N_A1_c_291_n N_A1_c_292_n N_A1_c_293_n A1 A1
+ PM_SKY130_FD_SC_HD__O2111AI_2%A1
x_PM_SKY130_FD_SC_HD__O2111AI_2%VPWR N_VPWR_M1005_d N_VPWR_M1017_d
+ N_VPWR_M1012_s N_VPWR_M1014_s N_VPWR_M1001_s N_VPWR_c_329_n N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n VPWR
+ N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_328_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n
+ PM_SKY130_FD_SC_HD__O2111AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O2111AI_2%Y N_Y_M1006_s N_Y_M1005_s N_Y_M1000_d
+ N_Y_M1002_d N_Y_M1003_s N_Y_c_416_n N_Y_c_452_n N_Y_c_429_n N_Y_c_456_n
+ N_Y_c_414_n N_Y_c_466_p N_Y_c_431_n N_Y_c_441_n Y Y Y Y Y N_Y_c_413_n Y
+ PM_SKY130_FD_SC_HD__O2111AI_2%Y
x_PM_SKY130_FD_SC_HD__O2111AI_2%A_664_297# N_A_664_297#_M1003_d
+ N_A_664_297#_M1011_d N_A_664_297#_M1008_d N_A_664_297#_c_474_n
+ N_A_664_297#_c_475_n N_A_664_297#_c_476_n N_A_664_297#_c_478_n
+ N_A_664_297#_c_480_n N_A_664_297#_c_482_n N_A_664_297#_c_499_n
+ PM_SKY130_FD_SC_HD__O2111AI_2%A_664_297#
x_PM_SKY130_FD_SC_HD__O2111AI_2%A_27_47# N_A_27_47#_M1006_d N_A_27_47#_M1007_d
+ N_A_27_47#_M1016_d N_A_27_47#_c_538_p N_A_27_47#_c_511_n N_A_27_47#_c_513_n
+ N_A_27_47#_c_508_n N_A_27_47#_c_509_n N_A_27_47#_c_510_n
+ PM_SKY130_FD_SC_HD__O2111AI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__O2111AI_2%A_298_47# N_A_298_47#_M1004_s
+ N_A_298_47#_M1013_s N_A_298_47#_c_548_n N_A_298_47#_c_551_n
+ N_A_298_47#_c_547_n PM_SKY130_FD_SC_HD__O2111AI_2%A_298_47#
x_PM_SKY130_FD_SC_HD__O2111AI_2%A_497_47# N_A_497_47#_M1013_d
+ N_A_497_47#_M1019_d N_A_497_47#_M1018_d N_A_497_47#_M1015_s
+ N_A_497_47#_c_573_n N_A_497_47#_c_604_p N_A_497_47#_c_580_n
+ N_A_497_47#_c_607_p N_A_497_47#_c_586_n N_A_497_47#_c_584_n
+ N_A_497_47#_c_585_n N_A_497_47#_c_574_n
+ PM_SKY130_FD_SC_HD__O2111AI_2%A_497_47#
x_PM_SKY130_FD_SC_HD__O2111AI_2%VGND N_VGND_M1009_s N_VGND_M1010_d
+ N_VGND_c_621_n N_VGND_c_622_n VGND N_VGND_c_623_n N_VGND_c_624_n
+ N_VGND_c_625_n N_VGND_c_626_n N_VGND_c_627_n N_VGND_c_628_n
+ PM_SKY130_FD_SC_HD__O2111AI_2%VGND
cc_1 VNB N_D1_c_93_n 0.0215964f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_2 VNB N_D1_c_94_n 0.0163088f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=0.995
cc_3 VNB N_D1_c_95_n 0.0327591f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_4 VNB N_D1_c_96_n 0.0266111f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_5 VNB D1 0.0100329f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_C1_M1004_g 0.017763f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_7 VNB N_C1_M1000_g 3.83102e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_C1_M1016_g 0.0240079f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.325
cc_9 VNB N_C1_M1012_g 4.33886e-19 $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_10 VNB N_C1_c_141_n 0.00822668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_C1_c_142_n 0.0131346f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_12 VNB N_C1_c_143_n 0.00964089f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB C1 0.00298086f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_14 VNB N_B1_M1002_g 3.83102e-19 $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_15 VNB N_B1_M1014_g 5.20615e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_M1013_g 0.0241107f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.325
cc_17 VNB N_B1_M1019_g 0.0180205f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_18 VNB N_B1_c_191_n 0.0127801f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_19 VNB N_B1_c_192_n 0.0147479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B1_c_193_n 0.0187557f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_21 VNB N_B1_c_194_n 0.0319228f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_22 VNB B1 0.00210397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A2_M1009_g 0.0178214f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_24 VNB N_A2_M1003_g 5.20615e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A2_M1018_g 0.0178214f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.325
cc_26 VNB N_A2_M1011_g 3.83102e-19 $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_27 VNB N_A2_c_246_n 0.00822936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A2_c_247_n 0.0132147f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_29 VNB N_A2_c_248_n 0.00822936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB A2 0.00932785f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_31 VNB N_A1_M1010_g 0.0178214f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_32 VNB N_A1_M1001_g 4.66859e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A1_M1015_g 0.0242965f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.325
cc_34 VNB N_A1_M1008_g 5.20615e-19 $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_35 VNB N_A1_c_291_n 0.00959742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A1_c_292_n 0.0132147f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_37 VNB N_A1_c_293_n 0.0133085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB A1 0.015006f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_39 VNB N_VPWR_c_328_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB Y 8.49635e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_413_n 6.30066e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_508_n 0.00273084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_c_509_n 0.00186829f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_44 VNB N_A_27_47#_c_510_n 0.00870418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_298_47#_c_547_n 0.00669637f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_46 VNB N_A_497_47#_c_573_n 0.00215605f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_47 VNB N_A_497_47#_c_574_n 0.01954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_621_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=0.56
cc_49 VNB N_VGND_c_622_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_50 VNB N_VGND_c_623_n 0.0891685f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.16
cc_51 VNB N_VGND_c_624_n 0.0118064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_625_n 0.0166039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_626_n 0.28004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_627_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_628_n 0.00436244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VPB N_D1_M1005_g 0.0247014f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_57 VPB N_D1_M1017_g 0.0187781f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_58 VPB N_D1_c_95_n 0.0126262f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_59 VPB N_D1_c_96_n 0.00434271f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.16
cc_60 VPB D1 0.007624f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_61 VPB N_C1_M1000_g 0.0197155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_C1_M1012_g 0.01985f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_63 VPB C1 0.00517544f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_64 VPB N_B1_M1002_g 0.0197428f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.56
cc_65 VPB N_B1_M1014_g 0.0264988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB B1 0.00663735f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A2_M1003_g 0.0273652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A2_M1011_g 0.0199855f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_69 VPB A2 0.0100179f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_70 VPB N_A1_M1001_g 0.0201624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A1_M1008_g 0.0271661f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_72 VPB A1 0.00924953f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_73 VPB N_VPWR_c_329_n 0.012566f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.16
cc_74 VPB N_VPWR_c_330_n 0.0406807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_331_n 3.22457e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_76 VPB N_VPWR_c_332_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_333_n 0.00932429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_334_n 0.00239351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_335_n 0.0157463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_336_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_337_n 0.0130339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_338_n 0.0388128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_339_n 0.0174443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_328_n 0.0580537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_341_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_342_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_343_n 0.00510842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_344_n 0.00375828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_Y_c_414_n 0.0121463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB Y 0.00151789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_664_297#_c_474_n 0.00168448f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=0.56
cc_92 VPB N_A_664_297#_c_475_n 0.00373754f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_93 N_D1_c_94_n N_C1_M1004_g 0.0217304f $X=0.985 $Y=0.995 $X2=0 $Y2=0
cc_94 N_D1_M1017_g N_C1_M1000_g 0.0217304f $X=0.985 $Y=1.985 $X2=0 $Y2=0
cc_95 N_D1_c_96_n N_C1_c_141_n 0.0217304f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_96 N_D1_c_96_n C1 0.00765539f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_97 N_D1_M1005_g N_VPWR_c_330_n 0.00675012f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_98 N_D1_c_95_n N_VPWR_c_330_n 0.00180829f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_99 D1 N_VPWR_c_330_n 0.0212679f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_100 N_D1_M1005_g N_VPWR_c_331_n 6.8852e-19 $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_101 N_D1_M1017_g N_VPWR_c_331_n 0.0108488f $X=0.985 $Y=1.985 $X2=0 $Y2=0
cc_102 N_D1_M1005_g N_VPWR_c_335_n 0.0054895f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_103 N_D1_M1017_g N_VPWR_c_335_n 0.00486043f $X=0.985 $Y=1.985 $X2=0 $Y2=0
cc_104 N_D1_M1005_g N_VPWR_c_328_n 0.0107517f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_105 N_D1_M1017_g N_VPWR_c_328_n 0.00822531f $X=0.985 $Y=1.985 $X2=0 $Y2=0
cc_106 N_D1_M1017_g N_Y_c_416_n 0.0176557f $X=0.985 $Y=1.985 $X2=0 $Y2=0
cc_107 N_D1_c_93_n Y 0.00453653f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_108 N_D1_M1005_g Y 0.00778359f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_109 N_D1_c_94_n Y 0.0023331f $X=0.985 $Y=0.995 $X2=0 $Y2=0
cc_110 N_D1_M1017_g Y 0.00421109f $X=0.985 $Y=1.985 $X2=0 $Y2=0
cc_111 N_D1_c_96_n Y 0.0244482f $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_112 D1 Y 0.019798f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_113 N_D1_M1005_g Y 0.00469133f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_114 N_D1_M1005_g Y 0.00961576f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_115 N_D1_c_93_n N_Y_c_413_n 0.00495465f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_116 N_D1_c_94_n N_Y_c_413_n 0.0041569f $X=0.985 $Y=0.995 $X2=0 $Y2=0
cc_117 N_D1_c_95_n N_A_27_47#_c_511_n 0.00640784f $X=0.48 $Y=1.16 $X2=0 $Y2=0
cc_118 D1 N_A_27_47#_c_511_n 0.0170321f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_119 N_D1_c_93_n N_A_27_47#_c_513_n 0.0119317f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_120 N_D1_c_94_n N_A_27_47#_c_513_n 0.0133103f $X=0.985 $Y=0.995 $X2=0 $Y2=0
cc_121 N_D1_c_96_n N_A_27_47#_c_513_n 3.20336e-19 $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_122 N_D1_c_94_n N_A_27_47#_c_509_n 4.56855e-19 $X=0.985 $Y=0.995 $X2=0 $Y2=0
cc_123 N_D1_c_93_n N_VGND_c_623_n 0.00358923f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_124 N_D1_c_94_n N_VGND_c_623_n 0.00358923f $X=0.985 $Y=0.995 $X2=0 $Y2=0
cc_125 N_D1_c_93_n N_VGND_c_626_n 0.00627986f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_126 N_D1_c_94_n N_VGND_c_626_n 0.00534612f $X=0.985 $Y=0.995 $X2=0 $Y2=0
cc_127 N_C1_M1012_g N_B1_M1002_g 0.0212779f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_128 N_C1_c_143_n N_B1_c_191_n 0.0212779f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_129 C1 N_B1_c_191_n 2.57295e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_130 N_C1_c_143_n B1 0.0011034f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_131 C1 B1 0.0102219f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_132 N_C1_M1000_g N_VPWR_c_331_n 0.0106688f $X=1.415 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C1_M1012_g N_VPWR_c_331_n 6.23052e-19 $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_134 N_C1_M1000_g N_VPWR_c_332_n 6.21637e-19 $X=1.415 $Y=1.985 $X2=0 $Y2=0
cc_135 N_C1_M1012_g N_VPWR_c_332_n 0.0106233f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_136 N_C1_M1000_g N_VPWR_c_336_n 0.00486043f $X=1.415 $Y=1.985 $X2=0 $Y2=0
cc_137 N_C1_M1012_g N_VPWR_c_336_n 0.00486043f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_138 N_C1_M1000_g N_VPWR_c_328_n 0.00822531f $X=1.415 $Y=1.985 $X2=0 $Y2=0
cc_139 N_C1_M1012_g N_VPWR_c_328_n 0.00822531f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_140 N_C1_M1000_g N_Y_c_416_n 0.0140805f $X=1.415 $Y=1.985 $X2=0 $Y2=0
cc_141 C1 N_Y_c_416_n 0.0305281f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_142 N_C1_M1012_g N_Y_c_429_n 0.015823f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_143 C1 N_Y_c_429_n 0.00319344f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_144 N_C1_c_142_n N_Y_c_431_n 7.32538e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_145 C1 N_Y_c_431_n 0.0150669f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_146 N_C1_M1004_g Y 3.82486e-19 $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_147 C1 Y 0.0185842f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_148 C1 N_A_27_47#_c_513_n 0.0012252f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_149 N_C1_M1004_g N_A_27_47#_c_508_n 0.01076f $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_150 N_C1_M1016_g N_A_27_47#_c_508_n 0.0110362f $X=1.845 $Y=0.56 $X2=0 $Y2=0
cc_151 N_C1_c_142_n N_A_27_47#_c_508_n 0.00228257f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_152 C1 N_A_27_47#_c_508_n 0.0354764f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_153 C1 N_A_27_47#_c_509_n 0.0159787f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_154 N_C1_M1016_g N_A_27_47#_c_510_n 4.70514e-19 $X=1.845 $Y=0.56 $X2=0 $Y2=0
cc_155 N_C1_M1004_g N_A_298_47#_c_548_n 0.00361103f $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_156 N_C1_M1016_g N_A_298_47#_c_548_n 0.0035946f $X=1.845 $Y=0.56 $X2=0 $Y2=0
cc_157 N_C1_M1016_g N_A_298_47#_c_547_n 0.0109617f $X=1.845 $Y=0.56 $X2=0 $Y2=0
cc_158 N_C1_M1004_g N_VGND_c_623_n 0.00428334f $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_159 N_C1_M1016_g N_VGND_c_623_n 0.0035787f $X=1.845 $Y=0.56 $X2=0 $Y2=0
cc_160 N_C1_M1004_g N_VGND_c_626_n 0.0060499f $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_161 N_C1_M1016_g N_VGND_c_626_n 0.00659231f $X=1.845 $Y=0.56 $X2=0 $Y2=0
cc_162 N_B1_M1019_g N_A2_M1009_g 0.0190118f $X=3.26 $Y=0.56 $X2=0 $Y2=0
cc_163 N_B1_c_194_n N_A2_c_246_n 0.0190118f $X=3.185 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B1_c_194_n A2 0.00232655f $X=3.185 $Y=1.16 $X2=0 $Y2=0
cc_165 B1 A2 0.0212995f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_166 N_B1_M1002_g N_VPWR_c_332_n 0.0106233f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_167 N_B1_M1014_g N_VPWR_c_332_n 6.21637e-19 $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_168 N_B1_M1002_g N_VPWR_c_333_n 6.32823e-19 $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_169 N_B1_M1014_g N_VPWR_c_333_n 0.0119128f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_170 N_B1_M1002_g N_VPWR_c_337_n 0.00486043f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B1_M1014_g N_VPWR_c_337_n 0.00486043f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_172 N_B1_M1002_g N_VPWR_c_328_n 0.00822531f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B1_M1014_g N_VPWR_c_328_n 0.00822531f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B1_M1002_g N_Y_c_429_n 0.0140854f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_175 B1 N_Y_c_429_n 0.0122739f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_176 N_B1_M1014_g N_Y_c_414_n 0.0161676f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B1_c_192_n N_Y_c_414_n 0.00247631f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B1_c_194_n N_Y_c_414_n 0.00450354f $X=3.185 $Y=1.16 $X2=0 $Y2=0
cc_179 B1 N_Y_c_414_n 0.041664f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_180 N_B1_c_193_n N_Y_c_441_n 7.32538e-19 $X=2.63 $Y=1.16 $X2=0 $Y2=0
cc_181 B1 N_Y_c_441_n 0.0146661f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_182 N_B1_M1013_g N_A_27_47#_c_510_n 0.00121964f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_183 N_B1_c_191_n N_A_27_47#_c_510_n 0.002092f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_184 B1 N_A_27_47#_c_510_n 0.00570112f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_185 N_B1_M1013_g N_A_298_47#_c_551_n 0.00266128f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_186 N_B1_M1019_g N_A_298_47#_c_551_n 0.00365488f $X=3.26 $Y=0.56 $X2=0 $Y2=0
cc_187 N_B1_M1013_g N_A_298_47#_c_547_n 0.00969765f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_188 N_B1_c_191_n N_A_298_47#_c_547_n 0.00374393f $X=2.35 $Y=1.16 $X2=0 $Y2=0
cc_189 B1 N_A_298_47#_c_547_n 0.00482211f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_190 N_B1_M1013_g N_A_497_47#_c_573_n 0.00940449f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_191 N_B1_M1019_g N_A_497_47#_c_573_n 0.0125951f $X=3.26 $Y=0.56 $X2=0 $Y2=0
cc_192 N_B1_c_193_n N_A_497_47#_c_573_n 0.00752369f $X=2.63 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B1_c_194_n N_A_497_47#_c_573_n 0.00219309f $X=3.185 $Y=1.16 $X2=0 $Y2=0
cc_194 B1 N_A_497_47#_c_573_n 0.0363106f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_195 N_B1_M1019_g N_VGND_c_621_n 0.00147382f $X=3.26 $Y=0.56 $X2=0 $Y2=0
cc_196 N_B1_M1013_g N_VGND_c_623_n 0.00357877f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_197 N_B1_M1019_g N_VGND_c_623_n 0.00416331f $X=3.26 $Y=0.56 $X2=0 $Y2=0
cc_198 N_B1_M1013_g N_VGND_c_626_n 0.00662861f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_199 N_B1_M1019_g N_VGND_c_626_n 0.00585646f $X=3.26 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A2_M1018_g N_A1_M1010_g 0.0178562f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A2_M1011_g N_A1_M1001_g 0.0178562f $X=4.12 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A2_c_248_n N_A1_c_291_n 0.0178562f $X=4.12 $Y=1.16 $X2=0 $Y2=0
cc_203 A2 N_A1_c_291_n 0.00256167f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_204 A2 A1 0.0212974f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_205 N_A2_M1003_g N_VPWR_c_333_n 0.00219786f $X=3.69 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A2_M1003_g N_VPWR_c_338_n 0.00357877f $X=3.69 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A2_M1011_g N_VPWR_c_338_n 0.00357877f $X=4.12 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A2_M1003_g N_VPWR_c_328_n 0.00657863f $X=3.69 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A2_M1011_g N_VPWR_c_328_n 0.00530427f $X=4.12 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A2_M1003_g N_Y_c_414_n 0.0141755f $X=3.69 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A2_c_247_n N_Y_c_414_n 7.21881e-19 $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_212 A2 N_Y_c_414_n 0.0444107f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_213 N_A2_M1003_g N_A_664_297#_c_476_n 0.0102895f $X=3.69 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A2_M1011_g N_A_664_297#_c_476_n 0.0128422f $X=4.12 $Y=1.985 $X2=0 $Y2=0
cc_215 A2 N_A_664_297#_c_478_n 0.0148233f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A2_M1009_g N_A_298_47#_c_551_n 3.52846e-19 $X=3.69 $Y=0.56 $X2=0 $Y2=0
cc_217 N_A2_M1009_g N_A_497_47#_c_580_n 0.0112467f $X=3.69 $Y=0.56 $X2=0 $Y2=0
cc_218 N_A2_M1018_g N_A_497_47#_c_580_n 0.0112467f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A2_c_247_n N_A_497_47#_c_580_n 0.00219309f $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_220 A2 N_A_497_47#_c_580_n 0.0316718f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_221 A2 N_A_497_47#_c_584_n 0.0116243f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_222 A2 N_A_497_47#_c_585_n 0.0116243f $X=4.285 $Y=1.105 $X2=0 $Y2=0
cc_223 N_A2_M1009_g N_VGND_c_621_n 0.00861335f $X=3.69 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A2_M1018_g N_VGND_c_621_n 0.00746783f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A2_M1018_g N_VGND_c_622_n 8.40876e-19 $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A2_M1009_g N_VGND_c_623_n 0.00355956f $X=3.69 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A2_M1018_g N_VGND_c_624_n 0.00355956f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A2_M1009_g N_VGND_c_626_n 0.00422417f $X=3.69 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A2_M1018_g N_VGND_c_626_n 0.00422417f $X=4.12 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A1_M1001_g N_VPWR_c_334_n 0.00285012f $X=4.55 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_M1008_g N_VPWR_c_334_n 0.0120017f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A1_M1001_g N_VPWR_c_338_n 0.00547432f $X=4.55 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_M1008_g N_VPWR_c_339_n 0.00486043f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A1_M1001_g N_VPWR_c_328_n 0.00971502f $X=4.55 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A1_M1008_g N_VPWR_c_328_n 0.00921385f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A1_M1001_g N_A_664_297#_c_478_n 0.00112604f $X=4.55 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A1_M1001_g N_A_664_297#_c_480_n 0.00950277f $X=4.55 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A1_M1008_g N_A_664_297#_c_480_n 4.50034e-19 $X=4.98 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A1_M1001_g N_A_664_297#_c_482_n 0.013047f $X=4.55 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A1_M1008_g N_A_664_297#_c_482_n 0.0144594f $X=4.98 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A1_c_292_n N_A_664_297#_c_482_n 6.38939e-19 $X=4.905 $Y=1.16 $X2=0
+ $Y2=0
cc_242 A1 N_A_664_297#_c_482_n 0.0466417f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_243 N_A1_M1010_g N_A_497_47#_c_586_n 0.0132299f $X=4.55 $Y=0.56 $X2=0 $Y2=0
cc_244 N_A1_M1015_g N_A_497_47#_c_586_n 0.0133929f $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_245 N_A1_c_292_n N_A_497_47#_c_586_n 0.0021949f $X=4.905 $Y=1.16 $X2=0 $Y2=0
cc_246 A1 N_A_497_47#_c_586_n 0.0218843f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_247 A1 N_A_497_47#_c_574_n 0.0214986f $X=5.205 $Y=1.105 $X2=0 $Y2=0
cc_248 N_A1_M1010_g N_VGND_c_621_n 8.4229e-19 $X=4.55 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A1_M1010_g N_VGND_c_622_n 0.00741718f $X=4.55 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A1_M1015_g N_VGND_c_622_n 0.0118588f $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_251 N_A1_M1010_g N_VGND_c_624_n 0.00355356f $X=4.55 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A1_M1015_g N_VGND_c_625_n 0.00355356f $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A1_M1010_g N_VGND_c_626_n 0.00421393f $X=4.55 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A1_M1015_g N_VGND_c_626_n 0.00521419f $X=4.98 $Y=0.56 $X2=0 $Y2=0
cc_255 N_VPWR_c_328_n N_Y_M1005_s 0.00379452f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_256 N_VPWR_c_328_n N_Y_M1000_d 0.00535672f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_257 N_VPWR_c_328_n N_Y_M1002_d 0.00570388f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_258 N_VPWR_c_328_n N_Y_M1003_s 0.00224864f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_259 N_VPWR_M1017_d N_Y_c_416_n 0.00353353f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_260 N_VPWR_c_331_n N_Y_c_416_n 0.0170777f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_261 N_VPWR_c_336_n N_Y_c_452_n 0.0124538f $X=1.895 $Y=2.72 $X2=0 $Y2=0
cc_262 N_VPWR_c_328_n N_Y_c_452_n 0.00724021f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_263 N_VPWR_M1012_s N_Y_c_429_n 0.00505842f $X=1.92 $Y=1.485 $X2=0 $Y2=0
cc_264 N_VPWR_c_332_n N_Y_c_429_n 0.0167051f $X=2.06 $Y=2 $X2=0 $Y2=0
cc_265 N_VPWR_c_337_n N_Y_c_456_n 0.012099f $X=2.755 $Y=2.72 $X2=0 $Y2=0
cc_266 N_VPWR_c_328_n N_Y_c_456_n 0.00684987f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_267 N_VPWR_M1014_s N_Y_c_414_n 0.00476073f $X=2.78 $Y=1.485 $X2=0 $Y2=0
cc_268 N_VPWR_c_333_n N_Y_c_414_n 0.0220026f $X=2.92 $Y=2 $X2=0 $Y2=0
cc_269 N_VPWR_c_335_n Y 0.0156896f $X=1.035 $Y=2.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_328_n Y 0.00975383f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_271 N_VPWR_c_328_n N_A_664_297#_M1003_d 0.00238016f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_272 N_VPWR_c_328_n N_A_664_297#_M1011_d 0.00223235f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_328_n N_A_664_297#_M1008_d 0.00513186f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_333_n N_A_664_297#_c_474_n 0.0138017f $X=2.92 $Y=2 $X2=0 $Y2=0
cc_275 N_VPWR_c_338_n N_A_664_297#_c_474_n 0.0177819f $X=4.67 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_328_n N_A_664_297#_c_474_n 0.00999318f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_333_n N_A_664_297#_c_475_n 0.0295518f $X=2.92 $Y=2 $X2=0 $Y2=0
cc_278 N_VPWR_c_338_n N_A_664_297#_c_476_n 0.0363338f $X=4.67 $Y=2.72 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_328_n N_A_664_297#_c_476_n 0.0235f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_338_n N_A_664_297#_c_480_n 0.0157932f $X=4.67 $Y=2.72 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_328_n N_A_664_297#_c_480_n 0.00982628f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_282 N_VPWR_M1001_s N_A_664_297#_c_482_n 0.00339101f $X=4.625 $Y=1.485 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_334_n N_A_664_297#_c_482_n 0.0152916f $X=4.765 $Y=2.02 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_339_n N_A_664_297#_c_499_n 0.0177595f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_328_n N_A_664_297#_c_499_n 0.00993603f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_286 N_Y_c_414_n N_A_664_297#_M1003_d 0.00650415f $X=3.815 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_287 N_Y_c_414_n N_A_664_297#_c_475_n 0.0199984f $X=3.815 $Y=1.58 $X2=0 $Y2=0
cc_288 N_Y_M1003_s N_A_664_297#_c_476_n 0.00333513f $X=3.765 $Y=1.485 $X2=0
+ $Y2=0
cc_289 N_Y_c_414_n N_A_664_297#_c_476_n 0.00354701f $X=3.815 $Y=1.58 $X2=0 $Y2=0
cc_290 N_Y_c_466_p N_A_664_297#_c_476_n 0.0126975f $X=3.905 $Y=1.9 $X2=0 $Y2=0
cc_291 N_Y_M1006_s N_A_27_47#_c_513_n 0.00324574f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_292 N_Y_c_413_n N_A_27_47#_c_513_n 0.0160586f $X=0.77 $Y=0.7 $X2=0 $Y2=0
cc_293 N_Y_c_429_n N_A_27_47#_c_508_n 0.00323264f $X=2.395 $Y=1.58 $X2=0 $Y2=0
cc_294 N_Y_c_413_n N_A_27_47#_c_509_n 0.00697079f $X=0.77 $Y=0.7 $X2=0 $Y2=0
cc_295 N_Y_c_429_n N_A_27_47#_c_510_n 0.00709456f $X=2.395 $Y=1.58 $X2=0 $Y2=0
cc_296 N_Y_c_414_n N_A_497_47#_c_573_n 0.00421852f $X=3.815 $Y=1.58 $X2=0 $Y2=0
cc_297 N_Y_M1006_s N_VGND_c_626_n 0.00225025f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_298 N_A_664_297#_c_478_n N_A_497_47#_c_586_n 5.9024e-19 $X=4.37 $Y=1.685
+ $X2=0 $Y2=0
cc_299 N_A_664_297#_c_482_n N_A_497_47#_c_586_n 0.00268557f $X=5.1 $Y=1.6 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_508_n N_A_298_47#_M1004_s 0.00172391f $X=1.925 $Y=0.82
+ $X2=-0.19 $Y2=-0.24
cc_301 N_A_27_47#_c_508_n N_A_298_47#_c_548_n 0.0138931f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1016_d N_A_298_47#_c_547_n 0.00599456f $X=1.92 $Y=0.235 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_508_n N_A_298_47#_c_547_n 0.00574729f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_510_n N_A_298_47#_c_547_n 0.0211074f $X=2.09 $Y=0.705 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_510_n N_A_497_47#_c_573_n 0.0159254f $X=2.09 $Y=0.705 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_538_p N_VGND_c_623_n 0.0171682f $X=0.305 $Y=0.445 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_513_n N_VGND_c_623_n 0.0474634f $X=1.115 $Y=0.352 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_508_n N_VGND_c_623_n 0.00200065f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_M1006_d N_VGND_c_626_n 0.00418036f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_M1007_d N_VGND_c_626_n 0.00245457f $X=1.06 $Y=0.235 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_M1016_d N_VGND_c_626_n 0.0023804f $X=1.92 $Y=0.235 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_538_p N_VGND_c_626_n 0.00995879f $X=0.305 $Y=0.445 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_513_n N_VGND_c_626_n 0.0309382f $X=1.115 $Y=0.352 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_508_n N_VGND_c_626_n 0.00461299f $X=1.925 $Y=0.82 $X2=0
+ $Y2=0
cc_315 N_A_298_47#_c_547_n N_A_497_47#_M1013_d 0.00520158f $X=2.88 $Y=0.37
+ $X2=-0.19 $Y2=-0.24
cc_316 N_A_298_47#_M1013_s N_A_497_47#_c_573_n 0.00348416f $X=2.905 $Y=0.235
+ $X2=0 $Y2=0
cc_317 N_A_298_47#_c_551_n N_A_497_47#_c_573_n 0.0150881f $X=3.045 $Y=0.36 $X2=0
+ $Y2=0
cc_318 N_A_298_47#_c_547_n N_A_497_47#_c_573_n 0.0212385f $X=2.88 $Y=0.37 $X2=0
+ $Y2=0
cc_319 N_A_298_47#_c_551_n N_VGND_c_621_n 0.0034179f $X=3.045 $Y=0.36 $X2=0
+ $Y2=0
cc_320 N_A_298_47#_c_548_n N_VGND_c_623_n 0.0166343f $X=1.775 $Y=0.35 $X2=0
+ $Y2=0
cc_321 N_A_298_47#_c_547_n N_VGND_c_623_n 0.084875f $X=2.88 $Y=0.37 $X2=0 $Y2=0
cc_322 N_A_298_47#_M1004_s N_VGND_c_626_n 0.00223231f $X=1.49 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_A_298_47#_M1013_s N_VGND_c_626_n 0.00223258f $X=2.905 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_A_298_47#_c_548_n N_VGND_c_626_n 0.0112629f $X=1.775 $Y=0.35 $X2=0
+ $Y2=0
cc_325 N_A_298_47#_c_547_n N_VGND_c_626_n 0.0520211f $X=2.88 $Y=0.37 $X2=0 $Y2=0
cc_326 N_A_497_47#_c_580_n N_VGND_M1009_s 0.00348016f $X=4.24 $Y=0.747 $X2=-0.19
+ $Y2=-0.24
cc_327 N_A_497_47#_c_586_n N_VGND_M1010_d 0.00348156f $X=5.1 $Y=0.745 $X2=0
+ $Y2=0
cc_328 N_A_497_47#_c_580_n N_VGND_c_621_n 0.0161999f $X=4.24 $Y=0.747 $X2=0
+ $Y2=0
cc_329 N_A_497_47#_c_586_n N_VGND_c_622_n 0.0162037f $X=5.1 $Y=0.745 $X2=0 $Y2=0
cc_330 N_A_497_47#_c_573_n N_VGND_c_623_n 0.00237525f $X=3.38 $Y=0.747 $X2=0
+ $Y2=0
cc_331 N_A_497_47#_c_604_p N_VGND_c_623_n 0.00711149f $X=3.47 $Y=0.575 $X2=0
+ $Y2=0
cc_332 N_A_497_47#_c_580_n N_VGND_c_623_n 0.00236596f $X=4.24 $Y=0.747 $X2=0
+ $Y2=0
cc_333 N_A_497_47#_c_580_n N_VGND_c_624_n 0.00236596f $X=4.24 $Y=0.747 $X2=0
+ $Y2=0
cc_334 N_A_497_47#_c_607_p N_VGND_c_624_n 0.00711149f $X=4.335 $Y=0.575 $X2=0
+ $Y2=0
cc_335 N_A_497_47#_c_586_n N_VGND_c_624_n 0.00239711f $X=5.1 $Y=0.745 $X2=0
+ $Y2=0
cc_336 N_A_497_47#_c_586_n N_VGND_c_625_n 0.00240362f $X=5.1 $Y=0.745 $X2=0
+ $Y2=0
cc_337 N_A_497_47#_c_574_n N_VGND_c_625_n 0.0131614f $X=5.255 $Y=0.58 $X2=0
+ $Y2=0
cc_338 N_A_497_47#_M1013_d N_VGND_c_626_n 0.00218346f $X=2.485 $Y=0.235 $X2=0
+ $Y2=0
cc_339 N_A_497_47#_M1019_d N_VGND_c_626_n 0.00267362f $X=3.335 $Y=0.235 $X2=0
+ $Y2=0
cc_340 N_A_497_47#_M1018_d N_VGND_c_626_n 0.00267034f $X=4.195 $Y=0.235 $X2=0
+ $Y2=0
cc_341 N_A_497_47#_M1015_s N_VGND_c_626_n 0.00297223f $X=5.055 $Y=0.235 $X2=0
+ $Y2=0
cc_342 N_A_497_47#_c_573_n N_VGND_c_626_n 0.00567289f $X=3.38 $Y=0.747 $X2=0
+ $Y2=0
cc_343 N_A_497_47#_c_604_p N_VGND_c_626_n 0.0067341f $X=3.47 $Y=0.575 $X2=0
+ $Y2=0
cc_344 N_A_497_47#_c_580_n N_VGND_c_626_n 0.00969868f $X=4.24 $Y=0.747 $X2=0
+ $Y2=0
cc_345 N_A_497_47#_c_607_p N_VGND_c_626_n 0.0067341f $X=4.335 $Y=0.575 $X2=0
+ $Y2=0
cc_346 N_A_497_47#_c_586_n N_VGND_c_626_n 0.00977124f $X=5.1 $Y=0.745 $X2=0
+ $Y2=0
cc_347 N_A_497_47#_c_574_n N_VGND_c_626_n 0.011928f $X=5.255 $Y=0.58 $X2=0 $Y2=0

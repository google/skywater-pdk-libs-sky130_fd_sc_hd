* File: sky130_fd_sc_hd__o211a_4.spice
* Created: Thu Aug 27 14:34:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o211a_4.spice.pex"
.subckt sky130_fd_sc_hd__o211a_4  VNB VPB B1 C1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_79_21#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_79_21#_M1013_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1013_d N_A_79_21#_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A_79_21#_M1021_g N_X_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.19175 AS=0.08775 PD=1.89 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 A_748_47# N_B1_M1000_g N_A_474_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.17225 PD=0.86 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1017 N_A_79_21#_M1017_d N_C1_M1017_g A_748_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.144625 AS=0.06825 PD=1.095 PS=0.86 NRD=12.912 NRS=9.228 M=1 R=4.33333
+ SA=75000.5 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1011 N_A_79_21#_M1017_d N_C1_M1011_g A_557_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.144625 AS=0.091 PD=1.095 PS=0.93 NRD=17.532 NRS=15.684 M=1 R=4.33333
+ SA=75001.1 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1022 A_557_47# N_B1_M1022_g N_A_474_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.104 PD=0.93 PS=0.97 NRD=15.684 NRS=4.608 M=1 R=4.33333
+ SA=75001.6 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A1_M1014_g N_A_474_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.104 PD=1.04 PS=0.97 NRD=7.38 NRS=2.76 M=1 R=4.33333 SA=75002
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1001 N_A_474_47#_M1001_d N_A2_M1001_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.12675 PD=0.93 PS=1.04 NRD=0 NRS=12.912 M=1 R=4.33333 SA=75002.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1002 N_A_474_47#_M1001_d N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1002_s N_A1_M1015_g N_A_474_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1004_d N_A_79_21#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1008 N_X_M1004_d N_A_79_21#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1018 N_X_M1018_d N_A_79_21#_M1018_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75004.4
+ A=0.15 P=2.3 MULT=1
MM1020 N_X_M1018_d N_A_79_21#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5 SB=75004
+ A=0.15 P=2.3 MULT=1
MM1006 N_A_79_21#_M1006_d N_B1_M1006_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2525 AS=0.14 PD=1.505 PS=1.28 NRD=19.7 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_79_21#_M1006_d N_C1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2525 AS=0.14 PD=1.505 PS=1.28 NRD=24.6053 NRS=0 M=1 R=6.66667 SA=75002.6
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1007 N_A_79_21#_M1007_d N_C1_M1007_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.14 PD=1.39 PS=1.28 NRD=13.7703 NRS=0 M=1 R=6.66667 SA=75003
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1009 N_A_79_21#_M1007_d N_B1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.16 PD=1.39 PS=1.32 NRD=7.8603 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1009_s N_A1_M1005_g A_950_297# VPB PHIGHVT L=0.15 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=7.8603 NRS=16.7253 M=1 R=6.66667 SA=75004
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1019 A_950_297# N_A2_M1019_g N_A_79_21#_M1019_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75004.4 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1023 A_1122_297# N_A2_M1023_g N_A_79_21#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75004.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g A_1122_297# VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=16.7253 M=1 R=6.66667 SA=75005.3 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.9461 P=16.85
c_707 A_950_297# 0 1.15267e-19 $X=4.75 $Y=1.485
*
.include "sky130_fd_sc_hd__o211a_4.spice.SKY130_FD_SC_HD__O211A_4.pxi"
*
.ends
*
*

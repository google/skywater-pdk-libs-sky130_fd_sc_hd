* NGSPICE file created from sky130_fd_sc_hd__and4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
M1000 VPWR a_27_47# X VPB phighvt w=1e+06u l=150000u
+  ad=1.43e+12p pd=1.286e+07u as=5.4e+11p ps=5.08e+06u
M1001 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=5.5575e+11p ps=5.61e+06u
M1002 a_285_47# C a_188_47# VNB nshort w=650000u l=150000u
+  ad=2.8275e+11p pd=2.17e+06u as=2.1775e+11p ps=1.97e+06u
M1003 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=7e+11p ps=5.4e+06u
M1006 VPWR a_27_47# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_188_47# B a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.5925e+11p ps=1.79e+06u
M1008 a_27_47# C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D a_285_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR D a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_109_47# A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1015 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__ha_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 1.075000 4.380000 1.245000 ;
        RECT 4.210000 1.245000 4.380000 1.505000 ;
        RECT 4.210000 1.505000 6.810000 1.675000 ;
        RECT 5.625000 0.995000 5.795000 1.505000 ;
        RECT 6.580000 0.995000 7.055000 1.325000 ;
        RECT 6.580000 1.325000 6.810000 1.505000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.550000 0.995000 5.455000 1.165000 ;
        RECT 4.550000 1.165000 4.720000 1.325000 ;
        RECT 5.285000 0.730000 6.315000 0.825000 ;
        RECT 5.285000 0.825000 5.535000 0.845000 ;
        RECT 5.285000 0.845000 5.495000 0.875000 ;
        RECT 5.285000 0.875000 5.455000 0.995000 ;
        RECT 5.295000 0.720000 6.315000 0.730000 ;
        RECT 5.310000 0.710000 6.315000 0.720000 ;
        RECT 5.320000 0.695000 6.315000 0.710000 ;
        RECT 5.335000 0.675000 6.315000 0.695000 ;
        RECT 5.345000 0.655000 6.315000 0.675000 ;
        RECT 6.085000 0.825000 6.315000 1.325000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595000 0.315000 7.845000 0.735000 ;
        RECT 7.595000 0.735000 8.685000 0.905000 ;
        RECT 7.595000 1.415000 8.685000 1.585000 ;
        RECT 7.595000 1.585000 7.765000 2.415000 ;
        RECT 8.405000 0.315000 8.685000 0.735000 ;
        RECT 8.405000 0.905000 8.685000 1.415000 ;
        RECT 8.405000 1.585000 8.685000 2.415000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.315000 0.845000 1.065000 ;
        RECT 0.515000 1.065000 1.550000 1.335000 ;
        RECT 0.515000 1.335000 0.845000 2.415000 ;
        RECT 1.355000 0.315000 1.685000 0.825000 ;
        RECT 1.355000 0.825000 1.550000 1.065000 ;
        RECT 1.355000 1.335000 1.550000 1.565000 ;
        RECT 1.355000 1.565000 1.685000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.200000 0.085000 ;
        RECT 0.135000  0.085000 0.345000 0.885000 ;
        RECT 1.015000  0.085000 1.185000 0.885000 ;
        RECT 1.855000  0.085000 2.095000 0.885000 ;
        RECT 3.555000  0.085000 3.910000 0.465000 ;
        RECT 4.420000  0.085000 4.750000 0.465000 ;
        RECT 5.385000  0.085000 5.715000 0.465000 ;
        RECT 7.055000  0.085000 7.385000 0.465000 ;
        RECT 8.015000  0.085000 8.225000 0.565000 ;
        RECT 8.855000  0.085000 9.065000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.200000 2.805000 ;
        RECT 0.135000 1.495000 0.345000 2.635000 ;
        RECT 1.015000 1.515000 1.185000 2.635000 ;
        RECT 1.855000 1.495000 2.365000 2.635000 ;
        RECT 3.190000 2.105000 3.360000 2.635000 ;
        RECT 5.240000 2.205000 5.570000 2.635000 ;
        RECT 6.175000 2.205000 6.505000 2.635000 ;
        RECT 7.055000 2.205000 7.385000 2.635000 ;
        RECT 7.935000 1.755000 8.225000 2.635000 ;
        RECT 8.855000 1.495000 9.065000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.720000 1.075000 2.750000 1.245000 ;
      RECT 2.270000 0.305000 3.385000 0.475000 ;
      RECT 2.580000 0.645000 3.045000 0.815000 ;
      RECT 2.580000 0.815000 2.750000 1.075000 ;
      RECT 2.580000 1.245000 2.750000 1.765000 ;
      RECT 2.580000 1.765000 3.700000 1.935000 ;
      RECT 2.770000 1.935000 2.940000 2.355000 ;
      RECT 2.920000 0.995000 3.090000 1.425000 ;
      RECT 2.920000 1.425000 4.040000 1.595000 ;
      RECT 3.215000 0.475000 3.385000 0.645000 ;
      RECT 3.215000 0.645000 5.115000 0.815000 ;
      RECT 3.530000 1.935000 3.700000 2.205000 ;
      RECT 3.530000 2.205000 4.330000 2.375000 ;
      RECT 3.870000 1.595000 4.040000 1.855000 ;
      RECT 3.870000 1.855000 7.395000 2.025000 ;
      RECT 4.080000 0.345000 4.250000 0.645000 ;
      RECT 4.920000 0.255000 5.190000 0.585000 ;
      RECT 4.920000 0.585000 5.115000 0.645000 ;
      RECT 5.835000 2.025000 6.005000 2.355000 ;
      RECT 6.175000 0.295000 6.875000 0.465000 ;
      RECT 6.675000 2.025000 6.845000 2.355000 ;
      RECT 6.705000 0.465000 6.875000 0.645000 ;
      RECT 6.705000 0.645000 7.395000 0.815000 ;
      RECT 7.225000 0.815000 7.395000 1.075000 ;
      RECT 7.225000 1.075000 8.225000 1.245000 ;
      RECT 7.225000 1.245000 7.395000 1.855000 ;
  END
END sky130_fd_sc_hd__ha_4

* File: sky130_fd_sc_hd__o22a_4.pxi.spice
* Created: Thu Aug 27 14:37:45 2020
* 
x_PM_SKY130_FD_SC_HD__O22A_4%A_96_21# N_A_96_21#_M1022_d N_A_96_21#_M1018_d
+ N_A_96_21#_M1009_s N_A_96_21#_M1011_s N_A_96_21#_c_110_n N_A_96_21#_M1000_g
+ N_A_96_21#_M1003_g N_A_96_21#_c_111_n N_A_96_21#_M1004_g N_A_96_21#_M1006_g
+ N_A_96_21#_c_112_n N_A_96_21#_M1005_g N_A_96_21#_M1007_g N_A_96_21#_c_113_n
+ N_A_96_21#_M1017_g N_A_96_21#_M1019_g N_A_96_21#_c_114_n N_A_96_21#_c_115_n
+ N_A_96_21#_c_116_n N_A_96_21#_c_117_n N_A_96_21#_c_132_p N_A_96_21#_c_168_p
+ N_A_96_21#_c_118_n N_A_96_21#_c_119_n N_A_96_21#_c_134_p N_A_96_21#_c_120_n
+ N_A_96_21#_c_121_n N_A_96_21#_c_139_p N_A_96_21#_c_163_p N_A_96_21#_c_122_n
+ PM_SKY130_FD_SC_HD__O22A_4%A_96_21#
x_PM_SKY130_FD_SC_HD__O22A_4%B1 N_B1_c_263_n N_B1_M1022_g N_B1_M1013_g
+ N_B1_c_264_n N_B1_M1023_g N_B1_M1021_g N_B1_c_271_n N_B1_c_265_n N_B1_c_266_n
+ B1 N_B1_c_267_n N_B1_c_268_n PM_SKY130_FD_SC_HD__O22A_4%B1
x_PM_SKY130_FD_SC_HD__O22A_4%B2 N_B2_c_349_n N_B2_M1001_g N_B2_M1009_g
+ N_B2_c_350_n N_B2_M1018_g N_B2_M1010_g B2 N_B2_c_352_n
+ PM_SKY130_FD_SC_HD__O22A_4%B2
x_PM_SKY130_FD_SC_HD__O22A_4%A1 N_A1_c_390_n N_A1_M1012_g N_A1_M1002_g
+ N_A1_c_391_n N_A1_M1016_g N_A1_M1008_g N_A1_c_392_n N_A1_c_393_n N_A1_c_402_n
+ N_A1_c_403_n N_A1_c_394_n N_A1_c_395_n A1 N_A1_c_397_n A1
+ PM_SKY130_FD_SC_HD__O22A_4%A1
x_PM_SKY130_FD_SC_HD__O22A_4%A2 N_A2_c_476_n N_A2_M1014_g N_A2_M1011_g
+ N_A2_c_477_n N_A2_M1015_g N_A2_M1020_g A2 N_A2_c_478_n
+ PM_SKY130_FD_SC_HD__O22A_4%A2
x_PM_SKY130_FD_SC_HD__O22A_4%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_M1019_d
+ N_VPWR_M1021_s N_VPWR_M1008_s N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n VPWR
+ N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_524_n N_VPWR_c_536_n
+ N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n PM_SKY130_FD_SC_HD__O22A_4%VPWR
x_PM_SKY130_FD_SC_HD__O22A_4%X N_X_M1000_d N_X_M1005_d N_X_M1003_s N_X_M1007_s
+ N_X_c_615_n N_X_c_616_n N_X_c_620_n N_X_c_621_n N_X_c_629_n N_X_c_663_n
+ N_X_c_622_n N_X_c_617_n N_X_c_645_n N_X_c_667_n N_X_c_618_n N_X_c_623_n X
+ PM_SKY130_FD_SC_HD__O22A_4%X
x_PM_SKY130_FD_SC_HD__O22A_4%A_566_297# N_A_566_297#_M1013_d
+ N_A_566_297#_M1010_d N_A_566_297#_c_690_n N_A_566_297#_c_694_n
+ N_A_566_297#_c_695_n PM_SKY130_FD_SC_HD__O22A_4%A_566_297#
x_PM_SKY130_FD_SC_HD__O22A_4%A_918_297# N_A_918_297#_M1002_d
+ N_A_918_297#_M1020_d N_A_918_297#_c_710_n N_A_918_297#_c_717_n
+ N_A_918_297#_c_713_n PM_SKY130_FD_SC_HD__O22A_4%A_918_297#
x_PM_SKY130_FD_SC_HD__O22A_4%VGND N_VGND_M1000_s N_VGND_M1004_s N_VGND_M1017_s
+ N_VGND_M1012_s N_VGND_M1015_s N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n
+ N_VGND_c_729_n N_VGND_c_730_n N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n
+ N_VGND_c_734_n N_VGND_c_735_n N_VGND_c_736_n VGND N_VGND_c_737_n
+ N_VGND_c_738_n N_VGND_c_739_n N_VGND_c_740_n N_VGND_c_741_n
+ PM_SKY130_FD_SC_HD__O22A_4%VGND
x_PM_SKY130_FD_SC_HD__O22A_4%A_484_47# N_A_484_47#_M1022_s N_A_484_47#_M1001_s
+ N_A_484_47#_M1023_s N_A_484_47#_M1014_d N_A_484_47#_M1016_d
+ N_A_484_47#_c_826_n N_A_484_47#_c_848_n N_A_484_47#_c_849_n
+ N_A_484_47#_c_827_n N_A_484_47#_c_828_n N_A_484_47#_c_857_n
+ N_A_484_47#_c_829_n N_A_484_47#_c_830_n N_A_484_47#_c_831_n
+ PM_SKY130_FD_SC_HD__O22A_4%A_484_47#
cc_1 VNB N_A_96_21#_c_110_n 0.0191784f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_2 VNB N_A_96_21#_c_111_n 0.0157977f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_3 VNB N_A_96_21#_c_112_n 0.0157964f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.995
cc_4 VNB N_A_96_21#_c_113_n 0.0190654f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=0.995
cc_5 VNB N_A_96_21#_c_114_n 6.30857e-19 $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.175
cc_6 VNB N_A_96_21#_c_115_n 6.59699e-19 $X=-0.19 $Y=-0.24 $X2=2.065 $Y2=1.785
cc_7 VNB N_A_96_21#_c_116_n 0.00475766f $X=-0.19 $Y=-0.24 $X2=2.085 $Y2=1.075
cc_8 VNB N_A_96_21#_c_117_n 0.00191669f $X=-0.19 $Y=-0.24 $X2=2.23 $Y2=0.82
cc_9 VNB N_A_96_21#_c_118_n 0.00259604f $X=-0.19 $Y=-0.24 $X2=2.545 $Y2=0.775
cc_10 VNB N_A_96_21#_c_119_n 0.00967441f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=0.73
cc_11 VNB N_A_96_21#_c_120_n 0.00424408f $X=-0.19 $Y=-0.24 $X2=2.065 $Y2=1.175
cc_12 VNB N_A_96_21#_c_121_n 0.00991332f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=0.775
cc_13 VNB N_A_96_21#_c_122_n 0.0689431f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=1.16
cc_14 VNB N_B1_c_263_n 0.0198931f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=0.235
cc_15 VNB N_B1_c_264_n 0.0170683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_c_265_n 0.00349127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B1_c_266_n 0.0196886f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_18 VNB N_B1_c_267_n 0.0241314f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_19 VNB N_B1_c_268_n 0.00590555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B2_c_349_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=0.235
cc_21 VNB N_B2_c_350_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB B2 0.00141292f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_23 VNB N_B2_c_352_n 0.0299865f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.56
cc_24 VNB N_A1_c_390_n 0.0169197f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=0.235
cc_25 VNB N_A1_c_391_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A1_c_392_n 0.00358781f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.985
cc_27 VNB N_A1_c_393_n 0.0192897f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.985
cc_28 VNB N_A1_c_394_n 2.72331e-19 $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.325
cc_29 VNB N_A1_c_395_n 0.00189758f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_30 VNB A1 0.0298833f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_31 VNB N_A1_c_397_n 0.0265824f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.56
cc_32 VNB N_A2_c_476_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=2.83 $Y2=0.235
cc_33 VNB N_A2_c_477_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A2_c_478_n 0.0313072f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.56
cc_35 VNB N_VPWR_c_524_n 0.269736f $X=-0.19 $Y=-0.24 $X2=5.02 $Y2=1.87
cc_36 VNB N_X_c_615_n 0.0014432f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_37 VNB N_X_c_616_n 0.00986769f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_38 VNB N_X_c_617_n 0.00440603f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.56
cc_39 VNB N_X_c_618_n 0.00222466f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_40 VNB X 0.0213229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_726_n 0.00419326f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.985
cc_42 VNB N_VGND_c_727_n 0.0169505f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.995
cc_43 VNB N_VGND_c_728_n 0.0130399f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=0.56
cc_44 VNB N_VGND_c_729_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_45 VNB N_VGND_c_730_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.56
cc_46 VNB N_VGND_c_731_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.985
cc_47 VNB N_VGND_c_732_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=0.56
cc_48 VNB N_VGND_c_733_n 0.0585747f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=1.985
cc_49 VNB N_VGND_c_734_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_735_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.175
cc_51 VNB N_VGND_c_736_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_52 VNB N_VGND_c_737_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=1.725 $Y2=1.175
cc_53 VNB N_VGND_c_738_n 0.0234308f $X=-0.19 $Y=-0.24 $X2=2.965 $Y2=0.73
cc_54 VNB N_VGND_c_739_n 0.326336f $X=-0.19 $Y=-0.24 $X2=3.805 $Y2=0.775
cc_55 VNB N_VGND_c_740_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_741_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_484_47#_c_826_n 0.00289463f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.325
cc_58 VNB N_A_484_47#_c_827_n 0.00332606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_484_47#_c_828_n 0.00807318f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=0.995
cc_60 VNB N_A_484_47#_c_829_n 0.0132865f $X=-0.19 $Y=-0.24 $X2=1.395 $Y2=1.985
cc_61 VNB N_A_484_47#_c_830_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=1.815 $Y2=0.56
cc_62 VNB N_A_484_47#_c_831_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VPB N_A_96_21#_M1003_g 0.0219695f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_64 VPB N_A_96_21#_M1006_g 0.0181176f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_65 VPB N_A_96_21#_M1007_g 0.0181312f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.985
cc_66 VPB N_A_96_21#_M1019_g 0.0218481f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.985
cc_67 VPB N_A_96_21#_c_115_n 0.0041539f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=1.785
cc_68 VPB N_A_96_21#_c_122_n 0.0103574f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.16
cc_69 VPB N_B1_M1013_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B1_M1021_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_71 VPB N_B1_c_271_n 0.00732858f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.56
cc_72 VPB N_B1_c_265_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B1_c_266_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.995
cc_74 VPB N_B1_c_267_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_75 VPB N_B1_c_268_n 0.00311667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_B2_M1009_g 0.0183531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_B2_M1010_g 0.0183545f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_78 VPB N_B2_c_352_n 0.00400363f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_79 VPB N_A1_M1002_g 0.0181129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A1_M1008_g 0.0245822f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_81 VPB N_A1_c_392_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_82 VPB N_A1_c_393_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_83 VPB N_A1_c_402_n 0.00689724f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.995
cc_84 VPB N_A1_c_403_n 2.50157e-19 $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_85 VPB N_A1_c_394_n 0.00130531f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.325
cc_86 VPB N_A1_c_397_n 0.00655427f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=0.56
cc_87 VPB N_A2_M1011_g 0.0183373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A2_M1020_g 0.0183337f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_89 VPB N_A2_c_478_n 0.00400351f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_90 VPB N_VPWR_c_525_n 0.0140014f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.325
cc_91 VPB N_VPWR_c_526_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.985
cc_92 VPB N_VPWR_c_527_n 0.0039289f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=0.56
cc_93 VPB N_VPWR_c_528_n 0.00561441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_529_n 0.00830908f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=1.325
cc_95 VPB N_VPWR_c_530_n 0.0363617f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=0.56
cc_96 VPB N_VPWR_c_531_n 0.00391723f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=0.56
cc_97 VPB N_VPWR_c_532_n 0.0163782f $X=-0.19 $Y=1.305 $X2=1.815 $Y2=1.985
cc_98 VPB N_VPWR_c_533_n 0.0349357f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=1.275
cc_99 VPB N_VPWR_c_534_n 0.0126445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_524_n 0.0565209f $X=-0.19 $Y=1.305 $X2=5.02 $Y2=1.87
cc_101 VPB N_VPWR_c_536_n 0.0047828f $X=-0.19 $Y=1.305 $X2=3.385 $Y2=1.96
cc_102 VPB N_VPWR_c_537_n 0.0163782f $X=-0.19 $Y=1.305 $X2=5.145 $Y2=1.96
cc_103 VPB N_VPWR_c_538_n 0.0222575f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.16
cc_104 VPB N_VPWR_c_539_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_105 VPB N_X_c_620_n 0.00152588f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.56
cc_106 VPB N_X_c_621_n 0.0124376f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.325
cc_107 VPB N_X_c_622_n 0.00471275f $X=-0.19 $Y=1.305 $X2=1.395 $Y2=0.995
cc_108 VPB N_X_c_623_n 0.00204415f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_109 VPB X 0.00756106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 N_A_96_21#_c_116_n N_B1_c_263_n 0.0024189f $X=2.085 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_96_21#_c_119_n N_B1_c_263_n 0.013778f $X=3.805 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_96_21#_c_115_n N_B1_M1013_g 0.00590249f $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_113 N_A_96_21#_c_132_p N_B1_M1013_g 0.0136543f $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_114 N_A_96_21#_c_119_n N_B1_c_264_n 0.00375446f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_115 N_A_96_21#_c_134_p N_B1_M1021_g 0.0119464f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_116 N_A_96_21#_M1009_s N_B1_c_271_n 0.00165831f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_117 N_A_96_21#_c_132_p N_B1_c_271_n 0.0165249f $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_118 N_A_96_21#_c_119_n N_B1_c_271_n 0.0116652f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_119 N_A_96_21#_c_134_p N_B1_c_271_n 0.0355123f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_120 N_A_96_21#_c_139_p N_B1_c_271_n 0.0120079f $X=3.385 $Y=1.87 $X2=0 $Y2=0
cc_121 N_A_96_21#_c_119_n N_B1_c_265_n 0.00964534f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_122 N_A_96_21#_c_119_n N_B1_c_266_n 0.00149384f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_123 N_A_96_21#_c_134_p N_B1_c_266_n 3.01349e-19 $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_124 N_A_96_21#_c_115_n N_B1_c_267_n 2.32165e-19 $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_125 N_A_96_21#_c_116_n N_B1_c_267_n 0.00245123f $X=2.085 $Y=1.075 $X2=0 $Y2=0
cc_126 N_A_96_21#_c_132_p N_B1_c_267_n 3.01349e-19 $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_127 N_A_96_21#_c_119_n N_B1_c_267_n 0.00298767f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_128 N_A_96_21#_c_120_n N_B1_c_267_n 0.00100933f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_129 N_A_96_21#_c_115_n N_B1_c_268_n 0.0267037f $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_130 N_A_96_21#_c_132_p N_B1_c_268_n 0.0326881f $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_131 N_A_96_21#_c_118_n N_B1_c_268_n 0.0436872f $X=2.545 $Y=0.775 $X2=0 $Y2=0
cc_132 N_A_96_21#_c_120_n N_B1_c_268_n 0.0169378f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_133 N_A_96_21#_c_122_n N_B1_c_268_n 0.00131745f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_96_21#_c_119_n N_B2_c_349_n 0.0112673f $X=3.805 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_96_21#_c_132_p N_B2_M1009_g 0.00924026f $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_136 N_A_96_21#_c_119_n N_B2_c_350_n 0.0109578f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_137 N_A_96_21#_c_134_p N_B2_M1010_g 0.00924026f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_138 N_A_96_21#_c_119_n B2 0.0405144f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_139 N_A_96_21#_c_119_n N_B2_c_352_n 0.00224214f $X=3.805 $Y=0.73 $X2=0 $Y2=0
cc_140 N_A_96_21#_c_134_p N_A1_M1002_g 0.0119464f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_141 N_A_96_21#_c_134_p N_A1_c_393_n 3.01349e-19 $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_142 N_A_96_21#_M1011_s N_A1_c_402_n 0.00165831f $X=5.01 $Y=1.485 $X2=0 $Y2=0
cc_143 N_A_96_21#_c_134_p N_A1_c_402_n 0.0190307f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_144 N_A_96_21#_c_163_p N_A1_c_402_n 0.0120079f $X=5.145 $Y=1.87 $X2=0 $Y2=0
cc_145 N_A_96_21#_c_134_p N_A1_c_403_n 0.0164816f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_146 N_A_96_21#_c_134_p N_A2_M1011_g 0.00924026f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_147 N_A_96_21#_c_115_n N_VPWR_M1019_d 0.00865609f $X=2.065 $Y=1.785 $X2=0
+ $Y2=0
cc_148 N_A_96_21#_c_132_p N_VPWR_M1019_d 0.0159609f $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_149 N_A_96_21#_c_168_p N_VPWR_M1019_d 0.00572923f $X=2.23 $Y=1.87 $X2=0 $Y2=0
cc_150 N_A_96_21#_c_134_p N_VPWR_M1021_s 0.0095835f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_151 N_A_96_21#_M1003_g N_VPWR_c_526_n 0.00338128f $X=0.555 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_96_21#_M1006_g N_VPWR_c_527_n 0.00157837f $X=0.975 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_96_21#_M1007_g N_VPWR_c_527_n 0.00157702f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_96_21#_c_134_p N_VPWR_c_528_n 0.0186532f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_155 N_A_96_21#_M1003_g N_VPWR_c_532_n 0.00585385f $X=0.555 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A_96_21#_M1006_g N_VPWR_c_532_n 0.00585385f $X=0.975 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_96_21#_M1009_s N_VPWR_c_524_n 0.00215227f $X=3.25 $Y=1.485 $X2=0
+ $Y2=0
cc_158 N_A_96_21#_M1011_s N_VPWR_c_524_n 0.0021603f $X=5.01 $Y=1.485 $X2=0 $Y2=0
cc_159 N_A_96_21#_M1003_g N_VPWR_c_524_n 0.0114631f $X=0.555 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_96_21#_M1006_g N_VPWR_c_524_n 0.0104367f $X=0.975 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_96_21#_M1007_g N_VPWR_c_524_n 0.0104367f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_96_21#_M1019_g N_VPWR_c_524_n 0.0117604f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_96_21#_c_132_p N_VPWR_c_524_n 0.00749156f $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_164 N_A_96_21#_c_168_p N_VPWR_c_524_n 0.00133688f $X=2.23 $Y=1.87 $X2=0 $Y2=0
cc_165 N_A_96_21#_c_134_p N_VPWR_c_524_n 0.0130817f $X=5.02 $Y=1.87 $X2=0 $Y2=0
cc_166 N_A_96_21#_M1007_g N_VPWR_c_537_n 0.00585385f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_96_21#_M1019_g N_VPWR_c_537_n 0.00585385f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_96_21#_M1019_g N_VPWR_c_538_n 0.00353572f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_96_21#_c_132_p N_VPWR_c_538_n 0.0308699f $X=3.26 $Y=1.87 $X2=0 $Y2=0
cc_170 N_A_96_21#_c_168_p N_VPWR_c_538_n 0.024545f $X=2.23 $Y=1.87 $X2=0 $Y2=0
cc_171 N_A_96_21#_c_110_n N_X_c_615_n 0.0111411f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_96_21#_c_114_n N_X_c_615_n 0.00410208f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_173 N_A_96_21#_M1003_g N_X_c_620_n 0.015729f $X=0.555 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_96_21#_c_114_n N_X_c_620_n 0.00686379f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_175 N_A_96_21#_c_110_n N_X_c_629_n 0.0108342f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_96_21#_c_111_n N_X_c_629_n 0.00621819f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_96_21#_c_112_n N_X_c_629_n 5.19281e-19 $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_96_21#_M1006_g N_X_c_622_n 0.0133439f $X=0.975 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_96_21#_M1007_g N_X_c_622_n 0.0133089f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_96_21#_M1019_g N_X_c_622_n 3.45391e-19 $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_96_21#_c_114_n N_X_c_622_n 0.0618991f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_182 N_A_96_21#_c_115_n N_X_c_622_n 0.00344747f $X=2.065 $Y=1.785 $X2=0 $Y2=0
cc_183 N_A_96_21#_c_122_n N_X_c_622_n 0.00436768f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_96_21#_c_111_n N_X_c_617_n 0.00870364f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_96_21#_c_112_n N_X_c_617_n 0.0098365f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_96_21#_c_113_n N_X_c_617_n 0.00273575f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_96_21#_c_114_n N_X_c_617_n 0.0626515f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_188 N_A_96_21#_c_117_n N_X_c_617_n 0.00808484f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_189 N_A_96_21#_c_118_n N_X_c_617_n 3.21899e-19 $X=2.545 $Y=0.775 $X2=0 $Y2=0
cc_190 N_A_96_21#_c_122_n N_X_c_617_n 0.00452472f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_96_21#_c_111_n N_X_c_645_n 5.22228e-19 $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_96_21#_c_112_n N_X_c_645_n 0.00630972f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_96_21#_c_113_n N_X_c_645_n 0.00924185f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_96_21#_c_118_n N_X_c_645_n 0.00241259f $X=2.545 $Y=0.775 $X2=0 $Y2=0
cc_195 N_A_96_21#_c_110_n N_X_c_618_n 0.00113258f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_96_21#_c_111_n N_X_c_618_n 0.00113258f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_96_21#_c_114_n N_X_c_618_n 0.0265057f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_198 N_A_96_21#_c_122_n N_X_c_618_n 0.00230227f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_96_21#_c_114_n N_X_c_623_n 0.0203891f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_200 N_A_96_21#_c_122_n N_X_c_623_n 0.00222737f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_96_21#_c_110_n X 0.0198998f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_96_21#_c_114_n X 0.0164324f $X=1.9 $Y=1.175 $X2=0 $Y2=0
cc_203 N_A_96_21#_c_132_p N_A_566_297#_M1013_d 0.00323325f $X=3.26 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_204 N_A_96_21#_c_134_p N_A_566_297#_M1010_d 0.00325521f $X=5.02 $Y=1.87 $X2=0
+ $Y2=0
cc_205 N_A_96_21#_M1009_s N_A_566_297#_c_690_n 0.00312348f $X=3.25 $Y=1.485
+ $X2=0 $Y2=0
cc_206 N_A_96_21#_c_132_p N_A_566_297#_c_690_n 0.00506389f $X=3.26 $Y=1.87 $X2=0
+ $Y2=0
cc_207 N_A_96_21#_c_134_p N_A_566_297#_c_690_n 0.00506389f $X=5.02 $Y=1.87 $X2=0
+ $Y2=0
cc_208 N_A_96_21#_c_139_p N_A_566_297#_c_690_n 0.0112811f $X=3.385 $Y=1.87 $X2=0
+ $Y2=0
cc_209 N_A_96_21#_c_132_p N_A_566_297#_c_694_n 0.0115714f $X=3.26 $Y=1.87 $X2=0
+ $Y2=0
cc_210 N_A_96_21#_c_134_p N_A_566_297#_c_695_n 0.0116461f $X=5.02 $Y=1.87 $X2=0
+ $Y2=0
cc_211 N_A_96_21#_c_134_p N_A_918_297#_M1002_d 0.00325521f $X=5.02 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_212 N_A_96_21#_M1011_s N_A_918_297#_c_710_n 0.00312348f $X=5.01 $Y=1.485
+ $X2=0 $Y2=0
cc_213 N_A_96_21#_c_134_p N_A_918_297#_c_710_n 0.00506389f $X=5.02 $Y=1.87 $X2=0
+ $Y2=0
cc_214 N_A_96_21#_c_163_p N_A_918_297#_c_710_n 0.0112811f $X=5.145 $Y=1.87 $X2=0
+ $Y2=0
cc_215 N_A_96_21#_c_134_p N_A_918_297#_c_713_n 0.0116461f $X=5.02 $Y=1.87 $X2=0
+ $Y2=0
cc_216 N_A_96_21#_c_117_n N_VGND_M1017_s 0.00426756f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_217 N_A_96_21#_c_110_n N_VGND_c_726_n 0.00316354f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_96_21#_c_110_n N_VGND_c_727_n 0.00423737f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_96_21#_c_111_n N_VGND_c_727_n 0.00423737f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_96_21#_c_111_n N_VGND_c_729_n 0.00146448f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_96_21#_c_112_n N_VGND_c_729_n 0.00146448f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_96_21#_c_113_n N_VGND_c_730_n 0.00316354f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_96_21#_c_117_n N_VGND_c_730_n 0.0133599f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_224 N_A_96_21#_c_117_n N_VGND_c_733_n 0.00195943f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_225 N_A_96_21#_c_121_n N_VGND_c_733_n 0.00223545f $X=2.415 $Y=0.775 $X2=0
+ $Y2=0
cc_226 N_A_96_21#_c_112_n N_VGND_c_737_n 0.00423334f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_96_21#_c_113_n N_VGND_c_737_n 0.00541359f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_96_21#_M1022_d N_VGND_c_739_n 0.00216833f $X=2.83 $Y=0.235 $X2=0
+ $Y2=0
cc_229 N_A_96_21#_M1018_d N_VGND_c_739_n 0.00216833f $X=3.67 $Y=0.235 $X2=0
+ $Y2=0
cc_230 N_A_96_21#_c_110_n N_VGND_c_739_n 0.00674307f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_96_21#_c_111_n N_VGND_c_739_n 0.00571669f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_96_21#_c_112_n N_VGND_c_739_n 0.0057163f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_96_21#_c_113_n N_VGND_c_739_n 0.0108276f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_96_21#_c_117_n N_VGND_c_739_n 0.00413086f $X=2.23 $Y=0.82 $X2=0 $Y2=0
cc_235 N_A_96_21#_c_121_n N_VGND_c_739_n 0.004011f $X=2.415 $Y=0.775 $X2=0 $Y2=0
cc_236 N_A_96_21#_c_118_n N_A_484_47#_M1022_s 0.00235892f $X=2.545 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_237 N_A_96_21#_c_119_n N_A_484_47#_M1022_s 8.01181e-19 $X=3.805 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_238 N_A_96_21#_c_119_n N_A_484_47#_M1001_s 0.00162317f $X=3.805 $Y=0.73 $X2=0
+ $Y2=0
cc_239 N_A_96_21#_M1022_d N_A_484_47#_c_826_n 0.00312026f $X=2.83 $Y=0.235 $X2=0
+ $Y2=0
cc_240 N_A_96_21#_M1018_d N_A_484_47#_c_826_n 0.00312026f $X=3.67 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_A_96_21#_c_118_n N_A_484_47#_c_826_n 0.0814184f $X=2.545 $Y=0.775 $X2=0
+ $Y2=0
cc_242 N_A_96_21#_c_121_n N_A_484_47#_c_826_n 0.0018027f $X=2.415 $Y=0.775 $X2=0
+ $Y2=0
cc_243 N_A_96_21#_c_119_n N_A_484_47#_c_828_n 0.00799569f $X=3.805 $Y=0.73 $X2=0
+ $Y2=0
cc_244 N_B1_c_263_n N_B2_c_349_n 0.0270078f $X=2.755 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_245 N_B1_M1013_g N_B2_M1009_g 0.0439608f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_246 N_B1_c_271_n N_B2_M1009_g 0.00991308f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_247 N_B1_c_264_n N_B2_c_350_n 0.0267413f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B1_M1021_g N_B2_M1010_g 0.0440009f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B1_c_271_n N_B2_M1010_g 0.0102793f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_250 N_B1_c_271_n B2 0.0391837f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_251 N_B1_c_265_n B2 0.0172311f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B1_c_266_n B2 6.66616e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_253 N_B1_c_267_n B2 2.07818e-19 $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_c_268_n B2 0.0169874f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B1_c_271_n N_B2_c_352_n 0.00214031f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_256 N_B1_c_265_n N_B2_c_352_n 0.00458063f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B1_c_266_n N_B2_c_352_n 0.0223771f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B1_c_267_n N_B2_c_352_n 0.0223106f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B1_c_268_n N_B2_c_352_n 0.00592594f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B1_c_264_n N_A1_c_390_n 0.00937759f $X=4.015 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_261 N_B1_M1021_g N_A1_M1002_g 0.0387452f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_262 N_B1_c_271_n N_A1_M1002_g 5.77655e-19 $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_263 N_B1_c_265_n N_A1_M1002_g 3.59226e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B1_M1021_g N_A1_c_392_n 3.59226e-19 $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B1_c_265_n N_A1_c_392_n 0.0307171f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_266 N_B1_c_266_n N_A1_c_392_n 7.80994e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B1_c_265_n N_A1_c_393_n 7.80994e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B1_c_266_n N_A1_c_393_n 0.0197715f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B1_M1021_g N_A1_c_403_n 5.77655e-19 $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_270 N_B1_c_271_n N_A1_c_403_n 0.0154679f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_271 N_B1_c_268_n N_VPWR_M1019_d 0.00407272f $X=2.755 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_c_271_n N_VPWR_M1021_s 0.00151212f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_273 N_B1_M1021_g N_VPWR_c_528_n 0.00323788f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B1_M1013_g N_VPWR_c_533_n 0.00585385f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B1_M1021_g N_VPWR_c_533_n 0.00585385f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B1_M1013_g N_VPWR_c_524_n 0.00723564f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B1_M1021_g N_VPWR_c_524_n 0.0061234f $X=4.015 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B1_M1013_g N_VPWR_c_538_n 0.00518337f $X=2.755 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B1_c_271_n N_A_566_297#_M1013_d 0.00124563f $X=3.85 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_280 N_B1_c_268_n N_A_566_297#_M1013_d 0.00104763f $X=2.755 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_281 N_B1_c_271_n N_A_566_297#_M1010_d 0.00165255f $X=3.85 $Y=1.53 $X2=0 $Y2=0
cc_282 N_B1_c_263_n N_VGND_c_730_n 0.0019578f $X=2.755 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B1_c_263_n N_VGND_c_733_n 0.00357877f $X=2.755 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B1_c_264_n N_VGND_c_733_n 0.00357877f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B1_c_263_n N_VGND_c_739_n 0.00657948f $X=2.755 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B1_c_264_n N_VGND_c_739_n 0.00546478f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B1_c_263_n N_A_484_47#_c_826_n 0.00886996f $X=2.755 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_B1_c_264_n N_A_484_47#_c_826_n 0.0105068f $X=4.015 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B1_c_265_n N_A_484_47#_c_826_n 0.00390962f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_290 N_B1_c_264_n N_A_484_47#_c_828_n 2.00828e-19 $X=4.015 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_B1_c_265_n N_A_484_47#_c_828_n 0.00353546f $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B1_c_266_n N_A_484_47#_c_828_n 2.55742e-19 $X=4.015 $Y=1.16 $X2=0 $Y2=0
cc_293 N_B2_M1009_g N_VPWR_c_533_n 0.00357877f $X=3.175 $Y=1.985 $X2=0 $Y2=0
cc_294 N_B2_M1010_g N_VPWR_c_533_n 0.00357877f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_295 N_B2_M1009_g N_VPWR_c_524_n 0.00525237f $X=3.175 $Y=1.985 $X2=0 $Y2=0
cc_296 N_B2_M1010_g N_VPWR_c_524_n 0.00525237f $X=3.595 $Y=1.985 $X2=0 $Y2=0
cc_297 N_B2_M1009_g N_A_566_297#_c_690_n 0.00851673f $X=3.175 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_B2_M1010_g N_A_566_297#_c_690_n 0.00851673f $X=3.595 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_B2_c_349_n N_VGND_c_733_n 0.00357877f $X=3.175 $Y=0.995 $X2=0 $Y2=0
cc_300 N_B2_c_350_n N_VGND_c_733_n 0.00357877f $X=3.595 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B2_c_349_n N_VGND_c_739_n 0.00525341f $X=3.175 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B2_c_350_n N_VGND_c_739_n 0.00525341f $X=3.595 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B2_c_349_n N_A_484_47#_c_826_n 0.00886996f $X=3.175 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_B2_c_350_n N_A_484_47#_c_826_n 0.00886996f $X=3.595 $Y=0.995 $X2=0
+ $Y2=0
cc_305 N_A1_c_390_n N_A2_c_476_n 0.0258191f $X=4.515 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_306 N_A1_M1002_g N_A2_M1011_g 0.0440009f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A1_c_402_n N_A2_M1011_g 0.0108086f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_308 N_A1_c_391_n N_A2_c_477_n 0.0258694f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A1_M1008_g N_A2_M1020_g 0.0270786f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A1_c_402_n N_A2_M1020_g 0.0153291f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_311 N_A1_c_392_n A2 0.0133594f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A1_c_393_n A2 2.2122e-19 $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A1_c_402_n A2 0.0349894f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_314 N_A1_c_395_n A2 0.0172564f $X=5.735 $Y=1.175 $X2=0 $Y2=0
cc_315 N_A1_c_397_n A2 2.00336e-19 $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A1_c_392_n N_A2_c_478_n 0.00527477f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A1_c_393_n N_A2_c_478_n 0.022397f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A1_c_402_n N_A2_c_478_n 0.00214031f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_319 N_A1_c_394_n N_A2_c_478_n 0.00362491f $X=5.65 $Y=1.445 $X2=0 $Y2=0
cc_320 N_A1_c_395_n N_A2_c_478_n 0.00144374f $X=5.735 $Y=1.175 $X2=0 $Y2=0
cc_321 N_A1_c_397_n N_A2_c_478_n 0.0222902f $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A1_c_403_n N_VPWR_M1021_s 0.00151212f $X=4.68 $Y=1.53 $X2=0 $Y2=0
cc_323 N_A1_M1002_g N_VPWR_c_528_n 0.00525229f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A1_M1008_g N_VPWR_c_529_n 0.00505805f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A1_c_402_n N_VPWR_c_529_n 0.00786716f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_326 A1 N_VPWR_c_529_n 0.0166332f $X=6.145 $Y=1.105 $X2=0 $Y2=0
cc_327 N_A1_M1002_g N_VPWR_c_530_n 0.00585385f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A1_M1008_g N_VPWR_c_530_n 0.00585385f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A1_M1002_g N_VPWR_c_524_n 0.00617642f $X=4.515 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A1_M1008_g N_VPWR_c_524_n 0.0116728f $X=5.775 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A1_c_402_n N_A_918_297#_M1002_d 0.00130005f $X=5.565 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_332 N_A1_c_403_n N_A_918_297#_M1002_d 3.52503e-19 $X=4.68 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_333 N_A1_c_402_n N_A_918_297#_M1020_d 0.00167564f $X=5.565 $Y=1.53 $X2=0
+ $Y2=0
cc_334 N_A1_c_402_n N_A_918_297#_c_717_n 0.0132239f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_335 N_A1_c_390_n N_VGND_c_731_n 0.00268723f $X=4.515 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A1_c_391_n N_VGND_c_732_n 0.00268723f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A1_c_390_n N_VGND_c_733_n 0.00422898f $X=4.515 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A1_c_391_n N_VGND_c_738_n 0.00423334f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A1_c_390_n N_VGND_c_739_n 0.00598371f $X=4.515 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A1_c_391_n N_VGND_c_739_n 0.00683939f $X=5.775 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A1_c_390_n N_A_484_47#_c_848_n 0.00255288f $X=4.515 $Y=0.995 $X2=0
+ $Y2=0
cc_342 N_A1_c_390_n N_A_484_47#_c_849_n 0.00393886f $X=4.515 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A1_c_390_n N_A_484_47#_c_827_n 0.00845282f $X=4.515 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A1_c_392_n N_A_484_47#_c_827_n 0.0160434f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A1_c_393_n N_A_484_47#_c_827_n 0.001478f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A1_c_402_n N_A_484_47#_c_827_n 0.0071189f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_347 N_A1_c_390_n N_A_484_47#_c_828_n 0.00111376f $X=4.515 $Y=0.995 $X2=0
+ $Y2=0
cc_348 N_A1_c_392_n N_A_484_47#_c_828_n 0.010391f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A1_c_393_n N_A_484_47#_c_828_n 0.00153445f $X=4.515 $Y=1.16 $X2=0 $Y2=0
cc_350 N_A1_c_390_n N_A_484_47#_c_857_n 5.22228e-19 $X=4.515 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A1_c_391_n N_A_484_47#_c_857_n 5.22228e-19 $X=5.775 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A1_c_391_n N_A_484_47#_c_829_n 0.00995081f $X=5.775 $Y=0.995 $X2=0
+ $Y2=0
cc_353 N_A1_c_402_n N_A_484_47#_c_829_n 0.00549032f $X=5.565 $Y=1.53 $X2=0 $Y2=0
cc_354 N_A1_c_395_n N_A_484_47#_c_829_n 0.0135931f $X=5.735 $Y=1.175 $X2=0 $Y2=0
cc_355 A1 N_A_484_47#_c_829_n 0.0333889f $X=6.145 $Y=1.105 $X2=0 $Y2=0
cc_356 N_A1_c_397_n N_A_484_47#_c_829_n 0.00301563f $X=5.775 $Y=1.16 $X2=0 $Y2=0
cc_357 N_A1_c_391_n N_A_484_47#_c_830_n 0.00630972f $X=5.775 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A2_M1011_g N_VPWR_c_530_n 0.00357877f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_359 N_A2_M1020_g N_VPWR_c_530_n 0.00357877f $X=5.355 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A2_M1011_g N_VPWR_c_524_n 0.00525237f $X=4.935 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A2_M1020_g N_VPWR_c_524_n 0.00525237f $X=5.355 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A2_M1011_g N_A_918_297#_c_710_n 0.00851673f $X=4.935 $Y=1.985 $X2=0
+ $Y2=0
cc_363 N_A2_M1020_g N_A_918_297#_c_710_n 0.0121306f $X=5.355 $Y=1.985 $X2=0
+ $Y2=0
cc_364 N_A2_c_476_n N_VGND_c_731_n 0.00146448f $X=4.935 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A2_c_477_n N_VGND_c_732_n 0.00146448f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A2_c_476_n N_VGND_c_735_n 0.00424416f $X=4.935 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A2_c_477_n N_VGND_c_735_n 0.00423334f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A2_c_476_n N_VGND_c_739_n 0.00576327f $X=4.935 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A2_c_477_n N_VGND_c_739_n 0.0057435f $X=5.355 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A2_c_476_n N_A_484_47#_c_849_n 4.86433e-19 $X=4.935 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A2_c_476_n N_A_484_47#_c_827_n 0.00894278f $X=4.935 $Y=0.995 $X2=0
+ $Y2=0
cc_372 A2 N_A_484_47#_c_827_n 0.00545718f $X=5.225 $Y=1.105 $X2=0 $Y2=0
cc_373 N_A2_c_476_n N_A_484_47#_c_857_n 0.00630972f $X=4.935 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_A2_c_477_n N_A_484_47#_c_857_n 0.00630972f $X=5.355 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A2_c_477_n N_A_484_47#_c_829_n 0.00908248f $X=5.355 $Y=0.995 $X2=0
+ $Y2=0
cc_376 A2 N_A_484_47#_c_829_n 0.00582553f $X=5.225 $Y=1.105 $X2=0 $Y2=0
cc_377 N_A2_c_477_n N_A_484_47#_c_830_n 5.22228e-19 $X=5.355 $Y=0.995 $X2=0
+ $Y2=0
cc_378 N_A2_c_476_n N_A_484_47#_c_831_n 0.00128009f $X=4.935 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A2_c_477_n N_A_484_47#_c_831_n 0.00113286f $X=5.355 $Y=0.995 $X2=0
+ $Y2=0
cc_380 A2 N_A_484_47#_c_831_n 0.0265405f $X=5.225 $Y=1.105 $X2=0 $Y2=0
cc_381 N_A2_c_478_n N_A_484_47#_c_831_n 0.00230339f $X=5.355 $Y=1.16 $X2=0 $Y2=0
cc_382 N_VPWR_c_524_n N_X_M1003_s 0.00284632f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_524_n N_X_M1007_s 0.00284632f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_M1003_d N_X_c_620_n 6.05749e-19 $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_385 N_VPWR_c_526_n N_X_c_620_n 0.00365338f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_386 N_VPWR_M1003_d N_X_c_621_n 0.00347536f $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_387 N_VPWR_c_526_n N_X_c_621_n 0.011469f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_388 N_VPWR_c_532_n N_X_c_663_n 0.0142343f $X=1.06 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_c_524_n N_X_c_663_n 0.00955092f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_M1006_d N_X_c_622_n 0.00169858f $X=1.05 $Y=1.485 $X2=0 $Y2=0
cc_391 N_VPWR_c_527_n N_X_c_622_n 0.0121607f $X=1.185 $Y=1.99 $X2=0 $Y2=0
cc_392 N_VPWR_c_524_n N_X_c_667_n 0.00955092f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_537_n N_X_c_667_n 0.0142343f $X=1.9 $Y=2.465 $X2=0 $Y2=0
cc_394 N_VPWR_c_524_n N_A_566_297#_M1013_d 0.00219968f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_395 N_VPWR_c_524_n N_A_566_297#_M1010_d 0.00219968f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_533_n N_A_566_297#_c_690_n 0.0330174f $X=4.1 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_524_n N_A_566_297#_c_690_n 0.0204707f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_533_n N_A_566_297#_c_694_n 0.0136719f $X=4.1 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_524_n N_A_566_297#_c_694_n 0.00938288f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_533_n N_A_566_297#_c_695_n 0.0137033f $X=4.1 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_c_524_n N_A_566_297#_c_695_n 0.00938745f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_524_n N_A_918_297#_M1002_d 0.00219968f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_403 N_VPWR_c_524_n N_A_918_297#_M1020_d 0.00246446f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_530_n N_A_918_297#_c_710_n 0.0473226f $X=5.905 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_524_n N_A_918_297#_c_710_n 0.0300947f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_530_n N_A_918_297#_c_713_n 0.0137033f $X=5.905 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_524_n N_A_918_297#_c_713_n 0.00938745f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_408 N_X_c_615_n N_VGND_M1000_s 5.40298e-19 $X=0.6 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_409 N_X_c_616_n N_VGND_M1000_s 0.00329182f $X=0.37 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_410 N_X_c_617_n N_VGND_M1004_s 0.00162089f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_411 N_X_c_615_n N_VGND_c_726_n 0.00402428f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_412 N_X_c_616_n N_VGND_c_726_n 0.00920832f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_413 N_X_c_629_n N_VGND_c_727_n 0.017716f $X=0.765 $Y=0.39 $X2=0 $Y2=0
cc_414 N_X_c_617_n N_VGND_c_727_n 0.00198695f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_415 N_X_c_615_n N_VGND_c_728_n 0.0019947f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_416 N_X_c_616_n N_VGND_c_728_n 0.00293744f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_417 N_X_c_617_n N_VGND_c_729_n 0.0122559f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_418 N_X_c_617_n N_VGND_c_737_n 0.00198695f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_419 N_X_c_645_n N_VGND_c_737_n 0.0188551f $X=1.605 $Y=0.39 $X2=0 $Y2=0
cc_420 N_X_M1000_d N_VGND_c_739_n 0.00215535f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_421 N_X_M1005_d N_VGND_c_739_n 0.00215201f $X=1.47 $Y=0.235 $X2=0 $Y2=0
cc_422 N_X_c_615_n N_VGND_c_739_n 0.00407016f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_423 N_X_c_616_n N_VGND_c_739_n 0.00542613f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_424 N_X_c_629_n N_VGND_c_739_n 0.0121406f $X=0.765 $Y=0.39 $X2=0 $Y2=0
cc_425 N_X_c_617_n N_VGND_c_739_n 0.00835832f $X=1.44 $Y=0.815 $X2=0 $Y2=0
cc_426 N_X_c_645_n N_VGND_c_739_n 0.0122069f $X=1.605 $Y=0.39 $X2=0 $Y2=0
cc_427 N_VGND_c_739_n N_A_484_47#_M1022_s 0.00209344f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_428 N_VGND_c_739_n N_A_484_47#_M1001_s 0.00215227f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_739_n N_A_484_47#_M1023_s 0.00279445f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_739_n N_A_484_47#_M1014_d 0.00215201f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_739_n N_A_484_47#_M1016_d 0.00209319f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_730_n N_A_484_47#_c_826_n 0.0130084f $X=2.025 $Y=0.39 $X2=0
+ $Y2=0
cc_433 N_VGND_c_733_n N_A_484_47#_c_826_n 0.0991765f $X=4.64 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_739_n N_A_484_47#_c_826_n 0.0628989f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_733_n N_A_484_47#_c_848_n 0.0208178f $X=4.64 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_739_n N_A_484_47#_c_848_n 0.0124843f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_M1012_s N_A_484_47#_c_827_n 0.00165819f $X=4.59 $Y=0.235 $X2=0
+ $Y2=0
cc_438 N_VGND_c_731_n N_A_484_47#_c_827_n 0.0116528f $X=4.725 $Y=0.39 $X2=0
+ $Y2=0
cc_439 N_VGND_c_733_n N_A_484_47#_c_827_n 0.00193763f $X=4.64 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_735_n N_A_484_47#_c_827_n 0.00193763f $X=5.48 $Y=0 $X2=0 $Y2=0
cc_441 N_VGND_c_739_n N_A_484_47#_c_827_n 0.00827287f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_442 N_VGND_c_735_n N_A_484_47#_c_857_n 0.0188551f $X=5.48 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_739_n N_A_484_47#_c_857_n 0.0122069f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_444 N_VGND_M1015_s N_A_484_47#_c_829_n 0.00162089f $X=5.43 $Y=0.235 $X2=0
+ $Y2=0
cc_445 N_VGND_c_732_n N_A_484_47#_c_829_n 0.0122559f $X=5.565 $Y=0.39 $X2=0
+ $Y2=0
cc_446 N_VGND_c_735_n N_A_484_47#_c_829_n 0.00198695f $X=5.48 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_c_738_n N_A_484_47#_c_829_n 0.00198695f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_448 N_VGND_c_739_n N_A_484_47#_c_829_n 0.00835832f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_738_n N_A_484_47#_c_830_n 0.0209752f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_739_n N_A_484_47#_c_830_n 0.0124119f $X=6.21 $Y=0 $X2=0 $Y2=0

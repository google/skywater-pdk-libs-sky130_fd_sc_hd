* File: sky130_fd_sc_hd__nand3_1.pex.spice
* Created: Tue Sep  1 19:16:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND3_1%C 1 3 6 8 9 16
r29 13 16 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r31 8 9 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=0.22 $Y=0.85 $X2=0.22
+ $Y2=1.16
r32 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r34 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_1%B 3 6 8 9 13 15
r34 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=1.325
r35 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.95 $Y2=0.995
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.16 $X2=0.95 $Y2=1.16
r37 9 14 0.921954 $w=3.73e-07 $l=3e-08 $layer=LI1_cond $X=1.052 $Y=1.19
+ $X2=1.052 $Y2=1.16
r38 8 14 9.52686 $w=3.73e-07 $l=3.1e-07 $layer=LI1_cond $X=1.052 $Y=0.85
+ $X2=1.052 $Y2=1.16
r39 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.985
+ $X2=0.89 $Y2=1.325
r40 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.56 $X2=0.89
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_1%A 1 3 6 8 13
r27 10 13 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.555 $Y2=1.16
r28 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.555
+ $Y=1.16 $X2=1.555 $Y2=1.16
r29 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.325
+ $X2=1.37 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.37 $Y=1.325 $X2=1.37
+ $Y2=1.985
r31 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=0.995
+ $X2=1.37 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.37 $Y=0.995 $X2=1.37
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_1%VPWR 1 2 7 9 15 17 19 26 27 33
r27 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r28 27 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 24 33 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.13 $Y2=2.72
r31 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.61 $Y2=2.72
r32 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r33 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r34 20 30 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r35 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r36 19 33 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.13 $Y2=2.72
r37 19 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r39 17 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r40 13 33 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.13 $Y2=2.72
r41 13 15 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.13 $Y=2.635
+ $X2=1.13 $Y2=2
r42 9 12 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r43 7 30 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r44 7 12 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r45 2 15 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r46 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r47 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_1%Y 1 2 3 12 14 16 18 20 22 24 27 31
r53 27 31 22.9811 $w=3.38e-07 $l=6.78e-07 $layer=LI1_cond $X=1.415 $Y=0.425
+ $X2=0.737 $Y2=0.425
r54 26 27 0.533618 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=0.425
+ $X2=1.415 $Y2=0.425
r55 24 26 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.58 $Y=0.38
+ $X2=1.58 $Y2=0.425
r56 20 31 40.3321 $w=2.63e-07 $l=9e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.605 $Y2=0.595
r57 20 22 3.64284 $w=2.55e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.605 $Y=1.495
+ $X2=0.68 $Y2=1.58
r58 16 30 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=1.665 $X2=1.58
+ $Y2=1.58
r59 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.58 $Y=1.665
+ $X2=1.58 $Y2=2.34
r60 15 22 2.83584 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.58
+ $X2=0.68 $Y2=1.58
r61 14 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=1.58
+ $X2=1.58 $Y2=1.58
r62 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.415 $Y=1.58
+ $X2=0.845 $Y2=1.58
r63 10 22 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=1.58
r64 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r65 3 30 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=1.485 $X2=1.58 $Y2=1.66
r66 3 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=1.485 $X2=1.58 $Y2=2.34
r67 2 22 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r68 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r69 1 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND3_1%VGND 1 4 6 8 15 16
r24 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r25 13 16 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r26 12 15 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r27 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r28 10 19 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r29 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r30 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r31 8 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r32 4 19 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r33 4 6 14.688 $w=2.53e-07 $l=3.25e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.41
r34 1 6 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.41
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 a_750_97# S0 a_757_363# VPB phighvt w=420000u l=150000u
+  ad=3.822e+11p pd=3.5e+06u as=2.171e+11p ps=2.72e+06u
M1001 a_1478_413# S1 a_277_47# VPB phighvt w=420000u l=150000u
+  ad=1.84175e+11p pd=1.98e+06u as=2.226e+11p ps=2.74e+06u
M1002 VPWR S0 a_247_21# VPB phighvt w=420000u l=150000u
+  ad=7.039e+11p pd=8e+06u as=1.083e+11p ps=1.36e+06u
M1003 a_750_97# a_1290_413# a_1478_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A3 a_923_363# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.8025e+11p ps=1.99e+06u
M1005 a_1478_413# S1 a_750_97# VNB nshort w=420000u l=150000u
+  ad=3.0205e+11p pd=2.57e+06u as=2.226e+11p ps=2.74e+06u
M1006 VGND S0 a_247_21# VNB nshort w=420000u l=150000u
+  ad=6.142e+11p pd=7.3e+06u as=1.092e+11p ps=1.36e+06u
M1007 a_277_47# a_1290_413# a_1478_413# VNB nshort w=420000u l=150000u
+  ad=2.7965e+11p pd=3.21e+06u as=0p ps=0u
M1008 a_923_363# a_247_21# a_750_97# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1290_413# S1 VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1010 VPWR A1 a_27_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.184e+11p ps=2.72e+06u
M1011 a_27_47# S0 a_277_47# VNB nshort w=420000u l=150000u
+  ad=2.184e+11p pd=2.72e+06u as=0p ps=0u
M1012 a_193_413# S0 a_277_47# VPB phighvt w=420000u l=150000u
+  ad=2.171e+11p pd=2.72e+06u as=0p ps=0u
M1013 a_193_47# A0 VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1014 a_277_47# a_247_21# a_27_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1290_413# S1 VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1016 X a_1478_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1017 a_277_47# a_247_21# a_193_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_750_97# S0 a_668_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.171e+11p ps=2.72e+06u
M1019 a_757_363# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_1478_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1021 VGND A1 a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_834_97# a_247_21# a_750_97# VNB nshort w=420000u l=150000u
+  ad=2.1715e+11p pd=2.72e+06u as=0p ps=0u
M1023 VGND A3 a_668_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_834_97# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_193_413# A0 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__clkdlybuf4s25_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.495000 1.615000 ;
    END
  END A
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  0.497000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.770000 0.285000 3.095000 0.615000 ;
        RECT 2.770000 1.625000 3.095000 2.460000 ;
        RECT 2.865000 0.615000 3.095000 0.765000 ;
        RECT 2.865000 0.765000 3.595000 1.275000 ;
        RECT 2.865000 1.275000 3.095000 1.625000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.305000 0.345000 0.640000 ;
      RECT 0.095000  0.640000 0.840000 0.810000 ;
      RECT 0.095000  1.785000 0.835000 1.955000 ;
      RECT 0.095000  1.955000 0.345000 2.465000 ;
      RECT 0.575000  0.085000 0.905000 0.470000 ;
      RECT 0.575000  2.125000 0.905000 2.635000 ;
      RECT 0.665000  0.810000 0.840000 0.995000 ;
      RECT 0.665000  0.995000 1.035000 1.325000 ;
      RECT 0.665000  1.325000 1.005000 1.750000 ;
      RECT 0.665000  1.750000 0.835000 1.785000 ;
      RECT 1.095000  0.255000 1.425000 0.780000 ;
      RECT 1.175000  1.425000 1.440000 2.465000 ;
      RECT 1.205000  0.780000 1.425000 0.995000 ;
      RECT 1.205000  0.995000 2.165000 1.325000 ;
      RECT 1.205000  1.325000 1.440000 1.425000 ;
      RECT 1.615000  0.255000 1.945000 0.635000 ;
      RECT 1.615000  0.635000 2.595000 0.805000 ;
      RECT 1.695000  1.500000 2.595000 1.745000 ;
      RECT 1.695000  1.745000 1.945000 2.465000 ;
      RECT 2.135000  0.085000 2.465000 0.465000 ;
      RECT 2.135000  1.915000 2.465000 2.635000 ;
      RECT 2.335000  0.805000 2.595000 1.500000 ;
      RECT 3.265000  0.085000 3.595000 0.550000 ;
      RECT 3.265000  1.635000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_2
END LIBRARY

* File: sky130_fd_sc_hd__nand4_4.spice
* Created: Thu Aug 27 14:30:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand4_4.spice.pex"
.subckt sky130_fd_sc_hd__nand4_4  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1009 N_A_27_47#_M1009_d N_D_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1014_d N_D_M1014_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1017 N_A_27_47#_M1014_d N_D_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1030 N_A_27_47#_M1030_d N_D_M1030_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1015 N_A_445_47#_M1015_d N_C_M1015_g N_A_27_47#_M1030_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1020 N_A_445_47#_M1015_d N_C_M1020_g N_A_27_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1025 N_A_445_47#_M1025_d N_C_M1025_g N_A_27_47#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1026 N_A_445_47#_M1025_d N_C_M1026_g N_A_27_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_445_47#_M1007_d N_B_M1007_g N_A_803_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_445_47#_M1007_d N_B_M1010_g N_A_803_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1016 N_A_445_47#_M1016_d N_B_M1016_g N_A_803_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1021 N_A_445_47#_M1016_d N_B_M1021_g N_A_803_47#_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=5.532 M=1 R=4.33333
+ SA=75001.4 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1011_d N_A_M1011_g N_A_803_47#_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75001.9
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1011_d N_A_M1013_g N_A_803_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1023 N_Y_M1023_d N_A_M1023_g N_A_803_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1024 N_Y_M1023_d N_A_M1024_g N_A_803_47#_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_D_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75007.1 A=0.15
+ P=2.3 MULT=1
MM1003 N_Y_M1002_d N_D_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75006.6
+ A=0.15 P=2.3 MULT=1
MM1018 N_Y_M1018_d N_D_M1018_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75006.2 A=0.15
+ P=2.3 MULT=1
MM1027 N_Y_M1018_d N_D_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75005.8
+ A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75005.4
+ A=0.15 P=2.3 MULT=1
MM1004 N_Y_M1000_d N_C_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75005 A=0.15
+ P=2.3 MULT=1
MM1022 N_Y_M1022_d N_C_M1022_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7 SB=75004.5
+ A=0.15 P=2.3 MULT=1
MM1028 N_Y_M1022_d N_C_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.395 PD=1.27 PS=1.79 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1 SB=75004.1
+ A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.395 PD=1.27 PS=1.79 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1 SB=75003.2
+ A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1001_d N_B_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5 SB=75002.8
+ A=0.15 P=2.3 MULT=1
MM1008 N_Y_M1008_d N_B_M1008_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.9 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1029 N_Y_M1008_d N_B_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.165 PD=1.27 PS=1.33 NRD=0 NRS=5.8903 M=1 R=6.66667 SA=75005.3 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1029_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.165 PD=1.27 PS=1.33 NRD=0 NRS=3.9203 M=1 R=6.66667 SA=75005.8 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1006_d N_A_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.2 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1019 N_Y_M1019_d N_A_M1019_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.6 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1031 N_Y_M1019_d N_A_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.1 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hd__nand4_4.spice.SKY130_FD_SC_HD__NAND4_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__dlxtp_1.spice
* Created: Tue Sep  1 19:06:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dlxtp_1.pex.spice"
.subckt sky130_fd_sc_hd__dlxtp_1  VNB VPB GATE D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_GATE_M1016_g N_A_27_47#_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_193_47#_M1012_d N_A_27_47#_M1012_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_D_M1005_g N_A_299_47#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 A_465_47# N_A_299_47#_M1010_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.0567 PD=0.802308 PS=0.69 NRD=32.628 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1015 N_A_560_47#_M1015_d N_A_193_47#_M1015_g A_465_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0621 AS=0.0609231 PD=0.705 PS=0.687692 NRD=21.66 NRS=38.076 M=1
+ R=2.4 SA=75001.1 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1007 A_659_47# N_A_27_47#_M1007_g N_A_560_47#_M1015_d VNB NSHORT L=0.15 W=0.36
+ AD=0.0486 AS=0.0621 PD=0.63 PS=0.705 NRD=26.664 NRS=0 M=1 R=2.4 SA=75001.6
+ SB=75000.6 A=0.054 P=1.02 MULT=1
MM1006 N_VGND_M1006_d N_A_713_21#_M1006_g A_659_47# VNB NSHORT L=0.15 W=0.36
+ AD=0.0936 AS=0.0486 PD=1.24 PS=0.63 NRD=0 NRS=26.664 M=1 R=2.4 SA=75002
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1008 N_VGND_M1008_d N_A_560_47#_M1008_g N_A_713_21#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.092625 AS=0.169 PD=0.935 PS=1.82 NRD=1.836 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_Q_M1017_d N_A_713_21#_M1017_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.092625 PD=1.87 PS=0.935 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_GATE_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_VPWR_M1014_d N_D_M1014_g N_A_299_47#_M1014_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1013 A_465_369# N_A_299_47#_M1013_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.115623 AS=0.0864 PD=1.16528 PS=0.91 NRD=38.6711 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 N_A_560_47#_M1004_d N_A_27_47#_M1004_g A_465_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0758774 PD=0.69 PS=0.764717 NRD=0 NRS=58.9227 M=1 R=2.8
+ SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_644_413# N_A_193_47#_M1002_g N_A_560_47#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07245 AS=0.0567 PD=0.765 PS=0.69 NRD=55.1009 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_713_21#_M1009_g A_644_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1134 AS=0.07245 PD=1.38 PS=0.765 NRD=2.3443 NRS=55.1009 M=1 R=2.8
+ SA=75002 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_560_47#_M1001_g N_A_713_21#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.1425 AS=0.26 PD=1.285 PS=2.52 NRD=1.9503 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_Q_M1003_d N_A_713_21#_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.1425 PD=2.57 PS=1.285 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.4695 P=15.01
c_126 VPB 0 1.54137e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dlxtp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nand4b_1.spice
* Created: Thu Aug 27 14:30:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand4b_1.pex.spice"
.subckt sky130_fd_sc_hd__nand4b_1  VNB VPB A_N D C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_N_M1009_g N_A_41_93#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.1113 PD=0.816449 PS=1.37 NRD=47.364 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 A_232_47# N_D_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.143516 PD=0.92 PS=1.26355 NRD=14.76 NRS=9.228 M=1 R=4.33333 SA=75000.6
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1000 A_316_47# N_C_M1000_g A_232_47# VNB NSHORT L=0.15 W=0.65 AD=0.125125
+ AS=0.08775 PD=1.035 PS=0.92 NRD=25.38 NRS=14.76 M=1 R=4.33333 SA=75001
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1007 A_423_47# N_B_M1007_g A_316_47# VNB NSHORT L=0.15 W=0.65 AD=0.12675
+ AS=0.125125 PD=1.04 PS=1.035 NRD=25.836 NRS=25.38 M=1 R=4.33333 SA=75001.5
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A_41_93#_M1004_g A_423_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.2275 AS=0.12675 PD=2 PS=1.04 NRD=11.988 NRS=25.836 M=1 R=4.33333
+ SA=75002.1 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_41_93#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.1092 PD=0.789718 PS=1.36 NRD=28.1316 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_D_M1008_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.205282 PD=1.27 PS=1.88028 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.4 SB=75001.7
+ A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g N_Y_M1008_d VPB PHIGHVT L=0.15 W=1 AD=0.1925
+ AS=0.135 PD=1.385 PS=1.27 NRD=10.8153 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.1925 PD=1.39 PS=1.385 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75001.3
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_41_93#_M1005_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.195 PD=2.56 PS=1.39 NRD=0 NRS=22.6353 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__nand4b_1.pxi.spice"
*
.ends
*
*

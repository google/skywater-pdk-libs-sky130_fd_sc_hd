* File: sky130_fd_sc_hd__o32a_1.spice.pex
* Created: Thu Aug 27 14:40:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O32A_1%A_77_199# 1 2 9 12 15 16 17 19 20 21 22 23 24
+ 27 29 30 39 42
c91 15 0 1.33587e-19 $X=0.725 $Y=1.495
r92 37 39 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=2.875 $Y=0.73
+ $X2=3.05 $Y2=0.73
r93 30 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.16
+ $X2=0.55 $Y2=1.325
r94 30 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.16
+ $X2=0.55 $Y2=0.995
r95 29 31 7.33677 $w=2.91e-07 $l=1.75e-07 $layer=LI1_cond $X=0.55 $Y=1.16
+ $X2=0.725 $Y2=1.16
r96 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.55
+ $Y=1.16 $X2=0.55 $Y2=1.16
r97 26 39 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.05 $Y=0.825 $X2=3.05
+ $Y2=0.73
r98 26 27 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.05 $Y=0.825
+ $X2=3.05 $Y2=1.835
r99 25 33 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.96
+ $X2=2.345 $Y2=1.96
r100 24 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.965 $Y=1.96
+ $X2=3.05 $Y2=1.835
r101 24 25 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=2.965 $Y=1.96
+ $X2=2.51 $Y2=1.96
r102 23 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=2.295
+ $X2=2.345 $Y2=2.38
r103 22 33 3.01144 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=2.345 $Y=2.085
+ $X2=2.345 $Y2=1.96
r104 22 23 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.345 $Y=2.085
+ $X2=2.345 $Y2=2.295
r105 20 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=2.38
+ $X2=2.345 $Y2=2.38
r106 20 21 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.18 $Y=2.38
+ $X2=1.315 $Y2=2.38
r107 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=2.295
+ $X2=1.315 $Y2=2.38
r108 18 19 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.23 $Y=1.665
+ $X2=1.23 $Y2=2.295
r109 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=1.58
+ $X2=1.23 $Y2=1.665
r110 16 17 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.145 $Y=1.58
+ $X2=0.81 $Y2=1.58
r111 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.725 $Y=1.495
+ $X2=0.81 $Y2=1.58
r112 14 31 3.88217 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.325
+ $X2=0.725 $Y2=1.16
r113 14 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.725 $Y=1.325
+ $X2=0.725 $Y2=1.495
r114 12 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.64 $Y=1.985
+ $X2=0.64 $Y2=1.325
r115 9 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.64 $Y=0.56
+ $X2=0.64 $Y2=0.995
r116 2 35 600 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.485 $X2=2.345 $Y2=2.34
r117 2 33 600 $w=1.7e-07 $l=6.02557e-07 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.485 $X2=2.345 $Y2=2
r118 1 37 182 $w=1.7e-07 $l=5.67913e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.235 $X2=2.875 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%A1 3 6 8 11 13
r33 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.16
+ $X2=1.09 $Y2=1.325
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.16
+ $X2=1.09 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.16 $X2=1.09 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.06 $Y=1.985
+ $X2=1.06 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.06 $Y=0.56 $X2=1.06
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%A2 3 6 8 9 10 15 17
c38 17 0 6.40318e-20 $X=1.63 $Y=0.995
c39 8 0 1.23066e-19 $X=1.605 $Y=1.19
r40 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=1.63 $Y2=1.325
r41 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=1.63 $Y2=0.995
r42 9 10 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.647 $Y=1.53
+ $X2=1.647 $Y2=1.87
r43 9 28 7.26926 $w=3.23e-07 $l=2.05e-07 $layer=LI1_cond $X=1.647 $Y=1.53
+ $X2=1.647 $Y2=1.325
r44 8 28 5.56418 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.637 $Y=1.16
+ $X2=1.637 $Y2=1.325
r45 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.16 $X2=1.63 $Y2=1.16
r46 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.54 $Y=1.985
+ $X2=1.54 $Y2=1.325
r47 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.54 $Y=0.56 $X2=1.54
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%A3 3 6 8 9 13 14 15
r37 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.16
+ $X2=2.17 $Y2=1.325
r38 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.16
+ $X2=2.17 $Y2=0.995
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.16 $X2=2.17 $Y2=1.16
r40 8 9 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=2.117 $Y=1.19
+ $X2=2.117 $Y2=1.53
r41 8 14 1.25721 $w=2.73e-07 $l=3e-08 $layer=LI1_cond $X=2.117 $Y=1.19 $X2=2.117
+ $Y2=1.16
r42 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.08 $Y=1.985
+ $X2=2.08 $Y2=1.325
r43 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.08 $Y=0.56 $X2=2.08
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%B2 3 6 8 9 13 14 15
c38 13 0 8.24349e-20 $X=2.71 $Y=1.16
r39 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.71 $Y2=1.325
r40 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=2.71 $Y2=0.995
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.16 $X2=2.71 $Y2=1.16
r42 8 9 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=2.617 $Y=1.19
+ $X2=2.617 $Y2=1.53
r43 8 14 0.973895 $w=3.53e-07 $l=3e-08 $layer=LI1_cond $X=2.617 $Y=1.19
+ $X2=2.617 $Y2=1.16
r44 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.62 $Y=1.985
+ $X2=2.62 $Y2=1.325
r45 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.62 $Y=0.56 $X2=2.62
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%B1 1 3 6 8 13
r27 10 13 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.18 $Y=1.16
+ $X2=3.405 $Y2=1.16
r28 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.405
+ $Y=1.16 $X2=3.405 $Y2=1.16
r29 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.18 $Y=1.325
+ $X2=3.18 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.18 $Y=1.325 $X2=3.18
+ $Y2=1.985
r31 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.18 $Y=0.995
+ $X2=3.18 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.18 $Y=0.995 $X2=3.18
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%X 1 2 9 10 11 12 13 18 25
r25 12 13 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.277 $Y=1.87
+ $X2=0.277 $Y2=2.21
r26 12 18 3.29269 $w=3.83e-07 $l=1.1e-07 $layer=LI1_cond $X=0.277 $Y=1.87
+ $X2=0.277 $Y2=1.76
r27 11 29 12.8932 $w=5.08e-07 $l=3.15e-07 $layer=LI1_cond $X=0.34 $Y=0.51
+ $X2=0.34 $Y2=0.825
r28 11 25 3.04883 $w=5.08e-07 $l=1.3e-07 $layer=LI1_cond $X=0.34 $Y=0.51
+ $X2=0.34 $Y2=0.38
r29 10 29 42.4623 $w=1.73e-07 $l=6.7e-07 $layer=LI1_cond $X=0.172 $Y=1.495
+ $X2=0.172 $Y2=0.825
r30 9 18 2.18515 $w=3.83e-07 $l=7.3e-08 $layer=LI1_cond $X=0.277 $Y=1.687
+ $X2=0.277 $Y2=1.76
r31 9 10 9.21419 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=0.277 $Y=1.687
+ $X2=0.277 $Y2=1.495
r32 2 18 300 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=2 $X=0.23
+ $Y=1.485 $X2=0.385 $Y2=1.76
r33 1 25 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.305
+ $Y=0.235 $X2=0.43 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%VPWR 1 2 11 13 15 19 21 30 34 38
c44 1 0 1.33587e-19 $X=0.715 $Y=1.485
r45 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 31 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r47 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r49 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 25 28 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 24 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 22 30 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=0.83 $Y2=2.72
r55 22 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.975 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 21 33 4.42954 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.305 $Y=2.72
+ $X2=3.492 $Y2=2.72
r57 21 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.305 $Y=2.72
+ $X2=2.99 $Y2=2.72
r58 19 38 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r59 15 18 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=3.45 $Y=1.66
+ $X2=3.45 $Y2=2.34
r60 13 33 3.0083 $w=2.9e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.45 $Y=2.635
+ $X2=3.492 $Y2=2.72
r61 13 18 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.45 $Y=2.635
+ $X2=3.45 $Y2=2.34
r62 9 30 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=2.635
+ $X2=0.83 $Y2=2.72
r63 9 11 25.2345 $w=2.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.83 $Y=2.635
+ $X2=0.83 $Y2=2
r64 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=1.485 $X2=3.39 $Y2=2.34
r65 2 15 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=1.485 $X2=3.39 $Y2=1.66
r66 1 11 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.715
+ $Y=1.485 $X2=0.85 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%VGND 1 2 9 13 16 17 19 20 21 34 35 40
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r45 32 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r46 31 34 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r47 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r48 29 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r49 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r50 25 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r51 25 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r52 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 21 40 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r54 19 28 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.61
+ $Y2=0
r55 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.81
+ $Y2=0
r56 18 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.07
+ $Y2=0
r57 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.81
+ $Y2=0
r58 16 24 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.69
+ $Y2=0
r59 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.85
+ $Y2=0
r60 15 28 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.61
+ $Y2=0
r61 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.85
+ $Y2=0
r62 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0
r63 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.38
r64 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=0.085 $X2=0.85
+ $Y2=0
r65 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.85 $Y=0.085 $X2=0.85
+ $Y2=0.38
r66 2 13 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.615
+ $Y=0.235 $X2=1.81 $Y2=0.38
r67 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.715
+ $Y=0.235 $X2=0.85 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O32A_1%A_227_47# 1 2 3 12 14 15 16 17 18
c35 18 0 8.24349e-20 $X=3.305 $Y=0.36
c36 15 0 6.40318e-20 $X=1.47 $Y=0.74
r37 19 21 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0.36
+ $X2=2.375 $Y2=0.36
r38 18 19 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=3.305 $Y=0.36
+ $X2=2.54 $Y2=0.36
r39 17 23 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0.655
+ $X2=2.375 $Y2=0.74
r40 16 21 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=2.375 $Y=0.465
+ $X2=2.375 $Y2=0.36
r41 16 17 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.375 $Y=0.465
+ $X2=2.375 $Y2=0.655
r42 14 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0.74
+ $X2=2.375 $Y2=0.74
r43 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.21 $Y=0.74
+ $X2=1.47 $Y2=0.74
r44 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.305 $Y=0.655
+ $X2=1.47 $Y2=0.74
r45 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.305 $Y=0.655
+ $X2=1.305 $Y2=0.38
r46 3 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.235 $X2=3.39 $Y2=0.38
r47 2 23 182 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.375 $Y2=0.72
r48 2 21 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.375 $Y2=0.38
r49 1 12 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=1.135
+ $Y=0.235 $X2=1.305 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__sdlclkp_4.pxi.spice
* Created: Tue Sep  1 19:31:48 2020
* 
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%SCE N_SCE_M1027_g N_SCE_M1014_g SCE SCE
+ N_SCE_c_165_n PM_SKY130_FD_SC_HD__SDLCLKP_4%SCE
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%GATE N_GATE_M1005_g N_GATE_M1011_g GATE GATE
+ N_GATE_c_191_n N_GATE_c_192_n PM_SKY130_FD_SC_HD__SDLCLKP_4%GATE
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%A_257_147# N_A_257_147#_M1025_d
+ N_A_257_147#_M1002_d N_A_257_147#_M1007_g N_A_257_147#_M1010_g
+ N_A_257_147#_M1020_g N_A_257_147#_M1012_g N_A_257_147#_c_234_n
+ N_A_257_147#_c_235_n N_A_257_147#_c_236_n N_A_257_147#_c_237_n
+ N_A_257_147#_c_244_n N_A_257_147#_c_238_n N_A_257_147#_c_239_n
+ N_A_257_147#_c_240_n N_A_257_147#_c_241_n N_A_257_147#_c_246_n
+ N_A_257_147#_c_258_n N_A_257_147#_c_247_n N_A_257_147#_c_248_n
+ N_A_257_147#_c_249_n N_A_257_147#_c_250_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_4%A_257_147#
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%A_257_243# N_A_257_243#_M1020_s
+ N_A_257_243#_M1012_s N_A_257_243#_M1026_g N_A_257_243#_c_405_n
+ N_A_257_243#_c_406_n N_A_257_243#_M1022_g N_A_257_243#_c_407_n
+ N_A_257_243#_c_408_n N_A_257_243#_c_409_n N_A_257_243#_c_421_n
+ N_A_257_243#_c_410_n N_A_257_243#_c_411_n N_A_257_243#_c_412_n
+ N_A_257_243#_c_413_n N_A_257_243#_c_414_n N_A_257_243#_c_415_n
+ N_A_257_243#_c_416_n PM_SKY130_FD_SC_HD__SDLCLKP_4%A_257_243#
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%A_465_315# N_A_465_315#_M1008_d
+ N_A_465_315#_M1000_d N_A_465_315#_M1023_g N_A_465_315#_M1016_g
+ N_A_465_315#_M1017_g N_A_465_315#_M1013_g N_A_465_315#_c_528_n
+ N_A_465_315#_c_521_n N_A_465_315#_c_541_n N_A_465_315#_c_530_n
+ N_A_465_315#_c_522_n N_A_465_315#_c_523_n N_A_465_315#_c_533_n
+ N_A_465_315#_c_553_n N_A_465_315#_c_554_n N_A_465_315#_c_524_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_4%A_465_315#
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%A_287_413# N_A_287_413#_M1007_d
+ N_A_287_413#_M1026_d N_A_287_413#_c_649_n N_A_287_413#_M1008_g
+ N_A_287_413#_M1000_g N_A_287_413#_c_660_n N_A_287_413#_c_664_n
+ N_A_287_413#_c_655_n N_A_287_413#_c_650_n N_A_287_413#_c_651_n
+ N_A_287_413#_c_652_n N_A_287_413#_c_653_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_4%A_287_413#
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%CLK N_CLK_M1025_g N_CLK_c_748_n N_CLK_M1002_g
+ N_CLK_M1019_g N_CLK_M1006_g N_CLK_c_749_n N_CLK_c_750_n CLK N_CLK_c_752_n
+ N_CLK_c_753_n N_CLK_c_754_n N_CLK_c_755_n N_CLK_c_763_n N_CLK_c_756_n
+ N_CLK_c_757_n N_CLK_c_758_n PM_SKY130_FD_SC_HD__SDLCLKP_4%CLK
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%A_1045_47# N_A_1045_47#_M1017_s
+ N_A_1045_47#_M1013_d N_A_1045_47#_M1003_g N_A_1045_47#_M1001_g
+ N_A_1045_47#_M1004_g N_A_1045_47#_M1018_g N_A_1045_47#_M1009_g
+ N_A_1045_47#_M1021_g N_A_1045_47#_M1015_g N_A_1045_47#_M1024_g
+ N_A_1045_47#_c_865_n N_A_1045_47#_c_902_p N_A_1045_47#_c_853_n
+ N_A_1045_47#_c_861_n N_A_1045_47#_c_862_n N_A_1045_47#_c_854_n
+ N_A_1045_47#_c_886_n N_A_1045_47#_c_855_n N_A_1045_47#_c_856_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_4%A_1045_47#
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%VPWR N_VPWR_M1014_s N_VPWR_M1023_d
+ N_VPWR_M1012_d N_VPWR_M1013_s N_VPWR_M1006_d N_VPWR_M1018_s N_VPWR_M1024_s
+ N_VPWR_c_982_n N_VPWR_c_983_n N_VPWR_c_984_n N_VPWR_c_985_n N_VPWR_c_986_n
+ N_VPWR_c_987_n N_VPWR_c_988_n N_VPWR_c_989_n VPWR N_VPWR_c_990_n
+ N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_993_n N_VPWR_c_994_n N_VPWR_c_995_n
+ N_VPWR_c_996_n N_VPWR_c_997_n N_VPWR_c_998_n N_VPWR_c_981_n
+ PM_SKY130_FD_SC_HD__SDLCLKP_4%VPWR
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%A_27_47# N_A_27_47#_M1027_s N_A_27_47#_M1011_d
+ N_A_27_47#_M1005_d N_A_27_47#_c_1101_n N_A_27_47#_c_1102_n N_A_27_47#_c_1103_n
+ N_A_27_47#_c_1104_n N_A_27_47#_c_1113_n N_A_27_47#_c_1121_n
+ N_A_27_47#_c_1126_n PM_SKY130_FD_SC_HD__SDLCLKP_4%A_27_47#
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%GCLK N_GCLK_M1003_s N_GCLK_M1009_s
+ N_GCLK_M1001_d N_GCLK_M1021_d N_GCLK_c_1162_n N_GCLK_c_1153_n N_GCLK_c_1169_n
+ N_GCLK_c_1157_n N_GCLK_c_1154_n N_GCLK_c_1158_n GCLK GCLK GCLK GCLK GCLK GCLK
+ GCLK GCLK GCLK GCLK GCLK N_GCLK_c_1156_n GCLK
+ PM_SKY130_FD_SC_HD__SDLCLKP_4%GCLK
x_PM_SKY130_FD_SC_HD__SDLCLKP_4%VGND N_VGND_M1027_d N_VGND_M1016_d
+ N_VGND_M1020_d N_VGND_M1019_d N_VGND_M1004_d N_VGND_M1015_d N_VGND_c_1227_n
+ N_VGND_c_1228_n N_VGND_c_1229_n N_VGND_c_1230_n N_VGND_c_1231_n
+ N_VGND_c_1232_n VGND N_VGND_c_1233_n N_VGND_c_1234_n N_VGND_c_1235_n
+ N_VGND_c_1236_n N_VGND_c_1237_n N_VGND_c_1238_n N_VGND_c_1239_n
+ N_VGND_c_1240_n N_VGND_c_1241_n N_VGND_c_1242_n N_VGND_c_1243_n
+ N_VGND_c_1244_n PM_SKY130_FD_SC_HD__SDLCLKP_4%VGND
cc_1 VNB N_SCE_M1027_g 0.0353274f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB SCE 0.0153259f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_SCE_c_165_n 0.0342729f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_GATE_M1011_g 0.0276674f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_5 VNB N_GATE_c_191_n 0.0274229f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_GATE_c_192_n 0.00458727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_257_147#_M1007_g 0.0195404f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_257_147#_M1020_g 0.0381097f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_9 VNB N_A_257_147#_c_234_n 0.00683453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_257_147#_c_235_n 0.026946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_257_147#_c_236_n 7.53315e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_257_147#_c_237_n 0.00836697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_257_147#_c_238_n 0.00238438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_257_147#_c_239_n 0.00353827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_257_147#_c_240_n 0.00214693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_257_147#_c_241_n 0.0238041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_257_243#_c_405_n 0.0152184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_257_243#_c_406_n 0.00503808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_257_243#_c_407_n 0.0111999f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_20 VNB N_A_257_243#_c_408_n 0.00775325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_257_243#_c_409_n 0.00739084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_257_243#_c_410_n 0.0088014f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_257_243#_c_411_n 0.00127255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_257_243#_c_412_n 0.00212966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_257_243#_c_413_n 0.00439228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_257_243#_c_414_n 0.0269987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_257_243#_c_415_n 0.00250527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_257_243#_c_416_n 0.0189173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_465_315#_M1016_g 0.044686f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_30 VNB N_A_465_315#_c_521_n 0.00919858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_465_315#_c_522_n 0.00483489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_465_315#_c_523_n 0.0278504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_465_315#_c_524_n 0.0192398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_287_413#_c_649_n 0.0210888f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_35 VNB N_A_287_413#_c_650_n 0.0018369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_287_413#_c_651_n 0.00624625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_287_413#_c_652_n 0.00187427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_287_413#_c_653_n 0.0292321f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_CLK_c_748_n 0.0205002f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_40 VNB N_CLK_c_749_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_CLK_c_750_n 0.0310005f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_42 VNB CLK 0.00153552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_CLK_c_752_n 0.00833113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_CLK_c_753_n 0.00270586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_CLK_c_754_n 9.30759e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_CLK_c_755_n 0.0147459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_CLK_c_756_n 0.0208982f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_CLK_c_757_n 0.00284829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_CLK_c_758_n 0.0158351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1045_47#_M1003_g 0.0179524f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_51 VNB N_A_1045_47#_M1001_g 3.73613e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_52 VNB N_A_1045_47#_M1004_g 0.0174082f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_53 VNB N_A_1045_47#_M1018_g 4.10048e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1045_47#_M1009_g 0.0171786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1045_47#_M1021_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1045_47#_M1015_g 0.0237792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1045_47#_M1024_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1045_47#_c_853_n 0.0014625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1045_47#_c_854_n 0.0120421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1045_47#_c_855_n 0.00131861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1045_47#_c_856_n 0.067157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VPWR_c_981_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_27_47#_c_1101_n 0.0141581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_27_47#_c_1102_n 0.00400734f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_65 VNB N_A_27_47#_c_1103_n 0.00595497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_27_47#_c_1104_n 0.0102139f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_67 VNB N_GCLK_c_1153_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_68 VNB N_GCLK_c_1154_n 0.0019351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB GCLK 0.0186676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_GCLK_c_1156_n 6.23889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1227_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1228_n 0.00566378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1229_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1230_n 0.00171783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1231_n 0.0107756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1232_n 0.0338712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1233_n 0.0142589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1234_n 0.0434128f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1235_n 0.0281079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1236_n 0.0169301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1237_n 0.0163097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1238_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1239_n 0.00663229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1240_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1241_n 0.0275285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1242_n 0.0129759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1243_n 0.00353477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1244_n 0.399563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VPB N_SCE_M1014_g 0.0419371f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_90 VPB SCE 0.0189103f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_91 VPB N_SCE_c_165_n 0.0109907f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_92 VPB N_GATE_M1005_g 0.036273f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_93 VPB GATE 0.00670128f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_94 VPB N_GATE_c_191_n 0.00607012f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_95 VPB N_GATE_c_192_n 8.45903e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_257_147#_M1010_g 0.0211245f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_97 VPB N_A_257_147#_c_236_n 0.00354288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_257_147#_c_244_n 0.00505794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_257_147#_c_241_n 0.00658814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_257_147#_c_246_n 0.0171138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_257_147#_c_247_n 0.00400932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_257_147#_c_248_n 7.50236e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_257_147#_c_249_n 0.0266048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_257_147#_c_250_n 0.0455237f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_257_243#_M1026_g 0.0505653f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_106 VPB N_A_257_243#_c_405_n 0.0163673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_257_243#_c_406_n 0.00221973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_257_243#_c_409_n 0.00468468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_257_243#_c_421_n 0.00295382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_465_315#_M1023_g 0.022326f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_111 VPB N_A_465_315#_M1016_g 0.0170562f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_112 VPB N_A_465_315#_M1013_g 0.0224813f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_465_315#_c_528_n 0.0033307f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_114 VPB N_A_465_315#_c_521_n 0.00400259f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_465_315#_c_530_n 0.0178401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_465_315#_c_522_n 0.00730657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_465_315#_c_523_n 0.00797286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_465_315#_c_533_n 0.0310341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_287_413#_M1000_g 0.0243607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_287_413#_c_655_n 0.0134653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_287_413#_c_651_n 0.00269176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_287_413#_c_652_n 0.00386605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_287_413#_c_653_n 0.00831864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_CLK_M1006_g 0.019688f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_125 VPB N_CLK_c_753_n 5.24179e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_CLK_c_754_n 0.00130257f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_CLK_c_755_n 0.00846978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_CLK_c_763_n 0.0473815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_CLK_c_756_n 0.0041594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_CLK_c_757_n 0.001598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_1045_47#_M1001_g 0.0191428f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_132 VPB N_A_1045_47#_M1018_g 0.0193742f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_1045_47#_M1021_g 0.0191015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_1045_47#_M1024_g 0.0267109f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_1045_47#_c_861_n 0.00159926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_1045_47#_c_862_n 0.00384171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_982_n 0.0098838f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_138 VPB N_VPWR_c_983_n 0.0318467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_984_n 0.00217662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_985_n 0.00165706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_986_n 0.0107497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_987_n 0.0480068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_988_n 0.013173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_989_n 0.0144538f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_990_n 0.0332603f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_991_n 0.0135857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_992_n 0.0158942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_993_n 0.0163094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_994_n 0.0487185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_995_n 0.0138172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_996_n 0.00455555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_997_n 0.00521963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_998_n 0.00353672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_981_n 0.0449635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_27_47#_c_1102_n 0.00313483f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_156 VPB N_GCLK_c_1157_n 0.00117749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_GCLK_c_1158_n 0.002754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB GCLK 0.00300463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB GCLK 0.00129449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB GCLK 0.00689571f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 N_SCE_M1014_g N_GATE_M1005_g 0.0495303f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_162 N_SCE_M1027_g N_GATE_M1011_g 0.0256093f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_163 N_SCE_c_165_n GATE 4.13543e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_164 N_SCE_c_165_n N_GATE_c_191_n 0.0495303f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_165 N_SCE_M1027_g N_GATE_c_192_n 4.13543e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_166 N_SCE_M1014_g N_VPWR_c_983_n 0.00472725f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_167 SCE N_VPWR_c_983_n 0.0242525f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_168 N_SCE_c_165_n N_VPWR_c_983_n 9.03791e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_169 N_SCE_M1014_g N_VPWR_c_994_n 0.00539841f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_170 N_SCE_M1014_g N_VPWR_c_981_n 0.0103231f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_171 N_SCE_M1027_g N_A_27_47#_c_1102_n 0.00889944f $X=0.47 $Y=0.445 $X2=0
+ $Y2=0
cc_172 N_SCE_M1014_g N_A_27_47#_c_1102_n 0.0181923f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_173 SCE N_A_27_47#_c_1102_n 0.0511821f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_174 N_SCE_c_165_n N_A_27_47#_c_1102_n 0.00719527f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_175 N_SCE_M1027_g N_A_27_47#_c_1104_n 0.0159826f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_176 SCE N_A_27_47#_c_1104_n 0.0218663f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_177 N_SCE_c_165_n N_A_27_47#_c_1104_n 0.00331025f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_178 N_SCE_M1014_g N_A_27_47#_c_1113_n 0.0070608f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_179 N_SCE_M1027_g N_VGND_c_1227_n 0.00809304f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_180 N_SCE_M1027_g N_VGND_c_1233_n 0.00337001f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_181 N_SCE_M1027_g N_VGND_c_1244_n 0.00485988f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_182 N_GATE_M1011_g N_A_257_147#_M1007_g 0.0143632f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_183 N_GATE_M1011_g N_A_257_147#_c_234_n 9.82505e-19 $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_184 N_GATE_c_191_n N_A_257_147#_c_234_n 0.00116699f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_GATE_c_192_n N_A_257_147#_c_234_n 0.0305181f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_186 N_GATE_M1011_g N_A_257_147#_c_235_n 0.0095729f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_187 N_GATE_c_191_n N_A_257_147#_c_235_n 6.18885e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_GATE_c_192_n N_A_257_147#_c_235_n 3.98477e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_189 GATE N_A_257_147#_c_258_n 0.00134565f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_190 N_GATE_c_192_n N_A_257_147#_c_258_n 2.00479e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_GATE_M1005_g N_A_257_147#_c_247_n 4.36779e-19 $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_192 GATE N_A_257_147#_c_247_n 0.0404082f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_193 N_GATE_c_192_n N_A_257_147#_c_247_n 0.00784692f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_194 GATE N_A_257_243#_M1026_g 0.00459698f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_195 N_GATE_M1005_g N_A_257_243#_c_406_n 0.0258836f $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_196 N_GATE_c_191_n N_A_257_243#_c_406_n 0.00719003f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_197 N_GATE_c_192_n N_A_257_243#_c_406_n 0.00194283f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_GATE_M1005_g N_VPWR_c_994_n 0.00357877f $X=0.83 $Y=2.165 $X2=0 $Y2=0
cc_199 N_GATE_M1005_g N_VPWR_c_981_n 0.00536442f $X=0.83 $Y=2.165 $X2=0 $Y2=0
cc_200 GATE N_A_27_47#_M1005_d 0.00345627f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_201 N_GATE_M1011_g N_A_27_47#_c_1102_n 0.00390472f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_GATE_c_191_n N_A_27_47#_c_1102_n 0.00960649f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_GATE_c_192_n N_A_27_47#_c_1102_n 0.0754313f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_204 N_GATE_M1011_g N_A_27_47#_c_1103_n 0.0123694f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_GATE_c_191_n N_A_27_47#_c_1103_n 0.00311345f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_206 N_GATE_c_192_n N_A_27_47#_c_1103_n 0.028952f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_207 N_GATE_M1005_g N_A_27_47#_c_1121_n 0.0145681f $X=0.83 $Y=2.165 $X2=0
+ $Y2=0
cc_208 GATE N_A_27_47#_c_1121_n 0.0261201f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_209 N_GATE_M1011_g N_VGND_c_1227_n 0.00763365f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_210 N_GATE_M1011_g N_VGND_c_1234_n 0.00337001f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_211 N_GATE_M1011_g N_VGND_c_1244_n 0.00408452f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_212 N_A_257_147#_M1010_g N_A_257_243#_M1026_g 0.0138034f $X=1.84 $Y=2.275
+ $X2=0 $Y2=0
cc_213 N_A_257_147#_c_247_n N_A_257_243#_M1026_g 0.0149237f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_214 N_A_257_147#_c_249_n N_A_257_243#_M1026_g 0.021304f $X=1.78 $Y=1.74 $X2=0
+ $Y2=0
cc_215 N_A_257_147#_c_240_n N_A_257_243#_c_405_n 0.0105586f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_216 N_A_257_147#_c_246_n N_A_257_243#_c_405_n 0.00213361f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_217 N_A_257_147#_c_247_n N_A_257_243#_c_405_n 0.00868281f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_218 N_A_257_147#_c_249_n N_A_257_243#_c_405_n 0.0180583f $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_219 N_A_257_147#_c_235_n N_A_257_243#_c_406_n 0.0227923f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_220 N_A_257_147#_c_240_n N_A_257_243#_c_406_n 0.0043361f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_221 N_A_257_147#_c_247_n N_A_257_243#_c_406_n 4.45536e-19 $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_222 N_A_257_147#_c_240_n N_A_257_243#_c_407_n 0.00150324f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_223 N_A_257_147#_M1020_g N_A_257_243#_c_408_n 0.00282429f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_224 N_A_257_147#_c_238_n N_A_257_243#_c_408_n 0.00771195f $X=4.72 $Y=0.615
+ $X2=0 $Y2=0
cc_225 N_A_257_147#_M1020_g N_A_257_243#_c_409_n 0.00236246f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_226 N_A_257_147#_c_236_n N_A_257_243#_c_409_n 0.0101973f $X=4.327 $Y=1.495
+ $X2=0 $Y2=0
cc_227 N_A_257_147#_c_237_n N_A_257_243#_c_409_n 0.0193569f $X=4.335 $Y=1.105
+ $X2=0 $Y2=0
cc_228 N_A_257_147#_c_241_n N_A_257_243#_c_409_n 0.00376938f $X=4.1 $Y=1.19
+ $X2=0 $Y2=0
cc_229 N_A_257_147#_c_246_n N_A_257_243#_c_409_n 0.0104083f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_230 N_A_257_147#_c_248_n N_A_257_243#_c_409_n 2.68226e-19 $X=4.395 $Y=1.53
+ $X2=0 $Y2=0
cc_231 N_A_257_147#_c_250_n N_A_257_243#_c_409_n 0.00385034f $X=4.1 $Y=1.325
+ $X2=0 $Y2=0
cc_232 N_A_257_147#_c_236_n N_A_257_243#_c_421_n 0.00660951f $X=4.327 $Y=1.495
+ $X2=0 $Y2=0
cc_233 N_A_257_147#_c_237_n N_A_257_243#_c_421_n 0.00185537f $X=4.335 $Y=1.105
+ $X2=0 $Y2=0
cc_234 N_A_257_147#_c_241_n N_A_257_243#_c_421_n 7.57315e-19 $X=4.1 $Y=1.19
+ $X2=0 $Y2=0
cc_235 N_A_257_147#_c_246_n N_A_257_243#_c_421_n 0.00988437f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_236 N_A_257_147#_c_248_n N_A_257_243#_c_421_n 2.78941e-19 $X=4.395 $Y=1.53
+ $X2=0 $Y2=0
cc_237 N_A_257_147#_c_250_n N_A_257_243#_c_421_n 0.00246207f $X=4.1 $Y=1.325
+ $X2=0 $Y2=0
cc_238 N_A_257_147#_c_246_n N_A_257_243#_c_410_n 0.0694573f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_239 N_A_257_147#_c_234_n N_A_257_243#_c_411_n 0.00155066f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_240 N_A_257_147#_c_246_n N_A_257_243#_c_411_n 0.0132091f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_241 N_A_257_147#_M1020_g N_A_257_243#_c_412_n 0.00504445f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_242 N_A_257_147#_c_237_n N_A_257_243#_c_412_n 0.00817201f $X=4.335 $Y=1.105
+ $X2=0 $Y2=0
cc_243 N_A_257_147#_c_238_n N_A_257_243#_c_412_n 0.00144026f $X=4.72 $Y=0.615
+ $X2=0 $Y2=0
cc_244 N_A_257_147#_c_241_n N_A_257_243#_c_412_n 7.14969e-19 $X=4.1 $Y=1.19
+ $X2=0 $Y2=0
cc_245 N_A_257_147#_c_246_n N_A_257_243#_c_412_n 0.0150763f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_246 N_A_257_147#_M1020_g N_A_257_243#_c_413_n 0.00636449f $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_247 N_A_257_147#_c_237_n N_A_257_243#_c_413_n 0.0148946f $X=4.335 $Y=1.105
+ $X2=0 $Y2=0
cc_248 N_A_257_147#_c_238_n N_A_257_243#_c_413_n 0.00132326f $X=4.72 $Y=0.615
+ $X2=0 $Y2=0
cc_249 N_A_257_147#_c_241_n N_A_257_243#_c_413_n 8.95761e-19 $X=4.1 $Y=1.19
+ $X2=0 $Y2=0
cc_250 N_A_257_147#_c_246_n N_A_257_243#_c_413_n 9.85771e-19 $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_251 N_A_257_147#_c_234_n N_A_257_243#_c_414_n 0.00708004f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_252 N_A_257_147#_c_235_n N_A_257_243#_c_414_n 0.0165261f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_253 N_A_257_147#_c_246_n N_A_257_243#_c_414_n 8.52878e-19 $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_254 N_A_257_147#_c_234_n N_A_257_243#_c_415_n 0.0242697f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_255 N_A_257_147#_c_235_n N_A_257_243#_c_415_n 2.60953e-19 $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_256 N_A_257_147#_c_246_n N_A_257_243#_c_415_n 0.00446365f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_257 N_A_257_147#_M1007_g N_A_257_243#_c_416_n 0.0107241f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_258 N_A_257_147#_c_246_n N_A_465_315#_M1000_d 3.75899e-19 $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_259 N_A_257_147#_M1010_g N_A_465_315#_M1023_g 0.0155568f $X=1.84 $Y=2.275
+ $X2=0 $Y2=0
cc_260 N_A_257_147#_c_246_n N_A_465_315#_M1016_g 0.00428067f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_261 N_A_257_147#_c_244_n N_A_465_315#_M1013_g 0.00101581f $X=4.81 $Y=1.66
+ $X2=0 $Y2=0
cc_262 N_A_257_147#_c_246_n N_A_465_315#_c_528_n 0.0228159f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_263 N_A_257_147#_M1020_g N_A_465_315#_c_521_n 4.88693e-19 $X=4.05 $Y=0.445
+ $X2=0 $Y2=0
cc_264 N_A_257_147#_c_246_n N_A_465_315#_c_521_n 0.0272857f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_265 N_A_257_147#_c_250_n N_A_465_315#_c_541_n 0.00465884f $X=4.1 $Y=1.325
+ $X2=0 $Y2=0
cc_266 N_A_257_147#_M1002_d N_A_465_315#_c_530_n 0.00477298f $X=4.675 $Y=1.515
+ $X2=0 $Y2=0
cc_267 N_A_257_147#_c_236_n N_A_465_315#_c_530_n 0.0210881f $X=4.327 $Y=1.495
+ $X2=0 $Y2=0
cc_268 N_A_257_147#_c_237_n N_A_465_315#_c_530_n 0.00128309f $X=4.335 $Y=1.105
+ $X2=0 $Y2=0
cc_269 N_A_257_147#_c_244_n N_A_465_315#_c_530_n 0.0282344f $X=4.81 $Y=1.66
+ $X2=0 $Y2=0
cc_270 N_A_257_147#_c_241_n N_A_465_315#_c_530_n 2.59847e-19 $X=4.1 $Y=1.19
+ $X2=0 $Y2=0
cc_271 N_A_257_147#_c_246_n N_A_465_315#_c_530_n 0.0139938f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_272 N_A_257_147#_c_248_n N_A_465_315#_c_530_n 0.00169866f $X=4.395 $Y=1.53
+ $X2=0 $Y2=0
cc_273 N_A_257_147#_c_250_n N_A_465_315#_c_530_n 0.0145602f $X=4.1 $Y=1.325
+ $X2=0 $Y2=0
cc_274 N_A_257_147#_c_244_n N_A_465_315#_c_522_n 0.0203633f $X=4.81 $Y=1.66
+ $X2=0 $Y2=0
cc_275 N_A_257_147#_c_246_n N_A_465_315#_c_533_n 0.0039188f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_276 N_A_257_147#_c_249_n N_A_465_315#_c_533_n 0.00753208f $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_277 N_A_257_147#_c_246_n N_A_465_315#_c_553_n 0.00517255f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_278 N_A_257_147#_c_250_n N_A_465_315#_c_554_n 0.00335885f $X=4.1 $Y=1.325
+ $X2=0 $Y2=0
cc_279 N_A_257_147#_c_246_n N_A_287_413#_M1000_g 0.00751079f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_280 N_A_257_147#_M1007_g N_A_287_413#_c_660_n 0.00581419f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_281 N_A_257_147#_c_234_n N_A_287_413#_c_660_n 0.0249382f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_282 N_A_257_147#_c_235_n N_A_287_413#_c_660_n 9.8177e-19 $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_283 N_A_257_147#_c_240_n N_A_287_413#_c_660_n 0.00398233f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_284 N_A_257_147#_M1010_g N_A_287_413#_c_664_n 0.0131252f $X=1.84 $Y=2.275
+ $X2=0 $Y2=0
cc_285 N_A_257_147#_c_246_n N_A_287_413#_c_664_n 0.00594058f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_286 N_A_257_147#_c_258_n N_A_287_413#_c_664_n 0.00121651f $X=1.76 $Y=1.53
+ $X2=0 $Y2=0
cc_287 N_A_257_147#_c_247_n N_A_287_413#_c_664_n 0.0302261f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_288 N_A_257_147#_c_249_n N_A_287_413#_c_664_n 6.45937e-19 $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_289 N_A_257_147#_c_246_n N_A_287_413#_c_655_n 0.0205826f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_290 N_A_257_147#_c_258_n N_A_287_413#_c_655_n 5.20192e-19 $X=1.76 $Y=1.53
+ $X2=0 $Y2=0
cc_291 N_A_257_147#_c_247_n N_A_287_413#_c_655_n 0.0436285f $X=1.615 $Y=1.53
+ $X2=0 $Y2=0
cc_292 N_A_257_147#_c_249_n N_A_287_413#_c_655_n 0.00709868f $X=1.78 $Y=1.74
+ $X2=0 $Y2=0
cc_293 N_A_257_147#_c_234_n N_A_287_413#_c_651_n 0.00602675f $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_294 N_A_257_147#_c_240_n N_A_287_413#_c_651_n 0.0146898f $X=1.615 $Y=1.325
+ $X2=0 $Y2=0
cc_295 N_A_257_147#_c_246_n N_A_287_413#_c_651_n 0.00783084f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_296 N_A_257_147#_c_246_n N_A_287_413#_c_652_n 0.00746407f $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_297 N_A_257_147#_c_246_n N_A_287_413#_c_653_n 3.55037e-19 $X=4.25 $Y=1.53
+ $X2=0 $Y2=0
cc_298 N_A_257_147#_M1020_g N_CLK_c_748_n 0.00386856f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_299 N_A_257_147#_c_237_n N_CLK_c_748_n 0.00634405f $X=4.335 $Y=1.105 $X2=0
+ $Y2=0
cc_300 N_A_257_147#_c_241_n N_CLK_c_748_n 0.0128434f $X=4.1 $Y=1.19 $X2=0 $Y2=0
cc_301 N_A_257_147#_M1020_g N_CLK_c_749_n 0.0199171f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_302 N_A_257_147#_c_238_n N_CLK_c_749_n 0.00705718f $X=4.72 $Y=0.615 $X2=0
+ $Y2=0
cc_303 N_A_257_147#_c_237_n N_CLK_c_750_n 0.00792429f $X=4.335 $Y=1.105 $X2=0
+ $Y2=0
cc_304 N_A_257_147#_c_244_n N_CLK_c_750_n 9.73222e-19 $X=4.81 $Y=1.66 $X2=0
+ $Y2=0
cc_305 N_A_257_147#_c_238_n N_CLK_c_750_n 0.0202151f $X=4.72 $Y=0.615 $X2=0
+ $Y2=0
cc_306 N_A_257_147#_c_239_n N_CLK_c_750_n 0.00148768f $X=4.68 $Y=0.465 $X2=0
+ $Y2=0
cc_307 N_A_257_147#_c_248_n N_CLK_c_750_n 0.00109922f $X=4.395 $Y=1.53 $X2=0
+ $Y2=0
cc_308 N_A_257_147#_c_236_n CLK 0.00244552f $X=4.327 $Y=1.495 $X2=0 $Y2=0
cc_309 N_A_257_147#_c_237_n CLK 0.0137996f $X=4.335 $Y=1.105 $X2=0 $Y2=0
cc_310 N_A_257_147#_c_244_n CLK 0.015439f $X=4.81 $Y=1.66 $X2=0 $Y2=0
cc_311 N_A_257_147#_c_238_n CLK 0.00653509f $X=4.72 $Y=0.615 $X2=0 $Y2=0
cc_312 N_A_257_147#_c_241_n CLK 2.84827e-19 $X=4.1 $Y=1.19 $X2=0 $Y2=0
cc_313 N_A_257_147#_c_236_n N_CLK_c_753_n 7.32681e-19 $X=4.327 $Y=1.495 $X2=0
+ $Y2=0
cc_314 N_A_257_147#_c_237_n N_CLK_c_753_n 0.00548008f $X=4.335 $Y=1.105 $X2=0
+ $Y2=0
cc_315 N_A_257_147#_c_244_n N_CLK_c_753_n 0.00376482f $X=4.81 $Y=1.66 $X2=0
+ $Y2=0
cc_316 N_A_257_147#_c_238_n N_CLK_c_753_n 0.00120125f $X=4.72 $Y=0.615 $X2=0
+ $Y2=0
cc_317 N_A_257_147#_c_236_n N_CLK_c_755_n 0.00491164f $X=4.327 $Y=1.495 $X2=0
+ $Y2=0
cc_318 N_A_257_147#_c_244_n N_CLK_c_755_n 0.00772226f $X=4.81 $Y=1.66 $X2=0
+ $Y2=0
cc_319 N_A_257_147#_c_244_n N_CLK_c_763_n 0.0159058f $X=4.81 $Y=1.66 $X2=0 $Y2=0
cc_320 N_A_257_147#_c_248_n N_CLK_c_763_n 0.00429027f $X=4.395 $Y=1.53 $X2=0
+ $Y2=0
cc_321 N_A_257_147#_c_250_n N_CLK_c_763_n 0.0381082f $X=4.1 $Y=1.325 $X2=0 $Y2=0
cc_322 N_A_257_147#_c_238_n N_A_1045_47#_c_854_n 0.0148333f $X=4.72 $Y=0.615
+ $X2=0 $Y2=0
cc_323 N_A_257_147#_c_239_n N_A_1045_47#_c_854_n 0.0299163f $X=4.68 $Y=0.465
+ $X2=0 $Y2=0
cc_324 N_A_257_147#_c_246_n N_VPWR_M1023_d 0.0020643f $X=4.25 $Y=1.53 $X2=0
+ $Y2=0
cc_325 N_A_257_147#_c_236_n N_VPWR_M1012_d 0.00511429f $X=4.327 $Y=1.495 $X2=0
+ $Y2=0
cc_326 N_A_257_147#_c_246_n N_VPWR_M1012_d 4.60476e-19 $X=4.25 $Y=1.53 $X2=0
+ $Y2=0
cc_327 N_A_257_147#_c_250_n N_VPWR_c_990_n 0.0230773f $X=4.1 $Y=1.325 $X2=0
+ $Y2=0
cc_328 N_A_257_147#_M1010_g N_VPWR_c_994_n 0.00357877f $X=1.84 $Y=2.275 $X2=0
+ $Y2=0
cc_329 N_A_257_147#_M1010_g N_VPWR_c_995_n 0.00145256f $X=1.84 $Y=2.275 $X2=0
+ $Y2=0
cc_330 N_A_257_147#_c_246_n N_VPWR_c_995_n 7.31718e-19 $X=4.25 $Y=1.53 $X2=0
+ $Y2=0
cc_331 N_A_257_147#_M1010_g N_VPWR_c_981_n 0.00579685f $X=1.84 $Y=2.275 $X2=0
+ $Y2=0
cc_332 N_A_257_147#_c_247_n N_VPWR_c_981_n 0.00150144f $X=1.615 $Y=1.53 $X2=0
+ $Y2=0
cc_333 N_A_257_147#_M1007_g N_A_27_47#_c_1103_n 0.0029712f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_334 N_A_257_147#_c_234_n N_A_27_47#_c_1103_n 0.0067219f $X=1.45 $Y=0.87 $X2=0
+ $Y2=0
cc_335 N_A_257_147#_c_235_n N_A_27_47#_c_1103_n 4.43441e-19 $X=1.45 $Y=0.87
+ $X2=0 $Y2=0
cc_336 N_A_257_147#_M1007_g N_A_27_47#_c_1126_n 0.00382934f $X=1.375 $Y=0.415
+ $X2=0 $Y2=0
cc_337 N_A_257_147#_c_238_n N_VGND_M1020_d 0.00192931f $X=4.72 $Y=0.615 $X2=0
+ $Y2=0
cc_338 N_A_257_147#_M1007_g N_VGND_c_1227_n 0.00109585f $X=1.375 $Y=0.415 $X2=0
+ $Y2=0
cc_339 N_A_257_147#_M1020_g N_VGND_c_1229_n 0.00853729f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_340 N_A_257_147#_c_237_n N_VGND_c_1229_n 0.00151747f $X=4.335 $Y=1.105 $X2=0
+ $Y2=0
cc_341 N_A_257_147#_c_238_n N_VGND_c_1229_n 0.0132365f $X=4.72 $Y=0.615 $X2=0
+ $Y2=0
cc_342 N_A_257_147#_c_241_n N_VGND_c_1229_n 8.45001e-19 $X=4.1 $Y=1.19 $X2=0
+ $Y2=0
cc_343 N_A_257_147#_M1007_g N_VGND_c_1234_n 0.00456464f $X=1.375 $Y=0.415 $X2=0
+ $Y2=0
cc_344 N_A_257_147#_c_235_n N_VGND_c_1234_n 2.64403e-19 $X=1.45 $Y=0.87 $X2=0
+ $Y2=0
cc_345 N_A_257_147#_M1020_g N_VGND_c_1235_n 0.0046653f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_346 N_A_257_147#_c_238_n N_VGND_c_1241_n 0.00258611f $X=4.72 $Y=0.615 $X2=0
+ $Y2=0
cc_347 N_A_257_147#_c_239_n N_VGND_c_1241_n 0.0165187f $X=4.68 $Y=0.465 $X2=0
+ $Y2=0
cc_348 N_A_257_147#_M1025_d N_VGND_c_1244_n 0.00227267f $X=4.545 $Y=0.235 $X2=0
+ $Y2=0
cc_349 N_A_257_147#_M1007_g N_VGND_c_1244_n 0.00806939f $X=1.375 $Y=0.415 $X2=0
+ $Y2=0
cc_350 N_A_257_147#_M1020_g N_VGND_c_1244_n 0.0060162f $X=4.05 $Y=0.445 $X2=0
+ $Y2=0
cc_351 N_A_257_147#_c_235_n N_VGND_c_1244_n 3.49206e-19 $X=1.45 $Y=0.87 $X2=0
+ $Y2=0
cc_352 N_A_257_147#_c_238_n N_VGND_c_1244_n 0.00544468f $X=4.72 $Y=0.615 $X2=0
+ $Y2=0
cc_353 N_A_257_147#_c_239_n N_VGND_c_1244_n 0.00940011f $X=4.68 $Y=0.465 $X2=0
+ $Y2=0
cc_354 N_A_257_243#_c_410_n N_A_465_315#_M1008_d 5.81953e-19 $X=3.79 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_355 N_A_257_243#_c_407_n N_A_465_315#_M1016_g 0.00692236f $X=1.9 $Y=1.215
+ $X2=0 $Y2=0
cc_356 N_A_257_243#_c_410_n N_A_465_315#_M1016_g 0.00342271f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_357 N_A_257_243#_c_414_n N_A_465_315#_M1016_g 0.0115616f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_358 N_A_257_243#_c_415_n N_A_465_315#_M1016_g 7.79891e-19 $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_359 N_A_257_243#_c_416_n N_A_465_315#_M1016_g 0.0139526f $X=1.96 $Y=0.705
+ $X2=0 $Y2=0
cc_360 N_A_257_243#_c_408_n N_A_465_315#_c_521_n 0.0925201f $X=3.84 $Y=0.465
+ $X2=0 $Y2=0
cc_361 N_A_257_243#_c_421_n N_A_465_315#_c_521_n 0.0041125f $X=3.84 $Y=1.66
+ $X2=0 $Y2=0
cc_362 N_A_257_243#_c_410_n N_A_465_315#_c_521_n 0.0209841f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_363 N_A_257_243#_c_412_n N_A_465_315#_c_521_n 2.94771e-19 $X=3.935 $Y=0.85
+ $X2=0 $Y2=0
cc_364 N_A_257_243#_M1012_s N_A_465_315#_c_530_n 0.00486982f $X=3.715 $Y=1.515
+ $X2=0 $Y2=0
cc_365 N_A_257_243#_c_421_n N_A_465_315#_c_530_n 0.0240477f $X=3.84 $Y=1.66
+ $X2=0 $Y2=0
cc_366 N_A_257_243#_c_421_n N_A_465_315#_c_554_n 0.00889195f $X=3.84 $Y=1.66
+ $X2=0 $Y2=0
cc_367 N_A_257_243#_c_410_n N_A_287_413#_c_649_n 0.00847687f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_368 N_A_257_243#_c_421_n N_A_287_413#_M1000_g 5.00151e-19 $X=3.84 $Y=1.66
+ $X2=0 $Y2=0
cc_369 N_A_257_243#_c_405_n N_A_287_413#_c_660_n 7.07243e-19 $X=1.825 $Y=1.29
+ $X2=0 $Y2=0
cc_370 N_A_257_243#_c_410_n N_A_287_413#_c_660_n 0.00173863f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_371 N_A_257_243#_c_411_n N_A_287_413#_c_660_n 0.0020338f $X=2.22 $Y=0.85
+ $X2=0 $Y2=0
cc_372 N_A_257_243#_c_414_n N_A_287_413#_c_660_n 0.00258224f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_373 N_A_257_243#_c_415_n N_A_287_413#_c_660_n 0.0175669f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_374 N_A_257_243#_c_416_n N_A_287_413#_c_660_n 0.0128508f $X=1.96 $Y=0.705
+ $X2=0 $Y2=0
cc_375 N_A_257_243#_M1026_g N_A_287_413#_c_664_n 0.00300964f $X=1.36 $Y=2.275
+ $X2=0 $Y2=0
cc_376 N_A_257_243#_M1026_g N_A_287_413#_c_655_n 6.3244e-19 $X=1.36 $Y=2.275
+ $X2=0 $Y2=0
cc_377 N_A_257_243#_c_410_n N_A_287_413#_c_650_n 0.0162752f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_378 N_A_257_243#_c_411_n N_A_287_413#_c_650_n 0.00275249f $X=2.22 $Y=0.85
+ $X2=0 $Y2=0
cc_379 N_A_257_243#_c_414_n N_A_287_413#_c_650_n 7.44567e-19 $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_380 N_A_257_243#_c_415_n N_A_287_413#_c_650_n 0.0205672f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_381 N_A_257_243#_c_416_n N_A_287_413#_c_650_n 0.00302624f $X=1.96 $Y=0.705
+ $X2=0 $Y2=0
cc_382 N_A_257_243#_c_407_n N_A_287_413#_c_651_n 0.00377955f $X=1.9 $Y=1.215
+ $X2=0 $Y2=0
cc_383 N_A_257_243#_c_410_n N_A_287_413#_c_651_n 0.00154998f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_384 N_A_257_243#_c_411_n N_A_287_413#_c_651_n 0.00160742f $X=2.22 $Y=0.85
+ $X2=0 $Y2=0
cc_385 N_A_257_243#_c_414_n N_A_287_413#_c_651_n 0.00153556f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_386 N_A_257_243#_c_415_n N_A_287_413#_c_651_n 0.0128543f $X=1.96 $Y=0.87
+ $X2=0 $Y2=0
cc_387 N_A_257_243#_c_410_n N_A_287_413#_c_652_n 0.0106635f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_388 N_A_257_243#_c_410_n N_A_287_413#_c_653_n 0.0044627f $X=3.79 $Y=0.85
+ $X2=0 $Y2=0
cc_389 N_A_257_243#_M1026_g N_VPWR_c_994_n 0.00577801f $X=1.36 $Y=2.275 $X2=0
+ $Y2=0
cc_390 N_A_257_243#_M1026_g N_VPWR_c_981_n 0.0103326f $X=1.36 $Y=2.275 $X2=0
+ $Y2=0
cc_391 N_A_257_243#_c_410_n N_VGND_M1016_d 4.25819e-19 $X=3.79 $Y=0.85 $X2=0
+ $Y2=0
cc_392 N_A_257_243#_c_410_n N_VGND_c_1228_n 0.0140576f $X=3.79 $Y=0.85 $X2=0
+ $Y2=0
cc_393 N_A_257_243#_c_416_n N_VGND_c_1234_n 0.00357877f $X=1.96 $Y=0.705 $X2=0
+ $Y2=0
cc_394 N_A_257_243#_c_408_n N_VGND_c_1235_n 0.0230197f $X=3.84 $Y=0.465 $X2=0
+ $Y2=0
cc_395 N_A_257_243#_M1020_s N_VGND_c_1244_n 0.0018314f $X=3.715 $Y=0.235 $X2=0
+ $Y2=0
cc_396 N_A_257_243#_c_408_n N_VGND_c_1244_n 0.00590194f $X=3.84 $Y=0.465 $X2=0
+ $Y2=0
cc_397 N_A_257_243#_c_410_n N_VGND_c_1244_n 0.0735105f $X=3.79 $Y=0.85 $X2=0
+ $Y2=0
cc_398 N_A_257_243#_c_411_n N_VGND_c_1244_n 0.014828f $X=2.22 $Y=0.85 $X2=0
+ $Y2=0
cc_399 N_A_257_243#_c_412_n N_VGND_c_1244_n 0.0153387f $X=3.935 $Y=0.85 $X2=0
+ $Y2=0
cc_400 N_A_257_243#_c_413_n N_VGND_c_1244_n 8.78282e-19 $X=3.935 $Y=0.85 $X2=0
+ $Y2=0
cc_401 N_A_257_243#_c_416_n N_VGND_c_1244_n 0.00589934f $X=1.96 $Y=0.705 $X2=0
+ $Y2=0
cc_402 N_A_465_315#_M1016_g N_A_287_413#_c_649_n 0.0188679f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_465_315#_c_521_n N_A_287_413#_c_649_n 0.0293052f $X=3.32 $Y=0.42
+ $X2=0 $Y2=0
cc_404 N_A_465_315#_M1023_g N_A_287_413#_M1000_g 0.0129074f $X=2.43 $Y=2.275
+ $X2=0 $Y2=0
cc_405 N_A_465_315#_M1016_g N_A_287_413#_M1000_g 0.00670688f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_406 N_A_465_315#_c_528_n N_A_287_413#_M1000_g 0.014093f $X=3.185 $Y=1.77
+ $X2=0 $Y2=0
cc_407 N_A_465_315#_c_533_n N_A_287_413#_M1000_g 0.00808806f $X=2.46 $Y=1.74
+ $X2=0 $Y2=0
cc_408 N_A_465_315#_c_553_n N_A_287_413#_M1000_g 2.06052e-19 $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_409 N_A_465_315#_c_554_n N_A_287_413#_M1000_g 0.00982347f $X=3.295 $Y=1.86
+ $X2=0 $Y2=0
cc_410 N_A_465_315#_M1016_g N_A_287_413#_c_660_n 0.00893118f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_411 N_A_465_315#_M1023_g N_A_287_413#_c_664_n 0.00282173f $X=2.43 $Y=2.275
+ $X2=0 $Y2=0
cc_412 N_A_465_315#_M1023_g N_A_287_413#_c_655_n 0.00426352f $X=2.43 $Y=2.275
+ $X2=0 $Y2=0
cc_413 N_A_465_315#_M1016_g N_A_287_413#_c_655_n 0.00550388f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_414 N_A_465_315#_c_533_n N_A_287_413#_c_655_n 0.00271662f $X=2.46 $Y=1.74
+ $X2=0 $Y2=0
cc_415 N_A_465_315#_c_553_n N_A_287_413#_c_655_n 0.0255746f $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_416 N_A_465_315#_M1016_g N_A_287_413#_c_650_n 0.0114396f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_465_315#_M1016_g N_A_287_413#_c_651_n 0.00791638f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_418 N_A_465_315#_c_533_n N_A_287_413#_c_651_n 0.00300149f $X=2.46 $Y=1.74
+ $X2=0 $Y2=0
cc_419 N_A_465_315#_c_553_n N_A_287_413#_c_651_n 0.00700208f $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_420 N_A_465_315#_M1016_g N_A_287_413#_c_652_n 0.00928658f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_421 N_A_465_315#_c_528_n N_A_287_413#_c_652_n 0.0171291f $X=3.185 $Y=1.77
+ $X2=0 $Y2=0
cc_422 N_A_465_315#_c_521_n N_A_287_413#_c_652_n 0.0310043f $X=3.32 $Y=0.42
+ $X2=0 $Y2=0
cc_423 N_A_465_315#_c_553_n N_A_287_413#_c_652_n 0.00230595f $X=2.545 $Y=1.74
+ $X2=0 $Y2=0
cc_424 N_A_465_315#_M1016_g N_A_287_413#_c_653_n 0.0213485f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_425 N_A_465_315#_c_528_n N_A_287_413#_c_653_n 0.00123339f $X=3.185 $Y=1.77
+ $X2=0 $Y2=0
cc_426 N_A_465_315#_c_522_n N_CLK_c_748_n 0.00112992f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_427 N_A_465_315#_c_523_n N_CLK_c_748_n 0.0131589f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_428 N_A_465_315#_M1013_g N_CLK_M1006_g 0.03873f $X=5.56 $Y=1.985 $X2=0 $Y2=0
cc_429 N_A_465_315#_c_522_n N_CLK_M1006_g 0.00115367f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_430 N_A_465_315#_c_524_n N_CLK_c_750_n 0.0072683f $X=5.445 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_A_465_315#_c_522_n CLK 0.0181504f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_432 N_A_465_315#_c_523_n CLK 4.91988e-19 $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_433 N_A_465_315#_c_522_n N_CLK_c_752_n 0.0317882f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_434 N_A_465_315#_c_523_n N_CLK_c_752_n 0.006986f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_435 N_A_465_315#_c_530_n N_CLK_c_753_n 8.29701e-19 $X=5.165 $Y=2 $X2=0 $Y2=0
cc_436 N_A_465_315#_c_522_n N_CLK_c_753_n 0.00271044f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_437 N_A_465_315#_c_522_n N_CLK_c_754_n 0.00267286f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_438 N_A_465_315#_c_523_n N_CLK_c_754_n 0.00154383f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_439 N_A_465_315#_c_530_n N_CLK_c_763_n 0.0130686f $X=5.165 $Y=2 $X2=0 $Y2=0
cc_440 N_A_465_315#_c_522_n N_CLK_c_763_n 0.00820469f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_441 N_A_465_315#_c_522_n N_CLK_c_756_n 3.15312e-19 $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_442 N_A_465_315#_c_523_n N_CLK_c_756_n 0.0390204f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A_465_315#_c_522_n N_CLK_c_757_n 0.0236254f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_444 N_A_465_315#_c_523_n N_CLK_c_757_n 0.00214976f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_445 N_A_465_315#_c_524_n N_CLK_c_758_n 0.0390204f $X=5.445 $Y=0.995 $X2=0
+ $Y2=0
cc_446 N_A_465_315#_c_522_n N_A_1045_47#_c_865_n 0.00348926f $X=5.39 $Y=1.16
+ $X2=0 $Y2=0
cc_447 N_A_465_315#_c_524_n N_A_1045_47#_c_865_n 0.0112508f $X=5.445 $Y=0.995
+ $X2=0 $Y2=0
cc_448 N_A_465_315#_c_522_n N_A_1045_47#_c_854_n 0.0180201f $X=5.39 $Y=1.16
+ $X2=0 $Y2=0
cc_449 N_A_465_315#_c_523_n N_A_1045_47#_c_854_n 0.00131961f $X=5.39 $Y=1.16
+ $X2=0 $Y2=0
cc_450 N_A_465_315#_c_528_n N_VPWR_M1023_d 0.00488989f $X=3.185 $Y=1.77 $X2=0
+ $Y2=0
cc_451 N_A_465_315#_c_530_n N_VPWR_M1012_d 0.00607953f $X=5.165 $Y=2 $X2=0 $Y2=0
cc_452 N_A_465_315#_c_530_n N_VPWR_M1013_s 0.00332048f $X=5.165 $Y=2 $X2=0 $Y2=0
cc_453 N_A_465_315#_c_522_n N_VPWR_M1013_s 0.00226383f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_454 N_A_465_315#_c_541_n N_VPWR_c_988_n 0.0163044f $X=3.32 $Y=2.205 $X2=0
+ $Y2=0
cc_455 N_A_465_315#_c_530_n N_VPWR_c_988_n 0.111679f $X=5.165 $Y=2 $X2=0 $Y2=0
cc_456 N_A_465_315#_c_541_n N_VPWR_c_989_n 0.0133789f $X=3.32 $Y=2.205 $X2=0
+ $Y2=0
cc_457 N_A_465_315#_c_530_n N_VPWR_c_989_n 0.00252001f $X=5.165 $Y=2 $X2=0 $Y2=0
cc_458 N_A_465_315#_c_530_n N_VPWR_c_990_n 0.0243297f $X=5.165 $Y=2 $X2=0 $Y2=0
cc_459 N_A_465_315#_M1013_g N_VPWR_c_991_n 0.0046653f $X=5.56 $Y=1.985 $X2=0
+ $Y2=0
cc_460 N_A_465_315#_M1023_g N_VPWR_c_994_n 7.6274e-19 $X=2.43 $Y=2.275 $X2=0
+ $Y2=0
cc_461 N_A_465_315#_M1023_g N_VPWR_c_995_n 0.0247949f $X=2.43 $Y=2.275 $X2=0
+ $Y2=0
cc_462 N_A_465_315#_c_533_n N_VPWR_c_995_n 0.0022365f $X=2.46 $Y=1.74 $X2=0
+ $Y2=0
cc_463 N_A_465_315#_c_553_n N_VPWR_c_995_n 0.044273f $X=2.545 $Y=1.74 $X2=0
+ $Y2=0
cc_464 N_A_465_315#_M1013_g N_VPWR_c_996_n 0.00835513f $X=5.56 $Y=1.985 $X2=0
+ $Y2=0
cc_465 N_A_465_315#_M1000_d N_VPWR_c_981_n 0.00223109f $X=3.185 $Y=1.485 $X2=0
+ $Y2=0
cc_466 N_A_465_315#_M1023_g N_VPWR_c_981_n 0.002381f $X=2.43 $Y=2.275 $X2=0
+ $Y2=0
cc_467 N_A_465_315#_M1013_g N_VPWR_c_981_n 0.00794739f $X=5.56 $Y=1.985 $X2=0
+ $Y2=0
cc_468 N_A_465_315#_c_528_n N_VPWR_c_981_n 0.00508158f $X=3.185 $Y=1.77 $X2=0
+ $Y2=0
cc_469 N_A_465_315#_c_541_n N_VPWR_c_981_n 0.00839556f $X=3.32 $Y=2.205 $X2=0
+ $Y2=0
cc_470 N_A_465_315#_c_530_n N_VPWR_c_981_n 0.0146489f $X=5.165 $Y=2 $X2=0 $Y2=0
cc_471 N_A_465_315#_c_533_n N_VPWR_c_981_n 6.86139e-19 $X=2.46 $Y=1.74 $X2=0
+ $Y2=0
cc_472 N_A_465_315#_c_553_n N_VPWR_c_981_n 0.00214472f $X=2.545 $Y=1.74 $X2=0
+ $Y2=0
cc_473 N_A_465_315#_M1016_g N_VGND_c_1228_n 0.00849127f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_474 N_A_465_315#_c_521_n N_VGND_c_1228_n 0.0156967f $X=3.32 $Y=0.42 $X2=0
+ $Y2=0
cc_475 N_A_465_315#_M1016_g N_VGND_c_1234_n 0.00486707f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_476 N_A_465_315#_c_521_n N_VGND_c_1235_n 0.0133789f $X=3.32 $Y=0.42 $X2=0
+ $Y2=0
cc_477 N_A_465_315#_c_524_n N_VGND_c_1241_n 0.00337001f $X=5.445 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_465_315#_c_524_n N_VGND_c_1242_n 0.00980361f $X=5.445 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_A_465_315#_M1008_d N_VGND_c_1244_n 0.00204319f $X=3.185 $Y=0.235 $X2=0
+ $Y2=0
cc_480 N_A_465_315#_M1016_g N_VGND_c_1244_n 0.00673447f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_481 N_A_465_315#_c_521_n N_VGND_c_1244_n 0.00399922f $X=3.32 $Y=0.42 $X2=0
+ $Y2=0
cc_482 N_A_465_315#_c_524_n N_VGND_c_1244_n 0.00531009f $X=5.445 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_287_413#_M1000_g N_VPWR_c_988_n 0.00237274f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_484 N_A_287_413#_M1000_g N_VPWR_c_989_n 0.00468308f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_A_287_413#_c_664_n N_VPWR_c_994_n 0.0463617f $X=2.035 $Y=2.295 $X2=0
+ $Y2=0
cc_486 N_A_287_413#_M1000_g N_VPWR_c_995_n 0.00517884f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_487 N_A_287_413#_c_664_n N_VPWR_c_995_n 0.0295853f $X=2.035 $Y=2.295 $X2=0
+ $Y2=0
cc_488 N_A_287_413#_c_655_n N_VPWR_c_995_n 0.00379592f $X=2.12 $Y=2.125 $X2=0
+ $Y2=0
cc_489 N_A_287_413#_M1026_d N_VPWR_c_981_n 0.00263412f $X=1.435 $Y=2.065 $X2=0
+ $Y2=0
cc_490 N_A_287_413#_M1000_g N_VPWR_c_981_n 0.00805978f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_491 N_A_287_413#_c_664_n N_VPWR_c_981_n 0.0285676f $X=2.035 $Y=2.295 $X2=0
+ $Y2=0
cc_492 N_A_287_413#_c_660_n N_A_27_47#_c_1126_n 0.0219377f $X=2.33 $Y=0.395
+ $X2=0 $Y2=0
cc_493 N_A_287_413#_c_664_n A_383_413# 0.00832946f $X=2.035 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_494 N_A_287_413#_c_655_n A_383_413# 0.00151526f $X=2.12 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_495 N_A_287_413#_c_649_n N_VGND_c_1228_n 0.00734556f $X=3.11 $Y=0.995 $X2=0
+ $Y2=0
cc_496 N_A_287_413#_c_660_n N_VGND_c_1228_n 0.0231479f $X=2.33 $Y=0.395 $X2=0
+ $Y2=0
cc_497 N_A_287_413#_c_650_n N_VGND_c_1228_n 0.0210362f $X=2.415 $Y=0.995 $X2=0
+ $Y2=0
cc_498 N_A_287_413#_c_652_n N_VGND_c_1228_n 0.022345f $X=2.93 $Y=1.16 $X2=0
+ $Y2=0
cc_499 N_A_287_413#_c_653_n N_VGND_c_1228_n 0.00484825f $X=3.11 $Y=1.16 $X2=0
+ $Y2=0
cc_500 N_A_287_413#_c_660_n N_VGND_c_1234_n 0.0673769f $X=2.33 $Y=0.395 $X2=0
+ $Y2=0
cc_501 N_A_287_413#_c_649_n N_VGND_c_1235_n 0.00585385f $X=3.11 $Y=0.995 $X2=0
+ $Y2=0
cc_502 N_A_287_413#_M1007_d N_VGND_c_1244_n 0.00299551f $X=1.45 $Y=0.235 $X2=0
+ $Y2=0
cc_503 N_A_287_413#_c_649_n N_VGND_c_1244_n 0.00794139f $X=3.11 $Y=0.995 $X2=0
+ $Y2=0
cc_504 N_A_287_413#_c_660_n N_VGND_c_1244_n 0.0299006f $X=2.33 $Y=0.395 $X2=0
+ $Y2=0
cc_505 N_A_287_413#_c_660_n A_395_47# 0.00874765f $X=2.33 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_506 N_A_287_413#_c_650_n A_395_47# 0.00160798f $X=2.415 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_507 N_CLK_c_756_n N_A_1045_47#_M1003_g 0.0149447f $X=5.98 $Y=1.16 $X2=0 $Y2=0
cc_508 N_CLK_c_757_n N_A_1045_47#_M1003_g 3.03588e-19 $X=5.98 $Y=1.16 $X2=0
+ $Y2=0
cc_509 N_CLK_c_758_n N_A_1045_47#_M1003_g 0.021131f $X=5.98 $Y=0.995 $X2=0 $Y2=0
cc_510 N_CLK_M1006_g N_A_1045_47#_M1001_g 0.0355284f $X=5.98 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_CLK_c_752_n N_A_1045_47#_c_865_n 0.00480193f $X=5.65 $Y=1.19 $X2=0
+ $Y2=0
cc_512 N_CLK_c_754_n N_A_1045_47#_c_865_n 0.00300199f $X=5.795 $Y=1.19 $X2=0
+ $Y2=0
cc_513 N_CLK_c_756_n N_A_1045_47#_c_865_n 0.00341374f $X=5.98 $Y=1.16 $X2=0
+ $Y2=0
cc_514 N_CLK_c_757_n N_A_1045_47#_c_865_n 0.0192296f $X=5.98 $Y=1.16 $X2=0 $Y2=0
cc_515 N_CLK_c_758_n N_A_1045_47#_c_865_n 0.0106654f $X=5.98 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_CLK_c_756_n N_A_1045_47#_c_853_n 3.98986e-19 $X=5.98 $Y=1.16 $X2=0
+ $Y2=0
cc_517 N_CLK_c_757_n N_A_1045_47#_c_853_n 0.00436902f $X=5.98 $Y=1.16 $X2=0
+ $Y2=0
cc_518 N_CLK_c_758_n N_A_1045_47#_c_853_n 0.00414454f $X=5.98 $Y=0.995 $X2=0
+ $Y2=0
cc_519 N_CLK_M1006_g N_A_1045_47#_c_861_n 0.0035261f $X=5.98 $Y=1.985 $X2=0
+ $Y2=0
cc_520 N_CLK_c_757_n N_A_1045_47#_c_861_n 6.35092e-19 $X=5.98 $Y=1.16 $X2=0
+ $Y2=0
cc_521 N_CLK_c_749_n N_A_1045_47#_c_854_n 3.56754e-19 $X=4.67 $Y=0.73 $X2=0
+ $Y2=0
cc_522 N_CLK_c_750_n N_A_1045_47#_c_854_n 7.25091e-19 $X=4.67 $Y=0.88 $X2=0
+ $Y2=0
cc_523 N_CLK_c_752_n N_A_1045_47#_c_854_n 0.00824021f $X=5.65 $Y=1.19 $X2=0
+ $Y2=0
cc_524 N_CLK_M1006_g N_A_1045_47#_c_886_n 0.0253822f $X=5.98 $Y=1.985 $X2=0
+ $Y2=0
cc_525 N_CLK_c_754_n N_A_1045_47#_c_886_n 0.00202388f $X=5.795 $Y=1.19 $X2=0
+ $Y2=0
cc_526 N_CLK_c_756_n N_A_1045_47#_c_886_n 0.00274158f $X=5.98 $Y=1.16 $X2=0
+ $Y2=0
cc_527 N_CLK_c_757_n N_A_1045_47#_c_886_n 0.0263899f $X=5.98 $Y=1.16 $X2=0 $Y2=0
cc_528 N_CLK_c_754_n N_A_1045_47#_c_855_n 0.00140401f $X=5.795 $Y=1.19 $X2=0
+ $Y2=0
cc_529 N_CLK_c_756_n N_A_1045_47#_c_855_n 0.0018984f $X=5.98 $Y=1.16 $X2=0 $Y2=0
cc_530 N_CLK_c_757_n N_A_1045_47#_c_855_n 0.0201661f $X=5.98 $Y=1.16 $X2=0 $Y2=0
cc_531 N_CLK_M1006_g N_VPWR_c_984_n 0.00166155f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_532 N_CLK_c_763_n N_VPWR_c_990_n 0.0240974f $X=4.735 $Y=1.325 $X2=0 $Y2=0
cc_533 N_CLK_M1006_g N_VPWR_c_991_n 0.00424386f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_534 N_CLK_M1006_g N_VPWR_c_996_n 5.79077e-19 $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_535 N_CLK_M1006_g N_VPWR_c_981_n 0.00576356f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_536 N_CLK_c_749_n N_VGND_c_1229_n 0.00809304f $X=4.67 $Y=0.73 $X2=0 $Y2=0
cc_537 N_CLK_c_749_n N_VGND_c_1241_n 0.00337001f $X=4.67 $Y=0.73 $X2=0 $Y2=0
cc_538 N_CLK_c_750_n N_VGND_c_1241_n 0.00230382f $X=4.67 $Y=0.88 $X2=0 $Y2=0
cc_539 N_CLK_c_758_n N_VGND_c_1242_n 0.0143705f $X=5.98 $Y=0.995 $X2=0 $Y2=0
cc_540 N_CLK_c_749_n N_VGND_c_1244_n 0.0053254f $X=4.67 $Y=0.73 $X2=0 $Y2=0
cc_541 N_CLK_c_750_n N_VGND_c_1244_n 0.00262886f $X=4.67 $Y=0.88 $X2=0 $Y2=0
cc_542 N_A_1045_47#_c_861_n N_VPWR_M1006_d 3.59643e-19 $X=6.325 $Y=1.495 $X2=0
+ $Y2=0
cc_543 N_A_1045_47#_c_886_n N_VPWR_M1006_d 0.00807023f $X=6.325 $Y=1.79 $X2=0
+ $Y2=0
cc_544 N_A_1045_47#_M1001_g N_VPWR_c_984_n 0.00547058f $X=6.455 $Y=1.985 $X2=0
+ $Y2=0
cc_545 N_A_1045_47#_M1018_g N_VPWR_c_984_n 6.13033e-19 $X=6.875 $Y=1.985 $X2=0
+ $Y2=0
cc_546 N_A_1045_47#_c_886_n N_VPWR_c_984_n 0.0177826f $X=6.325 $Y=1.79 $X2=0
+ $Y2=0
cc_547 N_A_1045_47#_M1018_g N_VPWR_c_985_n 0.00144921f $X=6.875 $Y=1.985 $X2=0
+ $Y2=0
cc_548 N_A_1045_47#_M1021_g N_VPWR_c_985_n 0.0113975f $X=7.295 $Y=1.985 $X2=0
+ $Y2=0
cc_549 N_A_1045_47#_M1024_g N_VPWR_c_985_n 7.74424e-19 $X=7.715 $Y=1.985 $X2=0
+ $Y2=0
cc_550 N_A_1045_47#_M1024_g N_VPWR_c_987_n 0.00588578f $X=7.715 $Y=1.985 $X2=0
+ $Y2=0
cc_551 N_A_1045_47#_c_902_p N_VPWR_c_991_n 0.0109464f $X=5.77 $Y=2.085 $X2=0
+ $Y2=0
cc_552 N_A_1045_47#_c_886_n N_VPWR_c_991_n 0.00315285f $X=6.325 $Y=1.79 $X2=0
+ $Y2=0
cc_553 N_A_1045_47#_M1001_g N_VPWR_c_992_n 0.00538448f $X=6.455 $Y=1.985 $X2=0
+ $Y2=0
cc_554 N_A_1045_47#_M1018_g N_VPWR_c_992_n 0.00541359f $X=6.875 $Y=1.985 $X2=0
+ $Y2=0
cc_555 N_A_1045_47#_c_886_n N_VPWR_c_992_n 4.25885e-19 $X=6.325 $Y=1.79 $X2=0
+ $Y2=0
cc_556 N_A_1045_47#_M1021_g N_VPWR_c_993_n 0.0046653f $X=7.295 $Y=1.985 $X2=0
+ $Y2=0
cc_557 N_A_1045_47#_M1024_g N_VPWR_c_993_n 0.00465454f $X=7.715 $Y=1.985 $X2=0
+ $Y2=0
cc_558 N_A_1045_47#_M1013_d N_VPWR_c_981_n 0.00408188f $X=5.635 $Y=1.485 $X2=0
+ $Y2=0
cc_559 N_A_1045_47#_M1001_g N_VPWR_c_981_n 0.00864801f $X=6.455 $Y=1.985 $X2=0
+ $Y2=0
cc_560 N_A_1045_47#_M1018_g N_VPWR_c_981_n 0.00954042f $X=6.875 $Y=1.985 $X2=0
+ $Y2=0
cc_561 N_A_1045_47#_M1021_g N_VPWR_c_981_n 0.00796766f $X=7.295 $Y=1.985 $X2=0
+ $Y2=0
cc_562 N_A_1045_47#_M1024_g N_VPWR_c_981_n 0.00884761f $X=7.715 $Y=1.985 $X2=0
+ $Y2=0
cc_563 N_A_1045_47#_c_902_p N_VPWR_c_981_n 0.00637602f $X=5.77 $Y=2.085 $X2=0
+ $Y2=0
cc_564 N_A_1045_47#_c_886_n N_VPWR_c_981_n 0.00754065f $X=6.325 $Y=1.79 $X2=0
+ $Y2=0
cc_565 N_A_1045_47#_M1004_g N_GCLK_c_1162_n 0.00930832f $X=6.875 $Y=0.56 $X2=0
+ $Y2=0
cc_566 N_A_1045_47#_M1009_g N_GCLK_c_1162_n 0.00161345f $X=7.295 $Y=0.56 $X2=0
+ $Y2=0
cc_567 N_A_1045_47#_c_862_n N_GCLK_c_1162_n 0.00346944f $X=6.41 $Y=1.185 $X2=0
+ $Y2=0
cc_568 N_A_1045_47#_c_856_n N_GCLK_c_1162_n 2.61826e-19 $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_569 N_A_1045_47#_M1004_g N_GCLK_c_1153_n 0.00238446f $X=6.875 $Y=0.56 $X2=0
+ $Y2=0
cc_570 N_A_1045_47#_c_862_n N_GCLK_c_1153_n 0.0172592f $X=6.41 $Y=1.185 $X2=0
+ $Y2=0
cc_571 N_A_1045_47#_c_856_n N_GCLK_c_1153_n 0.00208088f $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_572 N_A_1045_47#_M1018_g N_GCLK_c_1169_n 0.011586f $X=6.875 $Y=1.985 $X2=0
+ $Y2=0
cc_573 N_A_1045_47#_M1021_g N_GCLK_c_1169_n 0.00161345f $X=7.295 $Y=1.985 $X2=0
+ $Y2=0
cc_574 N_A_1045_47#_c_862_n N_GCLK_c_1169_n 0.00346944f $X=6.41 $Y=1.185 $X2=0
+ $Y2=0
cc_575 N_A_1045_47#_c_856_n N_GCLK_c_1169_n 2.45827e-19 $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_576 N_A_1045_47#_M1018_g N_GCLK_c_1157_n 0.00208253f $X=6.875 $Y=1.985 $X2=0
+ $Y2=0
cc_577 N_A_1045_47#_c_862_n N_GCLK_c_1157_n 0.0182275f $X=6.41 $Y=1.185 $X2=0
+ $Y2=0
cc_578 N_A_1045_47#_c_856_n N_GCLK_c_1157_n 6.77113e-19 $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_579 N_A_1045_47#_M1004_g N_GCLK_c_1154_n 0.00160474f $X=6.875 $Y=0.56 $X2=0
+ $Y2=0
cc_580 N_A_1045_47#_M1009_g N_GCLK_c_1154_n 0.00113977f $X=7.295 $Y=0.56 $X2=0
+ $Y2=0
cc_581 N_A_1045_47#_c_853_n N_GCLK_c_1154_n 0.0042649f $X=6.325 $Y=1.055 $X2=0
+ $Y2=0
cc_582 N_A_1045_47#_c_856_n N_GCLK_c_1154_n 0.00389977f $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_583 N_A_1045_47#_M1018_g N_GCLK_c_1158_n 0.0019548f $X=6.875 $Y=1.985 $X2=0
+ $Y2=0
cc_584 N_A_1045_47#_M1021_g N_GCLK_c_1158_n 0.00139033f $X=7.295 $Y=1.985 $X2=0
+ $Y2=0
cc_585 N_A_1045_47#_c_861_n N_GCLK_c_1158_n 0.00437861f $X=6.325 $Y=1.495 $X2=0
+ $Y2=0
cc_586 N_A_1045_47#_c_856_n N_GCLK_c_1158_n 0.00112702f $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_587 N_A_1045_47#_M1003_g GCLK 0.00301777f $X=6.455 $Y=0.56 $X2=0 $Y2=0
cc_588 N_A_1045_47#_M1004_g GCLK 0.00222143f $X=6.875 $Y=0.56 $X2=0 $Y2=0
cc_589 N_A_1045_47#_c_862_n GCLK 0.00132943f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_590 N_A_1045_47#_M1018_g GCLK 0.0110932f $X=6.875 $Y=1.985 $X2=0 $Y2=0
cc_591 N_A_1045_47#_M1021_g GCLK 4.73454e-19 $X=7.295 $Y=1.985 $X2=0 $Y2=0
cc_592 N_A_1045_47#_M1021_g GCLK 0.00696131f $X=7.295 $Y=1.985 $X2=0 $Y2=0
cc_593 N_A_1045_47#_M1024_g GCLK 5.88219e-19 $X=7.715 $Y=1.985 $X2=0 $Y2=0
cc_594 N_A_1045_47#_c_862_n GCLK 0.0217831f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_595 N_A_1045_47#_c_856_n GCLK 0.0311619f $X=7.715 $Y=1.16 $X2=0 $Y2=0
cc_596 N_A_1045_47#_M1021_g GCLK 0.00235666f $X=7.295 $Y=1.985 $X2=0 $Y2=0
cc_597 N_A_1045_47#_M1024_g GCLK 0.0267063f $X=7.715 $Y=1.985 $X2=0 $Y2=0
cc_598 N_A_1045_47#_c_856_n GCLK 0.00128432f $X=7.715 $Y=1.16 $X2=0 $Y2=0
cc_599 N_A_1045_47#_M1024_g GCLK 0.00371048f $X=7.715 $Y=1.985 $X2=0 $Y2=0
cc_600 N_A_1045_47#_c_856_n GCLK 0.00990909f $X=7.715 $Y=1.16 $X2=0 $Y2=0
cc_601 N_A_1045_47#_M1004_g GCLK 0.00559017f $X=6.875 $Y=0.56 $X2=0 $Y2=0
cc_602 N_A_1045_47#_M1009_g GCLK 4.51994e-19 $X=7.295 $Y=0.56 $X2=0 $Y2=0
cc_603 N_A_1045_47#_M1009_g N_GCLK_c_1156_n 0.00220005f $X=7.295 $Y=0.56 $X2=0
+ $Y2=0
cc_604 N_A_1045_47#_M1015_g N_GCLK_c_1156_n 0.0198692f $X=7.715 $Y=0.56 $X2=0
+ $Y2=0
cc_605 N_A_1045_47#_c_856_n N_GCLK_c_1156_n 0.00557847f $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_606 N_A_1045_47#_c_865_n N_VGND_M1019_d 0.00847186f $X=6.24 $Y=0.7 $X2=0
+ $Y2=0
cc_607 N_A_1045_47#_c_853_n N_VGND_M1019_d 0.00121461f $X=6.325 $Y=1.055 $X2=0
+ $Y2=0
cc_608 N_A_1045_47#_M1004_g N_VGND_c_1230_n 0.00151249f $X=6.875 $Y=0.56 $X2=0
+ $Y2=0
cc_609 N_A_1045_47#_M1009_g N_VGND_c_1230_n 0.00774463f $X=7.295 $Y=0.56 $X2=0
+ $Y2=0
cc_610 N_A_1045_47#_M1015_g N_VGND_c_1230_n 4.92355e-19 $X=7.715 $Y=0.56 $X2=0
+ $Y2=0
cc_611 N_A_1045_47#_c_856_n N_VGND_c_1230_n 3.5066e-19 $X=7.715 $Y=1.16 $X2=0
+ $Y2=0
cc_612 N_A_1045_47#_M1015_g N_VGND_c_1232_n 0.00487324f $X=7.715 $Y=0.56 $X2=0
+ $Y2=0
cc_613 N_A_1045_47#_M1003_g N_VGND_c_1236_n 0.00508675f $X=6.455 $Y=0.56 $X2=0
+ $Y2=0
cc_614 N_A_1045_47#_M1004_g N_VGND_c_1236_n 0.00422241f $X=6.875 $Y=0.56 $X2=0
+ $Y2=0
cc_615 N_A_1045_47#_c_865_n N_VGND_c_1236_n 0.00107125f $X=6.24 $Y=0.7 $X2=0
+ $Y2=0
cc_616 N_A_1045_47#_M1009_g N_VGND_c_1237_n 0.0046653f $X=7.295 $Y=0.56 $X2=0
+ $Y2=0
cc_617 N_A_1045_47#_M1015_g N_VGND_c_1237_n 0.00465454f $X=7.715 $Y=0.56 $X2=0
+ $Y2=0
cc_618 N_A_1045_47#_c_865_n N_VGND_c_1241_n 0.00255672f $X=6.24 $Y=0.7 $X2=0
+ $Y2=0
cc_619 N_A_1045_47#_c_854_n N_VGND_c_1241_n 0.0289373f $X=5.35 $Y=0.46 $X2=0
+ $Y2=0
cc_620 N_A_1045_47#_M1003_g N_VGND_c_1242_n 0.00299722f $X=6.455 $Y=0.56 $X2=0
+ $Y2=0
cc_621 N_A_1045_47#_c_865_n N_VGND_c_1242_n 0.0409497f $X=6.24 $Y=0.7 $X2=0
+ $Y2=0
cc_622 N_A_1045_47#_M1017_s N_VGND_c_1244_n 0.00226128f $X=5.225 $Y=0.235 $X2=0
+ $Y2=0
cc_623 N_A_1045_47#_M1003_g N_VGND_c_1244_n 0.00887252f $X=6.455 $Y=0.56 $X2=0
+ $Y2=0
cc_624 N_A_1045_47#_M1004_g N_VGND_c_1244_n 0.00569656f $X=6.875 $Y=0.56 $X2=0
+ $Y2=0
cc_625 N_A_1045_47#_M1009_g N_VGND_c_1244_n 0.00789179f $X=7.295 $Y=0.56 $X2=0
+ $Y2=0
cc_626 N_A_1045_47#_M1015_g N_VGND_c_1244_n 0.00880873f $X=7.715 $Y=0.56 $X2=0
+ $Y2=0
cc_627 N_A_1045_47#_c_865_n N_VGND_c_1244_n 0.00988208f $X=6.24 $Y=0.7 $X2=0
+ $Y2=0
cc_628 N_A_1045_47#_c_854_n N_VGND_c_1244_n 0.0159946f $X=5.35 $Y=0.46 $X2=0
+ $Y2=0
cc_629 N_A_1045_47#_c_865_n A_1127_47# 0.00202671f $X=6.24 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_630 N_VPWR_c_981_n A_109_369# 0.00168634f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_631 N_VPWR_c_981_n N_A_27_47#_M1005_d 0.00386882f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_632 N_VPWR_c_983_n N_A_27_47#_c_1102_n 0.0101554f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_633 N_VPWR_c_994_n N_A_27_47#_c_1113_n 0.0098369f $X=2.375 $Y=2.44 $X2=0
+ $Y2=0
cc_634 N_VPWR_c_981_n N_A_27_47#_c_1113_n 0.00639994f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_635 N_VPWR_c_994_n N_A_27_47#_c_1121_n 0.033302f $X=2.375 $Y=2.44 $X2=0 $Y2=0
cc_636 N_VPWR_c_981_n N_A_27_47#_c_1121_n 0.0209902f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_637 N_VPWR_c_981_n A_383_413# 0.00809303f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_638 N_VPWR_c_981_n N_GCLK_M1001_d 0.00393857f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_639 N_VPWR_c_981_n N_GCLK_M1021_d 0.00393857f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_640 N_VPWR_M1018_s N_GCLK_c_1169_n 0.00267387f $X=6.95 $Y=1.485 $X2=0 $Y2=0
cc_641 N_VPWR_c_985_n N_GCLK_c_1169_n 0.0131569f $X=7.085 $Y=2 $X2=0 $Y2=0
cc_642 N_VPWR_c_992_n GCLK 0.0151826f $X=7 $Y=2.72 $X2=0 $Y2=0
cc_643 N_VPWR_c_981_n GCLK 0.00941829f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_644 N_VPWR_c_985_n GCLK 9.45716e-19 $X=7.085 $Y=2 $X2=0 $Y2=0
cc_645 N_VPWR_c_987_n GCLK 0.0750802f $X=7.975 $Y=1.66 $X2=0 $Y2=0
cc_646 N_VPWR_c_993_n GCLK 0.0185916f $X=7.89 $Y=2.72 $X2=0 $Y2=0
cc_647 N_VPWR_c_981_n GCLK 0.0111152f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_648 N_VPWR_c_987_n GCLK 0.0259847f $X=7.975 $Y=1.66 $X2=0 $Y2=0
cc_649 A_109_369# N_A_27_47#_c_1102_n 0.00276145f $X=0.545 $Y=1.845 $X2=0 $Y2=0
cc_650 A_109_369# N_A_27_47#_c_1113_n 8.01918e-19 $X=0.545 $Y=1.845 $X2=0 $Y2=0
cc_651 A_109_369# N_A_27_47#_c_1121_n 6.12987e-19 $X=0.545 $Y=1.845 $X2=0 $Y2=0
cc_652 N_A_27_47#_c_1103_n N_VGND_M1027_d 7.33468e-19 $X=1.015 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_653 N_A_27_47#_c_1104_n N_VGND_M1027_d 8.45526e-19 $X=0.685 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_654 N_A_27_47#_c_1104_n N_VGND_c_1227_n 0.0158273f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_655 N_A_27_47#_c_1101_n N_VGND_c_1233_n 0.0172026f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_656 N_A_27_47#_c_1104_n N_VGND_c_1233_n 0.00258611f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_657 N_A_27_47#_c_1103_n N_VGND_c_1234_n 0.00256355f $X=1.015 $Y=0.7 $X2=0
+ $Y2=0
cc_658 N_A_27_47#_c_1126_n N_VGND_c_1234_n 0.0120906f $X=1.1 $Y=0.42 $X2=0 $Y2=0
cc_659 N_A_27_47#_M1027_s N_VGND_c_1244_n 0.00226128f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_660 N_A_27_47#_M1011_d N_VGND_c_1244_n 0.00617083f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_661 N_A_27_47#_c_1101_n N_VGND_c_1244_n 0.00977915f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_662 N_A_27_47#_c_1103_n N_VGND_c_1244_n 0.00427891f $X=1.015 $Y=0.7 $X2=0
+ $Y2=0
cc_663 N_A_27_47#_c_1104_n N_VGND_c_1244_n 0.00582244f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_664 N_A_27_47#_c_1126_n N_VGND_c_1244_n 0.00681108f $X=1.1 $Y=0.42 $X2=0
+ $Y2=0
cc_665 N_GCLK_c_1162_n N_VGND_M1004_d 0.0025724f $X=7.05 $Y=0.8 $X2=0 $Y2=0
cc_666 N_GCLK_c_1162_n N_VGND_c_1230_n 0.0126141f $X=7.05 $Y=0.8 $X2=0 $Y2=0
cc_667 GCLK N_VGND_c_1230_n 9.17352e-19 $X=7.55 $Y=1.105 $X2=0 $Y2=0
cc_668 GCLK N_VGND_c_1232_n 0.0259847f $X=8.01 $Y=1.105 $X2=0 $Y2=0
cc_669 N_GCLK_c_1156_n N_VGND_c_1232_n 0.0482658f $X=7.505 $Y=0.42 $X2=0 $Y2=0
cc_670 N_GCLK_c_1162_n N_VGND_c_1236_n 0.0020257f $X=7.05 $Y=0.8 $X2=0 $Y2=0
cc_671 GCLK N_VGND_c_1236_n 0.0186706f $X=6.63 $Y=0.425 $X2=0 $Y2=0
cc_672 N_GCLK_c_1156_n N_VGND_c_1237_n 0.0185589f $X=7.505 $Y=0.42 $X2=0 $Y2=0
cc_673 N_GCLK_M1003_s N_VGND_c_1244_n 0.00215201f $X=6.53 $Y=0.235 $X2=0 $Y2=0
cc_674 N_GCLK_M1009_s N_VGND_c_1244_n 0.0038878f $X=7.37 $Y=0.235 $X2=0 $Y2=0
cc_675 N_GCLK_c_1162_n N_VGND_c_1244_n 0.00476969f $X=7.05 $Y=0.8 $X2=0 $Y2=0
cc_676 GCLK N_VGND_c_1244_n 0.012115f $X=6.63 $Y=0.425 $X2=0 $Y2=0
cc_677 N_GCLK_c_1156_n N_VGND_c_1244_n 0.0110428f $X=7.505 $Y=0.42 $X2=0 $Y2=0
cc_678 N_VGND_c_1244_n A_395_47# 0.00299863f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_679 N_VGND_c_1242_n A_1127_47# 0.00105937f $X=6.33 $Y=0.18 $X2=-0.19
+ $Y2=-0.24

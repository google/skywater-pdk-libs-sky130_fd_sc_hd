* File: sky130_fd_sc_hd__sdlclkp_1.spice.pex
* Created: Thu Aug 27 14:47:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%SCE 3 7 9 10 17
r29 14 17 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.16
+ $X2=0.212 $Y2=1.53
r31 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r32 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r33 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.165
r34 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r35 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%GATE 3 7 9 10 14
c41 14 0 9.54602e-20 $X=0.935 $Y=1.16
c42 10 0 2.81292e-20 $X=1.15 $Y=1.87
r43 14 17 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.912 $Y=1.16
+ $X2=0.912 $Y2=1.325
r44 14 16 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.912 $Y=1.16
+ $X2=0.912 $Y2=0.995
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.935
+ $Y=1.16 $X2=0.935 $Y2=1.16
r46 9 10 12.0581 $w=3.44e-07 $l=3.4e-07 $layer=LI1_cond $X=1.042 $Y=1.53
+ $X2=1.042 $Y2=1.87
r47 9 15 13.1221 $w=3.44e-07 $l=3.7e-07 $layer=LI1_cond $X=1.042 $Y=1.53
+ $X2=1.042 $Y2=1.16
r48 7 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=0.995
r49 3 17 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.83 $Y=2.165
+ $X2=0.83 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%A_256_147# 1 2 9 13 17 21 24 25 28 30 33
+ 35 37 41 44 53 54 57 60 68 74
c171 68 0 1.23968e-19 $X=1.775 $Y=1.74
c172 60 0 1.37414e-19 $X=4.38 $Y=1.53
c173 57 0 3.38573e-20 $X=1.61 $Y=1.53
c174 44 0 1.86451e-19 $X=4.085 $Y=1.19
c175 41 0 2.00302e-19 $X=1.61 $Y=1.325
c176 24 0 3.18278e-20 $X=1.445 $Y=0.87
c177 9 0 2.35132e-20 $X=1.37 $Y=0.415
r178 68 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.74
+ $X2=1.775 $Y2=1.905
r179 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.775
+ $Y=1.74 $X2=1.775 $Y2=1.74
r180 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.38 $Y=1.53
+ $X2=4.38 $Y2=1.53
r181 57 69 5.52036 $w=4.53e-07 $l=2.1e-07 $layer=LI1_cond $X=1.632 $Y=1.53
+ $X2=1.632 $Y2=1.74
r182 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.53
+ $X2=1.61 $Y2=1.53
r183 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.53
+ $X2=1.61 $Y2=1.53
r184 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.235 $Y=1.53
+ $X2=4.38 $Y2=1.53
r185 53 54 3.0693 $w=1.4e-07 $l=2.48e-06 $layer=MET1_cond $X=4.235 $Y=1.53
+ $X2=1.755 $Y2=1.53
r186 44 74 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.085 $Y=1.19
+ $X2=4.085 $Y2=1.325
r187 44 73 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.085 $Y=1.19
+ $X2=4.085 $Y2=1.055
r188 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.085
+ $Y=1.19 $X2=4.085 $Y2=1.19
r189 41 57 5.38892 $w=4.53e-07 $l=2.05e-07 $layer=LI1_cond $X=1.632 $Y=1.325
+ $X2=1.632 $Y2=1.53
r190 40 41 3.94479 $w=4.53e-07 $l=1.2e-07 $layer=LI1_cond $X=1.61 $Y=1.205
+ $X2=1.61 $Y2=1.325
r191 35 37 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=4.705 $Y=0.615
+ $X2=4.705 $Y2=0.465
r192 31 61 3.79964 $w=2.5e-07 $l=1.53e-07 $layer=LI1_cond $X=4.465 $Y=1.62
+ $X2=4.312 $Y2=1.62
r193 31 33 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=4.465 $Y=1.62
+ $X2=4.795 $Y2=1.62
r194 29 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.32 $Y=0.7
+ $X2=4.705 $Y2=0.7
r195 29 30 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=4.32 $Y=0.785
+ $X2=4.32 $Y2=1.105
r196 28 61 3.10428 $w=3.05e-07 $l=1.25e-07 $layer=LI1_cond $X=4.312 $Y=1.495
+ $X2=4.312 $Y2=1.62
r197 27 30 0.521925 $w=1.68e-07 $l=8e-09 $layer=LI1_cond $X=4.312 $Y=1.19
+ $X2=4.32 $Y2=1.19
r198 27 43 14.8096 $w=1.68e-07 $l=2.27e-07 $layer=LI1_cond $X=4.312 $Y=1.19
+ $X2=4.085 $Y2=1.19
r199 27 28 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=4.312 $Y=1.275
+ $X2=4.312 $Y2=1.495
r200 25 63 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.445 $Y=0.87
+ $X2=1.37 $Y2=0.87
r201 24 40 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=1.53 $Y=0.87
+ $X2=1.53 $Y2=1.205
r202 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=0.87 $X2=1.445 $Y2=0.87
r203 21 74 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.035 $Y=1.835
+ $X2=4.035 $Y2=1.325
r204 17 73 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.035 $Y=0.445
+ $X2=4.035 $Y2=1.055
r205 13 71 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.835 $Y=2.275
+ $X2=1.835 $Y2=1.905
r206 7 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.37 $Y=0.735
+ $X2=1.37 $Y2=0.87
r207 7 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.37 $Y=0.735
+ $X2=1.37 $Y2=0.415
r208 2 33 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.66
+ $Y=1.515 $X2=4.795 $Y2=1.66
r209 1 37 182 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.235 $X2=4.665 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%A_256_243# 1 2 9 11 12 15 17 20 23 27 29
+ 30 36 37 40 41 42
c115 41 0 1.47482e-19 $X=1.955 $Y=0.87
c116 37 0 1.34642e-19 $X=3.92 $Y=0.85
c117 36 0 5.98268e-21 $X=3.92 $Y=0.85
c118 27 0 1.20845e-19 $X=3.825 $Y=1.66
c119 17 0 2.81292e-20 $X=1.895 $Y=1.215
c120 12 0 2.67301e-20 $X=1.43 $Y=1.29
c121 9 0 3.17216e-20 $X=1.355 $Y=2.275
r122 40 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=0.87
+ $X2=1.955 $Y2=1.035
r123 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=0.87
+ $X2=1.955 $Y2=0.705
r124 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=0.87 $X2=1.955 $Y2=0.87
r125 37 49 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.792 $Y=0.85
+ $X2=3.792 $Y2=0.935
r126 37 48 2.91128 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.792 $Y=0.85
+ $X2=3.792 $Y2=0.765
r127 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.92 $Y=0.85
+ $X2=3.92 $Y2=0.85
r128 32 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0.85
+ $X2=2.07 $Y2=0.85
r129 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.215 $Y=0.85
+ $X2=2.07 $Y2=0.85
r130 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.775 $Y=0.85
+ $X2=3.92 $Y2=0.85
r131 29 30 1.93069 $w=1.4e-07 $l=1.56e-06 $layer=MET1_cond $X=3.775 $Y=0.85
+ $X2=2.215 $Y2=0.85
r132 24 27 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.665 $Y=1.66
+ $X2=3.825 $Y2=1.66
r133 23 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=1.575
+ $X2=3.665 $Y2=1.66
r134 23 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.665 $Y=1.575
+ $X2=3.665 $Y2=0.935
r135 20 48 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.745 $Y=0.465
+ $X2=3.745 $Y2=0.765
r136 17 43 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.895 $Y=1.215
+ $X2=1.895 $Y2=1.035
r137 15 42 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.895 $Y=0.415
+ $X2=1.895 $Y2=0.705
r138 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.82 $Y=1.29
+ $X2=1.895 $Y2=1.215
r139 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.82 $Y=1.29
+ $X2=1.43 $Y2=1.29
r140 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.355 $Y=1.365
+ $X2=1.43 $Y2=1.29
r141 7 9 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.355 $Y=1.365
+ $X2=1.355 $Y2=2.275
r142 2 27 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=1.515 $X2=3.825 $Y2=1.66
r143 1 20 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=3.7
+ $Y=0.235 $X2=3.825 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%A_464_315# 1 2 9 13 17 21 23 27 31 33 36
+ 39 41 42 46 55
c132 46 0 1.8014e-19 $X=5.445 $Y=1.52
c133 39 0 1.77265e-19 $X=2.455 $Y=1.74
c134 36 0 1.82269e-19 $X=5.295 $Y=1.915
c135 13 0 1.38699e-19 $X=2.505 $Y=0.445
r136 47 55 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.445 $Y=1.52
+ $X2=5.535 $Y2=1.52
r137 47 52 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=5.445 $Y=1.52
+ $X2=5.395 $Y2=1.52
r138 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.445
+ $Y=1.52 $X2=5.445 $Y2=1.52
r139 39 51 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=1.74
+ $X2=2.455 $Y2=1.905
r140 39 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=1.74
+ $X2=2.455 $Y2=1.575
r141 38 41 3.38343 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=1.74
+ $X2=2.54 $Y2=1.74
r142 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.455
+ $Y=1.74 $X2=2.455 $Y2=1.74
r143 35 46 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.295 $Y=1.52
+ $X2=5.445 $Y2=1.52
r144 35 36 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=5.295 $Y=1.605
+ $X2=5.295 $Y2=1.915
r145 34 42 3.05 $w=1.7e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.4 $Y=2 $X2=3.29
+ $Y2=1.86
r146 33 36 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.14 $Y=2
+ $X2=5.295 $Y2=1.915
r147 33 34 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=5.14 $Y=2 $X2=3.4
+ $Y2=2
r148 29 42 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.29 $Y=2.085 $X2=3.29
+ $Y2=1.86
r149 29 31 11.2625 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=3.29 $Y=2.085
+ $X2=3.29 $Y2=2.3
r150 25 42 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.29 $Y=1.635 $X2=3.29
+ $Y2=1.86
r151 25 27 63.6463 $w=2.18e-07 $l=1.215e-06 $layer=LI1_cond $X=3.29 $Y=1.635
+ $X2=3.29 $Y2=0.42
r152 23 42 3.05 $w=2.7e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.18 $Y=1.77
+ $X2=3.29 $Y2=1.86
r153 23 41 27.3172 $w=2.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.18 $Y=1.77
+ $X2=2.54 $Y2=1.77
r154 19 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.535 $Y=1.655
+ $X2=5.535 $Y2=1.52
r155 19 21 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.535 $Y=1.655
+ $X2=5.535 $Y2=2.165
r156 15 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.395 $Y=1.385
+ $X2=5.395 $Y2=1.52
r157 15 17 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=5.395 $Y=1.385
+ $X2=5.395 $Y2=0.445
r158 13 50 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=2.505 $Y=0.445
+ $X2=2.505 $Y2=1.575
r159 9 51 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.425 $Y=2.275
+ $X2=2.425 $Y2=1.905
r160 2 31 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.485 $X2=3.315 $Y2=2.3
r161 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.235 $X2=3.305 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%A_286_413# 1 2 7 9 12 14 18 23 25 26 28 36
c100 28 0 1.77265e-19 $X=2.925 $Y=1.16
c101 26 0 3.17216e-20 $X=2.495 $Y=1.185
c102 25 0 3.18278e-20 $X=2.41 $Y=0.995
c103 14 0 2.67301e-20 $X=2.325 $Y=0.395
r104 35 36 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=3.095 $Y=1.16
+ $X2=3.105 $Y2=1.16
r105 31 32 14.6301 $w=2.46e-07 $l=2.95e-07 $layer=LI1_cond $X=2.115 $Y=1.205
+ $X2=2.41 $Y2=1.205
r106 29 35 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.925 $Y=1.16
+ $X2=3.095 $Y2=1.16
r107 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.925
+ $Y=1.16 $X2=2.925 $Y2=1.16
r108 26 32 4.2431 $w=3.8e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.495 $Y=1.185
+ $X2=2.41 $Y2=1.205
r109 26 28 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.495 $Y=1.185
+ $X2=2.925 $Y2=1.185
r110 25 32 2.90119 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.41 $Y=0.995
+ $X2=2.41 $Y2=1.205
r111 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.41 $Y=0.535
+ $X2=2.41 $Y2=0.995
r112 22 31 2.90119 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.115 $Y=1.375
+ $X2=2.115 $Y2=1.205
r113 22 23 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.115 $Y=1.375
+ $X2=2.115 $Y2=2.125
r114 18 23 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.03 $Y=2.295
+ $X2=2.115 $Y2=2.125
r115 18 20 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=2.03 $Y=2.295
+ $X2=1.595 $Y2=2.295
r116 14 24 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.325 $Y=0.395
+ $X2=2.41 $Y2=0.535
r117 14 16 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=2.325 $Y=0.395
+ $X2=1.63 $Y2=0.395
r118 10 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.325
+ $X2=3.105 $Y2=1.16
r119 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.105 $Y=1.325
+ $X2=3.105 $Y2=1.985
r120 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=0.995
+ $X2=3.095 $Y2=1.16
r121 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.095 $Y=0.995
+ $X2=3.095 $Y2=0.56
r122 2 20 600 $w=1.7e-07 $l=3.22102e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=2.065 $X2=1.595 $Y2=2.315
r123 1 16 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.63 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%CLK 3 5 8 11 15 17 18 21 22 24 27 29 36
c74 36 0 1.86451e-19 $X=4.93 $Y=1.14
c75 29 0 1.20845e-19 $X=4.72 $Y=1.325
c76 21 0 3.68683e-20 $X=5.845 $Y=1.05
c77 18 0 1.40624e-19 $X=4.655 $Y=0.88
c78 15 0 2.24995e-19 $X=5.955 $Y=2.165
r79 27 29 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.72 $Y=1.16
+ $X2=4.72 $Y2=1.325
r80 24 36 4.54172 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.795 $Y=1.14
+ $X2=4.93 $Y2=1.14
r81 24 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.795
+ $Y=1.16 $X2=4.795 $Y2=1.16
r82 22 32 41.4854 $w=3.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.855 $Y=1.05
+ $X2=5.855 $Y2=1.185
r83 22 31 41.4854 $w=3.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.855 $Y=1.05
+ $X2=5.855 $Y2=0.915
r84 21 36 34.0157 $w=3.08e-07 $l=9.15e-07 $layer=LI1_cond $X=5.845 $Y=1.11
+ $X2=4.93 $Y2=1.11
r85 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.845
+ $Y=1.05 $X2=5.845 $Y2=1.05
r86 17 18 44.1654 $w=4.2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.655 $Y=0.73
+ $X2=4.655 $Y2=0.88
r87 15 32 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=5.955 $Y=2.165
+ $X2=5.955 $Y2=1.185
r88 11 31 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.955 $Y=0.445 $X2=5.955
+ $Y2=0.915
r89 8 29 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.585 $Y=1.835
+ $X2=4.585 $Y2=1.325
r90 5 27 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=4.72 $Y=1.115
+ $X2=4.72 $Y2=1.16
r91 5 18 31.1181 $w=4.2e-07 $l=2.35e-07 $layer=POLY_cond $X=4.72 $Y=1.115
+ $X2=4.72 $Y2=0.88
r92 3 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.455 $Y=0.445
+ $X2=4.455 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%A_1012_47# 1 2 9 12 16 18 19 20 24 27 29
c58 29 0 3.68683e-20 $X=6.375 $Y=0.995
r59 27 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.375 $Y=1.16
+ $X2=6.375 $Y2=1.325
r60 27 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.375 $Y=1.16
+ $X2=6.375 $Y2=0.995
r61 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.375
+ $Y=1.16 $X2=6.375 $Y2=1.16
r62 24 26 9.57218 $w=4.78e-07 $l=2.09105e-07 $layer=LI1_cond $X=6.275 $Y=0.995
+ $X2=6.375 $Y2=1.16
r63 23 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.275 $Y=0.785
+ $X2=6.275 $Y2=0.995
r64 20 26 28.9697 $w=4.78e-07 $l=1.19932e-06 $layer=LI1_cond $X=5.745 $Y=2.085
+ $X2=6.375 $Y2=1.16
r65 20 22 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=5.745 $Y=2.085
+ $X2=5.745 $Y2=2.125
r66 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.19 $Y=0.7
+ $X2=6.275 $Y2=0.785
r67 18 19 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=6.19 $Y=0.7 $X2=5.27
+ $Y2=0.7
r68 14 19 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.14 $Y=0.615
+ $X2=5.27 $Y2=0.7
r69 14 16 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=5.14 $Y=0.615
+ $X2=5.14 $Y2=0.46
r70 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.985
+ $X2=6.43 $Y2=1.325
r71 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=0.56 $X2=6.43
+ $Y2=0.995
r72 2 22 600 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_PDIFF $count=1 $X=5.61
+ $Y=1.845 $X2=5.745 $Y2=2.125
r73 1 16 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.06
+ $Y=0.235 $X2=5.185 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%VPWR 1 2 3 4 5 16 18 22 24 26 27 41 47 54
+ 55 63 66 72 74
r90 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r91 71 72 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=2.53
+ $X2=5.49 $Y2=2.53
r92 68 71 0.761141 $w=5.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.29 $Y=2.53
+ $X2=5.325 $Y2=2.53
r93 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r94 65 66 11.8978 $w=7.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.79 $Y=2.44
+ $X2=3.01 $Y2=2.44
r95 61 65 4.26001 $w=7.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.79 $Y2=2.44
r96 61 63 10.9147 $w=7.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.37 $Y2=2.44
r97 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r98 55 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r99 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r100 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.195 $Y2=2.72
r101 52 54 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.36 $Y=2.72
+ $X2=6.67 $Y2=2.72
r102 51 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r103 51 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r104 50 72 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=5.49 $Y2=2.72
r105 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 47 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.03 $Y=2.72
+ $X2=6.195 $Y2=2.72
r107 47 50 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.03 $Y=2.72
+ $X2=5.75 $Y2=2.72
r108 44 69 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r109 43 46 8.69875 $w=5.48e-07 $l=4e-07 $layer=LI1_cond $X=3.91 $Y=2.53 $X2=4.31
+ $Y2=2.53
r110 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r111 41 68 1.63102 $w=5.48e-07 $l=7.5e-08 $layer=LI1_cond $X=5.215 $Y=2.53
+ $X2=5.29 $Y2=2.53
r112 41 46 19.6809 $w=5.48e-07 $l=9.05e-07 $layer=LI1_cond $X=5.215 $Y=2.53
+ $X2=4.31 $Y2=2.53
r113 40 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r114 40 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r115 39 66 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.01 $Y2=2.72
r116 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r117 36 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r118 35 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.07 $Y=2.72 $X2=2.37
+ $Y2=2.72
r119 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r120 33 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r121 32 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r122 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 30 58 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r124 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 27 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r126 27 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r127 26 39 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.58 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 24 43 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=3.855 $Y=2.53
+ $X2=3.91 $Y2=2.53
r129 24 26 12.2241 $w=5.48e-07 $l=2.75e-07 $layer=LI1_cond $X=3.855 $Y=2.53
+ $X2=3.58 $Y2=2.53
r130 20 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=2.635
+ $X2=6.195 $Y2=2.72
r131 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.195 $Y=2.635
+ $X2=6.195 $Y2=2.36
r132 16 58 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r133 16 18 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2
r134 5 22 600 $w=1.7e-07 $l=5.91777e-07 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=1.845 $X2=6.195 $Y2=2.36
r135 4 71 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.845 $X2=5.325 $Y2=2.34
r136 3 46 600 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=4.11
+ $Y=1.515 $X2=4.31 $Y2=2.34
r137 2 65 600 $w=1.7e-07 $l=4.15421e-07 $layer=licon1_PDIFF $count=1 $X=2.5
+ $Y=2.065 $X2=2.79 $Y2=2.36
r138 1 18 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%A_27_47# 1 2 3 12 17 18 19 20 22 26 31 32
r53 31 32 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.61 $Y=1.46
+ $X2=0.61 $Y2=1.755
r54 24 26 12.3584 $w=1.73e-07 $l=1.95e-07 $layer=LI1_cond $X=1.102 $Y=0.615
+ $X2=1.102 $Y2=0.42
r55 20 22 12.8802 $w=3.38e-07 $l=3.8e-07 $layer=LI1_cond $X=0.71 $Y=2.295
+ $X2=1.09 $Y2=2.295
r56 19 30 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.7
+ $X2=0.595 $Y2=0.7
r57 18 24 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.015 $Y=0.7
+ $X2=1.102 $Y2=0.615
r58 18 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.015 $Y=0.7
+ $X2=0.68 $Y2=0.7
r59 17 20 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.625 $Y=2.125
+ $X2=0.71 $Y2=2.295
r60 17 32 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.625 $Y=2.125
+ $X2=0.625 $Y2=1.755
r61 14 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0.785
+ $X2=0.595 $Y2=0.7
r62 14 31 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.595 $Y=0.785
+ $X2=0.595 $Y2=1.46
r63 10 30 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.215 $Y=0.7
+ $X2=0.595 $Y2=0.7
r64 10 12 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.43
r65 3 22 600 $w=1.7e-07 $l=5.29481e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.845 $X2=1.09 $Y2=2.29
r66 2 26 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.42
r67 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%GCLK 1 2 10 11 12 13 14 15 20
r17 14 15 15.9725 $w=2.83e-07 $l=3.95e-07 $layer=LI1_cond $X=6.672 $Y=1.815
+ $X2=6.672 $Y2=2.21
r18 13 20 3.63929 $w=2.83e-07 $l=9e-08 $layer=LI1_cond $X=6.672 $Y=0.51
+ $X2=6.672 $Y2=0.42
r19 11 14 7.19771 $w=2.83e-07 $l=1.78e-07 $layer=LI1_cond $X=6.672 $Y=1.637
+ $X2=6.672 $Y2=1.815
r20 11 12 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=6.672 $Y=1.637
+ $X2=6.672 $Y2=1.495
r21 10 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.73 $Y=0.825
+ $X2=6.73 $Y2=1.495
r22 9 13 6.99553 $w=2.83e-07 $l=1.73e-07 $layer=LI1_cond $X=6.672 $Y=0.683
+ $X2=6.672 $Y2=0.51
r23 9 10 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=6.672 $Y=0.683
+ $X2=6.672 $Y2=0.825
r24 2 14 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=6.505
+ $Y=1.485 $X2=6.64 $Y2=1.815
r25 1 20 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.505
+ $Y=0.235 $X2=6.64 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_1%VGND 1 2 3 4 15 19 23 25 27 32 40 52 53 56
+ 59 62 66 70
r104 68 70 9.36586 $w=5.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.21 $Y=0.18
+ $X2=6.36 $Y2=0.18
r105 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r106 65 68 1.01554 $w=5.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.165 $Y=0.18
+ $X2=6.21 $Y2=0.18
r107 65 66 20.8753 $w=5.28e-07 $l=6.6e-07 $layer=LI1_cond $X=6.165 $Y=0.18
+ $X2=5.505 $Y2=0.18
r108 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r109 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r110 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r111 53 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r112 52 70 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.36
+ $Y2=0
r113 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r114 49 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r115 49 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r116 48 66 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.505 $Y2=0
r117 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r118 46 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.245
+ $Y2=0
r119 46 48 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=5.29
+ $Y2=0
r120 44 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r121 44 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r122 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r123 41 59 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.837
+ $Y2=0
r124 41 43 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=3.91
+ $Y2=0
r125 40 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=4.245
+ $Y2=0
r126 40 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.91
+ $Y2=0
r127 39 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r128 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r129 36 39 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.53 $Y2=0
r130 36 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r131 35 38 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r132 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r133 33 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r134 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r135 32 59 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.665 $Y=0
+ $X2=2.837 $Y2=0
r136 32 38 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.665 $Y=0
+ $X2=2.53 $Y2=0
r137 27 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r138 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r139 25 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r140 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r141 21 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.085
+ $X2=4.245 $Y2=0
r142 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.245 $Y=0.085
+ $X2=4.245 $Y2=0.36
r143 17 59 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.837 $Y=0.085
+ $X2=2.837 $Y2=0
r144 17 19 14.1968 $w=3.43e-07 $l=4.25e-07 $layer=LI1_cond $X=2.837 $Y=0.085
+ $X2=2.837 $Y2=0.51
r145 13 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r146 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r147 4 65 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.03
+ $Y=0.235 $X2=6.165 $Y2=0.36
r148 3 23 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.11
+ $Y=0.235 $X2=4.245 $Y2=0.36
r149 2 19 182 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.235 $X2=2.81 $Y2=0.51
r150 1 15 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


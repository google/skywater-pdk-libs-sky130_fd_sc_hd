* File: sky130_fd_sc_hd__ha_2.pex.spice
* Created: Tue Sep  1 19:09:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__HA_2%A_79_21# 1 2 7 9 12 14 16 19 21 24 27 29 30 32
+ 37 39
c75 24 0 1.68161e-19 $X=1.115 $Y=1.16
r76 40 42 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.93 $Y2=1.16
r77 34 37 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.505 $Y=0.51
+ $X2=1.66 $Y2=0.51
r78 30 32 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.59 $Y=2.29
+ $X2=2.055 $Y2=2.29
r79 29 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=2.205
+ $X2=1.59 $Y2=2.29
r80 28 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=1.245
+ $X2=1.505 $Y2=1.16
r81 28 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.505 $Y=1.245
+ $X2=1.505 $Y2=2.205
r82 27 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=1.075
+ $X2=1.505 $Y2=1.16
r83 26 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=0.675
+ $X2=1.505 $Y2=0.51
r84 26 27 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.505 $Y=0.675
+ $X2=1.505 $Y2=1.075
r85 24 42 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.115 $Y=1.16
+ $X2=0.93 $Y2=1.16
r86 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.16 $X2=1.115 $Y2=1.16
r87 21 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=1.16
+ $X2=1.505 $Y2=1.16
r88 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.42 $Y=1.16
+ $X2=1.115 $Y2=1.16
r89 17 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.16
r90 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.93 $Y=1.325
+ $X2=0.93 $Y2=1.985
r91 14 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=1.16
r92 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.93 $Y=0.995
+ $X2=0.93 $Y2=0.56
r93 10 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r94 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r95 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r96 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
r97 2 32 600 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.845 $X2=2.055 $Y2=2.29
r98 1 37 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.66 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%A_342_199# 1 2 9 13 15 17 20 22 24 27 31 32 34
+ 35 38 40 41 44 46 48 49 50 60
c135 60 0 2.26883e-19 $X=5.05 $Y=1.16
c136 41 0 9.45908e-20 $X=3.63 $Y=0.8
c137 31 0 1.68161e-19 $X=1.845 $Y=1.16
c138 9 0 7.39302e-20 $X=1.845 $Y=2.165
r139 59 60 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=4.59 $Y=1.16
+ $X2=5.05 $Y2=1.16
r140 54 59 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.535 $Y=1.16
+ $X2=4.59 $Y2=1.16
r141 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=1.16 $X2=4.535 $Y2=1.16
r142 51 53 17.3597 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=4.457 $Y=0.8
+ $X2=4.457 $Y2=1.16
r143 48 53 9.27442 $w=2.53e-07 $l=1.99825e-07 $layer=LI1_cond $X=4.38 $Y=1.325
+ $X2=4.457 $Y2=1.16
r144 48 49 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.38 $Y=1.325
+ $X2=4.38 $Y2=1.855
r145 47 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=1.94
+ $X2=3.895 $Y2=1.94
r146 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.295 $Y=1.94
+ $X2=4.38 $Y2=1.855
r147 46 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.295 $Y=1.94
+ $X2=3.98 $Y2=1.94
r148 42 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=2.025
+ $X2=3.895 $Y2=1.94
r149 42 44 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=2.025
+ $X2=3.895 $Y2=2.19
r150 40 51 3.06467 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=4.295 $Y=0.8
+ $X2=4.457 $Y2=0.8
r151 40 41 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.295 $Y=0.8
+ $X2=3.63 $Y2=0.8
r152 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=0.715
+ $X2=3.63 $Y2=0.8
r153 36 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.545 $Y=0.715
+ $X2=3.545 $Y2=0.51
r154 34 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=1.94
+ $X2=3.895 $Y2=1.94
r155 34 35 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=3.81 $Y=1.94
+ $X2=1.93 $Y2=1.94
r156 32 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.16
+ $X2=1.845 $Y2=0.995
r157 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.16 $X2=1.845 $Y2=1.16
r158 29 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.845 $Y=1.855
+ $X2=1.93 $Y2=1.94
r159 29 31 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.845 $Y=1.855
+ $X2=1.845 $Y2=1.16
r160 25 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.16
r161 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.985
r162 22 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=1.16
r163 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=0.56
r164 18 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.16
r165 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.985
r166 15 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=1.16
r167 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=0.56
r168 13 56 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.87 $Y=0.445
+ $X2=1.87 $Y2=0.995
r169 7 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.16
r170 7 9 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=2.165
r171 2 44 600 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=1 $X=3.75
+ $Y=1.845 $X2=3.895 $Y2=2.19
r172 1 38 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.235 $X2=3.545 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%B 3 7 10 11 13 14 16 19 21 22 27 33 34 36
c77 27 0 1.24844e-19 $X=2.395 $Y=1.26
c78 21 0 7.39302e-20 $X=2.53 $Y=1.19
c79 19 0 6.64161e-20 $X=3.755 $Y=0.81
c80 7 0 3.18576e-20 $X=2.29 $Y=0.445
r81 32 34 10.4783 $w=2.76e-07 $l=6e-08 $layer=POLY_cond $X=3.43 $Y=1.55 $X2=3.49
+ $Y2=1.55
r82 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.52 $X2=3.43 $Y2=1.52
r83 28 36 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=2.462 $Y=1.26
+ $X2=2.462 $Y2=1.395
r84 27 30 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.26
+ $X2=2.36 $Y2=1.425
r85 27 29 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.26
+ $X2=2.36 $Y2=1.095
r86 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=1.26 $X2=2.395 $Y2=1.26
r87 22 36 3.26477 $w=3.05e-07 $l=1.4e-07 $layer=LI1_cond $X=2.462 $Y=1.535
+ $X2=2.462 $Y2=1.395
r88 22 33 23.3594 $w=4.48e-07 $l=8.15e-07 $layer=LI1_cond $X=2.615 $Y=1.535
+ $X2=3.43 $Y2=1.535
r89 21 28 2.64495 $w=3.03e-07 $l=7e-08 $layer=LI1_cond $X=2.462 $Y=1.19
+ $X2=2.462 $Y2=1.26
r90 17 19 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.49 $Y=0.81
+ $X2=3.755 $Y2=0.81
r91 14 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.755 $Y=0.735
+ $X2=3.755 $Y2=0.81
r92 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.755 $Y=0.735
+ $X2=3.755 $Y2=0.445
r93 11 34 32.308 $w=2.76e-07 $l=2.72213e-07 $layer=POLY_cond $X=3.675 $Y=1.745
+ $X2=3.49 $Y2=1.55
r94 11 13 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.675 $Y=1.745
+ $X2=3.675 $Y2=2.165
r95 10 34 17.0164 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.49 $Y=1.355
+ $X2=3.49 $Y2=1.55
r96 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.885
+ $X2=3.49 $Y2=0.81
r97 9 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.49 $Y=0.885 $X2=3.49
+ $Y2=1.355
r98 7 29 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.29 $Y=0.445
+ $X2=2.29 $Y2=1.095
r99 3 30 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.265 $Y=2.165
+ $X2=2.265 $Y2=1.425
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%A 1 3 4 6 10 14 16 17 29 31
c74 31 0 2.08591e-19 $X=3.932 $Y=1.225
c75 16 0 2.4141e-19 $X=3.905 $Y=1.19
c76 10 0 7.86312e-20 $X=4.115 $Y=0.445
c77 4 0 2.70336e-20 $X=2.815 $Y=1.305
c78 1 0 9.45908e-20 $X=2.71 $Y=0.735
r79 26 29 38.8804 $w=2.7e-07 $l=1.75e-07 $layer=POLY_cond $X=3.94 $Y=1.23
+ $X2=4.115 $Y2=1.23
r80 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.14 $X2=2.955 $Y2=1.14
r81 16 31 3.0159 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.932 $Y=1.14
+ $X2=3.932 $Y2=1.225
r82 16 24 36.3315 $w=2.88e-07 $l=8.65e-07 $layer=LI1_cond $X=3.82 $Y=1.14
+ $X2=2.955 $Y2=1.14
r83 16 17 15.3659 $w=2.23e-07 $l=3e-07 $layer=LI1_cond $X=3.932 $Y=1.23
+ $X2=3.932 $Y2=1.53
r84 16 31 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=3.932 $Y=1.23
+ $X2=3.932 $Y2=1.225
r85 16 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.23 $X2=3.94 $Y2=1.23
r86 12 29 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.115 $Y=1.365
+ $X2=4.115 $Y2=1.23
r87 12 14 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.115 $Y=1.365
+ $X2=4.115 $Y2=2.165
r88 8 29 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.115 $Y=1.095
+ $X2=4.115 $Y2=1.23
r89 8 10 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.115 $Y=1.095
+ $X2=4.115 $Y2=0.445
r90 4 23 38.5416 $w=3.03e-07 $l=1.87029e-07 $layer=POLY_cond $X=2.815 $Y=1.305
+ $X2=2.862 $Y2=1.14
r91 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.815 $Y=1.305
+ $X2=2.815 $Y2=2.165
r92 1 23 76.7198 $w=3.03e-07 $l=4.74958e-07 $layer=POLY_cond $X=2.71 $Y=0.735
+ $X2=2.862 $Y2=1.14
r93 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.71 $Y=0.735 $X2=2.71
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%VPWR 1 2 3 4 5 16 18 24 30 32 34 38 40 53 58 67
+ 71 75 77 81
r80 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r81 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r82 73 75 10.6544 $w=5.98e-07 $l=1.9e-07 $layer=LI1_cond $X=3.45 $Y=2.505
+ $X2=3.64 $Y2=2.505
r83 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r84 70 73 0.697712 $w=5.98e-07 $l=3.5e-08 $layer=LI1_cond $X=3.415 $Y=2.505
+ $X2=3.45 $Y2=2.505
r85 70 71 18.1299 $w=5.98e-07 $l=5.65e-07 $layer=LI1_cond $X=3.415 $Y=2.505
+ $X2=2.85 $Y2=2.505
r86 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r88 62 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r89 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r90 59 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.38 $Y2=2.72
r91 59 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.83 $Y2=2.72
r92 58 80 3.90446 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=5.145 $Y=2.72
+ $X2=5.332 $Y2=2.72
r93 58 61 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.145 $Y=2.72
+ $X2=4.83 $Y2=2.72
r94 57 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r95 57 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r96 56 75 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.91 $Y=2.72 $X2=3.64
+ $Y2=2.72
r97 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 53 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=2.72
+ $X2=4.38 $Y2=2.72
r99 53 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.215 $Y=2.72
+ $X2=3.91 $Y2=2.72
r100 52 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r101 51 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.85 $Y2=2.72
r102 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r104 49 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r105 48 51 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r106 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 46 67 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.25 $Y=2.72
+ $X2=1.152 $Y2=2.72
r108 46 48 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 44 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r110 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 41 64 3.90232 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.187 $Y2=2.72
r112 41 43 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 40 67 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=1.152 $Y2=2.72
r114 40 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r116 38 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r117 34 37 32.6526 $w=2.38e-07 $l=6.8e-07 $layer=LI1_cond $X=5.265 $Y=1.66
+ $X2=5.265 $Y2=2.34
r118 32 80 3.17368 $w=2.4e-07 $l=1.13666e-07 $layer=LI1_cond $X=5.265 $Y=2.635
+ $X2=5.332 $Y2=2.72
r119 32 37 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=5.265 $Y=2.635
+ $X2=5.265 $Y2=2.34
r120 28 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=2.635
+ $X2=4.38 $Y2=2.72
r121 28 30 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.38 $Y=2.635
+ $X2=4.38 $Y2=2.29
r122 24 27 38.676 $w=1.93e-07 $l=6.8e-07 $layer=LI1_cond $X=1.152 $Y=1.68
+ $X2=1.152 $Y2=2.36
r123 22 67 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.152 $Y=2.635
+ $X2=1.152 $Y2=2.72
r124 22 27 15.641 $w=1.93e-07 $l=2.75e-07 $layer=LI1_cond $X=1.152 $Y=2.635
+ $X2=1.152 $Y2=2.36
r125 18 21 32.6526 $w=2.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=2.34
r126 16 64 3.17582 $w=2.4e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.187 $Y2=2.72
r127 16 21 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.255 $Y2=2.34
r128 5 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.125
+ $Y=1.485 $X2=5.26 $Y2=2.34
r129 5 34 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.125
+ $Y=1.485 $X2=5.26 $Y2=1.66
r130 4 30 600 $w=1.7e-07 $l=5.31578e-07 $layer=licon1_PDIFF $count=1 $X=4.19
+ $Y=1.845 $X2=4.38 $Y2=2.29
r131 3 70 300 $w=1.7e-07 $l=7.13618e-07 $layer=licon1_PDIFF $count=2 $X=2.89
+ $Y=1.845 $X2=3.415 $Y2=2.29
r132 2 27 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.485 $X2=1.14 $Y2=2.36
r133 2 24 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.485 $X2=1.14 $Y2=1.68
r134 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r135 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%SUM 1 2 7 8 9 10 11 12 23 30 36
r20 36 48 1.79269 $w=2.23e-07 $l=3.5e-08 $layer=LI1_cond $X=0.667 $Y=1.53
+ $X2=0.667 $Y2=1.565
r21 30 46 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=0.667 $Y=0.85
+ $X2=0.667 $Y2=0.825
r22 12 43 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=2.21 $X2=0.72
+ $Y2=2.33
r23 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.72 $Y=1.87
+ $X2=0.72 $Y2=2.21
r24 11 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.72 $Y=1.87
+ $X2=0.72 $Y2=1.73
r25 10 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.72 $Y=1.59
+ $X2=0.72 $Y2=1.73
r26 10 48 2.04739 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.72 $Y=1.59
+ $X2=0.72 $Y2=1.565
r27 10 36 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=0.667 $Y=1.505
+ $X2=0.667 $Y2=1.53
r28 9 10 16.1342 $w=2.23e-07 $l=3.15e-07 $layer=LI1_cond $X=0.667 $Y=1.19
+ $X2=0.667 $Y2=1.505
r29 8 46 2.22201 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=0.795 $X2=0.72
+ $Y2=0.825
r30 8 21 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=0.795
+ $X2=0.72 $Y2=0.66
r31 8 9 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=0.667 $Y=0.88
+ $X2=0.667 $Y2=1.19
r32 8 30 1.53659 $w=2.23e-07 $l=3e-08 $layer=LI1_cond $X=0.667 $Y=0.88 $X2=0.667
+ $Y2=0.85
r33 7 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.72 $Y=0.51 $X2=0.72
+ $Y2=0.66
r34 7 23 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=0.51 $X2=0.72
+ $Y2=0.4
r35 2 10 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.72 $Y2=1.65
r36 2 43 400 $w=1.7e-07 $l=9.28386e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.72 $Y2=2.33
r37 1 23 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.72 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%COUT 1 2 10 11 12 13 14 15 20 25
c20 10 0 7.86312e-20 $X=4.8 $Y=0.825
r21 14 15 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.84 $Y=1.87
+ $X2=4.84 $Y2=2.21
r22 14 25 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=4.84 $Y=1.87
+ $X2=4.84 $Y2=1.71
r23 13 20 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.8 $Y=0.51 $X2=4.8
+ $Y2=0.4
r24 11 25 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=4.84 $Y=1.67 $X2=4.84
+ $Y2=1.71
r25 11 12 6.81244 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.84 $Y=1.67
+ $X2=4.84 $Y2=1.545
r26 10 12 45.6312 $w=1.73e-07 $l=7.2e-07 $layer=LI1_cond $X=4.877 $Y=0.825
+ $X2=4.877 $Y2=1.545
r27 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.8 $Y=0.66 $X2=4.8
+ $Y2=0.51
r28 9 10 8.29065 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.8 $Y=0.66 $X2=4.8
+ $Y2=0.825
r29 2 25 300 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=2 $X=4.665
+ $Y=1.485 $X2=4.8 $Y2=1.71
r30 1 20 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.665
+ $Y=0.235 $X2=4.8 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%VGND 1 2 3 4 5 16 18 22 26 30 32 34 36 38 43 48
+ 56 65 68 71 75
c83 75 0 2.70336e-20 $X=5.29 $Y=0
r84 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r85 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r86 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r87 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r88 60 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r89 60 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r90 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r91 57 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.34
+ $Y2=0
r92 57 59 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.83
+ $Y2=0
r93 56 74 3.90446 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=5.332
+ $Y2=0
r94 56 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=4.83
+ $Y2=0
r95 55 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r96 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r97 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r98 52 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r99 51 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r100 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r101 49 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=0 $X2=2.5
+ $Y2=0
r102 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.665 $Y=0
+ $X2=2.99 $Y2=0
r103 48 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.34
+ $Y2=0
r104 48 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.215 $Y=0
+ $X2=3.91 $Y2=0
r105 47 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r106 47 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r107 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r108 44 65 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.152
+ $Y2=0
r109 44 46 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=2.07
+ $Y2=0
r110 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.5
+ $Y2=0
r111 43 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=0
+ $X2=2.07 $Y2=0
r112 42 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r113 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r114 39 62 3.90232 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r115 39 41 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.69 $Y2=0
r116 38 65 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.152
+ $Y2=0
r117 38 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.69 $Y2=0
r118 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 36 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 32 74 3.17368 $w=2.4e-07 $l=1.13666e-07 $layer=LI1_cond $X=5.265 $Y=0.085
+ $X2=5.332 $Y2=0
r121 32 34 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=5.265 $Y=0.085
+ $X2=5.265 $Y2=0.38
r122 28 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.085
+ $X2=4.34 $Y2=0
r123 28 30 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.34 $Y=0.085
+ $X2=4.34 $Y2=0.38
r124 24 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=0.085 $X2=2.5
+ $Y2=0
r125 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.5 $Y=0.085
+ $X2=2.5 $Y2=0.38
r126 20 65 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.152 $Y=0.085
+ $X2=1.152 $Y2=0
r127 20 22 16.7786 $w=1.93e-07 $l=2.95e-07 $layer=LI1_cond $X=1.152 $Y=0.085
+ $X2=1.152 $Y2=0.38
r128 16 62 3.17582 $w=2.4e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.187 $Y2=0
r129 16 18 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.38
r130 5 34 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.125
+ $Y=0.235 $X2=5.26 $Y2=0.38
r131 4 30 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=4.19
+ $Y=0.235 $X2=4.38 $Y2=0.38
r132 3 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.235 $X2=2.5 $Y2=0.38
r133 2 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.235 $X2=1.14 $Y2=0.38
r134 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__HA_2%A_389_47# 1 2 9 11 12 15
r28 13 15 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.92 $Y=0.635
+ $X2=2.92 $Y2=0.51
r29 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.835 $Y=0.72
+ $X2=2.92 $Y2=0.635
r30 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.835 $Y=0.72
+ $X2=2.165 $Y2=0.72
r31 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.08 $Y=0.635
+ $X2=2.165 $Y2=0.72
r32 7 9 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.08 $Y=0.635
+ $X2=2.08 $Y2=0.51
r33 2 15 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.235 $X2=2.92 $Y2=0.51
r34 1 9 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.235 $X2=2.08 $Y2=0.51
.ends


* File: sky130_fd_sc_hd__a21boi_1.spice
* Created: Tue Sep  1 18:51:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21boi_1.pex.spice"
.subckt sky130_fd_sc_hd__a21boi_1  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_B1_N_M1007_g N_A_27_413#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0799766 AS=0.1113 PD=0.777196 PS=1.37 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_27_413#_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.143 AS=0.123773 PD=1.09 PS=1.2028 NRD=14.76 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1003 A_384_47# N_A1_M1003_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.143 PD=0.93 PS=1.09 NRD=15.684 NRS=14.76 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_384_47# VNB NSHORT L=0.15 W=0.65 AD=0.17225
+ AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75001.5 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_B1_N_M1001_g N_A_27_413#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_300_297#_M1006_d N_A_27_413#_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_300_297#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_300_297#_M1000_d N_A2_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
c_55 VPB 0 1.83237e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a21boi_1.pxi.spice"
*
.ends
*
*

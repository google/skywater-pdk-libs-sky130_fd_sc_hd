* File: sky130_fd_sc_hd__a2111oi_2.spice
* Created: Tue Sep  1 18:50:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2111oi_2.pex.spice"
.subckt sky130_fd_sc_hd__a2111oi_2  VNB VPB C1 D1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* D1	D1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1014 N_Y_M1014_d N_C1_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.091 PD=1.87 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1014_s N_D1_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75004.2
+ A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_D1_M1017_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.091 PD=1.04 PS=0.93 NRD=10.152 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1018_d N_C1_M1018_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.12675 PD=0.975 PS=1.04 NRD=2.76 NRS=10.152 M=1 R=4.33333
+ SA=75001.6 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1018_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.105625 PD=1.04 PS=0.975 NRD=7.38 NRS=5.532 M=1 R=4.33333
+ SA=75002.1 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1003_d N_B1_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.091 PD=1.04 PS=0.93 NRD=12.912 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1012_s N_A1_M1000_g A_684_47# VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.17875 PD=0.93 PS=1.2 NRD=0 NRS=40.608 M=1 R=4.33333 SA=75003.1 SB=75001.8
+ A=0.0975 P=1.6 MULT=1
MM1019 A_684_47# N_A2_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65 AD=0.17875
+ AS=0.112125 PD=1.2 PS=0.995 NRD=40.608 NRS=5.532 M=1 R=4.33333 SA=75003.8
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 A_923_47# N_A2_M1004_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.112125 PD=0.93 PS=0.995 NRD=15.684 NRS=6.456 M=1 R=4.33333 SA=75004.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1015_d N_A1_M1015_g A_923_47# VNB NSHORT L=0.15 W=0.65 AD=0.17225
+ AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75004.7 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1001 N_A_28_297#_M1001_d N_C1_M1001_g A_115_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=16.7253 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1007 A_115_297# N_D1_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1002 A_287_297# N_D1_M1002_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75001.1 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1013 N_A_28_297#_M1013_d N_C1_M1013_g A_287_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.14 PD=1.32 PS=1.28 NRD=0 NRS=16.7253 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 N_A_28_297#_M1013_d N_B1_M1005_g N_A_467_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.16 AS=0.14 PD=1.32 PS=1.28 NRD=7.8603 NRS=0 M=1 R=6.66667 SA=75002
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_28_297#_M1010_d N_B1_M1010_g N_A_467_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_467_297#_M1006_d N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1006_s N_A2_M1008_g N_A_467_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_A2_M1016_g N_A_467_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.14 PD=1.32 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1011 N_A_467_297#_M1011_d N_A1_M1011_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=1
+ AD=0.335 AS=0.16 PD=2.67 PS=1.32 NRD=9.8303 NRS=3.9203 M=1 R=6.66667
+ SA=75001.5 SB=75000.3 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__a2111oi_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdfstp_4.pex.spice
* Created: Thu Aug 27 14:46:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%SCD 1 2 3 5 6 8 11 13 14
r33 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r34 14 19 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.53
+ $X2=0.212 $Y2=1.16
r35 13 19 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.212 $Y=0.85
+ $X2=0.212 $Y2=1.16
r36 9 11 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.315 $Y=1.695
+ $X2=0.47 $Y2=1.695
r37 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=1.695
r38 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.77 $X2=0.47
+ $Y2=2.165
r39 3 18 87.63 $w=2.63e-07 $l=4.97242e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.325 $Y2=1.16
r40 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r41 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.315 $Y=1.62
+ $X2=0.315 $Y2=1.695
r42 1 18 39.0634 $w=2.63e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.325 $Y2=1.16
r43 1 2 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.315 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%SCE 3 5 7 11 15 17 19 20 26 33 34
c108 26 0 1.07953e-19 $X=2.53 $Y=1.19
c109 7 0 1.86564e-19 $X=0.89 $Y=2.165
r110 33 36 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.557 $Y=1.16
+ $X2=2.557 $Y2=1.325
r111 33 35 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.557 $Y=1.16
+ $X2=2.557 $Y2=0.995
r112 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=1.16 $X2=2.535 $Y2=1.16
r113 26 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r114 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.19
+ $X2=0.69 $Y2=1.19
r115 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r116 19 20 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.835 $Y2=1.19
r117 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.735
+ $Y=1.25 $X2=0.735 $Y2=1.25
r118 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.19
+ $X2=0.69 $Y2=1.19
r119 15 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.64 $Y=0.445
+ $X2=2.64 $Y2=0.995
r120 11 36 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.61 $Y=2.165
+ $X2=2.61 $Y2=1.325
r121 5 30 38.6139 $w=3.32e-07 $l=2.12238e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.782 $Y2=1.25
r122 5 7 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.89 $Y=1.415
+ $X2=0.89 $Y2=2.165
r123 1 30 38.6139 $w=3.32e-07 $l=1.8747e-07 $layer=POLY_cond $X=0.83 $Y=1.085
+ $X2=0.782 $Y2=1.25
r124 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.83 $Y=1.085 $X2=0.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%D 1 3 6 8 9 13
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=0.93 $X2=1.25 $Y2=0.93
r42 9 14 24.262 $w=2.83e-07 $l=6e-07 $layer=LI1_cond $X=1.192 $Y=1.53 $X2=1.192
+ $Y2=0.93
r43 8 14 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=1.192 $Y=0.85 $X2=1.192
+ $Y2=0.93
r44 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.095
+ $X2=1.25 $Y2=0.93
r45 4 6 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.25 $Y=1.095 $X2=1.25
+ $Y2=2.165
r46 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=0.765
+ $X2=1.25 $Y2=0.93
r47 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.25 $Y=0.765 $X2=1.25
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_319_21# 1 2 9 13 16 20 21 22 24 34 36
c76 21 0 1.4475e-19 $X=1.95 $Y=1.16
r77 34 36 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=2.395 $Y=1.927
+ $X2=2.4 $Y2=1.927
r78 22 24 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=2.39 $Y=0.715
+ $X2=2.39 $Y2=0.44
r79 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.16 $X2=1.95 $Y2=1.16
r80 18 34 13.2805 $w=3.13e-07 $l=3.63e-07 $layer=LI1_cond $X=2.032 $Y=1.927
+ $X2=2.395 $Y2=1.927
r81 18 20 20.9848 $w=3.33e-07 $l=6.1e-07 $layer=LI1_cond $X=2.032 $Y=1.77
+ $X2=2.032 $Y2=1.16
r82 17 22 20.8976 $w=1.88e-07 $l=3.58e-07 $layer=LI1_cond $X=2.032 $Y=0.81
+ $X2=2.39 $Y2=0.81
r83 17 20 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.032 $Y=0.905
+ $X2=2.032 $Y2=1.16
r84 15 21 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.745 $Y=1.16
+ $X2=1.95 $Y2=1.16
r85 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.745 $Y=1.16
+ $X2=1.67 $Y2=1.16
r86 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.325
+ $X2=1.67 $Y2=1.16
r87 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.67 $Y=1.325
+ $X2=1.67 $Y2=2.165
r88 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=0.995
+ $X2=1.67 $Y2=1.16
r89 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.67 $Y=0.995 $X2=1.67
+ $Y2=0.445
r90 2 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.845 $X2=2.4 $Y2=1.99
r91 1 24 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.235 $X2=2.43 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%CLK 7 8 10 13 15 16 17 18 19 20 26 28
c73 20 0 1.05862e-19 $X=3.45 $Y=1.19
c74 15 0 7.67918e-20 $X=3.52 $Y=1.62
c75 13 0 1.07242e-19 $X=3.58 $Y=0.805
r76 41 42 0.14951 $w=5.58e-07 $l=7e-09 $layer=LI1_cond $X=2.995 $Y=1.335
+ $X2=3.002 $Y2=1.335
r77 34 41 7.51078 $w=1.8e-07 $l=2.8e-07 $layer=LI1_cond $X=2.995 $Y=1.615
+ $X2=2.995 $Y2=1.335
r78 30 42 7.01796 $w=1.95e-07 $l=2.8e-07 $layer=LI1_cond $X=3.002 $Y=1.055
+ $X2=3.002 $Y2=1.335
r79 26 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.42
r80 26 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.255
+ $X2=3.43 $Y2=1.09
r81 20 42 9.14146 $w=5.58e-07 $l=4.28e-07 $layer=LI1_cond $X=3.43 $Y=1.335
+ $X2=3.002 $Y2=1.335
r82 20 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.255 $X2=3.43 $Y2=1.255
r83 19 34 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.995 $Y=1.87
+ $X2=2.995 $Y2=1.615
r84 18 41 0.106793 $w=5.58e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=1.335
+ $X2=2.995 $Y2=1.335
r85 17 30 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.002 $Y=0.85
+ $X2=3.002 $Y2=1.055
r86 15 16 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.52 $Y=1.62
+ $X2=3.52 $Y2=1.77
r87 15 29 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.49 $Y=1.62 $X2=3.49
+ $Y2=1.42
r88 11 13 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.49 $Y=0.805 $X2=3.58
+ $Y2=0.805
r89 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.58 $Y=0.73 $X2=3.58
+ $Y2=0.805
r90 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.58 $Y=0.73 $X2=3.58
+ $Y2=0.445
r91 7 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.55 $Y=2.165
+ $X2=3.55 $Y2=1.77
r92 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=0.88 $X2=3.49
+ $Y2=0.805
r93 1 28 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.49 $Y=0.88 $X2=3.49
+ $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_643_369# 1 2 9 13 15 16 18 20 23 27 31 33
+ 36 40 42 43 44 45 47 49 50 54 55 56 57 60 61 63 64 65 66 67 76 80 83 84
c285 84 0 1.78722e-19 $X=5.33 $Y=1.74
c286 80 0 3.22574e-20 $X=3.917 $Y=1.09
c287 76 0 1.95341e-19 $X=7.645 $Y=1.87
c288 66 0 1.36329e-19 $X=7.5 $Y=1.87
c289 64 0 1.42859e-19 $X=5.145 $Y=1.87
c290 61 0 6.7173e-20 $X=8.94 $Y=1.09
c291 60 0 3.87856e-19 $X=8.94 $Y=1.09
c292 49 0 7.67918e-20 $X=3.91 $Y=1.255
r293 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=1.74 $X2=5.33 $Y2=1.74
r294 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.645 $Y=1.87
+ $X2=7.645 $Y2=1.87
r295 73 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r296 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=1.87
+ $X2=3.91 $Y2=1.87
r297 67 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r298 66 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.5 $Y=1.87
+ $X2=7.645 $Y2=1.87
r299 66 67 2.55569 $w=1.4e-07 $l=2.065e-06 $layer=MET1_cond $X=7.5 $Y=1.87
+ $X2=5.435 $Y2=1.87
r300 65 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=1.87
+ $X2=3.91 $Y2=1.87
r301 64 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r302 64 65 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=4.055 $Y2=1.87
r303 63 77 9.70478 $w=2.83e-07 $l=2.4e-07 $layer=LI1_cond $X=7.885 $Y=1.812
+ $X2=7.645 $Y2=1.812
r304 61 90 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.94 $Y=1.09
+ $X2=8.94 $Y2=0.925
r305 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.94
+ $Y=1.09 $X2=8.94 $Y2=1.09
r306 58 60 7.48077 $w=2.83e-07 $l=1.85e-07 $layer=LI1_cond $X=8.962 $Y=0.905
+ $X2=8.962 $Y2=1.09
r307 56 58 7.22568 $w=1.85e-07 $l=1.82675e-07 $layer=LI1_cond $X=8.82 $Y=0.812
+ $X2=8.962 $Y2=0.905
r308 56 57 41.0663 $w=1.83e-07 $l=6.85e-07 $layer=LI1_cond $X=8.82 $Y=0.812
+ $X2=8.135 $Y2=0.812
r309 55 88 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.97 $Y=1.16
+ $X2=7.97 $Y2=1.325
r310 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.16 $X2=7.97 $Y2=1.16
r311 52 63 6.85451 $w=2.85e-07 $l=1.94715e-07 $layer=LI1_cond $X=8.01 $Y=1.67
+ $X2=7.885 $Y2=1.812
r312 52 54 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=8.01 $Y=1.67
+ $X2=8.01 $Y2=1.16
r313 51 57 7.01633 $w=1.85e-07 $l=1.65076e-07 $layer=LI1_cond $X=8.01 $Y=0.905
+ $X2=8.135 $Y2=0.812
r314 51 54 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.01 $Y=0.905
+ $X2=8.01 $Y2=1.16
r315 50 81 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.917 $Y=1.255
+ $X2=3.917 $Y2=1.42
r316 50 80 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.917 $Y=1.255
+ $X2=3.917 $Y2=1.09
r317 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.91
+ $Y=1.255 $X2=3.91 $Y2=1.255
r318 47 70 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=1.83
+ $X2=3.865 $Y2=1.915
r319 47 49 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.865 $Y=1.83
+ $X2=3.865 $Y2=1.255
r320 46 49 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.865 $Y=0.885
+ $X2=3.865 $Y2=1.255
r321 44 46 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.865 $Y2=0.885
r322 44 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.735 $Y=0.8
+ $X2=3.455 $Y2=0.8
r323 42 70 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.735 $Y=1.915
+ $X2=3.865 $Y2=1.915
r324 42 43 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.735 $Y=1.915
+ $X2=3.425 $Y2=1.915
r325 38 45 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.362 $Y=0.715
+ $X2=3.455 $Y2=0.8
r326 38 40 16.4865 $w=1.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.362 $Y=0.715
+ $X2=3.362 $Y2=0.44
r327 34 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.34 $Y=2
+ $X2=3.425 $Y2=1.915
r328 34 36 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.34 $Y=2 $X2=3.34
+ $Y2=2.16
r329 31 90 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9 $Y=0.445 $X2=9
+ $Y2=0.925
r330 27 88 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.91 $Y=2.065
+ $X2=7.91 $Y2=1.325
r331 21 83 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.33 $Y=1.905
+ $X2=5.33 $Y2=1.74
r332 21 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.33 $Y=1.905
+ $X2=5.33 $Y2=2.275
r333 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.94 $Y=0.73
+ $X2=4.94 $Y2=0.445
r334 17 33 5.30422 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=4.075 $Y=0.805
+ $X2=3.992 $Y2=0.805
r335 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.94 $Y2=0.73
r336 16 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.075 $Y2=0.805
r337 13 33 20.4101 $w=1.5e-07 $l=7.88987e-08 $layer=POLY_cond $X=4 $Y=0.73
+ $X2=3.992 $Y2=0.805
r338 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4 $Y=0.73 $X2=4
+ $Y2=0.445
r339 11 33 20.4101 $w=1.5e-07 $l=7.84219e-08 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=3.992 $Y2=0.805
r340 11 80 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.985 $Y=0.88
+ $X2=3.985 $Y2=1.09
r341 9 81 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.97 $Y=2.165
+ $X2=3.97 $Y2=1.42
r342 2 36 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.845 $X2=3.34 $Y2=2.16
r343 1 40 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.37 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_809_369# 1 2 8 9 11 13 16 20 22 24 28 35
+ 36 39 42 43 46 49 50 57 66
c179 66 0 8.01298e-20 $X=4.327 $Y=1.09
c180 46 0 3.47594e-20 $X=4.37 $Y=1.19
c181 22 0 5.6211e-20 $X=8.54 $Y=1.905
c182 16 0 9.48056e-20 $X=5.36 $Y=0.445
c183 9 0 1.42859e-19 $X=5.285 $Y=1.165
c184 8 0 1.78722e-19 $X=4.615 $Y=1.84
r185 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.56
+ $Y=1.74 $X2=8.56 $Y2=1.74
r186 56 57 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.615 $Y=1.255
+ $X2=4.69 $Y2=1.255
r187 53 56 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.405 $Y=1.255
+ $X2=4.615 $Y2=1.255
r188 50 60 28.1708 $w=2.23e-07 $l=5.5e-07 $layer=LI1_cond $X=8.537 $Y=1.19
+ $X2=8.537 $Y2=1.74
r189 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.565 $Y=1.19
+ $X2=8.565 $Y2=1.19
r190 46 67 8.46186 $w=3.23e-07 $l=2.3e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.42
r191 46 66 6.15528 $w=3.23e-07 $l=1e-07 $layer=LI1_cond $X=4.327 $Y=1.19
+ $X2=4.327 $Y2=1.09
r192 46 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.255 $X2=4.405 $Y2=1.255
r193 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=1.19
+ $X2=4.37 $Y2=1.19
r194 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=1.19
+ $X2=4.37 $Y2=1.19
r195 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.42 $Y=1.19
+ $X2=8.565 $Y2=1.19
r196 42 43 4.83291 $w=1.4e-07 $l=3.905e-06 $layer=MET1_cond $X=8.42 $Y=1.19
+ $X2=4.515 $Y2=1.19
r197 41 66 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.25 $Y=0.585
+ $X2=4.25 $Y2=1.09
r198 39 41 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0.42
+ $X2=4.23 $Y2=0.585
r199 36 67 29.9635 $w=2.73e-07 $l=7.15e-07 $layer=LI1_cond $X=4.302 $Y=2.135
+ $X2=4.302 $Y2=1.42
r200 35 36 6.01906 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.267 $Y=2.3
+ $X2=4.267 $Y2=2.135
r201 26 28 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=4.615 $Y=1.915
+ $X2=4.91 $Y2=1.915
r202 22 59 38.5495 $w=3.2e-07 $l=1.81659e-07 $layer=POLY_cond $X=8.54 $Y=1.905
+ $X2=8.505 $Y2=1.74
r203 22 24 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.54 $Y=1.905
+ $X2=8.54 $Y2=2.275
r204 18 59 38.5495 $w=3.2e-07 $l=2.14942e-07 $layer=POLY_cond $X=8.39 $Y=1.575
+ $X2=8.505 $Y2=1.74
r205 18 20 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=8.39 $Y=1.575
+ $X2=8.39 $Y2=0.555
r206 14 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.36 $Y=1.09
+ $X2=5.36 $Y2=0.445
r207 11 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.91 $Y=1.99
+ $X2=4.91 $Y2=1.915
r208 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.91 $Y=1.99
+ $X2=4.91 $Y2=2.275
r209 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.285 $Y=1.165
+ $X2=5.36 $Y2=1.09
r210 9 57 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.285 $Y=1.165
+ $X2=4.69 $Y2=1.165
r211 8 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.615 $Y=1.84
+ $X2=4.615 $Y2=1.915
r212 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.615 $Y=1.42
+ $X2=4.615 $Y2=1.255
r213 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.615 $Y=1.42
+ $X2=4.615 $Y2=1.84
r214 2 35 600 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.845 $X2=4.18 $Y2=2.3
r215 1 39 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.235 $X2=4.21 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_1129_21# 1 2 9 15 19 20 22 24 25 28 32 34
+ 38 44
c96 34 0 4.32543e-20 $X=5.81 $Y=0.72
c97 22 0 4.56917e-20 $X=6.285 $Y=0.72
c98 20 0 5.68782e-20 $X=6.01 $Y=1.74
r99 42 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.84 $Y=1.065
+ $X2=5.84 $Y2=1.575
r100 38 42 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=1.065
r101 38 41 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.81 $Y=0.93
+ $X2=5.81 $Y2=0.795
r102 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.81
+ $Y=0.93 $X2=5.81 $Y2=0.93
r103 34 37 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.81 $Y=0.72
+ $X2=5.81 $Y2=0.93
r104 30 32 9.64836 $w=2.13e-07 $l=1.8e-07 $layer=LI1_cond $X=6.712 $Y=2.105
+ $X2=6.712 $Y2=2.285
r105 26 28 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=0.635
+ $X2=6.41 $Y2=0.51
r106 24 30 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.712 $Y2=2.105
r107 24 25 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.095 $Y2=2.02
r108 23 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=0.72
+ $X2=5.81 $Y2=0.72
r109 22 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.285 $Y=0.72
+ $X2=6.41 $Y2=0.635
r110 22 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.285 $Y=0.72
+ $X2=5.975 $Y2=0.72
r111 20 45 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.74
+ $X2=5.955 $Y2=1.905
r112 20 44 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.74
+ $X2=5.955 $Y2=1.575
r113 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.01
+ $Y=1.74 $X2=6.01 $Y2=1.74
r114 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.01 $Y=1.935
+ $X2=6.095 $Y2=2.02
r115 17 19 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.01 $Y=1.935
+ $X2=6.01 $Y2=1.74
r116 15 45 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.84 $Y=2.275
+ $X2=5.84 $Y2=1.905
r117 9 41 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.72 $Y=0.445
+ $X2=5.72 $Y2=0.795
r118 2 32 600 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_PDIFF $count=1 $X=6.555
+ $Y=2.065 $X2=6.715 $Y2=2.285
r119 1 28 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.325
+ $Y=0.235 $X2=6.45 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_997_413# 1 2 11 13 15 18 21 25 29 31 36
+ 38 39 45 46 47 50 52 55
c145 52 0 4.32543e-20 $X=6.39 $Y=1.095
r146 50 56 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.465 $Y=1.16
+ $X2=7.465 $Y2=1.325
r147 50 55 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.465 $Y=1.16
+ $X2=7.465 $Y2=0.995
r148 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.44
+ $Y=1.16 $X2=7.44 $Y2=1.16
r149 45 53 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.39 $Y=1.23
+ $X2=6.39 $Y2=1.365
r150 45 52 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.39 $Y=1.23
+ $X2=6.39 $Y2=1.095
r151 44 47 3.29018 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.475 $Y2=1.185
r152 44 46 6.54147 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.185
+ $X2=6.305 $Y2=1.185
r153 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.39
+ $Y=1.23 $X2=6.39 $Y2=1.23
r154 39 49 3.24611 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.355 $Y=1.125
+ $X2=7.44 $Y2=1.125
r155 39 47 33.805 $w=2.98e-07 $l=8.8e-07 $layer=LI1_cond $X=7.355 $Y=1.125
+ $X2=6.475 $Y2=1.125
r156 38 42 6.20468 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=1.31
+ $X2=5.67 $Y2=1.31
r157 38 46 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.755 $Y=1.31
+ $X2=6.305 $Y2=1.31
r158 35 42 0.18542 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=1.395
+ $X2=5.67 $Y2=1.31
r159 35 36 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.67 $Y=1.395
+ $X2=5.67 $Y2=2.135
r160 31 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.585 $Y=2.3
+ $X2=5.67 $Y2=2.135
r161 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.585 $Y=2.3
+ $X2=5.12 $Y2=2.3
r162 27 42 35.1923 $w=1.56e-07 $l=4.5e-07 $layer=LI1_cond $X=5.22 $Y=1.31
+ $X2=5.67 $Y2=1.31
r163 27 29 21.0845 $w=4.38e-07 $l=8.05e-07 $layer=LI1_cond $X=5.22 $Y=1.225
+ $X2=5.22 $Y2=0.42
r164 23 25 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.48 $Y=0.805
+ $X2=6.66 $Y2=0.805
r165 21 56 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.55 $Y=2.065
+ $X2=7.55 $Y2=1.325
r166 18 55 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.495 $Y=0.555
+ $X2=7.495 $Y2=0.995
r167 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.66 $Y=0.73
+ $X2=6.66 $Y2=0.805
r168 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.66 $Y=0.73
+ $X2=6.66 $Y2=0.445
r169 11 53 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=6.48 $Y=2.275
+ $X2=6.48 $Y2=1.365
r170 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.48 $Y=0.88
+ $X2=6.48 $Y2=0.805
r171 7 52 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.48 $Y=0.88
+ $X2=6.48 $Y2=1.095
r172 2 33 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=2.065 $X2=5.12 $Y2=2.3
r173 1 29 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%SET_B 5 9 13 16 19 22 23 27 28 30 32 33 39
+ 40 44 45 46
c136 45 0 4.11784e-20 $X=6.9 $Y=1.68
c137 22 0 2.22391e-19 $X=9.715 $Y=1.985
c138 9 0 4.56917e-20 $X=7.02 $Y=0.445
c139 5 0 1.54163e-19 $X=6.97 $Y=2.275
r140 44 47 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=1.845
r141 44 46 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=1.515
r142 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.9
+ $Y=1.68 $X2=6.9 $Y2=1.68
r143 40 55 4.74535 $w=2.53e-07 $l=1.05e-07 $layer=LI1_cond $X=9.007 $Y=1.53
+ $X2=9.007 $Y2=1.635
r144 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.025 $Y=1.53
+ $X2=9.025 $Y2=1.53
r145 33 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.87 $Y=1.53
+ $X2=6.725 $Y2=1.53
r146 32 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.88 $Y=1.53
+ $X2=9.025 $Y2=1.53
r147 32 33 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=8.88 $Y=1.53
+ $X2=6.87 $Y2=1.53
r148 30 45 6.30242 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=6.725 $Y=1.605
+ $X2=6.9 $Y2=1.605
r149 30 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.725 $Y=1.53
+ $X2=6.725 $Y2=1.53
r150 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.63 $X2=9.78 $Y2=1.63
r151 25 55 2.77751 $w=1.8e-07 $l=1.28e-07 $layer=LI1_cond $X=9.135 $Y=1.635
+ $X2=9.007 $Y2=1.635
r152 25 27 39.7424 $w=1.78e-07 $l=6.45e-07 $layer=LI1_cond $X=9.135 $Y=1.635
+ $X2=9.78 $Y2=1.635
r153 23 28 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=9.78 $Y=1.6 $X2=9.78
+ $Y2=1.63
r154 23 24 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=9.78 $Y=1.6
+ $X2=9.78 $Y2=1.465
r155 21 28 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=9.78 $Y=1.835
+ $X2=9.78 $Y2=1.63
r156 21 22 45.0833 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=9.715 $Y=1.835
+ $X2=9.715 $Y2=1.985
r157 19 46 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.97 $Y=1.365
+ $X2=6.97 $Y2=1.515
r158 18 19 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.995 $Y=1.215
+ $X2=6.995 $Y2=1.365
r159 16 24 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=9.84 $Y=0.445
+ $X2=9.84 $Y2=1.465
r160 13 22 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.59 $Y=2.275
+ $X2=9.59 $Y2=1.985
r161 9 18 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.02 $Y=0.445
+ $X2=7.02 $Y2=1.215
r162 5 47 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.97 $Y=2.275
+ $X2=6.97 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_1781_295# 1 2 9 11 12 15 18 21 22 24 25
+ 28 31 33 36
c107 36 0 1.11257e-19 $X=10.785 $Y=1.28
c108 25 0 6.7173e-20 $X=9.53 $Y=1.28
c109 12 0 1.89883e-19 $X=9.055 $Y=1.55
c110 11 0 1.97973e-19 $X=9.285 $Y=1.55
r111 33 35 6.80499 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=0.42
+ $X2=10.745 $Y2=0.585
r112 31 36 3.77418 $w=2.45e-07 $l=9.21954e-08 $layer=LI1_cond $X=10.8 $Y=1.195
+ $X2=10.785 $Y2=1.28
r113 31 35 30.5648 $w=2.28e-07 $l=6.1e-07 $layer=LI1_cond $X=10.8 $Y=1.195
+ $X2=10.8 $Y2=0.585
r114 26 36 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.785 $Y=1.365
+ $X2=10.785 $Y2=1.28
r115 26 28 40.7788 $w=2.58e-07 $l=9.2e-07 $layer=LI1_cond $X=10.785 $Y=1.365
+ $X2=10.785 $Y2=2.285
r116 24 36 2.68609 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.655 $Y=1.28
+ $X2=10.785 $Y2=1.28
r117 24 25 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=10.655 $Y=1.28
+ $X2=9.53 $Y2=1.28
r118 22 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.42 $Y=1.02
+ $X2=9.42 $Y2=1.185
r119 22 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.42 $Y=1.02
+ $X2=9.42 $Y2=0.855
r120 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.42
+ $Y=1.02 $X2=9.42 $Y2=1.02
r121 19 25 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.425 $Y=1.195
+ $X2=9.53 $Y2=1.28
r122 19 21 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=9.425 $Y=1.195
+ $X2=9.425 $Y2=1.02
r123 18 39 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.36 $Y=1.475
+ $X2=9.36 $Y2=1.185
r124 15 38 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.36 $Y=0.445
+ $X2=9.36 $Y2=0.855
r125 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.285 $Y=1.55
+ $X2=9.36 $Y2=1.475
r126 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=9.285 $Y=1.55
+ $X2=9.055 $Y2=1.55
r127 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.98 $Y=1.625
+ $X2=9.055 $Y2=1.55
r128 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=8.98 $Y=1.625
+ $X2=8.98 $Y2=2.275
r129 2 28 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=2.065 $X2=10.74 $Y2=2.285
r130 1 33 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=10.485
+ $Y=0.235 $X2=10.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_1597_329# 1 2 3 14 17 19 23 27 29 30 32
+ 33 34 38 42 46 49 50 52 53 55 57 61 63 64 70
c155 63 0 1.3574e-19 $X=10.32 $Y=1.69
c156 57 0 1.42862e-19 $X=8.905 $Y=1.98
c157 23 0 1.64486e-19 $X=11.47 $Y=0.56
r158 64 71 43.2312 $w=4.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.38 $Y=1.69
+ $X2=10.38 $Y2=1.825
r159 64 70 17.8241 $w=4.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.38 $Y=1.69
+ $X2=10.38 $Y2=1.555
r160 63 66 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=10.32 $Y=1.69
+ $X2=10.32 $Y2=1.98
r161 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.32
+ $Y=1.69 $X2=10.32 $Y2=1.69
r162 56 61 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=9.965 $Y=1.98
+ $X2=9.812 $Y2=1.98
r163 55 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.155 $Y=1.98
+ $X2=10.32 $Y2=1.98
r164 55 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.155 $Y=1.98
+ $X2=9.965 $Y2=1.98
r165 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.35
+ $Y=0.93 $X2=10.35 $Y2=0.93
r166 50 52 22.0467 $w=2.28e-07 $l=4.4e-07 $layer=LI1_cond $X=9.91 $Y=0.9
+ $X2=10.35 $Y2=0.9
r167 49 50 6.85974 $w=2.3e-07 $l=1.57242e-07 $layer=LI1_cond $X=9.81 $Y=0.785
+ $X2=9.91 $Y2=0.9
r168 48 49 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=9.81 $Y=0.545
+ $X2=9.81 $Y2=0.785
r169 44 61 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.812 $Y=2.065
+ $X2=9.812 $Y2=1.98
r170 44 46 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=9.812 $Y=2.065
+ $X2=9.812 $Y2=2.285
r171 43 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=1.98
+ $X2=8.905 $Y2=1.98
r172 42 61 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.66 $Y=1.98
+ $X2=9.812 $Y2=1.98
r173 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.66 $Y=1.98
+ $X2=8.99 $Y2=1.98
r174 38 48 7.01501 $w=2.7e-07 $l=1.78115e-07 $layer=LI1_cond $X=9.71 $Y=0.41
+ $X2=9.81 $Y2=0.545
r175 38 40 46.0977 $w=2.68e-07 $l=1.08e-06 $layer=LI1_cond $X=9.71 $Y=0.41
+ $X2=8.63 $Y2=0.41
r176 34 57 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=8.905 $Y=2.292
+ $X2=8.905 $Y2=1.98
r177 34 36 18.9207 $w=3.33e-07 $l=5.5e-07 $layer=LI1_cond $X=8.82 $Y=2.292
+ $X2=8.27 $Y2=2.292
r178 31 53 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=10.35 $Y=1.205
+ $X2=10.35 $Y2=0.93
r179 31 32 10.1687 $w=3.3e-07 $l=1.00623e-07 $layer=POLY_cond $X=10.35 $Y=1.205
+ $X2=10.41 $Y2=1.28
r180 29 53 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=10.35 $Y=0.9
+ $X2=10.35 $Y2=0.93
r181 29 30 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=10.35 $Y=0.9
+ $X2=10.35 $Y2=0.765
r182 25 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.47 $Y=1.355
+ $X2=11.47 $Y2=1.28
r183 25 27 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.47 $Y=1.355
+ $X2=11.47 $Y2=1.985
r184 21 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.47 $Y=1.205
+ $X2=11.47 $Y2=1.28
r185 21 23 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=11.47 $Y=1.205
+ $X2=11.47 $Y2=0.56
r186 20 32 16.9349 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=10.605 $Y=1.28
+ $X2=10.41 $Y2=1.28
r187 19 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.395 $Y=1.28
+ $X2=11.47 $Y2=1.28
r188 19 20 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.395 $Y=1.28
+ $X2=10.605 $Y2=1.28
r189 17 71 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=10.53 $Y=2.275
+ $X2=10.53 $Y2=1.825
r190 14 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.41 $Y=0.445
+ $X2=10.41 $Y2=0.765
r191 10 32 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.41 $Y=1.355
+ $X2=10.41 $Y2=1.28
r192 10 70 28.5207 $w=3.9e-07 $l=2e-07 $layer=POLY_cond $X=10.41 $Y=1.355
+ $X2=10.41 $Y2=1.555
r193 3 46 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=2.065 $X2=9.8 $Y2=2.285
r194 2 36 600 $w=1.7e-07 $l=7.745e-07 $layer=licon1_PDIFF $count=1 $X=7.985
+ $Y=1.645 $X2=8.27 $Y2=2.29
r195 1 40 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=0.235 $X2=8.63 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_2227_47# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 37 41 45 48 54
r93 53 54 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.835 $Y=1.16
+ $X2=13.255 $Y2=1.16
r94 52 53 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=12.365 $Y=1.16
+ $X2=12.835 $Y2=1.16
r95 51 52 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=11.945 $Y=1.16
+ $X2=12.365 $Y2=1.16
r96 46 51 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=11.89 $Y=1.16
+ $X2=11.945 $Y2=1.16
r97 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.89
+ $Y=1.16 $X2=11.89 $Y2=1.16
r98 43 48 0.499868 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=11.345 $Y=1.16
+ $X2=11.215 $Y2=1.16
r99 43 45 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=11.345 $Y=1.16
+ $X2=11.89 $Y2=1.16
r100 39 48 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=11.215 $Y=1.325
+ $X2=11.215 $Y2=1.16
r101 39 41 27.9246 $w=2.58e-07 $l=6.3e-07 $layer=LI1_cond $X=11.215 $Y=1.325
+ $X2=11.215 $Y2=1.955
r102 35 48 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=11.215 $Y=0.995
+ $X2=11.215 $Y2=1.16
r103 35 37 25.2651 $w=2.58e-07 $l=5.7e-07 $layer=LI1_cond $X=11.215 $Y=0.995
+ $X2=11.215 $Y2=0.425
r104 31 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.255 $Y=1.325
+ $X2=13.255 $Y2=1.16
r105 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.255 $Y=1.325
+ $X2=13.255 $Y2=1.985
r106 28 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.255 $Y=0.995
+ $X2=13.255 $Y2=1.16
r107 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.255 $Y=0.995
+ $X2=13.255 $Y2=0.56
r108 24 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.835 $Y=1.325
+ $X2=12.835 $Y2=1.16
r109 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.835 $Y=1.325
+ $X2=12.835 $Y2=1.985
r110 21 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.835 $Y=0.995
+ $X2=12.835 $Y2=1.16
r111 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.835 $Y=0.995
+ $X2=12.835 $Y2=0.56
r112 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.365 $Y=1.325
+ $X2=12.365 $Y2=1.16
r113 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.365 $Y=1.325
+ $X2=12.365 $Y2=1.985
r114 14 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.365 $Y=0.995
+ $X2=12.365 $Y2=1.16
r115 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.365 $Y=0.995
+ $X2=12.365 $Y2=0.56
r116 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.945 $Y=1.325
+ $X2=11.945 $Y2=1.16
r117 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.945 $Y=1.325
+ $X2=11.945 $Y2=1.985
r118 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.945 $Y=0.995
+ $X2=11.945 $Y2=1.16
r119 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.945 $Y=0.995
+ $X2=11.945 $Y2=0.56
r120 2 41 300 $w=1.7e-07 $l=5.28819e-07 $layer=licon1_PDIFF $count=2 $X=11.135
+ $Y=1.485 $X2=11.26 $Y2=1.955
r121 1 37 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=11.135
+ $Y=0.235 $X2=11.26 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_27_369# 1 2 7 10 11 13 14 16
r41 14 16 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=1.125 $Y=2.36
+ $X2=1.88 $Y2=2.36
r42 13 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.04 $Y=2.255
+ $X2=1.125 $Y2=2.36
r43 12 13 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.04 $Y=2.025
+ $X2=1.04 $Y2=2.255
r44 10 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.955 $Y=1.935
+ $X2=1.04 $Y2=2.025
r45 10 11 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=0.955 $Y=1.935
+ $X2=0.345 $Y2=1.935
r46 7 11 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.345 $Y2=1.935
r47 7 9 2.11154 $w=2.6e-07 $l=4.5e-08 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.215 $Y2=2.07
r48 2 16 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=1.845 $X2=1.88 $Y2=2.34
r49 1 9 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 47 51 55
+ 61 65 67 72 73 75 76 78 79 80 82 94 98 110 114 123 128 131 134 143 149 151 154
+ 158
c207 158 0 5.68782e-20 $X=13.57 $Y=2.72
c208 37 0 3.22446e-20 $X=2.82 $Y=2.34
c209 5 0 1.36329e-19 $X=7.045 $Y=2.065
r210 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r211 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r212 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r213 147 149 15.2496 $w=6.78e-07 $l=4.25e-07 $layer=LI1_cond $X=7.59 $Y=2.465
+ $X2=8.015 $Y2=2.465
r214 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r215 145 147 6.42013 $w=6.78e-07 $l=3.65e-07 $layer=LI1_cond $X=7.225 $Y=2.465
+ $X2=7.59 $Y2=2.465
r216 142 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r217 141 145 1.67099 $w=6.78e-07 $l=9.5e-08 $layer=LI1_cond $X=7.13 $Y=2.465
+ $X2=7.225 $Y2=2.465
r218 141 143 9.00537 $w=6.78e-07 $l=7e-08 $layer=LI1_cond $X=7.13 $Y=2.465
+ $X2=7.06 $Y2=2.465
r219 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r220 138 142 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r221 131 132 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r222 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r223 126 158 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r224 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r225 123 157 4.85147 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=13.38 $Y=2.72
+ $X2=13.59 $Y2=2.72
r226 123 125 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=13.38 $Y=2.72
+ $X2=13.11 $Y2=2.72
r227 122 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=13.11 $Y2=2.72
r228 122 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r229 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r230 119 154 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=11.87 $Y=2.72
+ $X2=11.692 $Y2=2.72
r231 119 121 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.87 $Y=2.72
+ $X2=12.19 $Y2=2.72
r232 118 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r233 118 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=10.35 $Y2=2.72
r234 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r235 115 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=2.72
+ $X2=10.32 $Y2=2.72
r236 115 117 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=10.485 $Y=2.72
+ $X2=11.27 $Y2=2.72
r237 114 154 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=11.515 $Y=2.72
+ $X2=11.692 $Y2=2.72
r238 114 117 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.515 $Y=2.72
+ $X2=11.27 $Y2=2.72
r239 113 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r240 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r241 110 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.155 $Y=2.72
+ $X2=10.32 $Y2=2.72
r242 110 112 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.155 $Y=2.72
+ $X2=9.89 $Y2=2.72
r243 109 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r244 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r245 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r246 106 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r247 105 108 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r248 105 149 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.015 $Y2=2.72
r249 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r250 102 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r251 102 132 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=3.91 $Y2=2.72
r252 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r253 99 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=3.76 $Y2=2.72
r254 99 101 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r255 98 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r256 98 134 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=6.137 $Y=2.72
+ $X2=6.137 $Y2=2.36
r257 98 101 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=5.75 $Y2=2.72
r258 97 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r259 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r260 94 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.76 $Y2=2.72
r261 94 96 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.45 $Y2=2.72
r262 93 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r263 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r264 90 93 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r265 90 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r266 89 92 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r267 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r268 87 128 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.785 $Y=2.72
+ $X2=0.65 $Y2=2.72
r269 87 89 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=2.72
+ $X2=1.15 $Y2=2.72
r270 82 128 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.65 $Y2=2.72
r271 82 84 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r272 80 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r273 80 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r274 78 121 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.54 $Y=2.72
+ $X2=12.19 $Y2=2.72
r275 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.54 $Y=2.72
+ $X2=12.625 $Y2=2.72
r276 77 125 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=12.71 $Y=2.72
+ $X2=13.11 $Y2=2.72
r277 77 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.71 $Y=2.72
+ $X2=12.625 $Y2=2.72
r278 75 108 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.16 $Y=2.72
+ $X2=8.97 $Y2=2.72
r279 75 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.16 $Y=2.72
+ $X2=9.325 $Y2=2.72
r280 74 112 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.49 $Y=2.72
+ $X2=9.89 $Y2=2.72
r281 74 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.49 $Y=2.72
+ $X2=9.325 $Y2=2.72
r282 72 92 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r283 72 73 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.837 $Y2=2.72
r284 71 96 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.985 $Y=2.72
+ $X2=3.45 $Y2=2.72
r285 71 73 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.985 $Y=2.72
+ $X2=2.837 $Y2=2.72
r286 67 70 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=13.547 $Y=1.66
+ $X2=13.547 $Y2=2.34
r287 65 157 2.95709 $w=3.35e-07 $l=1.04307e-07 $layer=LI1_cond $X=13.547
+ $Y=2.635 $X2=13.59 $Y2=2.72
r288 65 70 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=13.547 $Y=2.635
+ $X2=13.547 $Y2=2.34
r289 61 64 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=12.625 $Y=1.66
+ $X2=12.625 $Y2=2.34
r290 59 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.625 $Y=2.635
+ $X2=12.625 $Y2=2.72
r291 59 64 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.625 $Y=2.635
+ $X2=12.625 $Y2=2.34
r292 55 58 22.075 $w=3.53e-07 $l=6.8e-07 $layer=LI1_cond $X=11.692 $Y=1.68
+ $X2=11.692 $Y2=2.36
r293 53 154 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.692 $Y=2.635
+ $X2=11.692 $Y2=2.72
r294 53 58 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=11.692 $Y=2.635
+ $X2=11.692 $Y2=2.36
r295 49 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.32 $Y=2.635
+ $X2=10.32 $Y2=2.72
r296 49 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.32 $Y=2.635
+ $X2=10.32 $Y2=2.34
r297 45 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=2.635
+ $X2=9.325 $Y2=2.72
r298 45 47 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.325 $Y=2.635
+ $X2=9.325 $Y2=2.36
r299 44 98 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=6.137 $Y2=2.72
r300 44 143 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=7.06 $Y2=2.72
r301 39 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=2.635
+ $X2=3.76 $Y2=2.72
r302 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.76 $Y=2.635
+ $X2=3.76 $Y2=2.36
r303 35 73 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.837 $Y=2.635
+ $X2=2.837 $Y2=2.72
r304 35 37 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=2.837 $Y=2.635
+ $X2=2.837 $Y2=2.34
r305 31 128 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=2.635
+ $X2=0.65 $Y2=2.72
r306 31 33 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.65 $Y=2.635
+ $X2=0.65 $Y2=2.36
r307 10 70 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=13.33
+ $Y=1.485 $X2=13.465 $Y2=2.34
r308 10 67 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=13.33
+ $Y=1.485 $X2=13.465 $Y2=1.66
r309 9 64 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=12.44
+ $Y=1.485 $X2=12.625 $Y2=2.34
r310 9 61 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=12.44
+ $Y=1.485 $X2=12.625 $Y2=1.66
r311 8 58 400 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=1.485 $X2=11.705 $Y2=2.36
r312 8 55 400 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=1.485 $X2=11.705 $Y2=1.68
r313 7 51 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=10.195
+ $Y=2.065 $X2=10.32 $Y2=2.34
r314 6 47 600 $w=1.7e-07 $l=4.08258e-07 $layer=licon1_PDIFF $count=1 $X=9.055
+ $Y=2.065 $X2=9.325 $Y2=2.36
r315 5 145 600 $w=1.7e-07 $l=3.74333e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=2.065 $X2=7.225 $Y2=2.36
r316 4 134 600 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_PDIFF $count=1 $X=5.915
+ $Y=2.065 $X2=6.11 $Y2=2.36
r317 3 41 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.845 $X2=3.76 $Y2=2.36
r318 2 37 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.845 $X2=2.82 $Y2=2.34
r319 1 33 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%A_181_47# 1 2 3 4 13 19 21 23 26 30 33 35
+ 36 37 40 43
c137 43 0 3.47594e-20 $X=4.83 $Y=1.53
c138 37 0 1.4475e-19 $X=1.755 $Y=1.53
c139 30 0 1.86564e-19 $X=1.6 $Y=1.965
c140 19 0 9.48056e-20 $X=4.73 $Y=0.42
r141 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.53
+ $X2=4.83 $Y2=1.53
r142 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.53
+ $X2=1.61 $Y2=1.53
r143 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.53
+ $X2=1.61 $Y2=1.53
r144 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.53
+ $X2=4.83 $Y2=1.53
r145 36 37 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=4.685 $Y=1.53
+ $X2=1.755 $Y2=1.53
r146 33 40 42.3206 $w=1.88e-07 $l=7.25e-07 $layer=LI1_cond $X=1.6 $Y=0.805
+ $X2=1.6 $Y2=1.53
r147 31 40 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=1.6 $Y=1.845
+ $X2=1.6 $Y2=1.53
r148 30 31 2.10789 $w=1.9e-07 $l=1.2e-07 $layer=LI1_cond $X=1.6 $Y=1.965 $X2=1.6
+ $Y2=1.845
r149 28 30 6.72258 $w=2.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.46 $Y=1.965
+ $X2=1.6 $Y2=1.965
r150 26 44 5.45457 $w=2.61e-07 $l=9.44722e-08 $layer=LI1_cond $X=4.745 $Y=1.445
+ $X2=4.765 $Y2=1.53
r151 26 35 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.745 $Y=1.445
+ $X2=4.745 $Y2=0.92
r152 21 44 4.38824 $w=2.61e-07 $l=1.04307e-07 $layer=LI1_cond $X=4.722 $Y=1.615
+ $X2=4.765 $Y2=1.53
r153 21 23 36.7174 $w=2.13e-07 $l=6.85e-07 $layer=LI1_cond $X=4.722 $Y=1.615
+ $X2=4.722 $Y2=2.3
r154 17 35 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=4.667 $Y=0.758
+ $X2=4.667 $Y2=0.92
r155 17 19 11.9854 $w=3.23e-07 $l=3.38e-07 $layer=LI1_cond $X=4.667 $Y=0.758
+ $X2=4.667 $Y2=0.42
r156 13 33 20.7082 $w=2.28e-07 $l=4.10293e-07 $layer=LI1_cond $X=1.537 $Y=0.425
+ $X2=1.6 $Y2=0.805
r157 13 15 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.38 $Y=0.425
+ $X2=1.04 $Y2=0.425
r158 4 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=4.575
+ $Y=2.065 $X2=4.7 $Y2=2.3
r159 3 28 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.325
+ $Y=1.845 $X2=1.46 $Y2=1.97
r160 2 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.605
+ $Y=0.235 $X2=4.73 $Y2=0.42
r161 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.905
+ $Y=0.235 $X2=1.04 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%Q 1 2 3 4 15 19 23 24 25 26 27 28 29 30 31
+ 44 51 72
c43 51 0 2.2939e-20 $X=12.285 $Y=0.85
c44 27 0 1.0279e-19 $X=12.285 $Y=1.19
r45 72 73 2.39662 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=12.205 $Y=1.53
+ $X2=12.205 $Y2=1.495
r46 51 68 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=12.257 $Y=0.85
+ $X2=12.257 $Y2=0.825
r47 30 62 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=12.205 $Y=2.21
+ $X2=12.205 $Y2=2.285
r48 29 30 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=12.205 $Y=1.87
+ $X2=12.205 $Y2=2.21
r49 29 56 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=12.205 $Y=1.87
+ $X2=12.205 $Y2=1.66
r50 28 56 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=12.205 $Y=1.555
+ $X2=12.205 $Y2=1.66
r51 28 72 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=12.205 $Y=1.555
+ $X2=12.205 $Y2=1.53
r52 28 73 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=12.257 $Y=1.47
+ $X2=12.257 $Y2=1.495
r53 28 53 7.42686 $w=2.23e-07 $l=1.45e-07 $layer=LI1_cond $X=12.257 $Y=1.47
+ $X2=12.257 $Y2=1.325
r54 27 49 5.99569 $w=2.25e-07 $l=1.35e-07 $layer=LI1_cond $X=12.257 $Y=1.19
+ $X2=12.257 $Y2=1.055
r55 27 53 5.99569 $w=2.25e-07 $l=1.35e-07 $layer=LI1_cond $X=12.257 $Y=1.19
+ $X2=12.257 $Y2=1.325
r56 27 31 11.5307 $w=4.38e-07 $l=3.75e-07 $layer=LI1_cond $X=12.37 $Y=1.19
+ $X2=12.745 $Y2=1.19
r57 26 68 2.22201 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=12.205 $Y=0.795
+ $X2=12.205 $Y2=0.825
r58 26 42 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=12.205 $Y=0.795
+ $X2=12.205 $Y2=0.66
r59 26 49 8.96345 $w=2.23e-07 $l=1.75e-07 $layer=LI1_cond $X=12.257 $Y=0.88
+ $X2=12.257 $Y2=1.055
r60 26 51 1.53659 $w=2.23e-07 $l=3e-08 $layer=LI1_cond $X=12.257 $Y=0.88
+ $X2=12.257 $Y2=0.85
r61 25 42 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=12.205 $Y=0.51
+ $X2=12.205 $Y2=0.66
r62 25 44 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=12.205 $Y=0.51
+ $X2=12.205 $Y2=0.44
r63 23 31 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=12.88 $Y=1.19
+ $X2=12.745 $Y2=1.19
r64 23 24 2.07418 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.88 $Y=1.19
+ $X2=13.045 $Y2=1.19
r65 19 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.045 $Y=1.675
+ $X2=13.045 $Y2=2.355
r66 17 24 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=13.045 $Y=1.325
+ $X2=13.045 $Y2=1.19
r67 17 19 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=13.045 $Y=1.325
+ $X2=13.045 $Y2=1.675
r68 13 24 4.35802 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=13.045 $Y=1.055
+ $X2=13.045 $Y2=1.19
r69 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=13.045 $Y=1.055
+ $X2=13.045 $Y2=0.36
r70 4 21 400 $w=1.7e-07 $l=9.35067e-07 $layer=licon1_PDIFF $count=1 $X=12.91
+ $Y=1.485 $X2=13.045 $Y2=2.355
r71 4 19 400 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_PDIFF $count=1 $X=12.91
+ $Y=1.485 $X2=13.045 $Y2=1.675
r72 3 62 600 $w=1.7e-07 $l=8.6487e-07 $layer=licon1_PDIFF $count=1 $X=12.02
+ $Y=1.485 $X2=12.155 $Y2=2.285
r73 2 15 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=12.91
+ $Y=0.235 $X2=13.045 $Y2=0.36
r74 1 44 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=12.02
+ $Y=0.235 $X2=12.155 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__SDFSTP_4%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 55 57 60 61 63 64 65 71 75 80 90 98 107 112 119 122 133 137 139 142 146
c190 146 0 2.71124e-20 $X=13.57 $Y=0
c191 37 0 4.13602e-20 $X=2.85 $Y=0.38
r192 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r193 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r194 139 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r195 135 137 11.6653 $w=8.88e-07 $l=1.25e-07 $layer=LI1_cond $X=7.59 $Y=0.36
+ $X2=7.715 $Y2=0.36
r196 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r197 132 135 4.79775 $w=8.88e-07 $l=3.5e-07 $layer=LI1_cond $X=7.24 $Y=0.36
+ $X2=7.59 $Y2=0.36
r198 132 133 17.2855 $w=8.88e-07 $l=5.35e-07 $layer=LI1_cond $X=7.24 $Y=0.36
+ $X2=6.705 $Y2=0.36
r199 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r200 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r201 112 117 8.24843 $w=6.36e-07 $l=4.3e-07 $layer=LI1_cond $X=0.35 $Y=0
+ $X2=0.35 $Y2=0.43
r202 112 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r203 110 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=13.57 $Y2=0
r204 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r205 107 145 4.85147 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=13.38 $Y=0
+ $X2=13.59 $Y2=0
r206 107 109 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=13.38 $Y=0
+ $X2=13.11 $Y2=0
r207 106 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=13.11 $Y2=0
r208 106 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r209 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r210 103 142 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=11.87 $Y=0
+ $X2=11.692 $Y2=0
r211 103 105 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.87 $Y=0
+ $X2=12.19 $Y2=0
r212 102 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r213 102 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=10.35 $Y2=0
r214 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r215 99 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=10.24 $Y2=0
r216 99 101 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=11.27 $Y2=0
r217 98 142 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=11.515 $Y=0
+ $X2=11.692 $Y2=0
r218 98 101 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.515 $Y=0
+ $X2=11.27 $Y2=0
r219 97 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r220 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r221 94 97 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=9.89 $Y2=0
r222 94 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r223 93 96 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=8.05 $Y=0 $X2=9.89
+ $Y2=0
r224 93 137 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=7.715 $Y2=0
r225 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r226 90 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.24 $Y2=0
r227 90 96 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.89 $Y2=0
r228 89 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r229 89 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=5.75 $Y2=0
r230 88 133 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=6.705 $Y2=0
r231 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r232 86 88 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.67 $Y2=0
r233 84 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r234 84 123 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=3.91 $Y2=0
r235 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r236 81 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=3.79 $Y2=0
r237 81 83 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=5.29 $Y2=0
r238 80 129 9.37134 $w=4.83e-07 $l=3.8e-07 $layer=LI1_cond $X=5.852 $Y=0
+ $X2=5.852 $Y2=0.38
r239 80 86 6.96588 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=5.852 $Y=0
+ $X2=6.095 $Y2=0
r240 80 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r241 80 83 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.29
+ $Y2=0
r242 79 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r243 79 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.99 $Y2=0
r244 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r245 76 119 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.895
+ $Y2=0
r246 76 78 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.45
+ $Y2=0
r247 75 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0
+ $X2=3.79 $Y2=0
r248 75 78 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.625 $Y=0
+ $X2=3.45 $Y2=0
r249 74 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.99 $Y2=0
r250 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r251 71 119 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.69 $Y=0
+ $X2=2.895 $Y2=0
r252 71 73 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.53
+ $Y2=0
r253 70 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r254 70 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=0.69 $Y2=0
r255 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r256 67 112 8.69404 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=0.7 $Y=0 $X2=0.35
+ $Y2=0
r257 67 69 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.7 $Y=0 $X2=1.61
+ $Y2=0
r258 65 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r259 65 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r260 63 105 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.54 $Y=0
+ $X2=12.19 $Y2=0
r261 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.54 $Y=0
+ $X2=12.625 $Y2=0
r262 62 109 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=12.71 $Y=0 $X2=13.11
+ $Y2=0
r263 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.71 $Y=0
+ $X2=12.625 $Y2=0
r264 60 69 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=1.61 $Y2=0
r265 60 61 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=1.825 $Y=0
+ $X2=1.957 $Y2=0
r266 59 73 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.53
+ $Y2=0
r267 59 61 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.957
+ $Y2=0
r268 55 145 2.95709 $w=3.35e-07 $l=1.04307e-07 $layer=LI1_cond $X=13.547
+ $Y=0.085 $X2=13.59 $Y2=0
r269 55 57 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=13.547 $Y=0.085
+ $X2=13.547 $Y2=0.38
r270 51 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.625 $Y=0.085
+ $X2=12.625 $Y2=0
r271 51 53 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.625 $Y=0.085
+ $X2=12.625 $Y2=0.38
r272 47 142 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.692 $Y=0.085
+ $X2=11.692 $Y2=0
r273 47 49 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=11.692 $Y=0.085
+ $X2=11.692 $Y2=0.36
r274 43 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.24 $Y=0.085
+ $X2=10.24 $Y2=0
r275 43 45 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=10.24 $Y=0.085
+ $X2=10.24 $Y2=0.36
r276 39 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0
r277 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0.36
r278 35 119 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0
r279 35 37 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0.38
r280 31 61 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.957 $Y=0.085
+ $X2=1.957 $Y2=0
r281 31 33 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.957 $Y=0.085
+ $X2=1.957 $Y2=0.38
r282 10 57 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=13.33
+ $Y=0.235 $X2=13.465 $Y2=0.38
r283 9 53 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=12.44
+ $Y=0.235 $X2=12.625 $Y2=0.38
r284 8 49 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=11.545
+ $Y=0.235 $X2=11.705 $Y2=0.36
r285 7 45 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=9.915
+ $Y=0.235 $X2=10.2 $Y2=0.36
r286 6 132 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.095
+ $Y=0.235 $X2=7.24 $Y2=0.36
r287 5 129 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.235 $X2=5.93 $Y2=0.38
r288 4 41 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.235 $X2=3.79 $Y2=0.36
r289 3 37 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.85 $Y2=0.38
r290 2 33 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=1.745
+ $Y=0.235 $X2=1.91 $Y2=0.38
r291 1 117 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__xor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 2.800000 1.275000 ;
        RECT 2.630000 1.275000 2.800000 1.445000 ;
        RECT 2.630000 1.445000 6.165000 1.615000 ;
        RECT 5.995000 1.075000 7.370000 1.275000 ;
        RECT 5.995000 1.275000 6.165000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.075000 5.000000 1.105000 ;
        RECT 2.970000 1.105000 5.740000 1.275000 ;
    END
  END B
  PIN X
    ANTENNAPARTIALMETALSIDEAREA  2.359000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 0.645000 5.580000 0.905000 ;
        RECT 5.150000 0.905000 5.580000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.850000 0.725000  8.630000 0.735000 ;
        RECT 7.850000 0.735000 10.035000 0.905000 ;
        RECT 7.850000 0.905000  8.305000 0.935000 ;
        RECT 7.880000 1.445000 10.035000 1.625000 ;
        RECT 7.880000 1.625000  9.010000 1.665000 ;
        RECT 7.880000 1.665000  8.170000 2.125000 ;
        RECT 8.300000 0.255000  8.630000 0.725000 ;
        RECT 8.760000 1.665000  9.010000 2.125000 ;
        RECT 9.140000 0.255000  9.470000 0.735000 ;
        RECT 9.600000 1.625000 10.035000 2.465000 ;
        RECT 9.735000 0.905000 10.035000 1.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.145000 0.735000 5.435000 0.780000 ;
        RECT 5.145000 0.780000 8.195000 0.920000 ;
        RECT 5.145000 0.920000 5.435000 0.965000 ;
        RECT 7.905000 0.735000 8.195000 0.780000 ;
        RECT 7.905000 0.920000 8.195000 0.965000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.085000  0.085000  0.360000 0.565000 ;
        RECT 1.030000  0.085000  1.200000 0.555000 ;
        RECT 1.870000  0.085000  2.040000 0.555000 ;
        RECT 2.710000  0.085000  2.880000 0.555000 ;
        RECT 3.550000  0.085000  3.820000 0.895000 ;
        RECT 6.170000  0.085000  6.340000 0.555000 ;
        RECT 7.010000  0.085000  7.180000 0.555000 ;
        RECT 7.960000  0.085000  8.130000 0.555000 ;
        RECT 8.800000  0.085000  8.970000 0.555000 ;
        RECT 9.640000  0.085000  9.810000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.570000 2.175000  0.820000 2.635000 ;
        RECT 1.410000 2.175000  1.660000 2.635000 ;
        RECT 4.450000 2.175000  4.700000 2.635000 ;
        RECT 5.290000 2.175000  5.540000 2.635000 ;
        RECT 6.130000 2.175000  6.380000 2.635000 ;
        RECT 6.970000 2.175000  7.220000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.735000 3.380000 0.905000 ;
      RECT 0.085000 0.905000 0.255000 1.445000 ;
      RECT 0.085000 1.445000 2.420000 1.615000 ;
      RECT 0.085000 1.785000 2.080000 2.005000 ;
      RECT 0.085000 2.005000 0.400000 2.465000 ;
      RECT 0.530000 0.255000 0.860000 0.725000 ;
      RECT 0.530000 0.725000 3.380000 0.735000 ;
      RECT 0.990000 2.005000 1.240000 2.465000 ;
      RECT 1.370000 0.255000 1.700000 0.725000 ;
      RECT 1.830000 2.005000 2.080000 2.295000 ;
      RECT 1.830000 2.295000 3.760000 2.465000 ;
      RECT 2.210000 0.255000 2.540000 0.725000 ;
      RECT 2.250000 1.615000 2.420000 1.785000 ;
      RECT 2.250000 1.785000 3.340000 1.955000 ;
      RECT 2.250000 1.955000 2.500000 2.125000 ;
      RECT 2.670000 2.125000 2.920000 2.295000 ;
      RECT 3.050000 0.255000 3.380000 0.725000 ;
      RECT 3.090000 1.955000 3.340000 2.125000 ;
      RECT 3.510000 1.795000 3.760000 2.295000 ;
      RECT 3.990000 0.255000 6.000000 0.475000 ;
      RECT 4.030000 1.785000 7.640000 2.005000 ;
      RECT 4.030000 2.005000 4.280000 2.465000 ;
      RECT 4.870000 2.005000 5.120000 2.465000 ;
      RECT 5.710000 2.005000 5.960000 2.465000 ;
      RECT 5.750000 0.475000 6.000000 0.725000 ;
      RECT 5.750000 0.725000 7.680000 0.905000 ;
      RECT 6.510000 0.255000 6.840000 0.725000 ;
      RECT 6.550000 1.455000 6.800000 1.785000 ;
      RECT 6.550000 2.005000 6.800000 2.465000 ;
      RECT 7.260000 1.445000 7.710000 1.615000 ;
      RECT 7.350000 0.255000 7.680000 0.725000 ;
      RECT 7.390000 2.005000 7.640000 2.295000 ;
      RECT 7.390000 2.295000 9.430000 2.465000 ;
      RECT 7.540000 1.105000 9.565000 1.275000 ;
      RECT 7.540000 1.275000 7.710000 1.445000 ;
      RECT 8.340000 1.835000 8.590000 2.295000 ;
      RECT 8.540000 1.075000 9.565000 1.105000 ;
      RECT 9.180000 1.795000 9.430000 2.295000 ;
    LAYER mcon ;
      RECT 1.985000 1.445000 2.155000 1.615000 ;
      RECT 7.505000 1.445000 7.675000 1.615000 ;
    LAYER met1 ;
      RECT 1.925000 1.415000 2.215000 1.460000 ;
      RECT 1.925000 1.460000 7.735000 1.600000 ;
      RECT 1.925000 1.600000 2.215000 1.645000 ;
      RECT 7.445000 1.415000 7.735000 1.460000 ;
      RECT 7.445000 1.600000 7.735000 1.645000 ;
  END
END sky130_fd_sc_hd__xor2_4

* File: sky130_fd_sc_hd__clkinv_1.pxi.spice
* Created: Tue Sep  1 19:01:21 2020
* 
x_PM_SKY130_FD_SC_HD__CLKINV_1%A N_A_M1000_g N_A_M1002_g N_A_M1001_g A A A
+ N_A_c_23_n PM_SKY130_FD_SC_HD__CLKINV_1%A
x_PM_SKY130_FD_SC_HD__CLKINV_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_c_52_n
+ N_VPWR_c_53_n N_VPWR_c_54_n N_VPWR_c_55_n VPWR N_VPWR_c_56_n N_VPWR_c_51_n
+ PM_SKY130_FD_SC_HD__CLKINV_1%VPWR
x_PM_SKY130_FD_SC_HD__CLKINV_1%Y N_Y_M1002_s N_Y_M1000_s N_Y_c_70_n Y Y Y
+ PM_SKY130_FD_SC_HD__CLKINV_1%Y
x_PM_SKY130_FD_SC_HD__CLKINV_1%VGND N_VGND_M1002_d N_VGND_c_92_n N_VGND_c_93_n
+ VGND N_VGND_c_94_n N_VGND_c_95_n PM_SKY130_FD_SC_HD__CLKINV_1%VGND
cc_1 VNB N_A_M1002_g 0.0412023f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=0.445
cc_2 VNB A 0.043896f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_3 VNB N_A_c_23_n 0.0736352f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.16
cc_4 VNB N_VPWR_c_51_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_Y_c_70_n 0.00995349f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.345
cc_6 VNB Y 0.0363467f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_7 VNB N_VGND_c_92_n 0.0103648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_VGND_c_93_n 0.0193136f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=0.445
cc_9 VNB N_VGND_c_94_n 0.0287474f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=2.065
cc_10 VNB N_VGND_c_95_n 0.113496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VPB N_A_M1000_g 0.0359234f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.065
cc_12 VPB N_A_M1001_g 0.0359234f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=2.065
cc_13 VPB A 0.00366f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.425
cc_14 VPB N_A_c_23_n 0.0188513f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=1.16
cc_15 VPB N_VPWR_c_52_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.885 $Y2=0.445
cc_16 VPB N_VPWR_c_53_n 0.0362093f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.345
cc_17 VPB N_VPWR_c_54_n 0.0102689f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=2.065
cc_18 VPB N_VPWR_c_55_n 0.036733f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.425
cc_19 VPB N_VPWR_c_56_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_51_n 0.0419516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_21 N_A_M1000_g N_VPWR_c_53_n 0.0055291f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_22 A N_VPWR_c_53_n 0.0123519f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_23 N_A_c_23_n N_VPWR_c_53_n 0.002208f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_24 N_A_M1001_g N_VPWR_c_55_n 0.00553885f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_25 N_A_M1000_g N_VPWR_c_56_n 0.00541359f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_26 N_A_M1001_g N_VPWR_c_56_n 0.00541359f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_27 N_A_M1000_g N_VPWR_c_51_n 0.0104557f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_28 N_A_M1001_g N_VPWR_c_51_n 0.0104744f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_29 N_A_M1002_g N_Y_c_70_n 0.0140555f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_30 A N_Y_c_70_n 0.0289142f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_31 N_A_c_23_n N_Y_c_70_n 0.00123281f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_32 N_A_M1000_g Y 0.0278674f $X=0.47 $Y=2.065 $X2=0 $Y2=0
cc_33 N_A_M1001_g Y 0.0278674f $X=0.89 $Y=2.065 $X2=0 $Y2=0
cc_34 A Y 0.00234543f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_35 N_A_c_23_n Y 0.0085603f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_36 N_A_M1002_g Y 0.0150252f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_37 A Y 0.0395886f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_38 N_A_c_23_n Y 0.0371028f $X=0.885 $Y=1.16 $X2=0 $Y2=0
cc_39 N_A_M1002_g N_VGND_c_93_n 0.00453359f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_40 N_A_M1002_g N_VGND_c_94_n 0.00426127f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_41 A N_VGND_c_94_n 0.00966373f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_42 N_A_M1002_g N_VGND_c_95_n 0.00818506f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_43 A N_VGND_c_95_n 0.00857725f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_44 N_VPWR_c_51_n N_Y_M1000_s 0.00215201f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_45 N_VPWR_c_56_n Y 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_46 N_VPWR_c_51_n Y 0.0122217f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_47 N_VPWR_c_55_n Y 0.0141111f $X=1.1 $Y=1.83 $X2=0 $Y2=0
cc_48 Y N_VGND_c_93_n 0.024392f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_49 N_Y_c_70_n N_VGND_c_94_n 0.02028f $X=0.675 $Y=0.435 $X2=0 $Y2=0
cc_50 Y N_VGND_c_94_n 0.00241655f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_51 N_Y_M1002_s N_VGND_c_95_n 0.00209319f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_52 N_Y_c_70_n N_VGND_c_95_n 0.01214f $X=0.675 $Y=0.435 $X2=0 $Y2=0
cc_53 Y N_VGND_c_95_n 0.005135f $X=1.065 $Y=0.765 $X2=0 $Y2=0

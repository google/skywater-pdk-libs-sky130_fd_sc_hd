* File: sky130_fd_sc_hd__mux4_1.spice
* Created: Thu Aug 27 14:28:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux4_1.pex.spice"
.subckt sky130_fd_sc_hd__mux4_1  VNB VPB A1 A0 S0 A3 A2 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A2	A2
* A3	A3
* S0	S0
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_A1_M1021_g N_A_27_47#_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1013 A_193_47# N_A0_M1013_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0567 PD=0.69 PS=0.69 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.9
+ A=0.063 P=1.14 MULT=1
MM1017 N_A_277_47#_M1017_d N_A_247_21#_M1017_g A_193_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.085225 AS=0.0567 PD=0.925 PS=0.69 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75001 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1011 N_A_27_47#_M1011_d N_S0_M1011_g N_A_277_47#_M1017_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.085225 PD=1.36 PS=0.925 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_S0_M1006_g N_A_247_21#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_750_97#_M1018_d N_S0_M1018_g N_A_668_97#_M1018_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_834_97#_M1022_d N_A_247_21#_M1022_g N_A_750_97#_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.10795 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A3_M1023_g N_A_668_97#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1079 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_834_97#_M1024_d N_A2_M1024_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_1290_413#_M1015_d N_S1_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_1478_413#_M1005_d N_S1_M1005_g N_A_750_97#_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.151025 AS=0.1092 PD=1.285 PS=1.36 NRD=78.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_277_47#_M1007_d N_A_1290_413#_M1007_g N_A_1478_413#_M1005_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.1092 AS=0.151025 PD=1.36 PS=1.285 NRD=0 NRS=87.012
+ M=1 R=2.8 SA=75000.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_X_M1020_d N_A_1478_413#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_27_413#_M1010_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_193_413#_M1025_d N_A0_M1025_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_277_47#_M1014_d N_A_247_21#_M1014_g N_A_27_413#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_193_413#_M1012_d N_S0_M1012_g N_A_277_47#_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1079 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_S0_M1002_g N_A_247_21#_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1079 AS=0.1083 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_750_97#_M1000_d N_S0_M1000_g N_A_757_363#_M1000_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.1079 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_923_363# N_A_247_21#_M1008_g N_A_750_97#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.090125 AS=0.0567 PD=0.995 PS=0.69 NRD=74.8403 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A3_M1004_g A_923_363# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.090125 PD=0.69 PS=0.995 NRD=0 NRS=74.8403 M=1 R=2.8 SA=75000.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_A_757_363#_M1019_d N_A2_M1019_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_1290_413#_M1009_d N_S1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_1478_413#_M1001_d N_S1_M1001_g N_A_277_47#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0920875 AS=0.1092 PD=0.99 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_750_97#_M1003_d N_A_1290_413#_M1003_g N_A_1478_413#_M1001_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.2688 AS=0.0920875 PD=2.12 PS=0.99 NRD=0 NRS=77.027
+ M=1 R=2.8 SA=75000.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_X_M1016_d N_A_1478_413#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_1606 A_193_47# 0 1.42804e-19 $X=0.965 $Y=0.235
*
.include "sky130_fd_sc_hd__mux4_1.pxi.spice"
*
.ends
*
*

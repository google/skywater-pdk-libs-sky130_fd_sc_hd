* File: sky130_fd_sc_hd__buf_6.pex.spice
* Created: Thu Aug 27 14:09:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUF_6%A 3 7 11 15 17 18 21 30
r51 28 30 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.15 $Y2=1.16
r52 26 28 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=0.73 $Y=1.16
+ $X2=1.02 $Y2=1.16
r53 21 26 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.73 $Y2=1.16
r54 21 23 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.545 $Y2=1.16
r55 18 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.02
+ $Y=1.16 $X2=1.02 $Y2=1.16
r56 17 18 24.0092 $w=2.38e-07 $l=5e-07 $layer=LI1_cond $X=0.475 $Y=1.195
+ $X2=0.975 $Y2=1.195
r57 17 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.545
+ $Y=1.16 $X2=0.545 $Y2=1.16
r58 13 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.16
r59 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.985
r60 9 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.15 $Y=1.025
+ $X2=1.15 $Y2=1.16
r61 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.15 $Y=1.025
+ $X2=1.15 $Y2=0.56
r62 5 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.73 $Y=1.295
+ $X2=0.73 $Y2=1.16
r63 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.73 $Y=1.295 $X2=0.73
+ $Y2=1.985
r64 1 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.73 $Y=1.025
+ $X2=0.73 $Y2=1.16
r65 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.73 $Y=1.025
+ $X2=0.73 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_6%A_161_47# 1 2 9 13 17 21 25 29 33 37 41 45 49
+ 53 57 59 61 63 64 65 68 70 73 78 86
c140 86 0 2.90279e-19 $X=3.67 $Y=1.16
r141 85 86 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.25 $Y=1.16
+ $X2=3.67 $Y2=1.16
r142 84 85 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.83 $Y=1.16
+ $X2=3.25 $Y2=1.16
r143 83 84 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.41 $Y=1.16
+ $X2=2.83 $Y2=1.16
r144 82 83 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.99 $Y=1.16
+ $X2=2.41 $Y2=1.16
r145 74 82 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=1.66 $Y=1.16
+ $X2=1.99 $Y2=1.16
r146 74 79 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.66 $Y=1.16 $X2=1.57
+ $Y2=1.16
r147 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.16 $X2=1.66 $Y2=1.16
r148 71 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=1.16
+ $X2=1.44 $Y2=1.16
r149 71 73 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.525 $Y=1.16
+ $X2=1.66 $Y2=1.16
r150 69 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=1.245
+ $X2=1.44 $Y2=1.16
r151 69 70 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.44 $Y=1.245
+ $X2=1.44 $Y2=1.485
r152 68 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=1.075
+ $X2=1.44 $Y2=1.16
r153 67 68 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.44 $Y=0.905
+ $X2=1.44 $Y2=1.075
r154 66 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=1.57
+ $X2=0.94 $Y2=1.57
r155 65 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.355 $Y=1.57
+ $X2=1.44 $Y2=1.485
r156 65 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.355 $Y=1.57
+ $X2=1.105 $Y2=1.57
r157 63 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.355 $Y=0.82
+ $X2=1.44 $Y2=0.905
r158 63 64 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.355 $Y=0.82
+ $X2=1.105 $Y2=0.82
r159 59 77 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=1.655
+ $X2=0.94 $Y2=1.57
r160 59 61 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.94 $Y=1.655
+ $X2=0.94 $Y2=2.31
r161 55 64 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.94 $Y=0.735
+ $X2=1.105 $Y2=0.82
r162 55 57 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.94 $Y=0.735
+ $X2=0.94 $Y2=0.38
r163 51 86 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.67 $Y=1.295
+ $X2=3.67 $Y2=1.16
r164 51 53 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.67 $Y=1.295
+ $X2=3.67 $Y2=1.985
r165 47 86 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.67 $Y=1.025
+ $X2=3.67 $Y2=1.16
r166 47 49 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.67 $Y=1.025
+ $X2=3.67 $Y2=0.56
r167 43 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.25 $Y=1.295
+ $X2=3.25 $Y2=1.16
r168 43 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.25 $Y=1.295
+ $X2=3.25 $Y2=1.985
r169 39 85 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.25 $Y=1.025
+ $X2=3.25 $Y2=1.16
r170 39 41 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.25 $Y=1.025
+ $X2=3.25 $Y2=0.56
r171 35 84 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.83 $Y=1.295
+ $X2=2.83 $Y2=1.16
r172 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.83 $Y=1.295
+ $X2=2.83 $Y2=1.985
r173 31 84 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.83 $Y=1.025
+ $X2=2.83 $Y2=1.16
r174 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.83 $Y=1.025
+ $X2=2.83 $Y2=0.56
r175 27 83 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.41 $Y=1.295
+ $X2=2.41 $Y2=1.16
r176 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.41 $Y=1.295
+ $X2=2.41 $Y2=1.985
r177 23 83 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.41 $Y=1.025
+ $X2=2.41 $Y2=1.16
r178 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.41 $Y=1.025
+ $X2=2.41 $Y2=0.56
r179 19 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.99 $Y=1.295
+ $X2=1.99 $Y2=1.16
r180 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.99 $Y=1.295
+ $X2=1.99 $Y2=1.985
r181 15 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.99 $Y=1.025
+ $X2=1.99 $Y2=1.16
r182 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.99 $Y=1.025
+ $X2=1.99 $Y2=0.56
r183 11 79 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.57 $Y=1.295
+ $X2=1.57 $Y2=1.16
r184 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.57 $Y=1.295
+ $X2=1.57 $Y2=1.985
r185 7 79 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.57 $Y=1.025
+ $X2=1.57 $Y2=1.16
r186 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.57 $Y=1.025
+ $X2=1.57 $Y2=0.56
r187 2 77 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.805
+ $Y=1.485 $X2=0.94 $Y2=1.63
r188 2 61 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.805
+ $Y=1.485 $X2=0.94 $Y2=2.31
r189 1 57 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.805
+ $Y=0.235 $X2=0.94 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_6%VPWR 1 2 3 4 5 18 24 26 30 34 36 38 43 44 45
+ 46 47 49 59 64 70 73 77
c71 30 0 1.4367e-19 $X=2.2 $Y=2
r72 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r74 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r75 68 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r76 68 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r77 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r78 65 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=3.04 $Y2=2.72
r79 65 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.205 $Y=2.72
+ $X2=3.45 $Y2=2.72
r80 64 76 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.927 $Y2=2.72
r81 64 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=2.72
+ $X2=3.45 $Y2=2.72
r82 63 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 63 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r84 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r85 60 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=2.72
+ $X2=2.2 $Y2=2.72
r86 60 62 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=2.72
+ $X2=2.53 $Y2=2.72
r87 59 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=3.04 $Y2=2.72
r88 59 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 58 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r90 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r91 49 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r92 47 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r93 45 57 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.275 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 45 46 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.275 $Y=2.72
+ $X2=1.395 $Y2=2.72
r95 43 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.23 $Y2=2.72
r96 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.52 $Y2=2.72
r97 42 57 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.52 $Y2=2.72
r99 38 41 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=1.66
+ $X2=3.88 $Y2=2.34
r100 36 76 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.927 $Y2=2.72
r101 36 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.88 $Y=2.635
+ $X2=3.88 $Y2=2.34
r102 32 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=2.635
+ $X2=3.04 $Y2=2.72
r103 32 34 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.04 $Y=2.635
+ $X2=3.04 $Y2=2
r104 28 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.635 $X2=2.2
+ $Y2=2.72
r105 28 30 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.2 $Y=2.635
+ $X2=2.2 $Y2=2
r106 27 46 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.395 $Y2=2.72
r107 26 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=2.72
+ $X2=2.2 $Y2=2.72
r108 26 27 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.035 $Y=2.72
+ $X2=1.515 $Y2=2.72
r109 22 46 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=2.635
+ $X2=1.395 $Y2=2.72
r110 22 24 30.4917 $w=2.38e-07 $l=6.35e-07 $layer=LI1_cond $X=1.395 $Y=2.635
+ $X2=1.395 $Y2=2
r111 18 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.52 $Y=1.66
+ $X2=0.52 $Y2=2.34
r112 16 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.52 $Y=2.635
+ $X2=0.52 $Y2=2.72
r113 16 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.52 $Y=2.635
+ $X2=0.52 $Y2=2.34
r114 5 41 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=2.34
r115 5 38 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=1.66
r116 4 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.905
+ $Y=1.485 $X2=3.04 $Y2=2
r117 3 30 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.065
+ $Y=1.485 $X2=2.2 $Y2=2
r118 2 24 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.225
+ $Y=1.485 $X2=1.36 $Y2=2
r119 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.485 $X2=0.52 $Y2=2.34
r120 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.485 $X2=0.52 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_6%X 1 2 3 4 5 6 21 25 29 33 37 41 43 44 45 61
r68 60 61 11.6455 $w=8.78e-07 $l=8.4e-07 $layer=LI1_cond $X=2.62 $Y=1.175
+ $X2=3.46 $Y2=1.175
r69 45 60 4.50568 $w=8.78e-07 $l=3.25e-07 $layer=LI1_cond $X=2.295 $Y=1.175
+ $X2=2.62 $Y2=1.175
r70 44 45 13.1335 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=1.865 $Y=1.53
+ $X2=2.21 $Y2=1.53
r71 43 45 14.1322 $w=3.08e-07 $l=3.45e-07 $layer=LI1_cond $X=1.865 $Y=0.82
+ $X2=2.21 $Y2=0.82
r72 39 61 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=3.46 $Y=1.615
+ $X2=3.46 $Y2=1.175
r73 39 41 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.46 $Y=1.615
+ $X2=3.46 $Y2=1.755
r74 35 61 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=3.46 $Y=0.735
+ $X2=3.46 $Y2=1.175
r75 35 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.46 $Y=0.735
+ $X2=3.46 $Y2=0.56
r76 31 60 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=2.62 $Y=1.615
+ $X2=2.62 $Y2=1.175
r77 31 33 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.62 $Y=1.615
+ $X2=2.62 $Y2=1.755
r78 27 60 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=2.62 $Y=0.735
+ $X2=2.62 $Y2=1.175
r79 27 29 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.62 $Y=0.735
+ $X2=2.62 $Y2=0.56
r80 23 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.78 $Y=1.615
+ $X2=1.865 $Y2=1.53
r81 23 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.78 $Y=1.615
+ $X2=1.78 $Y2=1.755
r82 19 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.78 $Y=0.735
+ $X2=1.865 $Y2=0.82
r83 19 21 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.78 $Y=0.735
+ $X2=1.78 $Y2=0.56
r84 6 41 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=1.485 $X2=3.46 $Y2=1.755
r85 5 33 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.485 $X2=2.62 $Y2=1.755
r86 4 25 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=1.645
+ $Y=1.485 $X2=1.78 $Y2=1.755
r87 3 37 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.46 $Y2=0.56
r88 2 29 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.62 $Y2=0.56
r89 1 21 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.78 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_6%VGND 1 2 3 4 5 18 22 24 28 32 34 36 39 40 41
+ 42 43 45 55 60 66 69 73
c77 28 0 1.46608e-19 $X=2.2 $Y=0.4
r78 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r79 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r80 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r81 64 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r82 64 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r83 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r84 61 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.04
+ $Y2=0
r85 61 63 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.45
+ $Y2=0
r86 60 72 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.927
+ $Y2=0
r87 60 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.45
+ $Y2=0
r88 59 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r89 59 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r90 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r91 56 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.2
+ $Y2=0
r92 56 58 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.53
+ $Y2=0
r93 55 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=3.04
+ $Y2=0
r94 55 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.53
+ $Y2=0
r95 54 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r96 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r97 45 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r98 43 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r99 41 53 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.15
+ $Y2=0
r100 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.36
+ $Y2=0
r101 39 43 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.435 $Y=0
+ $X2=0.23 $Y2=0
r102 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.52
+ $Y2=0
r103 38 53 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.605 $Y=0
+ $X2=1.15 $Y2=0
r104 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.52
+ $Y2=0
r105 34 72 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.927 $Y2=0
r106 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0.38
r107 30 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0
r108 30 32 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0.4
r109 26 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r110 26 28 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.2 $Y=0.085
+ $X2=2.2 $Y2=0.4
r111 25 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.36
+ $Y2=0
r112 24 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.2
+ $Y2=0
r113 24 25 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.445
+ $Y2=0
r114 20 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0
r115 20 22 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0.4
r116 16 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0
r117 16 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0.4
r118 5 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.38
r119 4 32 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.235 $X2=3.04 $Y2=0.4
r120 3 28 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.2 $Y2=0.4
r121 2 22 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.235 $X2=1.36 $Y2=0.4
r122 1 18 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.395
+ $Y=0.235 $X2=0.52 $Y2=0.4
.ends


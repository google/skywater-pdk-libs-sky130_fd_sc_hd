* File: sky130_fd_sc_hd__clkdlybuf4s15_1.spice
* Created: Tue Sep  1 19:00:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkdlybuf4s15_1.pex.spice"
.subckt sky130_fd_sc_hd__clkdlybuf4s15_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.174379 AS=0.1113 PD=1.06766 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_282_47#_M1007_d N_A_27_47#_M1007_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.65 AD=0.17225 AS=0.269871 PD=1.83 PS=1.65234 NRD=0 NRS=69.228 M=1
+ R=4.33333 SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_282_47#_M1005_g N_A_394_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.264981 AS=0.17225 PD=1.65234 PS=1.83 NRD=64.608 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_394_47#_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.171219 PD=1.37 PS=1.06766 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.38022 AS=0.265 PD=1.87912 PS=2.53 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1001 N_A_282_47#_M1001_d N_A_27_47#_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.82 AD=0.2173 AS=0.31178 PD=2.17 PS=1.54088 NRD=0 NRS=86.483 M=1 R=5.46667
+ SA=75001 SB=75000.2 A=0.123 P=1.94 MULT=1
MM1000 N_VPWR_M1000_d N_A_282_47#_M1000_g N_A_394_47#_M1000_s VPB PHIGHVT L=0.15
+ W=0.82 AD=0.306914 AS=0.2173 PD=1.54088 PS=2.17 NRD=84.0796 NRS=0 M=1
+ R=5.46667 SA=75000.2 SB=75001 A=0.123 P=1.94 MULT=1
MM1006 N_X_M1006_d N_A_394_47#_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.374286 PD=2.53 PS=1.87912 NRD=0 NRS=15.7403 M=1 R=6.66667
+ SA=75000.9 SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__clkdlybuf4s15_1.pxi.spice"
*
.ends
*
*

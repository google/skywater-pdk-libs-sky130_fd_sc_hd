* File: sky130_fd_sc_hd__lpflow_decapkapwr_4.pxi.spice
* Created: Thu Aug 27 14:24:36 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%VGND N_VGND_M1001_s VGND N_VGND_c_14_n
+ N_VGND_M1000_g N_VGND_c_15_n N_VGND_c_16_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%KAPWR N_KAPWR_M1000_s KAPWR
+ N_KAPWR_M1001_g N_KAPWR_c_26_n N_KAPWR_c_28_n N_KAPWR_c_29_n KAPWR
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%VPWR VPWR N_VPWR_c_40_n N_VPWR_c_39_n
+ PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_4%VPWR
cc_1 VNB N_VGND_c_14_n 0.0336337f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.29
cc_2 VNB N_VGND_c_15_n 0.115583f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=0.51
cc_3 VNB N_VGND_c_16_n 0.121884f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=0
cc_4 VNB N_KAPWR_M1001_g 0.151224f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=2.05
cc_5 VNB N_KAPWR_c_26_n 0.0137616f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=0.51
cc_6 VNB N_VPWR_c_39_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.775 $Y2=1.29
cc_7 VPB N_VGND_c_14_n 0.124937f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.29
cc_8 VPB N_VGND_c_15_n 0.00381416f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=0.51
cc_9 VPB N_KAPWR_c_26_n 0.0788122f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=0.51
cc_10 VPB N_KAPWR_c_28_n 0.0111567f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=0
cc_11 VPB N_KAPWR_c_29_n 0.0111567f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0
cc_12 VPB N_VPWR_c_40_n 0.0467232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_13 VPB N_VPWR_c_39_n 0.0419135f $X=-0.19 $Y=1.305 $X2=0.775 $Y2=1.29
cc_14 N_VGND_c_14_n N_KAPWR_M1001_g 0.0689775f $X=0.27 $Y=1.29 $X2=0 $Y2=0
cc_15 N_VGND_c_15_n N_KAPWR_M1001_g 0.142049f $X=1.58 $Y=0.51 $X2=0 $Y2=0
cc_16 N_VGND_c_14_n N_KAPWR_c_26_n 0.142595f $X=0.27 $Y=1.29 $X2=0 $Y2=0
cc_17 N_VGND_c_15_n N_KAPWR_c_26_n 0.16291f $X=1.58 $Y=0.51 $X2=0 $Y2=0
cc_18 N_VGND_c_14_n N_VPWR_c_40_n 0.0250367f $X=0.27 $Y=1.29 $X2=0 $Y2=0
cc_19 N_VGND_c_14_n N_VPWR_c_39_n 0.024908f $X=0.27 $Y=1.29 $X2=0 $Y2=0
cc_20 N_KAPWR_c_26_n N_VPWR_c_40_n 0.111288f $X=1.58 $Y=1.83 $X2=0 $Y2=0
cc_21 N_KAPWR_c_29_n N_VPWR_c_40_n 0.00121403f $X=0.215 $Y=2.21 $X2=0 $Y2=0
cc_22 N_KAPWR_M1000_s N_VPWR_c_39_n 0.0021408f $X=0.135 $Y=1.615 $X2=0 $Y2=0
cc_23 N_KAPWR_c_26_n N_VPWR_c_39_n 0.0143371f $X=1.58 $Y=1.83 $X2=0 $Y2=0
cc_24 N_KAPWR_c_29_n N_VPWR_c_39_n 0.173995f $X=0.215 $Y=2.21 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__dlymetal6s4s_1.spice.pex
* Created: Thu Aug 27 14:19:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%A 3 7 9 10 15 17
c31 17 0 1.57226e-19 $X=0.645 $Y=1.16
r32 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.42 $Y=1.16
+ $X2=0.645 $Y2=1.16
r33 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=1.16 $X2=0.42 $Y2=1.16
r34 9 10 8.38488 $w=4.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.327 $Y=1.19
+ $X2=0.327 $Y2=1.53
r35 9 15 0.739842 $w=4.83e-07 $l=3e-08 $layer=LI1_cond $X=0.327 $Y=1.19
+ $X2=0.327 $Y2=1.16
r36 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=1.325
+ $X2=0.645 $Y2=1.16
r37 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.645 $Y=1.325
+ $X2=0.645 $Y2=2.275
r38 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=0.995
+ $X2=0.645 $Y2=1.16
r39 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.645 $Y=0.995
+ $X2=0.645 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%A_62_47# 1 2 9 12 14 16 21 23 27 33
+ 34 35 38
c60 33 0 1.1704e-19 $X=1.065 $Y=1.16
c61 16 0 1.57226e-19 $X=0.74 $Y=1.955
r62 34 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.16
+ $X2=1.065 $Y2=1.325
r63 34 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.16
+ $X2=1.065 $Y2=0.995
r64 33 36 5.05753 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.16
+ $X2=0.945 $Y2=1.325
r65 33 35 5.05753 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.16
+ $X2=0.945 $Y2=0.995
r66 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.065
+ $Y=1.16 $X2=1.065 $Y2=1.16
r67 27 30 8.47774 $w=4.33e-07 $l=3.2e-07 $layer=LI1_cond $X=0.302 $Y=1.955
+ $X2=0.302 $Y2=2.275
r68 23 25 7.81542 $w=4.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.302 $Y=0.445
+ $X2=0.302 $Y2=0.74
r69 21 36 18.7487 $w=3.33e-07 $l=5.45e-07 $layer=LI1_cond $X=0.907 $Y=1.87
+ $X2=0.907 $Y2=1.325
r70 18 35 5.84822 $w=3.33e-07 $l=1.7e-07 $layer=LI1_cond $X=0.907 $Y=0.825
+ $X2=0.907 $Y2=0.995
r71 17 27 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.52 $Y=1.955
+ $X2=0.302 $Y2=1.955
r72 16 21 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=0.74 $Y=1.955
+ $X2=0.907 $Y2=1.87
r73 16 17 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.74 $Y=1.955
+ $X2=0.52 $Y2=1.955
r74 15 25 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.52 $Y=0.74
+ $X2=0.302 $Y2=0.74
r75 14 18 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=0.74 $Y=0.74
+ $X2=0.907 $Y2=0.825
r76 14 15 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.74 $Y=0.74
+ $X2=0.52 $Y2=0.74
r77 12 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.12 $Y=1.985
+ $X2=1.12 $Y2=1.325
r78 9 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.12 $Y=0.56 $X2=1.12
+ $Y2=0.995
r79 2 30 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.31
+ $Y=2.065 $X2=0.435 $Y2=2.275
r80 1 23 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.235 $X2=0.435 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%A_239_47# 1 2 9 13 17 19 21 24 25 31
r55 28 31 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.835 $Y=1.16
+ $X2=2.06 $Y2=1.16
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=1.16 $X2=1.835 $Y2=1.16
r57 24 27 9.80533 $w=6.69e-07 $l=2.59711e-07 $layer=LI1_cond $X=1.417 $Y=0.995
+ $X2=1.607 $Y2=1.16
r58 24 25 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=1.417 $Y=0.995
+ $X2=1.417 $Y2=0.825
r59 19 27 13.8675 $w=6.69e-07 $l=6.18167e-07 $layer=LI1_cond $X=1.38 $Y=1.675
+ $X2=1.607 $Y2=1.16
r60 19 21 12.1647 $w=2.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.38 $Y=1.675
+ $X2=1.38 $Y2=1.96
r61 15 25 6.67067 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.38 $Y=0.69
+ $X2=1.38 $Y2=0.825
r62 15 17 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.38 $Y=0.69
+ $X2=1.38 $Y2=0.44
r63 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.325
+ $X2=2.06 $Y2=1.16
r64 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.06 $Y=1.325
+ $X2=2.06 $Y2=2.275
r65 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=0.995
+ $X2=2.06 $Y2=1.16
r66 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.06 $Y=0.995 $X2=2.06
+ $Y2=0.445
r67 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.195
+ $Y=1.485 $X2=1.33 $Y2=1.96
r68 1 17 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.235 $X2=1.33 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%A_345_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c67 26 0 1.27733e-19 $X=2.315 $Y=1.325
r68 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.48 $Y=1.16
+ $X2=2.48 $Y2=1.325
r69 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.48 $Y=1.16
+ $X2=2.48 $Y2=0.995
r70 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.16 $X2=2.48 $Y2=1.16
r71 28 30 13.2746 $w=3.86e-07 $l=4.2e-07 $layer=LI1_cond $X=2.352 $Y=0.74
+ $X2=2.352 $Y2=1.16
r72 26 30 5.34605 $w=3.86e-07 $l=1.82565e-07 $layer=LI1_cond $X=2.315 $Y=1.325
+ $X2=2.352 $Y2=1.16
r73 26 27 17.122 $w=3.48e-07 $l=5.2e-07 $layer=LI1_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.845
r74 24 27 7.55928 $w=1.95e-07 $l=2.18174e-07 $layer=LI1_cond $X=2.14 $Y=1.942
+ $X2=2.315 $Y2=1.845
r75 24 25 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=2.14 $Y=1.942
+ $X2=1.935 $Y2=1.942
r76 22 28 5.5624 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.14 $Y=0.74
+ $X2=2.352 $Y2=0.74
r77 22 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.14 $Y=0.74
+ $X2=1.935 $Y2=0.74
r78 18 25 6.9528 $w=1.95e-07 $l=1.66958e-07 $layer=LI1_cond $X=1.81 $Y=2.04
+ $X2=1.935 $Y2=1.942
r79 18 20 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=1.81 $Y=2.04
+ $X2=1.81 $Y2=2.275
r80 14 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.81 $Y=0.655
+ $X2=1.935 $Y2=0.74
r81 14 16 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.81 $Y=0.655
+ $X2=1.81 $Y2=0.44
r82 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.535 $Y=1.985
+ $X2=2.535 $Y2=1.325
r83 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.535 $Y=0.56
+ $X2=2.535 $Y2=0.995
r84 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=2.065 $X2=1.85 $Y2=2.275
r85 1 16 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.235 $X2=1.85 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%X 1 2 9 13 15 16 17 18 19 20 21 22 35
+ 37
r48 32 35 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.43 $Y=1.16
+ $X2=3.655 $Y2=1.16
r49 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.16 $X2=3.43 $Y2=1.16
r50 20 41 6.4744 $w=4.43e-07 $l=2.5e-07 $layer=LI1_cond $X=2.882 $Y=2.21
+ $X2=2.882 $Y2=1.96
r51 19 41 2.33078 $w=4.43e-07 $l=9e-08 $layer=LI1_cond $X=2.882 $Y=1.87
+ $X2=2.882 $Y2=1.96
r52 19 37 5.05003 $w=4.43e-07 $l=1.95e-07 $layer=LI1_cond $X=2.882 $Y=1.87
+ $X2=2.882 $Y2=1.675
r53 18 37 3.87245 $w=6.29e-07 $l=2.86468e-07 $layer=LI1_cond $X=3.105 $Y=1.53
+ $X2=2.882 $Y2=1.675
r54 18 22 8.62214 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=3.105 $Y=1.53
+ $X2=3.445 $Y2=1.53
r55 17 18 6.59459 $w=6.29e-07 $l=3.4e-07 $layer=LI1_cond $X=3.105 $Y=1.19
+ $X2=3.105 $Y2=1.53
r56 17 21 8.62214 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=3.105 $Y=1.19
+ $X2=3.445 $Y2=1.19
r57 17 33 0.581876 $w=6.29e-07 $l=3e-08 $layer=LI1_cond $X=3.105 $Y=1.19
+ $X2=3.105 $Y2=1.16
r58 16 33 6.01272 $w=6.29e-07 $l=3.1e-07 $layer=LI1_cond $X=3.105 $Y=0.85
+ $X2=3.105 $Y2=1.16
r59 15 16 6.59459 $w=6.29e-07 $l=3.4e-07 $layer=LI1_cond $X=3.105 $Y=0.51
+ $X2=3.105 $Y2=0.85
r60 15 46 1.35771 $w=6.29e-07 $l=7e-08 $layer=LI1_cond $X=3.105 $Y=0.51
+ $X2=3.105 $Y2=0.44
r61 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.325
+ $X2=3.655 $Y2=1.16
r62 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.655 $Y=1.325
+ $X2=3.655 $Y2=2.275
r63 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=0.995
+ $X2=3.655 $Y2=1.16
r64 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.655 $Y=0.995
+ $X2=3.655 $Y2=0.445
r65 2 41 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.61
+ $Y=1.485 $X2=2.745 $Y2=1.96
r66 1 46 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=2.61
+ $Y=0.235 $X2=2.745 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%A_664_47# 1 2 9 12 16 20 22 23 24 25
+ 26 27 31 33
c64 26 0 1.27733e-19 $X=3.91 $Y=1.325
r65 31 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.16
+ $X2=4.075 $Y2=1.325
r66 31 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.16
+ $X2=4.075 $Y2=0.995
r67 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.075
+ $Y=1.16 $X2=4.075 $Y2=1.16
r68 28 30 13.2746 $w=3.86e-07 $l=4.2e-07 $layer=LI1_cond $X=3.947 $Y=0.74
+ $X2=3.947 $Y2=1.16
r69 26 30 5.34605 $w=3.86e-07 $l=1.82565e-07 $layer=LI1_cond $X=3.91 $Y=1.325
+ $X2=3.947 $Y2=1.16
r70 26 27 17.122 $w=3.48e-07 $l=5.2e-07 $layer=LI1_cond $X=3.91 $Y=1.325
+ $X2=3.91 $Y2=1.845
r71 24 27 7.55928 $w=1.95e-07 $l=2.18174e-07 $layer=LI1_cond $X=3.735 $Y=1.942
+ $X2=3.91 $Y2=1.845
r72 24 25 11.6597 $w=1.93e-07 $l=2.05e-07 $layer=LI1_cond $X=3.735 $Y=1.942
+ $X2=3.53 $Y2=1.942
r73 22 28 5.5624 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.735 $Y=0.74
+ $X2=3.947 $Y2=0.74
r74 22 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.735 $Y=0.74
+ $X2=3.53 $Y2=0.74
r75 18 25 6.9753 $w=1.95e-07 $l=1.70082e-07 $layer=LI1_cond $X=3.402 $Y=2.04
+ $X2=3.53 $Y2=1.942
r76 18 20 10.6206 $w=2.53e-07 $l=2.35e-07 $layer=LI1_cond $X=3.402 $Y=2.04
+ $X2=3.402 $Y2=2.275
r77 14 23 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=3.402 $Y=0.655
+ $X2=3.53 $Y2=0.74
r78 14 16 9.71668 $w=2.53e-07 $l=2.15e-07 $layer=LI1_cond $X=3.402 $Y=0.655
+ $X2=3.402 $Y2=0.44
r79 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.13 $Y=1.985
+ $X2=4.13 $Y2=1.325
r80 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.56 $X2=4.13
+ $Y2=0.995
r81 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=2.065 $X2=3.445 $Y2=2.275
r82 1 16 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.235 $X2=3.445 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%VPWR 1 2 3 14 18 22 25 26 27 36 45 46
+ 49 52 57
r62 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 50 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 46 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r66 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r67 43 52 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=3.892 $Y2=2.72
r68 43 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=2.72
+ $X2=4.37 $Y2=2.72
r69 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r71 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r73 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r74 36 52 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.7 $Y=2.72
+ $X2=3.892 $Y2=2.72
r75 36 41 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.45
+ $Y2=2.72
r76 35 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r77 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r78 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r79 32 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 31 34 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r81 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r82 29 49 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=0.882 $Y2=2.72
r83 29 31 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=1.15 $Y2=2.72
r84 27 57 0.00711354 $w=4.8e-07 $l=2.5e-08 $layer=MET1_cond $X=0.205 $Y=2.72
+ $X2=0.23 $Y2=2.72
r85 25 34 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r86 25 26 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.297 $Y2=2.72
r87 24 38 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.49 $Y=2.72 $X2=2.53
+ $Y2=2.72
r88 24 26 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.49 $Y=2.72
+ $X2=2.297 $Y2=2.72
r89 20 52 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.892 $Y2=2.72
r90 20 22 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.892 $Y2=2.36
r91 16 26 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.297 $Y=2.635
+ $X2=2.297 $Y2=2.72
r92 16 18 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=2.297 $Y=2.635
+ $X2=2.297 $Y2=2.36
r93 12 49 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.882 $Y=2.635
+ $X2=0.882 $Y2=2.72
r94 12 14 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=0.882 $Y=2.635
+ $X2=0.882 $Y2=2.36
r95 3 22 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=2.065 $X2=3.895 $Y2=2.36
r96 2 18 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=2.065 $X2=2.3 $Y2=2.36
r97 1 14 600 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=2.065 $X2=0.885 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%A_841_47# 1 2 9 11 13 17 18
r17 17 18 40.1671 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=4.422 $Y=0.825
+ $X2=4.422 $Y2=1.495
r18 11 18 6.73749 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=4.385 $Y=1.625
+ $X2=4.385 $Y2=1.495
r19 11 13 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=4.385 $Y=1.625
+ $X2=4.385 $Y2=1.96
r20 7 17 6.73749 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=4.385 $Y=0.695
+ $X2=4.385 $Y2=0.825
r21 7 9 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=4.385 $Y=0.695
+ $X2=4.385 $Y2=0.44
r22 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.205
+ $Y=1.485 $X2=4.34 $Y2=1.96
r23 1 9 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.235 $X2=4.34 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HD__DLYMETAL6S4S_1%VGND 1 2 3 14 18 22 25 26 27 36 45 46
+ 49 52 57
r65 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r66 50 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r67 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r68 46 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r69 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r70 43 52 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=3.892
+ $Y2=0
r71 43 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.37
+ $Y2=0
r72 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r73 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r74 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r75 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r76 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r77 36 52 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.892
+ $Y2=0
r78 36 41 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.45
+ $Y2=0
r79 35 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r80 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r81 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r82 32 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r83 31 34 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r84 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r85 29 49 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.882
+ $Y2=0
r86 29 31 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.15
+ $Y2=0
r87 27 57 0.00711354 $w=4.8e-07 $l=2.5e-08 $layer=MET1_cond $X=0.205 $Y=0
+ $X2=0.23 $Y2=0
r88 25 34 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.07
+ $Y2=0
r89 25 26 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.297
+ $Y2=0
r90 24 38 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.49 $Y=0 $X2=2.53
+ $Y2=0
r91 24 26 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.49 $Y=0 $X2=2.297
+ $Y2=0
r92 20 52 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.892 $Y2=0
r93 20 22 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.892 $Y2=0.38
r94 16 26 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.297 $Y=0.085
+ $X2=2.297 $Y2=0
r95 16 18 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=2.297 $Y=0.085
+ $X2=2.297 $Y2=0.38
r96 12 49 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.882 $Y=0.085
+ $X2=0.882 $Y2=0
r97 12 14 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.882 $Y=0.085
+ $X2=0.882 $Y2=0.38
r98 3 22 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.89 $Y2=0.38
r99 2 18 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.235 $X2=2.295 $Y2=0.38
r100 1 14 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.72
+ $Y=0.235 $X2=0.88 $Y2=0.38
.ends


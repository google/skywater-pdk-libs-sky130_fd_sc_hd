* File: sky130_fd_sc_hd__fahcon_1.spice.pex
* Created: Thu Aug 27 14:21:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_67_199# 1 2 3 4 5 18 21 23 24 25 27 28 29
+ 32 33 37 39 44 47 55 56 59 62 63 66
c175 44 0 3.27481e-19 $X=0.51 $Y=1.16
r176 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.295 $Y=1.87
+ $X2=4.295 $Y2=1.87
r177 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.365 $Y=1.87
+ $X2=1.365 $Y2=1.87
r178 56 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.51 $Y=1.87
+ $X2=1.365 $Y2=1.87
r179 55 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.15 $Y=1.87
+ $X2=4.295 $Y2=1.87
r180 55 56 3.26732 $w=1.4e-07 $l=2.64e-06 $layer=MET1_cond $X=4.15 $Y=1.87
+ $X2=1.51 $Y2=1.87
r181 50 59 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.365 $Y=1.875
+ $X2=1.365 $Y2=1.87
r182 47 59 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.365 $Y=1.67
+ $X2=1.365 $Y2=1.87
r183 47 49 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=1.67
+ $X2=1.365 $Y2=1.585
r184 44 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.16
+ $X2=0.5 $Y2=1.325
r185 44 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.16
+ $X2=0.5 $Y2=0.995
r186 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r187 37 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=1.96
+ $X2=1.365 $Y2=1.875
r188 37 39 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=1.45 $Y=1.96
+ $X2=2.725 $Y2=1.96
r189 34 46 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=0.36
+ $X2=1.16 $Y2=0.36
r190 34 36 29.5758 $w=2.08e-07 $l=5.6e-07 $layer=LI1_cond $X=1.325 $Y=0.36
+ $X2=1.885 $Y2=0.36
r191 33 36 71.5628 $w=2.08e-07 $l=1.355e-06 $layer=LI1_cond $X=3.24 $Y=0.36
+ $X2=1.885 $Y2=0.36
r192 30 32 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.16 $Y=0.735
+ $X2=1.16 $Y2=0.72
r193 29 46 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.36
r194 29 32 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.72
r195 27 49 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.585
+ $X2=1.365 $Y2=1.585
r196 27 28 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.28 $Y=1.585
+ $X2=0.78 $Y2=1.585
r197 26 43 15.1941 $w=2.73e-07 $l=4.19667e-07 $layer=LI1_cond $X=0.78 $Y=0.82
+ $X2=0.602 $Y2=1.16
r198 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.995 $Y=0.82
+ $X2=1.16 $Y2=0.735
r199 25 26 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.995 $Y=0.82
+ $X2=0.78 $Y2=0.82
r200 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.695 $Y=1.5
+ $X2=0.78 $Y2=1.585
r201 23 43 9.1003 $w=2.73e-07 $l=2.06325e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.602 $Y2=1.16
r202 23 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.695 $Y2=1.5
r203 21 67 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.325
r204 18 66 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.475 $Y=0.555
+ $X2=0.475 $Y2=0.995
r205 5 63 600 $w=1.7e-07 $l=3.81576e-07 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.61 $X2=4.295 $Y2=1.93
r206 4 39 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.725 $Y2=1.96
r207 3 49 600 $w=1.7e-07 $l=3.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.485 $X2=1.365 $Y2=1.665
r208 2 33 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.235 $X2=3.325 $Y2=0.42
r209 1 46 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.16 $Y2=0.38
r210 1 36 182 $w=1.7e-07 $l=9.29677e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.885 $Y2=0.38
r211 1 32 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.16 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A 1 3 6 8 14
c44 8 0 1.76755e-19 $X=1.15 $Y=1.19
c45 1 0 5.07203e-20 $X=0.95 $Y=0.995
r46 12 14 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.975 $Y=1.16
+ $X2=1.175 $Y2=1.16
r47 10 12 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.975 $Y2=1.16
r48 8 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=1.16 $X2=1.175 $Y2=1.16
r49 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.16
r50 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.985
r51 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=1.16
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.95 $Y=0.995 $X2=0.95
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%B 1 3 6 10 14 17 19 21 22 24 26 29 31 32 34
+ 35 37 38 39 40 42 43 45 51 52
c179 52 0 1.03294e-19 $X=4.395 $Y=0.85
c180 40 0 1.31043e-19 $X=1.61 $Y=0.85
c181 32 0 1.94707e-19 $X=2.095 $Y=1.16
c182 10 0 1.51029e-19 $X=4.085 $Y=2.03
r183 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.35
+ $Y=1.16 $X2=4.35 $Y2=1.16
r184 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.16 $X2=1.655 $Y2=1.16
r185 52 60 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=4.39 $Y=0.85
+ $X2=4.39 $Y2=1.16
r186 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.395 $Y=0.85
+ $X2=4.395 $Y2=0.85
r187 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=0.85
+ $X2=1.61 $Y2=0.85
r188 42 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.25 $Y=0.85
+ $X2=4.395 $Y2=0.85
r189 42 43 3.08787 $w=1.4e-07 $l=2.495e-06 $layer=MET1_cond $X=4.25 $Y=0.85
+ $X2=1.755 $Y2=0.85
r190 40 56 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.645 $Y=0.85
+ $X2=1.645 $Y2=1.16
r191 40 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0.85
+ $X2=1.61 $Y2=0.85
r192 37 59 124.152 $w=3.3e-07 $l=7.1e-07 $layer=POLY_cond $X=5.06 $Y=1.16
+ $X2=4.35 $Y2=1.16
r193 37 38 4.10278 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.06 $Y=1.16
+ $X2=5.145 $Y2=1.16
r194 34 59 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.295 $Y=1.16
+ $X2=4.35 $Y2=1.16
r195 34 36 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=4.152 $Y=1.16
+ $X2=4.152 $Y2=1.325
r196 34 35 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=4.152 $Y=1.16
+ $X2=4.152 $Y2=0.995
r197 31 55 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.02 $Y=1.16
+ $X2=1.655 $Y2=1.16
r198 31 32 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.02 $Y=1.16
+ $X2=2.095 $Y2=1.16
r199 27 39 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.645 $Y=1.325
+ $X2=5.645 $Y2=1.16
r200 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.645 $Y=1.325
+ $X2=5.645 $Y2=1.985
r201 24 39 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.645 $Y=0.995
+ $X2=5.645 $Y2=1.16
r202 24 26 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.645 $Y=0.995
+ $X2=5.645 $Y2=0.565
r203 23 38 4.10278 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.23 $Y=1.16
+ $X2=5.145 $Y2=1.16
r204 22 39 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.57 $Y=1.16
+ $X2=5.645 $Y2=1.16
r205 22 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.57 $Y=1.16
+ $X2=5.23 $Y2=1.16
r206 19 38 22.6206 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=5.155 $Y=0.995
+ $X2=5.145 $Y2=1.16
r207 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.155 $Y=0.995
+ $X2=5.155 $Y2=0.56
r208 15 38 22.6206 $w=1.5e-07 $l=1.69926e-07 $layer=POLY_cond $X=5.135 $Y=1.325
+ $X2=5.145 $Y2=1.16
r209 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.135 $Y=1.325
+ $X2=5.135 $Y2=1.985
r210 14 35 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.22 $Y=0.565
+ $X2=4.22 $Y2=0.995
r211 10 36 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=4.085 $Y=2.03
+ $X2=4.085 $Y2=1.325
r212 4 32 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.325
+ $X2=2.095 $Y2=1.16
r213 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.095 $Y=1.325
+ $X2=2.095 $Y2=1.905
r214 1 32 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.095 $Y2=1.16
r215 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.095 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_488_21# 1 2 7 9 12 14 16 19 22 23 24 27
+ 29 32 33 39 40 44 48
c120 44 0 1.94707e-19 $X=2.81 $Y=1.16
c121 24 0 1.61409e-19 $X=3.582 $Y=1.16
c122 22 0 1.31043e-19 $X=2.515 $Y=1.16
c123 14 0 4.61014e-20 $X=3.555 $Y=0.995
r124 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=1.16 $X2=2.81 $Y2=1.16
r125 40 48 4.64666 $w=4.78e-07 $l=1.45e-07 $layer=LI1_cond $X=4.94 $Y=1.53
+ $X2=4.94 $Y2=1.385
r126 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.855 $Y=1.53
+ $X2=4.855 $Y2=1.53
r127 36 44 10.2591 $w=4.4e-07 $l=3.7e-07 $layer=LI1_cond $X=2.87 $Y=1.53
+ $X2=2.87 $Y2=1.16
r128 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.53
+ $X2=3.015 $Y2=1.53
r129 33 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.16 $Y=1.53
+ $X2=3.015 $Y2=1.53
r130 32 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.71 $Y=1.53
+ $X2=4.855 $Y2=1.53
r131 32 33 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=4.71 $Y=1.53
+ $X2=3.16 $Y2=1.53
r132 29 31 7.98749 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=5.01 $Y=1.165
+ $X2=5.01 $Y2=0.995
r133 29 48 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=5.01 $Y=1.165
+ $X2=5.01 $Y2=1.385
r134 27 31 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=4.935 $Y=0.73
+ $X2=4.935 $Y2=0.995
r135 23 43 117.157 $w=3.3e-07 $l=6.7e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=2.81 $Y2=1.16
r136 23 24 5.03009 $w=3.3e-07 $l=1.02e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=3.582 $Y2=1.16
r137 21 43 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.81 $Y2=1.16
r138 21 22 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=2.515 $Y2=1.16
r139 17 24 37.0704 $w=1.5e-07 $l=1.73767e-07 $layer=POLY_cond $X=3.6 $Y=1.325
+ $X2=3.582 $Y2=1.16
r140 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.6 $Y=1.325
+ $X2=3.6 $Y2=1.905
r141 14 24 37.0704 $w=1.5e-07 $l=1.77989e-07 $layer=POLY_cond $X=3.555 $Y=0.995
+ $X2=3.582 $Y2=1.16
r142 14 16 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.555 $Y=0.995
+ $X2=3.555 $Y2=0.555
r143 10 22 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=1.325
+ $X2=2.515 $Y2=1.16
r144 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.515 $Y=1.325
+ $X2=2.515 $Y2=1.905
r145 7 22 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.515 $Y2=1.16
r146 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.515 $Y2=0.565
r147 2 40 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=1.485 $X2=4.925 $Y2=1.64
r148 1 27 182 $w=1.7e-07 $l=1.76777e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.605 $X2=4.945 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_434_49# 1 2 9 11 13 16 19 21 22 23 24 31
+ 33 41 44 45 46 49
c176 41 0 2.59669e-19 $X=6.64 $Y=1.16
c177 33 0 3.03414e-19 $X=8.995 $Y=1.19
c178 11 0 1.78045e-19 $X=6.64 $Y=0.995
c179 2 0 8.07134e-20 $X=2.17 $Y=1.485
r180 44 47 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.96 $Y=1.16
+ $X2=8.96 $Y2=1.325
r181 44 46 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.96 $Y=1.16
+ $X2=8.96 $Y2=0.995
r182 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.945
+ $Y=1.16 $X2=8.945 $Y2=1.16
r183 40 41 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.585 $Y=1.16
+ $X2=6.64 $Y2=1.16
r184 37 40 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=6.35 $Y=1.16
+ $X2=6.585 $Y2=1.16
r185 33 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.995 $Y=1.19
+ $X2=8.995 $Y2=1.19
r186 31 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.35
+ $Y=1.16 $X2=6.35 $Y2=1.16
r187 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.235 $Y=1.19
+ $X2=6.235 $Y2=1.19
r188 27 53 10.1844 $w=5.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.217 $Y=1.19
+ $X2=2.217 $Y2=1.62
r189 27 49 11.1318 $w=5.03e-07 $l=4.7e-07 $layer=LI1_cond $X=2.217 $Y=1.19
+ $X2=2.217 $Y2=0.72
r190 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=1.19
+ $X2=2.07 $Y2=1.19
r191 24 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.38 $Y=1.19
+ $X2=6.235 $Y2=1.19
r192 23 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.85 $Y=1.19
+ $X2=8.995 $Y2=1.19
r193 23 24 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=8.85 $Y=1.19
+ $X2=6.38 $Y2=1.19
r194 22 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.215 $Y=1.19
+ $X2=2.07 $Y2=1.19
r195 21 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.09 $Y=1.19
+ $X2=6.235 $Y2=1.19
r196 21 22 4.79578 $w=1.4e-07 $l=3.875e-06 $layer=MET1_cond $X=6.09 $Y=1.19
+ $X2=2.215 $Y2=1.19
r197 19 47 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.945 $Y=1.995
+ $X2=8.945 $Y2=1.325
r198 16 46 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.915 $Y=0.565
+ $X2=8.915 $Y2=0.995
r199 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.64 $Y=0.995
+ $X2=6.64 $Y2=1.16
r200 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.64 $Y=0.995
+ $X2=6.64 $Y2=0.565
r201 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.585 $Y=1.325
+ $X2=6.585 $Y2=1.16
r202 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.585 $Y=1.325
+ $X2=6.585 $Y2=1.905
r203 2 53 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.17
+ $Y=1.485 $X2=2.305 $Y2=1.62
r204 1 49 182 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.245 $X2=2.305 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_726_47# 1 2 9 11 13 14 16 17 19 21 22 23
+ 28 29 30 33 36 37 38 40 41 42 44 47 52 55
c191 28 0 5.81156e-20 $X=3.81 $Y=1.7
c192 9 0 1.73441e-19 $X=7.005 $Y=1.905
r193 54 55 7.68295 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=7.917 $Y=1.55
+ $X2=7.917 $Y2=1.72
r194 50 52 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.81 $Y=1.235
+ $X2=4.01 $Y2=1.235
r195 47 54 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.96 $Y=1.16
+ $X2=7.96 $Y2=1.55
r196 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.96
+ $Y=1.16 $X2=7.96 $Y2=1.16
r197 44 55 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.875 $Y=2.295
+ $X2=7.875 $Y2=1.72
r198 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.79 $Y=2.38
+ $X2=7.875 $Y2=2.295
r199 41 42 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=7.79 $Y=2.38
+ $X2=6.005 $Y2=2.38
r200 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.92 $Y=2.295
+ $X2=6.005 $Y2=2.38
r201 39 40 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.92 $Y=2.065
+ $X2=5.92 $Y2=2.295
r202 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.835 $Y=1.98
+ $X2=5.92 $Y2=2.065
r203 37 38 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.835 $Y=1.98
+ $X2=5.1 $Y2=1.98
r204 35 38 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=4.987 $Y=2.065
+ $X2=5.1 $Y2=1.98
r205 35 36 11.7805 $w=2.23e-07 $l=2.3e-07 $layer=LI1_cond $X=4.987 $Y=2.065
+ $X2=4.987 $Y2=2.295
r206 31 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.01 $Y=1.15
+ $X2=4.01 $Y2=1.235
r207 31 33 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.01 $Y=1.15
+ $X2=4.01 $Y2=0.76
r208 29 36 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.875 $Y=2.38
+ $X2=4.987 $Y2=2.295
r209 29 30 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.875 $Y=2.38
+ $X2=3.895 $Y2=2.38
r210 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=2.295
+ $X2=3.895 $Y2=2.38
r211 26 28 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.81 $Y=2.295
+ $X2=3.81 $Y2=1.7
r212 25 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=1.32
+ $X2=3.81 $Y2=1.235
r213 25 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.81 $Y=1.32
+ $X2=3.81 $Y2=1.7
r214 23 24 5.07368 $w=4.75e-07 $l=5e-08 $layer=POLY_cond $X=8.475 $Y=1.247
+ $X2=8.525 $Y2=1.247
r215 22 48 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=8.005 $Y=1.16
+ $X2=7.96 $Y2=1.16
r216 22 23 52.2322 $w=4.75e-07 $l=5.11654e-07 $layer=POLY_cond $X=8.005 $Y=1.16
+ $X2=8.475 $Y2=1.247
r217 20 48 143.386 $w=3.3e-07 $l=8.2e-07 $layer=POLY_cond $X=7.14 $Y=1.16
+ $X2=7.96 $Y2=1.16
r218 20 21 5.03009 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=7.14 $Y=1.16
+ $X2=7.035 $Y2=1.16
r219 17 24 30.117 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=8.525 $Y=1.5
+ $X2=8.525 $Y2=1.247
r220 17 19 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.525 $Y=1.5
+ $X2=8.525 $Y2=1.995
r221 14 23 30.117 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=8.475 $Y=0.995
+ $X2=8.475 $Y2=1.247
r222 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.475 $Y=0.995
+ $X2=8.475 $Y2=0.565
r223 11 21 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=7.065 $Y=0.995
+ $X2=7.035 $Y2=1.16
r224 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.065 $Y=0.995
+ $X2=7.065 $Y2=0.565
r225 7 21 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=7.005 $Y=1.325
+ $X2=7.035 $Y2=1.16
r226 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.005 $Y=1.325
+ $X2=7.005 $Y2=1.905
r227 2 28 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.485 $X2=3.81 $Y2=1.7
r228 1 33 182 $w=1.7e-07 $l=6.89293e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.235 $X2=4.01 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_1589_49# 1 2 3 4 15 18 22 25 26 30 32 34
+ 37 38 39 45 49 51 53
c148 49 0 1.96825e-19 $X=10.075 $Y=1.16
c149 32 0 1.49929e-19 $X=10.73 $Y=2.045
r150 50 57 12.9309 $w=4.34e-07 $l=4.6e-07 $layer=LI1_cond $X=10.36 $Y=1.16
+ $X2=10.36 $Y2=1.62
r151 49 51 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.075 $Y=1.16
+ $X2=10.075 $Y2=0.995
r152 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.075
+ $Y=1.16 $X2=10.075 $Y2=1.16
r153 46 57 7.02765 $w=4.34e-07 $l=2.5e-07 $layer=LI1_cond $X=10.36 $Y=1.87
+ $X2=10.36 $Y2=1.62
r154 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.275 $Y=1.87
+ $X2=10.275 $Y2=1.87
r155 41 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.365 $Y=1.87
+ $X2=9.365 $Y2=1.87
r156 39 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.51 $Y=1.87
+ $X2=9.365 $Y2=1.87
r157 38 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.13 $Y=1.87
+ $X2=10.275 $Y2=1.87
r158 38 39 0.767325 $w=1.4e-07 $l=6.2e-07 $layer=MET1_cond $X=10.13 $Y=1.87
+ $X2=9.51 $Y2=1.87
r159 32 46 8.17867 $w=4.34e-07 $l=4.49055e-07 $layer=LI1_cond $X=10.73 $Y=2.045
+ $X2=10.36 $Y2=1.87
r160 32 34 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=10.73 $Y=2.045
+ $X2=10.73 $Y2=2.3
r161 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.73 $Y=0.735
+ $X2=10.73 $Y2=0.4
r162 27 50 9.5576 $w=4.34e-07 $l=3.4e-07 $layer=LI1_cond $X=10.36 $Y=0.82
+ $X2=10.36 $Y2=1.16
r163 26 28 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=10.54 $Y=0.82
+ $X2=10.73 $Y2=0.735
r164 26 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.54 $Y=0.82
+ $X2=10.36 $Y2=0.82
r165 25 53 9.2186 $w=3.75e-07 $l=2.16217e-07 $layer=LI1_cond $X=9.365 $Y=1.53
+ $X2=9.26 $Y2=1.7
r166 24 25 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=9.365 $Y=0.425
+ $X2=9.365 $Y2=1.53
r167 23 37 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.27 $Y=0.34
+ $X2=8.102 $Y2=0.34
r168 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.28 $Y=0.34
+ $X2=9.365 $Y2=0.425
r169 22 23 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.28 $Y=0.34
+ $X2=8.27 $Y2=0.34
r170 16 49 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.075 $Y=1.325
+ $X2=10.075 $Y2=1.16
r171 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.075 $Y=1.325
+ $X2=10.075 $Y2=1.985
r172 15 51 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.045 $Y=0.565
+ $X2=10.045 $Y2=0.995
r173 4 57 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=10.57
+ $Y=1.485 $X2=10.71 $Y2=1.62
r174 4 34 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=10.57
+ $Y=1.485 $X2=10.71 $Y2=2.3
r175 3 53 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=9.02
+ $Y=1.575 $X2=9.235 $Y2=1.7
r176 2 30 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=10.595
+ $Y=0.235 $X2=10.73 $Y2=0.4
r177 1 37 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=7.945
+ $Y=0.245 $X2=8.105 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%CI 3 5 7 8 10 13 16 17 18 19
c65 19 0 1.5713e-19 $X=10.835 $Y=1.19
c66 5 0 8.35847e-20 $X=10.52 $Y=0.995
r67 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.775
+ $Y=1.16 $X2=10.775 $Y2=1.16
r68 17 22 106.665 $w=3.3e-07 $l=6.1e-07 $layer=POLY_cond $X=11.385 $Y=1.16
+ $X2=10.775 $Y2=1.16
r69 17 18 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.385 $Y=1.16
+ $X2=11.46 $Y2=1.16
r70 15 22 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=10.595 $Y=1.16
+ $X2=10.775 $Y2=1.16
r71 15 16 5.03009 $w=3.3e-07 $l=8.8e-08 $layer=POLY_cond $X=10.595 $Y=1.16
+ $X2=10.507 $Y2=1.16
r72 11 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.46 $Y=1.325
+ $X2=11.46 $Y2=1.16
r73 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.46 $Y=1.325
+ $X2=11.46 $Y2=1.985
r74 8 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.46 $Y=0.995
+ $X2=11.46 $Y2=1.16
r75 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.46 $Y=0.995
+ $X2=11.46 $Y2=0.565
r76 5 16 37.0704 $w=1.5e-07 $l=1.71377e-07 $layer=POLY_cond $X=10.52 $Y=0.995
+ $X2=10.507 $Y2=1.16
r77 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.52 $Y=0.995
+ $X2=10.52 $Y2=0.56
r78 1 16 37.0704 $w=1.5e-07 $l=1.70895e-07 $layer=POLY_cond $X=10.495 $Y=1.325
+ $X2=10.507 $Y2=1.16
r79 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.495 $Y=1.325
+ $X2=10.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_1710_49# 1 2 9 13 15 16 18 20 22 24 25 31
+ 35 36 37
c118 35 0 1.52424e-19 $X=11.88 $Y=1.16
c119 16 0 1.91615e-19 $X=8.735 $Y=1.615
r120 35 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.88 $Y=1.16
+ $X2=11.88 $Y2=0.995
r121 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.88
+ $Y=1.16 $X2=11.88 $Y2=1.16
r122 32 36 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=11.81 $Y=1.53
+ $X2=11.81 $Y2=1.16
r123 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.775 $Y=1.53
+ $X2=11.775 $Y2=1.53
r124 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.535 $Y=1.53
+ $X2=8.535 $Y2=1.53
r125 25 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.68 $Y=1.53
+ $X2=8.535 $Y2=1.53
r126 24 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.63 $Y=1.53
+ $X2=11.775 $Y2=1.53
r127 24 25 3.65098 $w=1.4e-07 $l=2.95e-06 $layer=MET1_cond $X=11.63 $Y=1.53
+ $X2=8.68 $Y2=1.53
r128 20 22 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.61 $Y=0.68
+ $X2=8.705 $Y2=0.68
r129 16 28 2.97297 $w=3.8e-07 $l=1.12916e-07 $layer=LI1_cond $X=8.735 $Y=1.615
+ $X2=8.67 $Y2=1.53
r130 16 18 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=1.615
+ $X2=8.735 $Y2=1.7
r131 15 28 6.50522 $w=3.8e-07 $l=1.8262e-07 $layer=LI1_cond $X=8.525 $Y=1.445
+ $X2=8.67 $Y2=1.53
r132 14 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.525 $Y=0.765
+ $X2=8.61 $Y2=0.68
r133 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.525 $Y=0.765
+ $X2=8.525 $Y2=1.445
r134 13 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.935 $Y=0.56
+ $X2=11.935 $Y2=0.995
r135 7 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.88 $Y=1.325
+ $X2=11.88 $Y2=1.16
r136 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.88 $Y=1.325
+ $X2=11.88 $Y2=1.985
r137 2 18 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=8.6
+ $Y=1.575 $X2=8.735 $Y2=1.7
r138 1 22 182 $w=1.7e-07 $l=5.06606e-07 $layer=licon1_NDIFF $count=1 $X=8.55
+ $Y=0.245 $X2=8.705 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_28_47# 1 2 3 4 5 6 23 27 29 32 34 37 40
+ 42 44 46 48 50 51 54 55 58 63 64
c152 63 0 4.61014e-20 $X=4.43 $Y=0.39
c153 55 0 8.07134e-20 $X=2.545 $Y=2.34
c154 50 0 1.3431e-19 $X=0.265 $Y=1.63
c155 48 0 5.07203e-20 $X=0.257 $Y=0.805
c156 40 0 1.51029e-19 $X=3.355 $Y=2.295
r157 63 64 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=0.365
+ $X2=4.265 $Y2=0.365
r158 57 58 33.7186 $w=1.99e-07 $l=5.5e-07 $layer=LI1_cond $X=2.805 $Y=0.79
+ $X2=3.355 $Y2=0.79
r159 54 55 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.375 $Y=2.34
+ $X2=2.545 $Y2=2.34
r160 52 53 2.75937 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=0.262 $Y=1.925
+ $X2=0.262 $Y2=2.01
r161 50 52 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=1.63
+ $X2=0.262 $Y2=1.925
r162 50 51 7.36284 $w=3.53e-07 $l=1.3e-07 $layer=LI1_cond $X=0.262 $Y=1.63
+ $X2=0.262 $Y2=1.5
r163 48 51 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.17 $Y=0.805
+ $X2=0.17 $Y2=1.5
r164 47 48 5.14454 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.805
r165 46 64 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=3.75 $Y=0.34
+ $X2=4.265 $Y2=0.34
r166 44 58 19.005 $w=1.99e-07 $l=3.1e-07 $layer=LI1_cond $X=3.665 $Y=0.79
+ $X2=3.355 $Y2=0.79
r167 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.665 $Y=0.425
+ $X2=3.75 $Y2=0.34
r168 43 44 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.665 $Y=0.425
+ $X2=3.665 $Y2=0.755
r169 40 61 3.40825 $w=1.7e-07 $l=1.07121e-07 $layer=LI1_cond $X=3.355 $Y=2.295
+ $X2=3.405 $Y2=2.38
r170 40 42 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.355 $Y=2.295
+ $X2=3.355 $Y2=1.62
r171 39 58 1.66034 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.355 $Y=0.925
+ $X2=3.355 $Y2=0.79
r172 39 42 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.355 $Y=0.925
+ $X2=3.355 $Y2=1.62
r173 37 61 3.40825 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.27 $Y=2.38
+ $X2=3.405 $Y2=2.38
r174 37 55 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.27 $Y=2.38
+ $X2=2.545 $Y2=2.38
r175 36 54 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.805 $Y=2.3
+ $X2=2.375 $Y2=2.3
r176 34 36 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.11 $Y=2.3
+ $X2=1.805 $Y2=2.3
r177 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.025 $Y=2.215
+ $X2=1.11 $Y2=2.3
r178 31 32 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.025 $Y=2.01
+ $X2=1.025 $Y2=2.215
r179 30 52 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.44 $Y=1.925
+ $X2=0.262 $Y2=1.925
r180 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.94 $Y=1.925
+ $X2=1.025 $Y2=2.01
r181 29 30 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=0.94 $Y=1.925
+ $X2=0.44 $Y2=1.925
r182 27 47 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.265 $Y=0.38
+ $X2=0.265 $Y2=0.735
r183 23 53 10.0212 $w=3.43e-07 $l=3e-07 $layer=LI1_cond $X=0.257 $Y=2.31
+ $X2=0.257 $Y2=2.01
r184 6 61 600 $w=1.7e-07 $l=9.55458e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.485 $X2=3.315 $Y2=2.38
r185 6 42 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.485 $X2=3.355 $Y2=1.62
r186 5 36 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.66
+ $Y=2.155 $X2=1.805 $Y2=2.3
r187 4 50 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.63
r188 4 23 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=2.31
r189 3 63 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.295
+ $Y=0.245 $X2=4.43 $Y2=0.39
r190 2 57 182 $w=1.7e-07 $l=5.92832e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.245 $X2=2.805 $Y2=0.74
r191 1 27 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%VPWR 1 2 3 4 15 17 21 25 29 31 33 38 46 53
+ 54 57 60 63 66
c129 33 0 1.3431e-19 $X=0.6 $Y=2.72
c130 29 0 1.52424e-19 $X=11.67 $Y=1.95
r131 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r132 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r133 60 61 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 58 61 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=5.29 $Y2=2.72
r135 57 58 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 54 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r137 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r138 51 66 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=11.84 $Y=2.72
+ $X2=11.712 $Y2=2.72
r139 51 53 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=11.84 $Y=2.72
+ $X2=12.19 $Y2=2.72
r140 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r141 50 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=10.35 $Y2=2.72
r142 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r143 47 63 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=10.455 $Y=2.72
+ $X2=10.287 $Y2=2.72
r144 47 49 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=10.455 $Y=2.72
+ $X2=11.27 $Y2=2.72
r145 46 66 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=11.585 $Y=2.72
+ $X2=11.712 $Y2=2.72
r146 46 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=11.585 $Y=2.72
+ $X2=11.27 $Y2=2.72
r147 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r148 44 45 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r149 42 45 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=9.89 $Y2=2.72
r150 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r151 41 44 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=9.89 $Y2=2.72
r152 41 42 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r153 39 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=2.72
+ $X2=5.435 $Y2=2.72
r154 39 41 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.6 $Y=2.72 $X2=5.75
+ $Y2=2.72
r155 38 63 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=10.12 $Y=2.72
+ $X2=10.287 $Y2=2.72
r156 38 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=10.12 $Y=2.72
+ $X2=9.89 $Y2=2.72
r157 33 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.685 $Y2=2.72
r158 33 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r159 31 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r160 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r161 27 66 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.712 $Y=2.635
+ $X2=11.712 $Y2=2.72
r162 27 29 30.9578 $w=2.53e-07 $l=6.85e-07 $layer=LI1_cond $X=11.712 $Y=2.635
+ $X2=11.712 $Y2=1.95
r163 23 63 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=10.287 $Y=2.635
+ $X2=10.287 $Y2=2.72
r164 23 25 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=10.287 $Y=2.635
+ $X2=10.287 $Y2=2.36
r165 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=2.635
+ $X2=5.435 $Y2=2.72
r166 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.435 $Y=2.635
+ $X2=5.435 $Y2=2.32
r167 18 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=2.72
+ $X2=0.685 $Y2=2.72
r168 17 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=2.72
+ $X2=5.435 $Y2=2.72
r169 17 18 293.583 $w=1.68e-07 $l=4.5e-06 $layer=LI1_cond $X=5.27 $Y=2.72
+ $X2=0.77 $Y2=2.72
r170 13 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.72
r171 13 15 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.685 $Y=2.635
+ $X2=0.685 $Y2=2.345
r172 4 29 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=11.535
+ $Y=1.485 $X2=11.67 $Y2=1.95
r173 3 25 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=10.15
+ $Y=1.485 $X2=10.285 $Y2=2.36
r174 2 21 600 $w=1.7e-07 $l=9.40798e-07 $layer=licon1_PDIFF $count=1 $X=5.21
+ $Y=1.485 $X2=5.435 $Y2=2.32
r175 1 15 600 $w=1.7e-07 $l=9.25041e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.485 $X2=0.685 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_1144_49# 1 2 3 12 15 16 19 20 22 23 26 30
c73 30 0 1.73441e-19 $X=6.54 $Y=2.01
c74 23 0 8.41027e-20 $X=7.135 $Y=1.955
c75 22 0 3.53612e-19 $X=7.135 $Y=1.23
r76 29 30 13.0837 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.295 $Y=2.01
+ $X2=6.54 $Y2=2.01
r77 22 32 26.0563 $w=2.27e-07 $l=5.03786e-07 $layer=LI1_cond $X=7.135 $Y=1.23
+ $X2=7.205 $Y2=0.76
r78 22 23 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.135 $Y=1.23
+ $X2=7.135 $Y2=1.955
r79 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=2.04
+ $X2=7.135 $Y2=1.955
r80 20 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.05 $Y=2.04
+ $X2=6.54 $Y2=2.04
r81 19 29 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.295 $Y=1.895
+ $X2=6.295 $Y2=2.01
r82 18 19 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.295 $Y=1.725
+ $X2=6.295 $Y2=1.895
r83 17 25 3.40825 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=5.98 $Y=1.64
+ $X2=5.812 $Y2=1.64
r84 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.21 $Y=1.64
+ $X2=6.295 $Y2=1.725
r85 16 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.21 $Y=1.64
+ $X2=5.98 $Y2=1.64
r86 15 25 3.40825 $w=1.7e-07 $l=1.19499e-07 $layer=LI1_cond $X=5.895 $Y=1.555
+ $X2=5.812 $Y2=1.64
r87 15 26 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.895 $Y=1.555
+ $X2=5.895 $Y2=0.815
r88 10 26 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=5.84 $Y=0.675
+ $X2=5.84 $Y2=0.815
r89 10 12 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=5.84 $Y=0.675
+ $X2=5.84 $Y2=0.58
r90 3 29 600 $w=1.7e-07 $l=8.679e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.485 $X2=6.375 $Y2=1.98
r91 3 25 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.485 $X2=5.855 $Y2=1.64
r92 2 32 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=7.14
+ $Y=0.245 $X2=7.275 $Y2=0.76
r93 1 12 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=5.72
+ $Y=0.245 $X2=5.855 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%COUT_N 1 2 7 8 13 18
r28 14 18 0.426831 $w=2.68e-07 $l=1e-08 $layer=LI1_cond $X=6.745 $Y=1.54
+ $X2=6.745 $Y2=1.53
r29 8 24 2.33156 $w=2.25e-07 $l=4.3e-08 $layer=LI1_cond $X=6.745 $Y=1.577
+ $X2=6.745 $Y2=1.62
r30 8 14 2.0467 $w=2.7e-07 $l=3.7e-08 $layer=LI1_cond $X=6.745 $Y=1.577
+ $X2=6.745 $Y2=1.54
r31 8 18 1.62196 $w=2.68e-07 $l=3.8e-08 $layer=LI1_cond $X=6.745 $Y=1.492
+ $X2=6.745 $Y2=1.53
r32 7 13 3.70924 $w=2.7e-07 $l=9.25203e-08 $layer=LI1_cond $X=6.772 $Y=0.845
+ $X2=6.745 $Y2=0.925
r33 7 20 4.16466 $w=2.49e-07 $l=8.5e-08 $layer=LI1_cond $X=6.772 $Y=0.845
+ $X2=6.772 $Y2=0.76
r34 7 8 23.9879 $w=2.68e-07 $l=5.62e-07 $layer=LI1_cond $X=6.745 $Y=0.93
+ $X2=6.745 $Y2=1.492
r35 7 13 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=6.745 $Y=0.93
+ $X2=6.745 $Y2=0.925
r36 2 24 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.66
+ $Y=1.485 $X2=6.795 $Y2=1.62
r37 1 20 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=6.715
+ $Y=0.245 $X2=6.85 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_1261_49# 1 2 3 4 13 17 19 21 27 29 34 38
+ 40 41 44 47 48
r131 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.315 $Y=0.85
+ $X2=11.315 $Y2=0.85
r132 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.615 $Y=0.85
+ $X2=7.615 $Y2=0.85
r133 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.76 $Y=0.85
+ $X2=7.615 $Y2=0.85
r134 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.17 $Y=0.85
+ $X2=11.315 $Y2=0.85
r135 40 41 4.22029 $w=1.4e-07 $l=3.41e-06 $layer=MET1_cond $X=11.17 $Y=0.85
+ $X2=7.76 $Y2=0.85
r136 38 48 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=11.29 $Y=0.805
+ $X2=11.29 $Y2=0.85
r137 38 39 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.29 $Y=0.805
+ $X2=11.29 $Y2=0.68
r138 37 48 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=11.29 $Y=1.455
+ $X2=11.29 $Y2=0.85
r139 35 44 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.615 $Y=0.425
+ $X2=7.615 $Y2=0.85
r140 34 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.615 $Y=1.105
+ $X2=7.615 $Y2=0.85
r141 29 32 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.43 $Y=0.34
+ $X2=6.43 $Y2=0.485
r142 27 39 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=11.25 $Y=0.55
+ $X2=11.25 $Y2=0.68
r143 21 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.25 $Y=1.635
+ $X2=11.25 $Y2=2.315
r144 19 37 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.25 $Y=1.62
+ $X2=11.25 $Y2=1.455
r145 19 21 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.25 $Y=1.62
+ $X2=11.25 $Y2=1.635
r146 15 34 22.7412 $w=2.28e-07 $l=4.90026e-07 $layer=LI1_cond $X=7.475 $Y=1.53
+ $X2=7.615 $Y2=1.105
r147 15 17 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.475 $Y=1.53
+ $X2=7.475 $Y2=1.62
r148 14 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=0.34
+ $X2=6.43 $Y2=0.34
r149 13 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.53 $Y=0.34
+ $X2=7.615 $Y2=0.425
r150 13 14 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=7.53 $Y=0.34 $X2=6.595
+ $Y2=0.34
r151 4 23 400 $w=1.7e-07 $l=8.90309e-07 $layer=licon1_PDIFF $count=1 $X=11.125
+ $Y=1.485 $X2=11.25 $Y2=2.315
r152 4 21 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=11.125
+ $Y=1.485 $X2=11.25 $Y2=1.635
r153 3 17 300 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_PDIFF $count=2 $X=7.08
+ $Y=1.485 $X2=7.475 $Y2=1.62
r154 2 27 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=11.125
+ $Y=0.245 $X2=11.25 $Y2=0.55
r155 1 32 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=6.305
+ $Y=0.245 $X2=6.43 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%A_1634_315# 1 2 3 12 14 15 18 22 25 26 27
c58 26 0 8.35847e-20 $X=9.835 $Y=0.825
r59 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=9.735 $Y=0.825
+ $X2=9.735 $Y2=1.535
r60 23 25 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=9.8 $Y=2.215
+ $X2=9.8 $Y2=1.86
r61 22 27 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=9.8 $Y=1.685 $X2=9.8
+ $Y2=1.535
r62 22 25 6.72258 $w=2.98e-07 $l=1.75e-07 $layer=LI1_cond $X=9.8 $Y=1.685
+ $X2=9.8 $Y2=1.86
r63 16 26 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.835 $Y=0.64
+ $X2=9.835 $Y2=0.825
r64 16 18 7.47531 $w=3.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.835 $Y=0.64
+ $X2=9.835 $Y2=0.4
r65 14 23 7.51767 $w=1.7e-07 $l=2.49199e-07 $layer=LI1_cond $X=9.62 $Y=2.38
+ $X2=9.8 $Y2=2.215
r66 14 15 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=9.62 $Y=2.38
+ $X2=8.4 $Y2=2.38
r67 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.315 $Y=2.295
+ $X2=8.4 $Y2=2.38
r68 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.315 $Y=2.295
+ $X2=8.315 $Y2=1.95
r69 3 25 300 $w=1.7e-07 $l=4.66369e-07 $layer=licon1_PDIFF $count=2 $X=9.65
+ $Y=1.485 $X2=9.855 $Y2=1.86
r70 2 12 300 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_PDIFF $count=2 $X=8.17
+ $Y=1.575 $X2=8.315 $Y2=1.95
r71 1 18 91 $w=1.7e-07 $l=9.09203e-07 $layer=licon1_NDIFF $count=2 $X=8.99
+ $Y=0.245 $X2=9.825 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%SUM 1 2 7 8 9 10 11 12 24
r19 12 36 8.86495 $w=3.23e-07 $l=2.5e-07 $layer=LI1_cond $X=12.172 $Y=2.21
+ $X2=12.172 $Y2=1.96
r20 11 33 2.87224 $w=3.23e-07 $l=8.1e-08 $layer=LI1_cond $X=12.172 $Y=1.866
+ $X2=12.172 $Y2=1.947
r21 11 36 0.319138 $w=3.23e-07 $l=9e-09 $layer=LI1_cond $X=12.172 $Y=1.951
+ $X2=12.172 $Y2=1.96
r22 11 33 0.141839 $w=3.23e-07 $l=4e-09 $layer=LI1_cond $X=12.172 $Y=1.951
+ $X2=12.172 $Y2=1.947
r23 10 11 10.3592 $w=3.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.235 $Y=1.53
+ $X2=12.235 $Y2=1.785
r24 9 10 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=12.235 $Y=1.19
+ $X2=12.235 $Y2=1.53
r25 8 40 2.95469 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=12.165 $Y=0.795
+ $X2=12.165 $Y2=0.825
r26 8 22 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=12.165 $Y=0.795
+ $X2=12.165 $Y2=0.655
r27 8 9 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=12.235 $Y=0.88
+ $X2=12.235 $Y2=1.19
r28 8 40 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=12.235 $Y=0.88
+ $X2=12.235 $Y2=0.825
r29 7 22 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=12.165 $Y=0.51
+ $X2=12.165 $Y2=0.655
r30 7 24 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=12.165 $Y=0.51
+ $X2=12.165 $Y2=0.39
r31 2 36 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=11.955
+ $Y=1.485 $X2=12.095 $Y2=1.96
r32 1 24 91 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_NDIFF $count=2 $X=12.01
+ $Y=0.235 $X2=12.16 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__FAHCON_1%VGND 1 2 3 4 17 21 25 29 31 33 41 49 56 57
+ 60 63 66 69
c131 41 0 1.49929e-19 $X=10.2 $Y=0
c132 25 0 3.96944e-20 $X=10.285 $Y=0.4
c133 17 0 1.50726e-19 $X=0.715 $Y=0.38
r134 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r135 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r136 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r137 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r138 57 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r139 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r140 54 69 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=11.68 $Y2=0
r141 54 56 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.825 $Y=0
+ $X2=12.19 $Y2=0
r142 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r143 53 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=10.35 $Y2=0
r144 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r145 50 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.37 $Y=0
+ $X2=10.285 $Y2=0
r146 50 52 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=10.37 $Y=0 $X2=11.27
+ $Y2=0
r147 49 69 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.535 $Y=0
+ $X2=11.68 $Y2=0
r148 49 52 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.535 $Y=0
+ $X2=11.27 $Y2=0
r149 48 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r150 47 48 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r151 45 48 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=9.89
+ $Y2=0
r152 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r153 44 47 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=9.89
+ $Y2=0
r154 44 45 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r155 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.365
+ $Y2=0
r156 42 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.75
+ $Y2=0
r157 41 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.2 $Y=0 $X2=10.285
+ $Y2=0
r158 41 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.2 $Y=0 $X2=9.89
+ $Y2=0
r159 40 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r160 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r161 37 40 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r162 37 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r163 36 39 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r164 36 37 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r165 34 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0 $X2=0.715
+ $Y2=0
r166 34 36 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.8 $Y=0 $X2=1.15
+ $Y2=0
r167 33 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.2 $Y=0 $X2=5.365
+ $Y2=0
r168 33 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.2 $Y=0 $X2=4.83
+ $Y2=0
r169 31 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r170 27 69 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0
r171 27 29 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0.39
r172 23 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0
r173 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.4
r174 19 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0
r175 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0.38
r176 15 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r177 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.38
r178 4 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=11.535
+ $Y=0.245 $X2=11.67 $Y2=0.39
r179 3 25 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=10.12
+ $Y=0.245 $X2=10.285 $Y2=0.4
r180 2 21 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.23
+ $Y=0.235 $X2=5.365 $Y2=0.38
r181 1 17 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.715 $Y2=0.38
.ends


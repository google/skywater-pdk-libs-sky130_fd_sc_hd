* File: sky130_fd_sc_hd__einvn_2.spice.pex
* Created: Thu Aug 27 14:20:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVN_2%TE_B 3 5 7 9 11 13 14 16 18 19 20
c42 16 0 1.87565e-19 $X=1.365 $Y=1.47
c43 14 0 1.73709e-19 $X=1.29 $Y=1.395
r44 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r45 16 18 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.365 $Y=1.47
+ $X2=1.365 $Y2=2.015
r46 15 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.395
+ $X2=0.945 $Y2=1.395
r47 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.29 $Y=1.395
+ $X2=1.365 $Y2=1.47
r48 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.29 $Y=1.395
+ $X2=1.02 $Y2=1.395
r49 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.945 $Y=1.47
+ $X2=0.945 $Y2=1.395
r50 11 13 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.945 $Y=1.47
+ $X2=0.945 $Y2=2.015
r51 10 23 32.2707 $w=3.51e-07 $l=3.26994e-07 $layer=POLY_cond $X=0.545 $Y=1.395
+ $X2=0.325 $Y2=1.16
r52 9 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.395
+ $X2=0.945 $Y2=1.395
r53 9 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.87 $Y=1.395
+ $X2=0.545 $Y2=1.395
r54 5 10 26.4367 $w=3.51e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.47 $Y=1.47
+ $X2=0.545 $Y2=1.395
r55 5 7 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.47 $Y=1.47 $X2=0.47
+ $Y2=2.165
r56 1 23 38.7956 $w=3.51e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.325 $Y2=1.16
r57 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_2%A_27_47# 1 2 7 9 10 11 12 14 17 21 24 25 27
+ 36
c64 24 0 1.87565e-19 $X=0.695 $Y=1.555
r65 28 36 19.8845 $w=3.03e-07 $l=1.25e-07 $layer=POLY_cond $X=1.87 $Y=1.16
+ $X2=1.87 $Y2=1.035
r66 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.87
+ $Y=1.16 $X2=1.87 $Y2=1.16
r67 25 31 7.35142 $w=3.69e-07 $l=2.38747e-07 $layer=LI1_cond $X=0.895 $Y=1.135
+ $X2=0.695 $Y2=1.05
r68 25 27 40.1297 $w=2.78e-07 $l=9.75e-07 $layer=LI1_cond $X=0.895 $Y=1.135
+ $X2=1.87 $Y2=1.135
r69 23 31 0.218444 $w=4e-07 $l=2.25e-07 $layer=LI1_cond $X=0.695 $Y=1.275
+ $X2=0.695 $Y2=1.05
r70 23 24 8.0671 $w=3.98e-07 $l=2.8e-07 $layer=LI1_cond $X=0.695 $Y=1.275
+ $X2=0.695 $Y2=1.555
r71 19 24 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.215 $Y=1.64
+ $X2=0.695 $Y2=1.64
r72 19 21 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=0.215 $Y=1.725
+ $X2=0.215 $Y2=2.165
r73 15 31 15.8699 $w=3.69e-07 $l=6.48074e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.695 $Y2=1.05
r74 15 17 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r75 12 36 24.2248 $w=3.03e-07 $l=9.48683e-08 $layer=POLY_cond $X=1.825 $Y=0.96
+ $X2=1.87 $Y2=1.035
r76 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.825 $Y=0.96
+ $X2=1.825 $Y2=0.56
r77 10 36 19.2026 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.035
+ $X2=1.87 $Y2=1.035
r78 10 11 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.705 $Y=1.035
+ $X2=1.48 $Y2=1.035
r79 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.405 $Y=0.96
+ $X2=1.48 $Y2=1.035
r80 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.405 $Y=0.96 $X2=1.405
+ $Y2=0.56
r81 2 21 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.165
r82 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_2%A 3 7 11 15 17 20 23
r47 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r48 17 23 27.9249 $w=2.9e-07 $l=1.35e-07 $layer=POLY_cond $X=2.815 $Y=1.16
+ $X2=2.95 $Y2=1.16
r49 17 19 12.6442 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=2.815 $Y=1.16
+ $X2=2.74 $Y2=1.16
r50 13 19 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.74 $Y=1.305
+ $X2=2.74 $Y2=1.16
r51 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.74 $Y=1.305
+ $X2=2.74 $Y2=1.985
r52 9 19 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.74 $Y=1.015
+ $X2=2.74 $Y2=1.16
r53 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.74 $Y=1.015
+ $X2=2.74 $Y2=0.56
r54 1 19 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=2.32 $Y=1.16
+ $X2=2.74 $Y2=1.16
r55 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.32 $Y=1.295 $X2=2.32
+ $Y2=1.985
r56 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.32 $Y=1.025
+ $X2=2.32 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_2%VPWR 1 2 9 11 12 16 17 19 30 31 34 39
c49 11 0 5.07009e-20 $X=2 $Y=2.53
r50 37 39 10.7019 $w=5.48e-07 $l=2.05e-07 $layer=LI1_cond $X=2.07 $Y=2.53
+ $X2=2.275 $Y2=2.53
r51 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 31 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 30 39 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.275 $Y2=2.72
r55 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 27 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 27 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r58 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 24 34 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r60 24 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 19 34 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r62 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 17 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 16 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 15 16 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=2.53
+ $X2=1.41 $Y2=2.53
r67 12 15 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.685 $Y=2.53
+ $X2=1.575 $Y2=2.53
r68 11 37 1.52228 $w=5.48e-07 $l=7e-08 $layer=LI1_cond $X=2 $Y=2.53 $X2=2.07
+ $Y2=2.53
r69 11 12 6.85027 $w=5.48e-07 $l=3.15e-07 $layer=LI1_cond $X=2 $Y=2.53 $X2=1.685
+ $Y2=2.53
r70 7 34 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r71 7 9 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.02
r72 2 15 600 $w=1.7e-07 $l=8.59855e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.545 $X2=1.575 $Y2=2.34
r73 1 9 300 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.845 $X2=0.705 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_2%A_204_309# 1 2 9 11 15 20
c31 9 0 1.73709e-19 $X=1.155 $Y=2.265
r32 18 20 17.0802 $w=6.38e-07 $l=6.2e-07 $layer=LI1_cond $X=1.155 $Y=1.765
+ $X2=1.775 $Y2=1.765
r33 13 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.53 $Y=2.085
+ $X2=2.53 $Y2=2.265
r34 11 13 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.445 $Y=1.975
+ $X2=2.53 $Y2=2.085
r35 11 20 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=2.445 $Y=1.975
+ $X2=1.775 $Y2=1.975
r36 7 18 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=1.155 $Y=2.085
+ $X2=1.155 $Y2=1.765
r37 7 9 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.155 $Y=2.085
+ $X2=1.155 $Y2=2.265
r38 2 15 600 $w=1.7e-07 $l=8.44808e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.485 $X2=2.53 $Y2=2.265
r39 1 18 600 $w=1.7e-07 $l=4.4238e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.545 $X2=1.155 $Y2=1.925
r40 1 9 600 $w=1.7e-07 $l=7.84602e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.545 $X2=1.155 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_2%Z 1 2 3 10 11 12 13 14 15 16 26 34
c39 2 0 5.07009e-20 $X=1.965 $Y=1.485
r40 34 49 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.49 $Y=0.85 $X2=2.49
+ $Y2=0.845
r41 26 50 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.365 $Y=1.57
+ $X2=2.49 $Y2=1.57
r42 15 16 13.0061 $w=3.48e-07 $l=3.95e-07 $layer=LI1_cond $X=2.96 $Y=1.815
+ $X2=2.96 $Y2=2.21
r43 15 39 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=2.96 $Y=1.815
+ $X2=2.96 $Y2=1.695
r44 14 39 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=2.99 $Y=1.57 $X2=2.96
+ $Y2=1.57
r45 13 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.53 $Y=1.57 $X2=2.96
+ $Y2=1.57
r46 13 50 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=2.53 $Y=1.57 $X2=2.49
+ $Y2=1.57
r47 13 50 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=2.49 $Y=1.445
+ $X2=2.49 $Y2=1.57
r48 12 13 8.86994 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.49 $Y=1.19
+ $X2=2.49 $Y2=1.445
r49 11 49 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=0.76
+ $X2=2.53 $Y2=0.845
r50 11 12 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=2.49 $Y=0.89 $X2=2.49
+ $Y2=1.19
r51 11 34 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=2.49 $Y=0.89 $X2=2.49
+ $Y2=0.85
r52 10 26 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.07 $Y=1.57
+ $X2=2.365 $Y2=1.57
r53 3 15 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=2.815
+ $Y=1.485 $X2=2.95 $Y2=1.815
r54 2 10 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.485 $X2=2.11 $Y2=1.61
r55 1 11 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.53 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r46 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r47 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r49 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r50 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r51 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r52 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r53 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.615
+ $Y2=0
r54 27 29 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=2.07
+ $Y2=0
r55 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r56 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r57 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r59 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r60 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.615
+ $Y2=0
r61 22 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.15
+ $Y2=0
r62 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r63 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r64 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r65 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0
r67 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.36
r68 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r69 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r70 2 13 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.235 $X2=1.615 $Y2=0.36
r71 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__EINVN_2%A_214_120# 1 2 3 12 18 19 22 25
r35 20 22 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3 $Y=0.425 $X2=3
+ $Y2=0.56
r36 18 20 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.865 $Y=0.34
+ $X2=3 $Y2=0.425
r37 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.865 $Y=0.34
+ $X2=2.195 $Y2=0.34
r38 15 17 4.46866 $w=2.43e-07 $l=9.5e-08 $layer=LI1_cond $X=2.072 $Y=0.655
+ $X2=2.072 $Y2=0.56
r39 14 19 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=2.072 $Y=0.425
+ $X2=2.195 $Y2=0.34
r40 14 17 6.3502 $w=2.43e-07 $l=1.35e-07 $layer=LI1_cond $X=2.072 $Y=0.425
+ $X2=2.072 $Y2=0.56
r41 13 25 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.28 $Y=0.74
+ $X2=1.147 $Y2=0.74
r42 12 15 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=1.95 $Y=0.74
+ $X2=2.072 $Y2=0.655
r43 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.95 $Y=0.74
+ $X2=1.28 $Y2=0.74
r44 3 22 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.235 $X2=2.95 $Y2=0.56
r45 2 17 182 $w=1.7e-07 $l=4.03113e-07 $layer=licon1_NDIFF $count=1 $X=1.9
+ $Y=0.235 $X2=2.075 $Y2=0.56
r46 1 25 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.6 $X2=1.195 $Y2=0.74
.ends


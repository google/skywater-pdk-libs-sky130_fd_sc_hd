* File: sky130_fd_sc_hd__einvp_8.spice.pex
* Created: Thu Aug 27 14:20:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVP_8%TE 1 3 6 8 9 10 12 13 15 17 18 20 22 23 25
+ 27 28 30 32 33 35 37 38 40 42 43 45 47 48 49 50 51 52 53 54 55 56
c136 54 0 9.62962e-20 $X=3.43 $Y=1.035
c137 53 0 9.62962e-20 $X=3.01 $Y=1.035
c138 52 0 9.62962e-20 $X=2.59 $Y=1.035
c139 51 0 9.62962e-20 $X=2.17 $Y=1.035
c140 50 0 9.62962e-20 $X=1.75 $Y=1.035
c141 49 0 9.62962e-20 $X=1.33 $Y=1.035
c142 43 0 4.50788e-20 $X=3.775 $Y=1.035
c143 38 0 1.96823e-19 $X=3.355 $Y=1.035
c144 28 0 1.96823e-19 $X=2.515 $Y=1.035
c145 18 0 1.96823e-19 $X=1.675 $Y=1.035
r146 60 62 31.7105 $w=3.42e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.142
+ $X2=0.47 $Y2=1.142
r147 55 56 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r148 55 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r149 45 47 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.85 $Y=0.96 $X2=3.85
+ $Y2=0.56
r150 44 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=1.035
+ $X2=3.43 $Y2=1.035
r151 43 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.775 $Y=1.035
+ $X2=3.85 $Y2=0.96
r152 43 44 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.775 $Y=1.035
+ $X2=3.505 $Y2=1.035
r153 40 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.43 $Y=0.96
+ $X2=3.43 $Y2=1.035
r154 40 42 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.43 $Y=0.96 $X2=3.43
+ $Y2=0.56
r155 39 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.085 $Y=1.035
+ $X2=3.01 $Y2=1.035
r156 38 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.355 $Y=1.035
+ $X2=3.43 $Y2=1.035
r157 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.355 $Y=1.035
+ $X2=3.085 $Y2=1.035
r158 35 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.01 $Y=0.96
+ $X2=3.01 $Y2=1.035
r159 35 37 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.01 $Y=0.96 $X2=3.01
+ $Y2=0.56
r160 34 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.665 $Y=1.035
+ $X2=2.59 $Y2=1.035
r161 33 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.935 $Y=1.035
+ $X2=3.01 $Y2=1.035
r162 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.935 $Y=1.035
+ $X2=2.665 $Y2=1.035
r163 30 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.59 $Y=0.96
+ $X2=2.59 $Y2=1.035
r164 30 32 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.59 $Y=0.96 $X2=2.59
+ $Y2=0.56
r165 29 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.245 $Y=1.035
+ $X2=2.17 $Y2=1.035
r166 28 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.515 $Y=1.035
+ $X2=2.59 $Y2=1.035
r167 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.515 $Y=1.035
+ $X2=2.245 $Y2=1.035
r168 25 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.17 $Y=0.96
+ $X2=2.17 $Y2=1.035
r169 25 27 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.17 $Y=0.96 $X2=2.17
+ $Y2=0.56
r170 24 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.035
+ $X2=1.75 $Y2=1.035
r171 23 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.095 $Y=1.035
+ $X2=2.17 $Y2=1.035
r172 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.095 $Y=1.035
+ $X2=1.825 $Y2=1.035
r173 20 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=0.96
+ $X2=1.75 $Y2=1.035
r174 20 22 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.75 $Y=0.96 $X2=1.75
+ $Y2=0.56
r175 19 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.405 $Y=1.035
+ $X2=1.33 $Y2=1.035
r176 18 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.035
+ $X2=1.75 $Y2=1.035
r177 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.675 $Y=1.035
+ $X2=1.405 $Y2=1.035
r178 15 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.33 $Y=0.96
+ $X2=1.33 $Y2=1.035
r179 15 17 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.33 $Y=0.96 $X2=1.33
+ $Y2=0.56
r180 14 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.965 $Y=1.035
+ $X2=0.89 $Y2=1.035
r181 13 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.255 $Y=1.035
+ $X2=1.33 $Y2=1.035
r182 13 14 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.255 $Y=1.035
+ $X2=0.965 $Y2=1.035
r183 10 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=0.96
+ $X2=0.89 $Y2=1.035
r184 10 12 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.89 $Y=0.96 $X2=0.89
+ $Y2=0.56
r185 9 62 26.0143 $w=3.42e-07 $l=1.39549e-07 $layer=POLY_cond $X=0.545 $Y=1.035
+ $X2=0.47 $Y2=1.142
r186 8 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.815 $Y=1.035
+ $X2=0.89 $Y2=1.035
r187 8 9 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.815 $Y=1.035
+ $X2=0.545 $Y2=1.035
r188 4 62 22.0749 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.142
r189 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r190 1 62 22.0749 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.47 $Y=0.96
+ $X2=0.47 $Y2=1.142
r191 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.47 $Y=0.96 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_8%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 25 27 29 30 32 34 35 37 39 40 42 43 44 45 46 47 51 55 59 61 62 64 67 68 78
c163 78 0 1.9418e-19 $X=0.687 $Y=1.16
c164 47 0 1.50055e-19 $X=3.51 $Y=1.395
c165 46 0 1.51809e-19 $X=3.09 $Y=1.395
c166 45 0 1.50055e-19 $X=2.67 $Y=1.395
c167 44 0 1.51809e-19 $X=2.25 $Y=1.395
c168 43 0 1.50055e-19 $X=1.83 $Y=1.395
c169 40 0 2.25041e-19 $X=4.35 $Y=1.47
c170 35 0 7.37964e-20 $X=3.855 $Y=1.395
c171 30 0 7.37964e-20 $X=3.435 $Y=1.395
c172 25 0 7.37964e-20 $X=3.015 $Y=1.395
c173 20 0 7.37964e-20 $X=2.595 $Y=1.395
c174 15 0 7.37964e-20 $X=2.175 $Y=1.395
c175 11 0 1.86371e-19 $X=1.485 $Y=1.395
c176 10 0 7.37964e-20 $X=1.755 $Y=1.395
r177 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.29
+ $Y=1.16 $X2=4.29 $Y2=1.16
r178 65 78 0.820356 $w=3.3e-07 $l=1.88e-07 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=0.687 $Y2=1.16
r179 65 67 119.26 $w=3.28e-07 $l=3.415e-06 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=4.29 $Y2=1.16
r180 63 78 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=0.687 $Y=1.325
+ $X2=0.687 $Y2=1.16
r181 63 64 14.1366 $w=3.73e-07 $l=4.6e-07 $layer=LI1_cond $X=0.687 $Y=1.325
+ $X2=0.687 $Y2=1.785
r182 62 78 5.82594 $w=2.85e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.597 $Y=0.995
+ $X2=0.687 $Y2=1.16
r183 61 62 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.597 $Y=0.825
+ $X2=0.597 $Y2=0.995
r184 57 64 30.7936 $w=1.68e-07 $l=4.72e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.687 $Y2=1.87
r185 57 59 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=1.955
+ $X2=0.215 $Y2=2.165
r186 53 61 24.9219 $w=1.68e-07 $l=3.82e-07 $layer=LI1_cond $X=0.215 $Y=0.74
+ $X2=0.597 $Y2=0.74
r187 53 55 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r188 50 68 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=4.29 $Y=1.32
+ $X2=4.29 $Y2=1.16
r189 50 51 30.766 $w=1.5e-07 $l=6e-08 $layer=POLY_cond $X=4.29 $Y=1.395 $X2=4.35
+ $Y2=1.395
r190 48 50 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.93 $Y=1.395
+ $X2=4.29 $Y2=1.395
r191 40 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.35 $Y=1.47
+ $X2=4.35 $Y2=1.395
r192 40 42 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.35 $Y=1.47
+ $X2=4.35 $Y2=2.015
r193 37 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.93 $Y=1.47
+ $X2=3.93 $Y2=1.395
r194 37 39 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.93 $Y=1.47
+ $X2=3.93 $Y2=2.015
r195 36 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=1.395
+ $X2=3.51 $Y2=1.395
r196 35 48 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.855 $Y=1.395
+ $X2=3.93 $Y2=1.395
r197 35 36 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.855 $Y=1.395
+ $X2=3.585 $Y2=1.395
r198 32 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=1.47
+ $X2=3.51 $Y2=1.395
r199 32 34 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.51 $Y=1.47
+ $X2=3.51 $Y2=2.015
r200 31 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.395
+ $X2=3.09 $Y2=1.395
r201 30 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.435 $Y=1.395
+ $X2=3.51 $Y2=1.395
r202 30 31 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.435 $Y=1.395
+ $X2=3.165 $Y2=1.395
r203 27 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.09 $Y=1.47
+ $X2=3.09 $Y2=1.395
r204 27 29 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.09 $Y=1.47
+ $X2=3.09 $Y2=2.015
r205 26 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=1.395
+ $X2=2.67 $Y2=1.395
r206 25 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=1.395
+ $X2=3.09 $Y2=1.395
r207 25 26 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.015 $Y=1.395
+ $X2=2.745 $Y2=1.395
r208 22 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=1.47
+ $X2=2.67 $Y2=1.395
r209 22 24 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.67 $Y=1.47
+ $X2=2.67 $Y2=2.015
r210 21 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.325 $Y=1.395
+ $X2=2.25 $Y2=1.395
r211 20 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.595 $Y=1.395
+ $X2=2.67 $Y2=1.395
r212 20 21 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.595 $Y=1.395
+ $X2=2.325 $Y2=1.395
r213 17 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=1.47
+ $X2=2.25 $Y2=1.395
r214 17 19 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.25 $Y=1.47
+ $X2=2.25 $Y2=2.015
r215 16 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.395
+ $X2=1.83 $Y2=1.395
r216 15 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.175 $Y=1.395
+ $X2=2.25 $Y2=1.395
r217 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.175 $Y=1.395
+ $X2=1.905 $Y2=1.395
r218 12 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.47
+ $X2=1.83 $Y2=1.395
r219 12 14 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.83 $Y=1.47
+ $X2=1.83 $Y2=2.015
r220 10 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=1.395
+ $X2=1.83 $Y2=1.395
r221 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.755 $Y=1.395
+ $X2=1.485 $Y2=1.395
r222 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.47
+ $X2=1.485 $Y2=1.395
r223 7 9 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.41 $Y=1.47
+ $X2=1.41 $Y2=2.015
r224 2 59 600 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.165
r225 1 55 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_8%A 1 3 6 8 10 13 17 21 25 29 31 33 36 38 40
+ 43 47 51 53 55 59 61 62 63 64 65 66
r133 100 101 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.965
+ $Y=1.16 $X2=7.965 $Y2=1.16
r134 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.285
+ $Y=1.16 $X2=7.285 $Y2=1.16
r135 89 92 56.1233 $w=2.92e-07 $l=3.4e-07 $layer=POLY_cond $X=6.945 $Y=1.16
+ $X2=7.285 $Y2=1.16
r136 89 90 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.945
+ $Y=1.16 $X2=6.945 $Y2=1.16
r137 87 89 3.30137 $w=2.92e-07 $l=2e-08 $layer=POLY_cond $X=6.925 $Y=1.16
+ $X2=6.945 $Y2=1.16
r138 86 87 69.3288 $w=2.92e-07 $l=4.2e-07 $layer=POLY_cond $X=6.505 $Y=1.16
+ $X2=6.925 $Y2=1.16
r139 84 86 39.6164 $w=2.92e-07 $l=2.4e-07 $layer=POLY_cond $X=6.265 $Y=1.16
+ $X2=6.505 $Y2=1.16
r140 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.925
+ $Y=1.16 $X2=5.925 $Y2=1.16
r141 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.585
+ $Y=1.16 $X2=5.585 $Y2=1.16
r142 74 76 56.1233 $w=2.92e-07 $l=3.4e-07 $layer=POLY_cond $X=5.245 $Y=1.16
+ $X2=5.585 $Y2=1.16
r143 73 74 69.3288 $w=2.92e-07 $l=4.2e-07 $layer=POLY_cond $X=4.825 $Y=1.16
+ $X2=5.245 $Y2=1.16
r144 66 101 4.97132 $w=2.53e-07 $l=1.1e-07 $layer=LI1_cond $X=8.075 $Y=1.147
+ $X2=7.965 $Y2=1.147
r145 65 101 15.8178 $w=2.53e-07 $l=3.5e-07 $layer=LI1_cond $X=7.615 $Y=1.147
+ $X2=7.965 $Y2=1.147
r146 65 93 14.914 $w=2.53e-07 $l=3.3e-07 $layer=LI1_cond $X=7.615 $Y=1.147
+ $X2=7.285 $Y2=1.147
r147 65 96 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.625
+ $Y=1.16 $X2=7.625 $Y2=1.16
r148 64 93 5.8752 $w=2.53e-07 $l=1.3e-07 $layer=LI1_cond $X=7.155 $Y=1.147
+ $X2=7.285 $Y2=1.147
r149 64 90 9.49071 $w=2.53e-07 $l=2.1e-07 $layer=LI1_cond $X=7.155 $Y=1.147
+ $X2=6.945 $Y2=1.147
r150 63 90 11.2985 $w=2.53e-07 $l=2.5e-07 $layer=LI1_cond $X=6.695 $Y=1.147
+ $X2=6.945 $Y2=1.147
r151 62 63 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=6.235 $Y=1.147
+ $X2=6.695 $Y2=1.147
r152 62 81 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=6.235 $Y=1.147
+ $X2=5.925 $Y2=1.147
r153 62 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.265
+ $Y=1.16 $X2=6.265 $Y2=1.16
r154 61 81 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=5.775 $Y=1.147
+ $X2=5.925 $Y2=1.147
r155 61 77 8.58683 $w=2.53e-07 $l=1.9e-07 $layer=LI1_cond $X=5.775 $Y=1.147
+ $X2=5.585 $Y2=1.147
r156 53 100 33.0137 $w=2.92e-07 $l=2e-07 $layer=POLY_cond $X=7.765 $Y=1.16
+ $X2=7.965 $Y2=1.16
r157 53 96 23.1096 $w=2.92e-07 $l=1.4e-07 $layer=POLY_cond $X=7.765 $Y=1.16
+ $X2=7.625 $Y2=1.16
r158 53 59 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.765 $Y=1.305
+ $X2=7.765 $Y2=1.985
r159 53 55 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.765 $Y=1.015
+ $X2=7.765 $Y2=0.56
r160 45 96 46.2192 $w=2.92e-07 $l=2.8e-07 $layer=POLY_cond $X=7.345 $Y=1.16
+ $X2=7.625 $Y2=1.16
r161 45 92 9.90411 $w=2.92e-07 $l=6e-08 $layer=POLY_cond $X=7.345 $Y=1.16
+ $X2=7.285 $Y2=1.16
r162 45 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.345 $Y=1.295
+ $X2=7.345 $Y2=1.985
r163 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.345 $Y=1.025
+ $X2=7.345 $Y2=0.56
r164 41 87 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=1.16
r165 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=1.985
r166 38 87 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=0.995
+ $X2=6.925 $Y2=1.16
r167 38 40 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.925 $Y=0.995
+ $X2=6.925 $Y2=0.56
r168 34 86 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=1.325
+ $X2=6.505 $Y2=1.16
r169 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.505 $Y=1.325
+ $X2=6.505 $Y2=1.985
r170 31 86 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=0.995
+ $X2=6.505 $Y2=1.16
r171 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.505 $Y=0.995
+ $X2=6.505 $Y2=0.56
r172 23 84 29.7123 $w=2.92e-07 $l=1.8e-07 $layer=POLY_cond $X=6.085 $Y=1.16
+ $X2=6.265 $Y2=1.16
r173 23 80 26.411 $w=2.92e-07 $l=1.6e-07 $layer=POLY_cond $X=6.085 $Y=1.16
+ $X2=5.925 $Y2=1.16
r174 23 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.085 $Y=1.295
+ $X2=6.085 $Y2=1.985
r175 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.085 $Y=1.025
+ $X2=6.085 $Y2=0.56
r176 15 80 42.9178 $w=2.92e-07 $l=2.6e-07 $layer=POLY_cond $X=5.665 $Y=1.16
+ $X2=5.925 $Y2=1.16
r177 15 76 13.2055 $w=2.92e-07 $l=8e-08 $layer=POLY_cond $X=5.665 $Y=1.16
+ $X2=5.585 $Y2=1.16
r178 15 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.665 $Y=1.295
+ $X2=5.665 $Y2=1.985
r179 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.665 $Y=1.025
+ $X2=5.665 $Y2=0.56
r180 11 74 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.325
+ $X2=5.245 $Y2=1.16
r181 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.245 $Y=1.325
+ $X2=5.245 $Y2=1.985
r182 8 74 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=0.995
+ $X2=5.245 $Y2=1.16
r183 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.245 $Y=0.995
+ $X2=5.245 $Y2=0.56
r184 4 73 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.825 $Y=1.325
+ $X2=4.825 $Y2=1.16
r185 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.825 $Y=1.325
+ $X2=4.825 $Y2=1.985
r186 1 73 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.825 $Y=0.995
+ $X2=4.825 $Y2=1.16
r187 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.825 $Y=0.995
+ $X2=4.825 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_8%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 42
+ 44 49 54 70 71 74 77 80
r121 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r122 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r123 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r125 68 71 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=8.05 $Y2=2.72
r126 67 70 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=8.05 $Y2=2.72
r127 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r128 65 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r129 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r130 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r131 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r132 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r133 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=2.72
+ $X2=2.46 $Y2=2.72
r134 59 61 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.625 $Y=2.72
+ $X2=2.99 $Y2=2.72
r135 58 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r136 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r138 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r139 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r140 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.46 $Y2=2.72
r141 54 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 53 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r143 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r144 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r145 50 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.695 $Y2=2.72
r146 50 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r147 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r148 49 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r149 44 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.695 $Y2=2.72
r150 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r151 42 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r152 42 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r153 40 64 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=3.91 $Y2=2.72
r154 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=4.14 $Y2=2.72
r155 39 67 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.37 $Y2=2.72
r156 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=2.72
+ $X2=4.14 $Y2=2.72
r157 37 61 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=2.99 $Y2=2.72
r158 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.3 $Y2=2.72
r159 36 64 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.91 $Y2=2.72
r160 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.3 $Y2=2.72
r161 32 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.72
r162 32 34 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=4.14 $Y=2.635
+ $X2=4.14 $Y2=2.02
r163 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.635 $X2=3.3
+ $Y2=2.72
r164 28 30 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.3 $Y=2.635
+ $X2=3.3 $Y2=2.02
r165 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.72
r166 24 26 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.46 $Y=2.635
+ $X2=2.46 $Y2=2.02
r167 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r168 20 22 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.02
r169 16 74 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r170 16 18 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.34
r171 5 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.005
+ $Y=1.545 $X2=4.14 $Y2=2.02
r172 4 30 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.545 $X2=3.3 $Y2=2.02
r173 3 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.325
+ $Y=1.545 $X2=2.46 $Y2=2.02
r174 2 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.545 $X2=1.62 $Y2=2.02
r175 1 18 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_8%A_215_309# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 56 57 60 62 66 68 72 74 76 79 80 81 82 83 84
c102 50 0 4.50788e-20 $X=4.475 $Y=1.64
c103 44 0 3.89415e-19 $X=3.635 $Y=1.64
c104 38 0 3.89415e-19 $X=2.795 $Y=1.64
c105 32 0 3.89415e-19 $X=1.955 $Y=1.64
r106 76 78 13.4 $w=3.05e-07 $l=3.35e-07 $layer=LI1_cond $X=8.042 $Y=2.295
+ $X2=8.042 $Y2=1.96
r107 75 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.38
+ $X2=7.135 $Y2=2.38
r108 74 76 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=7.89 $Y=2.38
+ $X2=8.042 $Y2=2.295
r109 74 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.89 $Y=2.38
+ $X2=7.22 $Y2=2.38
r110 70 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.135 $Y=2.295
+ $X2=7.135 $Y2=2.38
r111 70 72 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.135 $Y=2.295
+ $X2=7.135 $Y2=1.96
r112 69 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=2.38
+ $X2=6.295 $Y2=2.38
r113 68 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.05 $Y=2.38
+ $X2=7.135 $Y2=2.38
r114 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.05 $Y=2.38
+ $X2=6.38 $Y2=2.38
r115 64 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.295
+ $X2=6.295 $Y2=2.38
r116 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.295 $Y=2.295
+ $X2=6.295 $Y2=1.96
r117 63 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.54 $Y=2.38
+ $X2=5.455 $Y2=2.38
r118 62 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=2.38
+ $X2=6.295 $Y2=2.38
r119 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.21 $Y=2.38
+ $X2=5.54 $Y2=2.38
r120 58 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.455 $Y2=2.38
r121 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.455 $Y2=1.96
r122 56 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.37 $Y=2.38
+ $X2=5.455 $Y2=2.38
r123 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.37 $Y=2.38
+ $X2=4.7 $Y2=2.38
r124 53 57 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=4.587 $Y=2.295
+ $X2=4.7 $Y2=2.38
r125 53 55 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=4.587 $Y=2.295
+ $X2=4.587 $Y2=1.96
r126 52 55 12.0366 $w=2.23e-07 $l=2.35e-07 $layer=LI1_cond $X=4.587 $Y=1.725
+ $X2=4.587 $Y2=1.96
r127 51 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=1.64
+ $X2=3.72 $Y2=1.64
r128 50 52 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.475 $Y=1.64
+ $X2=4.587 $Y2=1.725
r129 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.475 $Y=1.64
+ $X2=3.805 $Y2=1.64
r130 46 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.725
+ $X2=3.72 $Y2=1.64
r131 46 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.72 $Y=1.725
+ $X2=3.72 $Y2=1.96
r132 45 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=1.64
+ $X2=2.88 $Y2=1.64
r133 44 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=1.64
+ $X2=3.72 $Y2=1.64
r134 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.635 $Y=1.64
+ $X2=2.965 $Y2=1.64
r135 40 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=1.725
+ $X2=2.88 $Y2=1.64
r136 40 42 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.88 $Y=1.725
+ $X2=2.88 $Y2=1.96
r137 39 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=1.64
+ $X2=2.04 $Y2=1.64
r138 38 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=1.64
+ $X2=2.88 $Y2=1.64
r139 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.795 $Y=1.64
+ $X2=2.125 $Y2=1.64
r140 34 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=1.725
+ $X2=2.04 $Y2=1.64
r141 34 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.04 $Y=1.725
+ $X2=2.04 $Y2=1.96
r142 32 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.64
+ $X2=2.04 $Y2=1.64
r143 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=1.64
+ $X2=1.285 $Y2=1.64
r144 28 33 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.18 $Y=1.725
+ $X2=1.285 $Y2=1.64
r145 28 30 27.1991 $w=2.08e-07 $l=5.15e-07 $layer=LI1_cond $X=1.18 $Y=1.725
+ $X2=1.18 $Y2=2.24
r146 9 78 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.84
+ $Y=1.485 $X2=7.975 $Y2=1.96
r147 8 72 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7
+ $Y=1.485 $X2=7.135 $Y2=1.96
r148 7 66 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.16
+ $Y=1.485 $X2=6.295 $Y2=1.96
r149 6 60 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.32
+ $Y=1.485 $X2=5.455 $Y2=1.96
r150 5 55 300 $w=1.7e-07 $l=4.90612e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.545 $X2=4.59 $Y2=1.96
r151 4 48 300 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=1.545 $X2=3.72 $Y2=1.96
r152 3 42 300 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.545 $X2=2.88 $Y2=1.96
r153 2 36 300 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.545 $X2=2.04 $Y2=1.96
r154 1 30 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.545 $X2=1.2 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_8%Z 1 2 3 4 5 6 7 8 33 35 38 39 40 41 42 43 44
+ 45 60 63 66 75 88
c97 38 0 2.25041e-19 $X=5.23 $Y=1.445
r98 88 89 3.28461 $w=3.3e-07 $l=2.55e-07 $layer=LI1_cond $X=5.875 $Y=1.87
+ $X2=5.875 $Y2=1.615
r99 86 88 2.11073 $w=5.08e-07 $l=9e-08 $layer=LI1_cond $X=5.785 $Y=1.87
+ $X2=5.875 $Y2=1.87
r100 61 63 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.25 $Y=1.53
+ $X2=5.315 $Y2=1.53
r101 44 75 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.555 $Y=1.53
+ $X2=7.39 $Y2=1.53
r102 44 45 7.48369 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=7.555 $Y=1.615
+ $X2=7.555 $Y2=1.87
r103 43 75 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.155 $Y=1.53
+ $X2=7.39 $Y2=1.53
r104 43 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.155 $Y=1.53
+ $X2=6.88 $Y2=1.53
r105 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=1.53
+ $X2=6.55 $Y2=1.53
r106 41 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=1.53
+ $X2=6.88 $Y2=1.53
r107 41 42 7.48369 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=6.715 $Y=1.615
+ $X2=6.715 $Y2=1.87
r108 40 66 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.235 $Y=1.53
+ $X2=6.55 $Y2=1.53
r109 40 67 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.235 $Y=1.53
+ $X2=6.04 $Y2=1.53
r110 39 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=1.53
+ $X2=5.875 $Y2=1.615
r111 39 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=1.53
+ $X2=5.71 $Y2=1.53
r112 39 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=1.53
+ $X2=6.04 $Y2=1.53
r113 39 86 8.07657 $w=1.5e-07 $l=2.55e-07 $layer=LI1_cond $X=5.785 $Y=1.615
+ $X2=5.785 $Y2=1.87
r114 39 60 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.7 $Y=1.53 $X2=5.71
+ $Y2=1.53
r115 38 61 4.08752 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.06 $Y=1.53
+ $X2=5.25 $Y2=1.53
r116 38 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.325 $Y=1.53
+ $X2=5.7 $Y2=1.53
r117 38 63 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.325 $Y=1.53
+ $X2=5.315 $Y2=1.53
r118 35 38 17.1828 $w=3.98e-07 $l=5.95e-07 $layer=LI1_cond $X=5.06 $Y=0.85
+ $X2=5.06 $Y2=1.445
r119 35 37 2.72589 $w=3.8e-07 $l=1.08e-07 $layer=LI1_cond $X=5.06 $Y=0.85
+ $X2=5.06 $Y2=0.742
r120 31 33 45.0257 $w=2.13e-07 $l=8.4e-07 $layer=LI1_cond $X=6.715 $Y=0.742
+ $X2=7.555 $Y2=0.742
r121 29 31 45.0257 $w=2.13e-07 $l=8.4e-07 $layer=LI1_cond $X=5.875 $Y=0.742
+ $X2=6.715 $Y2=0.742
r122 27 37 4.79554 $w=2.15e-07 $l=1.9e-07 $layer=LI1_cond $X=5.25 $Y=0.742
+ $X2=5.06 $Y2=0.742
r123 27 29 33.5013 $w=2.13e-07 $l=6.25e-07 $layer=LI1_cond $X=5.25 $Y=0.742
+ $X2=5.875 $Y2=0.742
r124 8 44 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=7.42
+ $Y=1.485 $X2=7.555 $Y2=1.61
r125 7 41 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=6.58
+ $Y=1.485 $X2=6.715 $Y2=1.61
r126 6 39 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=5.74
+ $Y=1.485 $X2=5.875 $Y2=1.61
r127 5 38 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=4.9
+ $Y=1.485 $X2=5.035 $Y2=1.61
r128 4 33 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=7.42
+ $Y=0.235 $X2=7.555 $Y2=0.76
r129 3 31 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.235 $X2=6.715 $Y2=0.76
r130 2 29 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=5.74
+ $Y=0.235 $X2=5.875 $Y2=0.76
r131 1 37 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=4.9
+ $Y=0.235 $X2=5.035 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_8%VGND 1 2 3 4 5 18 22 26 30 32 36 39 40 41 42
+ 43 45 50 67 68 71 74 77
r127 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r128 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r129 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r130 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r131 65 68 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=8.05
+ $Y2=0
r132 65 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r133 64 67 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=8.05
+ $Y2=0
r134 64 65 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r135 62 77 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.235 $Y=0 $X2=4.065
+ $Y2=0
r136 62 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.235 $Y=0
+ $X2=4.37 $Y2=0
r137 61 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r138 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r139 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r140 58 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r141 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r142 55 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.54
+ $Y2=0
r143 55 57 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r144 54 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r145 54 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r146 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r147 51 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r148 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r149 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.54
+ $Y2=0
r150 50 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.15 $Y2=0
r151 45 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r152 45 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r153 43 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r154 43 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r155 41 60 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.99
+ $Y2=0
r156 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.22
+ $Y2=0
r157 39 57 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.215 $Y=0
+ $X2=2.07 $Y2=0
r158 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=0 $X2=2.38
+ $Y2=0
r159 38 60 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=0
+ $X2=2.99 $Y2=0
r160 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.38
+ $Y2=0
r161 34 77 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0
r162 34 36 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0.36
r163 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.22
+ $Y2=0
r164 32 77 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.065
+ $Y2=0
r165 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=3.385 $Y2=0
r166 28 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0
r167 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0.36
r168 24 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=0.085
+ $X2=2.38 $Y2=0
r169 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.38 $Y=0.085
+ $X2=2.38 $Y2=0.36
r170 20 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0
r171 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.54 $Y=0.085
+ $X2=1.54 $Y2=0.36
r172 16 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r173 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r174 5 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.925
+ $Y=0.235 $X2=4.06 $Y2=0.36
r175 4 30 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.36
r176 3 26 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.36
r177 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.36
r178 1 18 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_8%A_193_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 55 56 64 66 67 68
c95 68 0 1.50055e-19 $X=3.64 $Y=0.74
c96 67 0 1.50055e-19 $X=2.8 $Y=0.74
c97 66 0 1.50055e-19 $X=1.96 $Y=0.74
c98 50 0 7.37964e-20 $X=4.405 $Y=0.74
c99 44 0 2.99402e-19 $X=3.555 $Y=0.74
c100 38 0 2.99402e-19 $X=2.715 $Y=0.74
c101 32 0 2.60168e-19 $X=1.875 $Y=0.74
r102 62 64 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=7.135 $Y=0.36
+ $X2=7.975 $Y2=0.36
r103 60 62 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=6.295 $Y=0.36
+ $X2=7.135 $Y2=0.36
r104 58 60 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=5.455 $Y=0.36
+ $X2=6.295 $Y2=0.36
r105 56 58 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=4.7 $Y=0.36
+ $X2=5.455 $Y2=0.36
r106 53 55 4.6879 $w=2.93e-07 $l=1.2e-07 $layer=LI1_cond $X=4.552 $Y=0.655
+ $X2=4.552 $Y2=0.535
r107 52 56 7.07071 $w=2.1e-07 $l=1.93505e-07 $layer=LI1_cond $X=4.552 $Y=0.465
+ $X2=4.7 $Y2=0.36
r108 52 55 2.73461 $w=2.93e-07 $l=7e-08 $layer=LI1_cond $X=4.552 $Y=0.465
+ $X2=4.552 $Y2=0.535
r109 51 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.74
+ $X2=3.64 $Y2=0.74
r110 50 53 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=4.405 $Y=0.74
+ $X2=4.552 $Y2=0.655
r111 50 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.405 $Y=0.74
+ $X2=3.725 $Y2=0.74
r112 46 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.655
+ $X2=3.64 $Y2=0.74
r113 46 48 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.64 $Y=0.655
+ $X2=3.64 $Y2=0.535
r114 45 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0.74
+ $X2=2.8 $Y2=0.74
r115 44 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0.74
+ $X2=3.64 $Y2=0.74
r116 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.555 $Y=0.74
+ $X2=2.885 $Y2=0.74
r117 40 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.655 $X2=2.8
+ $Y2=0.74
r118 40 42 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.8 $Y=0.655
+ $X2=2.8 $Y2=0.535
r119 39 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.74
+ $X2=1.96 $Y2=0.74
r120 38 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.74
+ $X2=2.8 $Y2=0.74
r121 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.715 $Y=0.74
+ $X2=2.045 $Y2=0.74
r122 34 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.655
+ $X2=1.96 $Y2=0.74
r123 34 36 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.96 $Y=0.655
+ $X2=1.96 $Y2=0.535
r124 32 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.96 $Y2=0.74
r125 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.205 $Y2=0.74
r126 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.655
+ $X2=1.205 $Y2=0.74
r127 28 30 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.12 $Y=0.655
+ $X2=1.12 $Y2=0.535
r128 9 64 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.84
+ $Y=0.235 $X2=7.975 $Y2=0.36
r129 8 62 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7
+ $Y=0.235 $X2=7.135 $Y2=0.36
r130 7 60 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.16
+ $Y=0.235 $X2=6.295 $Y2=0.36
r131 6 58 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.235 $X2=5.455 $Y2=0.36
r132 5 55 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.235 $X2=4.615 $Y2=0.535
r133 4 48 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.535
r134 3 42 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.535
r135 2 36 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.535
r136 1 30 182 $w=1.7e-07 $l=3.69459e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.12 $Y2=0.535
.ends


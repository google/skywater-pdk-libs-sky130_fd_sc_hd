* File: sky130_fd_sc_hd__o2bb2a_4.pxi.spice
* Created: Thu Aug 27 14:38:27 2020
* 
x_PM_SKY130_FD_SC_HD__O2BB2A_4%B1 N_B1_M1016_g N_B1_M1019_g N_B1_c_128_n
+ N_B1_M1027_g N_B1_M1025_g N_B1_c_136_n N_B1_c_129_n N_B1_c_130_n B1
+ N_B1_c_131_n N_B1_c_132_n N_B1_c_133_n PM_SKY130_FD_SC_HD__O2BB2A_4%B1
x_PM_SKY130_FD_SC_HD__O2BB2A_4%B2 N_B2_c_208_n N_B2_M1013_g N_B2_M1001_g
+ N_B2_c_209_n N_B2_M1018_g N_B2_M1003_g B2 N_B2_c_211_n
+ PM_SKY130_FD_SC_HD__O2BB2A_4%B2
x_PM_SKY130_FD_SC_HD__O2BB2A_4%A_415_21# N_A_415_21#_M1007_d N_A_415_21#_M1009_s
+ N_A_415_21#_M1015_d N_A_415_21#_c_256_n N_A_415_21#_M1020_g
+ N_A_415_21#_M1004_g N_A_415_21#_c_257_n N_A_415_21#_M1024_g
+ N_A_415_21#_M1022_g N_A_415_21#_c_258_n N_A_415_21#_c_259_n
+ N_A_415_21#_c_260_n N_A_415_21#_c_261_n N_A_415_21#_c_262_n
+ N_A_415_21#_c_276_p N_A_415_21#_c_330_p N_A_415_21#_c_288_p
+ N_A_415_21#_c_263_n N_A_415_21#_c_289_p N_A_415_21#_c_264_n
+ N_A_415_21#_c_265_n N_A_415_21#_c_291_p PM_SKY130_FD_SC_HD__O2BB2A_4%A_415_21#
x_PM_SKY130_FD_SC_HD__O2BB2A_4%A1_N N_A1_N_M1008_g N_A1_N_M1009_g N_A1_N_c_378_n
+ N_A1_N_M1021_g N_A1_N_M1023_g N_A1_N_c_385_n N_A1_N_c_379_n N_A1_N_c_387_n
+ N_A1_N_c_388_n A1_N N_A1_N_c_381_n N_A1_N_c_382_n
+ PM_SKY130_FD_SC_HD__O2BB2A_4%A1_N
x_PM_SKY130_FD_SC_HD__O2BB2A_4%A2_N N_A2_N_c_468_n N_A2_N_M1007_g N_A2_N_M1012_g
+ N_A2_N_c_469_n N_A2_N_M1014_g N_A2_N_M1015_g A2_N N_A2_N_c_470_n
+ N_A2_N_c_471_n PM_SKY130_FD_SC_HD__O2BB2A_4%A2_N
x_PM_SKY130_FD_SC_HD__O2BB2A_4%A_193_297# N_A_193_297#_M1020_s
+ N_A_193_297#_M1001_s N_A_193_297#_M1004_s N_A_193_297#_c_513_n
+ N_A_193_297#_M1006_g N_A_193_297#_M1000_g N_A_193_297#_c_514_n
+ N_A_193_297#_M1010_g N_A_193_297#_M1002_g N_A_193_297#_c_515_n
+ N_A_193_297#_M1011_g N_A_193_297#_M1005_g N_A_193_297#_c_516_n
+ N_A_193_297#_M1017_g N_A_193_297#_M1026_g N_A_193_297#_c_531_n
+ N_A_193_297#_c_517_n N_A_193_297#_c_572_n N_A_193_297#_c_619_p
+ N_A_193_297#_c_536_n N_A_193_297#_c_548_n N_A_193_297#_c_524_n
+ N_A_193_297#_c_525_n N_A_193_297#_c_526_n N_A_193_297#_c_527_n
+ N_A_193_297#_c_518_n N_A_193_297#_c_519_n
+ PM_SKY130_FD_SC_HD__O2BB2A_4%A_193_297#
x_PM_SKY130_FD_SC_HD__O2BB2A_4%VPWR N_VPWR_M1019_s N_VPWR_M1025_s N_VPWR_M1022_d
+ N_VPWR_M1012_s N_VPWR_M1023_d N_VPWR_M1002_s N_VPWR_M1026_s N_VPWR_c_671_n
+ N_VPWR_c_672_n N_VPWR_c_673_n N_VPWR_c_674_n N_VPWR_c_675_n N_VPWR_c_676_n
+ N_VPWR_c_677_n N_VPWR_c_678_n N_VPWR_c_679_n N_VPWR_c_680_n N_VPWR_c_681_n
+ N_VPWR_c_682_n N_VPWR_c_683_n N_VPWR_c_684_n VPWR N_VPWR_c_685_n
+ N_VPWR_c_686_n N_VPWR_c_670_n N_VPWR_c_688_n N_VPWR_c_689_n N_VPWR_c_690_n
+ N_VPWR_c_691_n PM_SKY130_FD_SC_HD__O2BB2A_4%VPWR
x_PM_SKY130_FD_SC_HD__O2BB2A_4%A_109_297# N_A_109_297#_M1019_d
+ N_A_109_297#_M1003_d N_A_109_297#_c_792_n N_A_109_297#_c_793_n
+ N_A_109_297#_c_804_n N_A_109_297#_c_799_n
+ PM_SKY130_FD_SC_HD__O2BB2A_4%A_109_297#
x_PM_SKY130_FD_SC_HD__O2BB2A_4%X N_X_M1006_d N_X_M1011_d N_X_M1000_d N_X_M1005_d
+ N_X_c_817_n N_X_c_856_n N_X_c_820_n N_X_c_824_n N_X_c_808_n N_X_c_809_n
+ N_X_c_838_n N_X_c_861_n N_X_c_810_n N_X_c_811_n X X
+ PM_SKY130_FD_SC_HD__O2BB2A_4%X
x_PM_SKY130_FD_SC_HD__O2BB2A_4%A_27_47# N_A_27_47#_M1016_d N_A_27_47#_M1013_d
+ N_A_27_47#_M1027_d N_A_27_47#_M1024_d N_A_27_47#_c_882_n N_A_27_47#_c_883_n
+ N_A_27_47#_c_884_n N_A_27_47#_c_895_n N_A_27_47#_c_885_n N_A_27_47#_c_901_n
+ N_A_27_47#_c_902_n N_A_27_47#_c_886_n N_A_27_47#_c_887_n
+ PM_SKY130_FD_SC_HD__O2BB2A_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O2BB2A_4%VGND N_VGND_M1016_s N_VGND_M1018_s N_VGND_M1008_s
+ N_VGND_M1021_s N_VGND_M1010_s N_VGND_M1017_s N_VGND_c_946_n N_VGND_c_947_n
+ N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n N_VGND_c_952_n
+ N_VGND_c_953_n N_VGND_c_954_n N_VGND_c_955_n N_VGND_c_956_n N_VGND_c_957_n
+ N_VGND_c_958_n N_VGND_c_959_n N_VGND_c_960_n N_VGND_c_961_n N_VGND_c_962_n
+ VGND N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n
+ PM_SKY130_FD_SC_HD__O2BB2A_4%VGND
x_PM_SKY130_FD_SC_HD__O2BB2A_4%A_717_47# N_A_717_47#_M1008_d N_A_717_47#_M1014_s
+ N_A_717_47#_c_1066_n N_A_717_47#_c_1071_n N_A_717_47#_c_1064_n
+ PM_SKY130_FD_SC_HD__O2BB2A_4%A_717_47#
cc_1 VNB N_B1_c_128_n 0.0162167f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_2 VNB N_B1_c_129_n 0.00357799f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_3 VNB N_B1_c_130_n 0.0190067f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_4 VNB N_B1_c_131_n 0.0267423f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_5 VNB N_B1_c_132_n 0.0131186f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_6 VNB N_B1_c_133_n 0.021688f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_7 VNB N_B2_c_208_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_B2_c_209_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_9 VNB B2 0.0015816f $X=-0.19 $Y=-0.24 $X2=1.565 $Y2=1.53
cc_10 VNB N_B2_c_211_n 0.0308136f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_11 VNB N_A_415_21#_c_256_n 0.01577f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_12 VNB N_A_415_21#_c_257_n 0.0194896f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.445
cc_13 VNB N_A_415_21#_c_258_n 6.87055e-19 $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_14 VNB N_A_415_21#_c_259_n 0.0496516f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_15 VNB N_A_415_21#_c_260_n 0.00338858f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_16 VNB N_A_415_21#_c_261_n 9.04747e-19 $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.19
cc_17 VNB N_A_415_21#_c_262_n 0.0057395f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.53
cc_18 VNB N_A_415_21#_c_263_n 0.00115914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_415_21#_c_264_n 0.00206877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_415_21#_c_265_n 0.00710224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A1_N_c_378_n 0.016414f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_22 VNB N_A1_N_c_379_n 0.027267f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_23 VNB A1_N 0.00383212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A1_N_c_381_n 0.0196192f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_25 VNB N_A1_N_c_382_n 0.0204331f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_26 VNB N_A2_N_c_468_n 0.0160171f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_27 VNB N_A2_N_c_469_n 0.0161504f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_28 VNB N_A2_N_c_470_n 0.00334158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A2_N_c_471_n 0.0286689f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_30 VNB N_A_193_297#_c_513_n 0.0161462f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_31 VNB N_A_193_297#_c_514_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.445
cc_32 VNB N_A_193_297#_c_515_n 0.0157971f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_33 VNB N_A_193_297#_c_516_n 0.0191578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_193_297#_c_517_n 9.40276e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_193_297#_c_518_n 0.0657138f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_193_297#_c_519_n 0.00158183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_670_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_808_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_809_n 0.00211281f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_40 VNB N_X_c_810_n 0.0110739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_X_c_811_n 0.00222406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB X 0.0214978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_c_882_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=1.565 $Y2=1.53
cc_44 VNB N_A_27_47#_c_883_n 0.00382625f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.445
cc_45 VNB N_A_27_47#_c_884_n 0.0100021f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_46 VNB N_A_27_47#_c_885_n 0.00938439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_27_47#_c_886_n 0.00298253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_27_47#_c_887_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_946_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_947_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_51 VNB N_VGND_c_948_n 0.00469239f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_52 VNB N_VGND_c_949_n 0.00682968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_950_n 0.0176493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_951_n 0.00359433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_952_n 0.00416791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_953_n 0.0172255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_954_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_955_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_956_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_957_n 0.0382271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_958_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_959_n 0.0373934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_960_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_961_n 0.017009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_962_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_963_n 0.0211037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_964_n 0.371806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_965_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_717_47#_c_1064_n 0.00249478f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_70 VPB N_B1_M1019_g 0.0223957f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_71 VPB N_B1_M1025_g 0.0172429f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_72 VPB N_B1_c_136_n 0.008734f $X=-0.19 $Y=1.305 $X2=1.565 $Y2=1.53
cc_73 VPB N_B1_c_129_n 0.00229153f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_74 VPB N_B1_c_130_n 0.00441099f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_75 VPB N_B1_c_131_n 0.00483422f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_76 VPB N_B1_c_132_n 0.0160332f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_77 VPB N_B2_M1001_g 0.0183629f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_78 VPB N_B2_M1003_g 0.0183559f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_79 VPB N_B2_c_211_n 0.00405369f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_80 VPB N_A_415_21#_M1004_g 0.0172006f $X=-0.19 $Y=1.305 $X2=1.565 $Y2=1.53
cc_81 VPB N_A_415_21#_M1022_g 0.0227001f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_82 VPB N_A_415_21#_c_259_n 0.0154948f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=0.995
cc_83 VPB N_A_415_21#_c_261_n 0.00306758f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.19
cc_84 VPB N_A1_N_M1009_g 0.0223541f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_85 VPB N_A1_N_M1023_g 0.0172429f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_86 VPB N_A1_N_c_385_n 0.00220361f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.445
cc_87 VPB N_A1_N_c_379_n 0.00655096f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_88 VPB N_A1_N_c_387_n 0.00871758f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_89 VPB N_A1_N_c_388_n 2.03604e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB A1_N 0.00232127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A1_N_c_382_n 0.00441099f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_92 VPB N_A2_N_M1012_g 0.0183412f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_93 VPB N_A2_N_M1015_g 0.0183385f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_94 VPB N_A2_N_c_471_n 0.00400439f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_95 VPB N_A_193_297#_M1000_g 0.0179782f $X=-0.19 $Y=1.305 $X2=1.565 $Y2=1.53
cc_96 VPB N_A_193_297#_M1002_g 0.0184574f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_97 VPB N_A_193_297#_M1005_g 0.0184765f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_98 VPB N_A_193_297#_M1026_g 0.0220575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_193_297#_c_524_n 0.00686111f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_193_297#_c_525_n 0.00119374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_193_297#_c_526_n 0.00106182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_193_297#_c_527_n 0.00152765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_193_297#_c_518_n 0.0111791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_193_297#_c_519_n 0.00235068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_671_n 0.010584f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_106 VPB N_VPWR_c_672_n 0.00492706f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_107 VPB N_VPWR_c_673_n 0.00459443f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.325
cc_108 VPB N_VPWR_c_674_n 0.0039289f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.19
cc_109 VPB N_VPWR_c_675_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_676_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_677_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_678_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_679_n 0.0362026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_680_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_681_n 0.0163086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_682_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_683_n 0.0157745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_684_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_685_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_686_n 0.0204409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_670_n 0.0650773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_688_n 0.0168209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_689_n 0.0206381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_690_n 0.00478125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_691_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB X 0.00591752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB X 0.0201413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 N_B1_c_133_n N_B2_c_208_n 0.0234927f $X=0.41 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_129 N_B1_M1019_g N_B2_M1001_g 0.0234927f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_130 N_B1_c_136_n N_B2_M1001_g 0.0145375f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_131 N_B1_c_128_n N_B2_c_209_n 0.0258191f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_M1025_g N_B2_M1003_g 0.043521f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_133 N_B1_c_136_n N_B2_M1003_g 0.0107644f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_134 N_B1_c_136_n B2 0.0381541f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_135 N_B1_c_129_n B2 0.0134455f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B1_c_130_n B2 2.20976e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_137 N_B1_c_131_n B2 7.59344e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_138 N_B1_c_132_n B2 0.0143152f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B1_c_136_n N_B2_c_211_n 0.00214031f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_140 N_B1_c_129_n N_B2_c_211_n 0.00527477f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B1_c_130_n N_B2_c_211_n 0.022397f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B1_c_131_n N_B2_c_211_n 0.0234927f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_143 N_B1_c_132_n N_B2_c_211_n 0.00483648f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B1_c_128_n N_A_415_21#_c_256_n 0.0118576f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B1_M1025_g N_A_415_21#_M1004_g 0.0429632f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_146 N_B1_c_136_n N_A_415_21#_M1004_g 6.60451e-19 $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_147 N_B1_c_129_n N_A_415_21#_c_259_n 0.00120189f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B1_c_130_n N_A_415_21#_c_259_n 0.0220852f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_149 N_B1_c_136_n N_A_193_297#_M1001_s 0.00165831f $X=1.565 $Y=1.53 $X2=0
+ $Y2=0
cc_150 N_B1_M1025_g N_A_193_297#_c_531_n 0.0115072f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B1_c_136_n N_A_193_297#_c_531_n 0.0355123f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_152 N_B1_c_130_n N_A_193_297#_c_531_n 3.01349e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_153 N_B1_c_128_n N_A_193_297#_c_517_n 4.41707e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_B1_c_130_n N_A_193_297#_c_517_n 4.25752e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B1_c_136_n N_A_193_297#_c_536_n 0.0120079f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B1_c_136_n N_A_193_297#_c_525_n 7.23574e-19 $X=1.565 $Y=1.53 $X2=0
+ $Y2=0
cc_157 N_B1_M1025_g N_A_193_297#_c_519_n 5.62413e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_B1_c_136_n N_A_193_297#_c_519_n 0.00895055f $X=1.565 $Y=1.53 $X2=0
+ $Y2=0
cc_159 N_B1_c_129_n N_A_193_297#_c_519_n 0.0312176f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B1_c_130_n N_A_193_297#_c_519_n 7.85686e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_161 N_B1_c_132_n N_VPWR_M1019_s 0.00296816f $X=0.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_162 N_B1_c_136_n N_VPWR_M1025_s 0.00145947f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_163 N_B1_M1019_g N_VPWR_c_672_n 0.00443865f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_164 N_B1_c_131_n N_VPWR_c_672_n 2.81509e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_132_n N_VPWR_c_672_n 0.0167281f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_166 N_B1_M1025_g N_VPWR_c_673_n 0.00302074f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_167 N_B1_M1019_g N_VPWR_c_679_n 0.00585385f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_168 N_B1_M1025_g N_VPWR_c_679_n 0.00585385f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_169 N_B1_M1019_g N_VPWR_c_670_n 0.0115185f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_170 N_B1_M1025_g N_VPWR_c_670_n 0.00593924f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_171 N_B1_c_136_n N_A_109_297#_M1019_d 0.00165831f $X=1.565 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_172 N_B1_c_136_n N_A_109_297#_M1003_d 0.00165255f $X=1.565 $Y=1.53 $X2=0
+ $Y2=0
cc_173 N_B1_c_136_n N_A_109_297#_c_792_n 0.0126919f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_174 N_B1_c_133_n N_A_27_47#_c_882_n 0.00630972f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B1_c_136_n N_A_27_47#_c_883_n 0.00780885f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_176 N_B1_c_132_n N_A_27_47#_c_883_n 0.0113814f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_177 N_B1_c_133_n N_A_27_47#_c_883_n 0.00865195f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B1_c_131_n N_A_27_47#_c_884_n 0.0030689f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B1_c_132_n N_A_27_47#_c_884_n 0.0294933f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B1_c_133_n N_A_27_47#_c_884_n 0.00129412f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B1_c_128_n N_A_27_47#_c_895_n 5.22228e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B1_c_133_n N_A_27_47#_c_895_n 5.22228e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B1_c_128_n N_A_27_47#_c_885_n 0.00951765f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B1_c_136_n N_A_27_47#_c_885_n 0.0071189f $X=1.565 $Y=1.53 $X2=0 $Y2=0
cc_185 N_B1_c_129_n N_A_27_47#_c_885_n 0.0264344f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_186 N_B1_c_130_n N_A_27_47#_c_885_n 0.00301245f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_187 N_B1_c_128_n N_A_27_47#_c_901_n 0.00255288f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_128_n N_A_27_47#_c_902_n 0.00393886f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_133_n N_VGND_c_946_n 0.00268723f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B1_c_128_n N_VGND_c_947_n 0.00268723f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_191 N_B1_c_133_n N_VGND_c_953_n 0.00423334f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_192 N_B1_c_128_n N_VGND_c_957_n 0.00422898f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B1_c_128_n N_VGND_c_964_n 0.00579955f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B1_c_133_n N_VGND_c_964_n 0.00669771f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B2_M1003_g N_A_193_297#_c_531_n 0.00924026f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_B2_M1001_g N_VPWR_c_679_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B2_M1003_g N_VPWR_c_679_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B2_M1001_g N_VPWR_c_670_n 0.00525237f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B2_M1003_g N_VPWR_c_670_n 0.00525237f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B2_M1001_g N_A_109_297#_c_793_n 0.0121306f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_201 N_B2_M1003_g N_A_109_297#_c_793_n 0.00851673f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_202 N_B2_c_208_n N_A_27_47#_c_882_n 5.22228e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B2_c_208_n N_A_27_47#_c_883_n 0.00865686f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_204 B2 N_A_27_47#_c_883_n 0.00900407f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_205 N_B2_c_208_n N_A_27_47#_c_895_n 0.00630972f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B2_c_209_n N_A_27_47#_c_895_n 0.00630972f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B2_c_209_n N_A_27_47#_c_885_n 0.00894278f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_208 B2 N_A_27_47#_c_885_n 0.00545718f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_209 N_B2_c_209_n N_A_27_47#_c_902_n 4.87589e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B2_c_208_n N_A_27_47#_c_887_n 0.00113286f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B2_c_209_n N_A_27_47#_c_887_n 0.00128009f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_212 B2 N_A_27_47#_c_887_n 0.0265405f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_213 N_B2_c_211_n N_A_27_47#_c_887_n 0.00230339f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_214 N_B2_c_208_n N_VGND_c_946_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B2_c_209_n N_VGND_c_947_n 0.00146448f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B2_c_208_n N_VGND_c_955_n 0.00423334f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B2_c_209_n N_VGND_c_955_n 0.00424416f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B2_c_208_n N_VGND_c_964_n 0.0057435f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B2_c_209_n N_VGND_c_964_n 0.00576327f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_415_21#_c_261_n N_A1_N_M1009_g 0.00665142f $X=3.05 $Y=1.785 $X2=0
+ $Y2=0
cc_221 N_A_415_21#_c_276_p N_A1_N_M1009_g 0.0123266f $X=3.595 $Y=1.875 $X2=0
+ $Y2=0
cc_222 N_A_415_21#_c_261_n N_A1_N_c_385_n 0.0155745f $X=3.05 $Y=1.785 $X2=0
+ $Y2=0
cc_223 N_A_415_21#_c_263_n N_A1_N_c_385_n 0.0140485f $X=3.05 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_415_21#_c_265_n N_A1_N_c_385_n 0.0245987f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_225 N_A_415_21#_c_259_n N_A1_N_c_379_n 0.00912582f $X=2.78 $Y=1.16 $X2=0
+ $Y2=0
cc_226 N_A_415_21#_c_260_n N_A1_N_c_379_n 0.00182346f $X=3.05 $Y=1.075 $X2=0
+ $Y2=0
cc_227 N_A_415_21#_c_261_n N_A1_N_c_379_n 5.95846e-19 $X=3.05 $Y=1.785 $X2=0
+ $Y2=0
cc_228 N_A_415_21#_c_276_p N_A1_N_c_379_n 3.71138e-19 $X=3.595 $Y=1.875 $X2=0
+ $Y2=0
cc_229 N_A_415_21#_c_263_n N_A1_N_c_379_n 0.00137346f $X=3.05 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_415_21#_c_265_n N_A1_N_c_379_n 0.00447326f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_231 N_A_415_21#_M1009_s N_A1_N_c_387_n 0.00161579f $X=3.585 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_415_21#_M1015_d N_A1_N_c_387_n 0.00164852f $X=4.425 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_A_415_21#_c_288_p N_A1_N_c_387_n 0.0288156f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_234 N_A_415_21#_c_289_p N_A1_N_c_387_n 0.0106118f $X=3.72 $Y=1.875 $X2=0
+ $Y2=0
cc_235 N_A_415_21#_c_265_n N_A1_N_c_387_n 0.00458181f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_236 N_A_415_21#_c_291_p N_A1_N_c_387_n 0.0116235f $X=4.56 $Y=1.96 $X2=0 $Y2=0
cc_237 N_A_415_21#_c_261_n N_A1_N_c_388_n 0.0124042f $X=3.05 $Y=1.785 $X2=0
+ $Y2=0
cc_238 N_A_415_21#_c_276_p N_A1_N_c_388_n 0.0149193f $X=3.595 $Y=1.875 $X2=0
+ $Y2=0
cc_239 N_A_415_21#_c_289_p N_A1_N_c_388_n 2.32234e-19 $X=3.72 $Y=1.875 $X2=0
+ $Y2=0
cc_240 N_A_415_21#_c_260_n N_A1_N_c_381_n 0.00271538f $X=3.05 $Y=1.075 $X2=0
+ $Y2=0
cc_241 N_A_415_21#_c_264_n N_A1_N_c_381_n 3.91234e-19 $X=4.14 $Y=0.73 $X2=0
+ $Y2=0
cc_242 N_A_415_21#_c_265_n N_A1_N_c_381_n 0.0140908f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_243 N_A_415_21#_c_264_n N_A2_N_c_468_n 0.00298393f $X=4.14 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_415_21#_c_265_n N_A2_N_c_468_n 0.00762189f $X=3.975 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_245 N_A_415_21#_c_288_p N_A2_N_M1012_g 0.0103689f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_246 N_A_415_21#_c_264_n N_A2_N_c_469_n 0.00381491f $X=4.14 $Y=0.73 $X2=0
+ $Y2=0
cc_247 N_A_415_21#_c_288_p N_A2_N_M1015_g 0.0103689f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_248 N_A_415_21#_c_265_n N_A2_N_c_470_n 0.034704f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_249 N_A_415_21#_c_264_n N_A2_N_c_471_n 0.00224214f $X=4.14 $Y=0.73 $X2=0
+ $Y2=0
cc_250 N_A_415_21#_c_256_n N_A_193_297#_c_517_n 0.00347918f $X=2.15 $Y=0.995
+ $X2=0 $Y2=0
cc_251 N_A_415_21#_c_257_n N_A_193_297#_c_517_n 0.00131112f $X=2.57 $Y=0.995
+ $X2=0 $Y2=0
cc_252 N_A_415_21#_c_259_n N_A_193_297#_c_517_n 0.00666811f $X=2.78 $Y=1.16
+ $X2=0 $Y2=0
cc_253 N_A_415_21#_c_260_n N_A_193_297#_c_517_n 0.00580513f $X=3.05 $Y=1.075
+ $X2=0 $Y2=0
cc_254 N_A_415_21#_c_262_n N_A_193_297#_c_517_n 0.00230097f $X=3.145 $Y=0.815
+ $X2=0 $Y2=0
cc_255 N_A_415_21#_c_256_n N_A_193_297#_c_548_n 0.00217268f $X=2.15 $Y=0.995
+ $X2=0 $Y2=0
cc_256 N_A_415_21#_c_257_n N_A_193_297#_c_548_n 0.00618959f $X=2.57 $Y=0.995
+ $X2=0 $Y2=0
cc_257 N_A_415_21#_c_262_n N_A_193_297#_c_548_n 0.00379909f $X=3.145 $Y=0.815
+ $X2=0 $Y2=0
cc_258 N_A_415_21#_c_258_n N_A_193_297#_c_524_n 0.0111482f $X=2.955 $Y=1.16
+ $X2=0 $Y2=0
cc_259 N_A_415_21#_c_259_n N_A_193_297#_c_524_n 0.00639596f $X=2.78 $Y=1.16
+ $X2=0 $Y2=0
cc_260 N_A_415_21#_c_261_n N_A_193_297#_c_524_n 0.0201205f $X=3.05 $Y=1.785
+ $X2=0 $Y2=0
cc_261 N_A_415_21#_c_276_p N_A_193_297#_c_524_n 0.0096537f $X=3.595 $Y=1.875
+ $X2=0 $Y2=0
cc_262 N_A_415_21#_c_288_p N_A_193_297#_c_524_n 0.00428749f $X=4.435 $Y=1.875
+ $X2=0 $Y2=0
cc_263 N_A_415_21#_c_289_p N_A_193_297#_c_524_n 0.00195811f $X=3.72 $Y=1.875
+ $X2=0 $Y2=0
cc_264 N_A_415_21#_c_265_n N_A_193_297#_c_524_n 0.00835128f $X=3.975 $Y=0.775
+ $X2=0 $Y2=0
cc_265 N_A_415_21#_c_291_p N_A_193_297#_c_524_n 0.00209035f $X=4.56 $Y=1.96
+ $X2=0 $Y2=0
cc_266 N_A_415_21#_M1022_g N_A_193_297#_c_525_n 0.00894358f $X=2.57 $Y=1.985
+ $X2=0 $Y2=0
cc_267 N_A_415_21#_c_258_n N_A_193_297#_c_525_n 0.00252139f $X=2.955 $Y=1.16
+ $X2=0 $Y2=0
cc_268 N_A_415_21#_c_259_n N_A_193_297#_c_525_n 8.13808e-19 $X=2.78 $Y=1.16
+ $X2=0 $Y2=0
cc_269 N_A_415_21#_c_261_n N_A_193_297#_c_525_n 0.00248394f $X=3.05 $Y=1.785
+ $X2=0 $Y2=0
cc_270 N_A_415_21#_M1004_g N_A_193_297#_c_519_n 0.0174919f $X=2.15 $Y=1.985
+ $X2=0 $Y2=0
cc_271 N_A_415_21#_M1022_g N_A_193_297#_c_519_n 0.0286386f $X=2.57 $Y=1.985
+ $X2=0 $Y2=0
cc_272 N_A_415_21#_c_258_n N_A_193_297#_c_519_n 0.0133541f $X=2.955 $Y=1.16
+ $X2=0 $Y2=0
cc_273 N_A_415_21#_c_259_n N_A_193_297#_c_519_n 0.0189574f $X=2.78 $Y=1.16 $X2=0
+ $Y2=0
cc_274 N_A_415_21#_c_261_n N_A_193_297#_c_519_n 0.0193649f $X=3.05 $Y=1.785
+ $X2=0 $Y2=0
cc_275 N_A_415_21#_c_330_p N_A_193_297#_c_519_n 0.00913982f $X=3.145 $Y=1.875
+ $X2=0 $Y2=0
cc_276 N_A_415_21#_c_261_n N_VPWR_M1022_d 0.00909039f $X=3.05 $Y=1.785 $X2=0
+ $Y2=0
cc_277 N_A_415_21#_c_276_p N_VPWR_M1022_d 0.0062656f $X=3.595 $Y=1.875 $X2=0
+ $Y2=0
cc_278 N_A_415_21#_c_330_p N_VPWR_M1022_d 0.00612176f $X=3.145 $Y=1.875 $X2=0
+ $Y2=0
cc_279 N_A_415_21#_c_288_p N_VPWR_M1012_s 0.00303737f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_280 N_A_415_21#_M1004_g N_VPWR_c_673_n 0.00162987f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_A_415_21#_c_288_p N_VPWR_c_674_n 0.0119173f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_282 N_A_415_21#_c_276_p N_VPWR_c_681_n 0.0020229f $X=3.595 $Y=1.875 $X2=0
+ $Y2=0
cc_283 N_A_415_21#_c_288_p N_VPWR_c_681_n 0.0020229f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_284 N_A_415_21#_c_289_p N_VPWR_c_681_n 0.00414246f $X=3.72 $Y=1.875 $X2=0
+ $Y2=0
cc_285 N_A_415_21#_c_288_p N_VPWR_c_683_n 0.0020229f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_286 N_A_415_21#_c_291_p N_VPWR_c_683_n 0.0142343f $X=4.56 $Y=1.96 $X2=0 $Y2=0
cc_287 N_A_415_21#_M1009_s N_VPWR_c_670_n 0.00302071f $X=3.585 $Y=1.485 $X2=0
+ $Y2=0
cc_288 N_A_415_21#_M1015_d N_VPWR_c_670_n 0.00253991f $X=4.425 $Y=1.485 $X2=0
+ $Y2=0
cc_289 N_A_415_21#_M1004_g N_VPWR_c_670_n 0.00590957f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_A_415_21#_M1022_g N_VPWR_c_670_n 0.00799454f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_291 N_A_415_21#_c_276_p N_VPWR_c_670_n 0.00460674f $X=3.595 $Y=1.875 $X2=0
+ $Y2=0
cc_292 N_A_415_21#_c_330_p N_VPWR_c_670_n 7.8019e-19 $X=3.145 $Y=1.875 $X2=0
+ $Y2=0
cc_293 N_A_415_21#_c_288_p N_VPWR_c_670_n 0.00806641f $X=4.435 $Y=1.875 $X2=0
+ $Y2=0
cc_294 N_A_415_21#_c_289_p N_VPWR_c_670_n 0.00745459f $X=3.72 $Y=1.875 $X2=0
+ $Y2=0
cc_295 N_A_415_21#_c_291_p N_VPWR_c_670_n 0.00955092f $X=4.56 $Y=1.96 $X2=0
+ $Y2=0
cc_296 N_A_415_21#_M1004_g N_VPWR_c_688_n 0.00585385f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_A_415_21#_M1022_g N_VPWR_c_688_n 0.00455174f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_415_21#_M1022_g N_VPWR_c_689_n 0.00331225f $X=2.57 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A_415_21#_c_276_p N_VPWR_c_689_n 0.0176659f $X=3.595 $Y=1.875 $X2=0
+ $Y2=0
cc_300 N_A_415_21#_c_330_p N_VPWR_c_689_n 0.015863f $X=3.145 $Y=1.875 $X2=0
+ $Y2=0
cc_301 N_A_415_21#_c_256_n N_A_27_47#_c_886_n 0.010549f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_415_21#_c_257_n N_A_27_47#_c_886_n 0.0122128f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_415_21#_c_258_n N_A_27_47#_c_886_n 0.00797286f $X=2.955 $Y=1.16 $X2=0
+ $Y2=0
cc_304 N_A_415_21#_c_259_n N_A_27_47#_c_886_n 0.00525812f $X=2.78 $Y=1.16 $X2=0
+ $Y2=0
cc_305 N_A_415_21#_c_265_n N_VGND_M1008_s 0.00315681f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_306 N_A_415_21#_c_257_n N_VGND_c_948_n 0.0019578f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_415_21#_c_265_n N_VGND_c_948_n 0.0127273f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_308 N_A_415_21#_c_256_n N_VGND_c_957_n 0.00357877f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_415_21#_c_257_n N_VGND_c_957_n 0.00357877f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_A_415_21#_c_262_n N_VGND_c_957_n 0.00323451f $X=3.145 $Y=0.815 $X2=0
+ $Y2=0
cc_311 N_A_415_21#_c_265_n N_VGND_c_957_n 0.00102539f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_312 N_A_415_21#_c_265_n N_VGND_c_959_n 0.00199263f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_313 N_A_415_21#_M1007_d N_VGND_c_964_n 0.00220248f $X=4.005 $Y=0.235 $X2=0
+ $Y2=0
cc_314 N_A_415_21#_c_256_n N_VGND_c_964_n 0.00525237f $X=2.15 $Y=0.995 $X2=0
+ $Y2=0
cc_315 N_A_415_21#_c_257_n N_VGND_c_964_n 0.00655123f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_316 N_A_415_21#_c_262_n N_VGND_c_964_n 0.00534938f $X=3.145 $Y=0.815 $X2=0
+ $Y2=0
cc_317 N_A_415_21#_c_265_n N_VGND_c_964_n 0.00733587f $X=3.975 $Y=0.775 $X2=0
+ $Y2=0
cc_318 N_A_415_21#_c_265_n N_A_717_47#_M1008_d 0.00191752f $X=3.975 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_319 N_A_415_21#_M1007_d N_A_717_47#_c_1066_n 0.00318958f $X=4.005 $Y=0.235
+ $X2=0 $Y2=0
cc_320 N_A_415_21#_c_264_n N_A_717_47#_c_1066_n 0.015032f $X=4.14 $Y=0.73 $X2=0
+ $Y2=0
cc_321 N_A_415_21#_c_265_n N_A_717_47#_c_1066_n 0.014624f $X=3.975 $Y=0.775
+ $X2=0 $Y2=0
cc_322 N_A_415_21#_c_264_n N_A_717_47#_c_1064_n 0.0105027f $X=4.14 $Y=0.73 $X2=0
+ $Y2=0
cc_323 N_A1_N_c_381_n N_A2_N_c_468_n 0.0269138f $X=3.48 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_324 N_A1_N_M1009_g N_A2_N_M1012_g 0.0420013f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A1_N_c_385_n N_A2_N_M1012_g 0.00265828f $X=3.48 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A1_N_c_387_n N_A2_N_M1012_g 0.0103235f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_327 N_A1_N_c_378_n N_A2_N_c_469_n 0.012379f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A1_N_M1023_g N_A2_N_M1015_g 0.0277801f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A1_N_c_387_n N_A2_N_M1015_g 0.0103235f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_330 N_A1_N_c_385_n N_A2_N_c_470_n 0.0165706f $X=3.48 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A1_N_c_379_n N_A2_N_c_470_n 0.00119401f $X=3.48 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A1_N_c_387_n N_A2_N_c_470_n 0.0399588f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_333 A1_N N_A2_N_c_470_n 0.0174911f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_334 N_A1_N_c_382_n N_A2_N_c_470_n 6.80324e-19 $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A1_N_c_385_n N_A2_N_c_471_n 6.0934e-19 $X=3.48 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A1_N_c_379_n N_A2_N_c_471_n 0.0222728f $X=3.48 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A1_N_c_387_n N_A2_N_c_471_n 0.00214031f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_338 A1_N N_A2_N_c_471_n 0.00465908f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_339 N_A1_N_c_382_n N_A2_N_c_471_n 0.0223771f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A1_N_c_378_n N_A_193_297#_c_513_n 0.0123221f $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A1_N_M1023_g N_A_193_297#_M1000_g 0.0279096f $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A1_N_c_387_n N_A_193_297#_M1000_g 9.45935e-19 $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_343 A1_N N_A_193_297#_c_572_n 0.0126993f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_344 N_A1_N_c_387_n N_A_193_297#_c_524_n 0.0657556f $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_345 N_A1_N_c_388_n N_A_193_297#_c_524_n 0.0162437f $X=3.645 $Y=1.53 $X2=0
+ $Y2=0
cc_346 N_A1_N_c_387_n N_A_193_297#_c_526_n 7.58576e-19 $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_347 A1_N N_A_193_297#_c_526_n 7.39655e-19 $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_348 N_A1_N_M1023_g N_A_193_297#_c_527_n 3.87046e-19 $X=4.77 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A1_N_c_387_n N_A_193_297#_c_527_n 0.00983194f $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_350 A1_N N_A_193_297#_c_527_n 0.0134769f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_351 A1_N N_A_193_297#_c_518_n 0.00251711f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_352 N_A1_N_c_382_n N_A_193_297#_c_518_n 0.02273f $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A1_N_c_388_n N_VPWR_M1022_d 0.00138147f $X=3.645 $Y=1.53 $X2=0 $Y2=0
cc_354 N_A1_N_c_387_n N_VPWR_M1012_s 0.00166235f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_355 N_A1_N_c_387_n N_VPWR_M1023_d 0.0014624f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_356 N_A1_N_M1023_g N_VPWR_c_675_n 0.00157837f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_357 N_A1_N_c_387_n N_VPWR_c_675_n 0.0048223f $X=4.605 $Y=1.53 $X2=0 $Y2=0
cc_358 N_A1_N_M1009_g N_VPWR_c_681_n 0.00441875f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_359 N_A1_N_M1023_g N_VPWR_c_683_n 0.00585385f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A1_N_M1009_g N_VPWR_c_670_n 0.00725698f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A1_N_M1023_g N_VPWR_c_670_n 0.0104912f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A1_N_M1009_g N_VPWR_c_689_n 0.00353572f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A1_N_c_381_n N_VGND_c_948_n 0.00438629f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A1_N_c_378_n N_VGND_c_949_n 0.00275369f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_365 A1_N N_VGND_c_949_n 0.0057781f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_366 N_A1_N_c_382_n N_VGND_c_949_n 2.29798e-19 $X=4.77 $Y=1.16 $X2=0 $Y2=0
cc_367 N_A1_N_c_378_n N_VGND_c_959_n 0.00541892f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A1_N_c_381_n N_VGND_c_959_n 0.00423906f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A1_N_c_378_n N_VGND_c_964_n 0.00952298f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A1_N_c_381_n N_VGND_c_964_n 0.0070828f $X=3.48 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A1_N_c_381_n N_A_717_47#_c_1066_n 0.00265651f $X=3.48 $Y=0.995 $X2=0
+ $Y2=0
cc_372 N_A1_N_c_378_n N_A_717_47#_c_1071_n 0.00208315f $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_373 N_A1_N_c_378_n N_A_717_47#_c_1064_n 0.00487681f $X=4.77 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_A1_N_c_387_n N_A_717_47#_c_1064_n 0.00368291f $X=4.605 $Y=1.53 $X2=0
+ $Y2=0
cc_375 A1_N N_A_717_47#_c_1064_n 0.00947365f $X=4.765 $Y=1.105 $X2=0 $Y2=0
cc_376 N_A1_N_c_382_n N_A_717_47#_c_1064_n 0.00152217f $X=4.77 $Y=1.16 $X2=0
+ $Y2=0
cc_377 N_A2_N_c_470_n N_A_193_297#_c_524_n 0.00443567f $X=4.145 $Y=1.16 $X2=0
+ $Y2=0
cc_378 N_A2_N_M1012_g N_VPWR_c_674_n 0.00157702f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A2_N_M1015_g N_VPWR_c_674_n 0.00157837f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A2_N_M1012_g N_VPWR_c_681_n 0.00441875f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A2_N_M1015_g N_VPWR_c_683_n 0.00441875f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_382 N_A2_N_M1012_g N_VPWR_c_670_n 0.00593338f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_383 N_A2_N_M1015_g N_VPWR_c_670_n 0.00588739f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_384 N_A2_N_c_468_n N_VGND_c_959_n 0.00368123f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_385 N_A2_N_c_469_n N_VGND_c_959_n 0.00368123f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A2_N_c_468_n N_VGND_c_964_n 0.00527354f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A2_N_c_469_n N_VGND_c_964_n 0.00527354f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_388 N_A2_N_c_468_n N_A_717_47#_c_1066_n 0.0083291f $X=3.93 $Y=0.995 $X2=0
+ $Y2=0
cc_389 N_A2_N_c_469_n N_A_717_47#_c_1066_n 0.00957565f $X=4.35 $Y=0.995 $X2=0
+ $Y2=0
cc_390 N_A2_N_c_470_n N_A_717_47#_c_1066_n 0.00305114f $X=4.145 $Y=1.16 $X2=0
+ $Y2=0
cc_391 N_A_193_297#_c_531_n N_VPWR_M1025_s 0.00663764f $X=2.065 $Y=1.87 $X2=0
+ $Y2=0
cc_392 N_A_193_297#_c_524_n N_VPWR_M1022_d 0.00582483f $X=5.165 $Y=1.53 $X2=0
+ $Y2=0
cc_393 N_A_193_297#_c_525_n N_VPWR_M1022_d 0.00162949f $X=2.675 $Y=1.53 $X2=0
+ $Y2=0
cc_394 N_A_193_297#_c_524_n N_VPWR_M1023_d 0.00154493f $X=5.165 $Y=1.53 $X2=0
+ $Y2=0
cc_395 N_A_193_297#_c_531_n N_VPWR_c_673_n 0.0123301f $X=2.065 $Y=1.87 $X2=0
+ $Y2=0
cc_396 N_A_193_297#_M1000_g N_VPWR_c_675_n 0.00157837f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_397 N_A_193_297#_c_524_n N_VPWR_c_675_n 0.00805046f $X=5.165 $Y=1.53 $X2=0
+ $Y2=0
cc_398 N_A_193_297#_M1000_g N_VPWR_c_676_n 0.00585385f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_399 N_A_193_297#_M1002_g N_VPWR_c_676_n 0.00585385f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_400 N_A_193_297#_M1002_g N_VPWR_c_677_n 0.00157837f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_401 N_A_193_297#_M1005_g N_VPWR_c_677_n 0.00157837f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_402 N_A_193_297#_M1026_g N_VPWR_c_678_n 0.00338128f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_403 N_A_193_297#_M1005_g N_VPWR_c_685_n 0.00585385f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_404 N_A_193_297#_M1026_g N_VPWR_c_685_n 0.00585385f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_405 N_A_193_297#_M1001_s N_VPWR_c_670_n 0.0021603f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_406 N_A_193_297#_M1004_s N_VPWR_c_670_n 0.00219397f $X=2.225 $Y=1.485 $X2=0
+ $Y2=0
cc_407 N_A_193_297#_M1000_g N_VPWR_c_670_n 0.010464f $X=5.19 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_A_193_297#_M1002_g N_VPWR_c_670_n 0.00588483f $X=5.61 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A_193_297#_M1005_g N_VPWR_c_670_n 0.00588483f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_410 N_A_193_297#_M1026_g N_VPWR_c_670_n 0.0117628f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_411 N_A_193_297#_c_531_n N_VPWR_c_670_n 0.00682229f $X=2.065 $Y=1.87 $X2=0
+ $Y2=0
cc_412 N_A_193_297#_c_519_n N_VPWR_c_670_n 0.0186938f $X=2.36 $Y=1.96 $X2=0
+ $Y2=0
cc_413 N_A_193_297#_c_519_n N_VPWR_c_688_n 0.0177981f $X=2.36 $Y=1.96 $X2=0
+ $Y2=0
cc_414 N_A_193_297#_c_524_n N_VPWR_c_689_n 0.0108145f $X=5.165 $Y=1.53 $X2=0
+ $Y2=0
cc_415 N_A_193_297#_c_531_n N_A_109_297#_M1003_d 0.00325521f $X=2.065 $Y=1.87
+ $X2=0 $Y2=0
cc_416 N_A_193_297#_M1001_s N_A_109_297#_c_793_n 0.00312348f $X=0.965 $Y=1.485
+ $X2=0 $Y2=0
cc_417 N_A_193_297#_c_531_n N_A_109_297#_c_793_n 0.00506389f $X=2.065 $Y=1.87
+ $X2=0 $Y2=0
cc_418 N_A_193_297#_c_536_n N_A_109_297#_c_793_n 0.0112811f $X=1.1 $Y=1.87 $X2=0
+ $Y2=0
cc_419 N_A_193_297#_c_531_n N_A_109_297#_c_799_n 0.0116461f $X=2.065 $Y=1.87
+ $X2=0 $Y2=0
cc_420 N_A_193_297#_c_526_n N_X_M1000_d 0.00466631f $X=5.31 $Y=1.53 $X2=0 $Y2=0
cc_421 N_A_193_297#_c_527_n N_X_M1000_d 0.00237412f $X=5.31 $Y=1.53 $X2=0 $Y2=0
cc_422 N_A_193_297#_c_513_n N_X_c_817_n 0.00494802f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_423 N_A_193_297#_c_514_n N_X_c_817_n 0.00612654f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_424 N_A_193_297#_c_515_n N_X_c_817_n 5.16334e-19 $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_425 N_A_193_297#_M1002_g N_X_c_820_n 0.0113688f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_426 N_A_193_297#_M1005_g N_X_c_820_n 0.0113688f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_427 N_A_193_297#_c_619_p N_X_c_820_n 0.0140663f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_428 N_A_193_297#_c_518_n N_X_c_820_n 0.00166652f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_429 N_A_193_297#_c_619_p N_X_c_824_n 0.00134408f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_430 N_A_193_297#_c_526_n N_X_c_824_n 0.0053154f $X=5.31 $Y=1.53 $X2=0 $Y2=0
cc_431 N_A_193_297#_c_527_n N_X_c_824_n 0.0103526f $X=5.31 $Y=1.53 $X2=0 $Y2=0
cc_432 N_A_193_297#_c_518_n N_X_c_824_n 3.77487e-19 $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_433 N_A_193_297#_c_514_n N_X_c_808_n 0.00870364f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A_193_297#_c_515_n N_X_c_808_n 0.00870364f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_435 N_A_193_297#_c_619_p N_X_c_808_n 0.0356734f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_436 N_A_193_297#_c_518_n N_X_c_808_n 0.00222133f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_193_297#_c_513_n N_X_c_809_n 0.00261784f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_438 N_A_193_297#_c_514_n N_X_c_809_n 0.00113229f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_439 N_A_193_297#_c_572_n N_X_c_809_n 0.0183805f $X=5.455 $Y=1.16 $X2=0 $Y2=0
cc_440 N_A_193_297#_c_619_p N_X_c_809_n 0.00865078f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_441 N_A_193_297#_c_526_n N_X_c_809_n 9.14672e-19 $X=5.31 $Y=1.53 $X2=0 $Y2=0
cc_442 N_A_193_297#_c_518_n N_X_c_809_n 0.00229945f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A_193_297#_c_514_n N_X_c_838_n 5.16334e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_444 N_A_193_297#_c_515_n N_X_c_838_n 0.00612654f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_445 N_A_193_297#_c_516_n N_X_c_838_n 0.0107369f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_446 N_A_193_297#_c_516_n N_X_c_810_n 0.0113812f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_447 N_A_193_297#_c_619_p N_X_c_810_n 0.00200821f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_448 N_A_193_297#_c_515_n N_X_c_811_n 0.00113229f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_449 N_A_193_297#_c_516_n N_X_c_811_n 0.00113229f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_450 N_A_193_297#_c_619_p N_X_c_811_n 0.0261859f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_451 N_A_193_297#_c_518_n N_X_c_811_n 0.00230115f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_452 N_A_193_297#_c_516_n X 0.0200556f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_453 N_A_193_297#_c_619_p X 0.014013f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_454 N_A_193_297#_M1005_g X 0.0012299f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_455 N_A_193_297#_M1026_g X 0.019019f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_456 N_A_193_297#_c_619_p X 0.0251128f $X=6.21 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_193_297#_c_527_n X 0.0025429f $X=5.31 $Y=1.53 $X2=0 $Y2=0
cc_458 N_A_193_297#_c_518_n X 0.00231083f $X=6.45 $Y=1.16 $X2=0 $Y2=0
cc_459 N_A_193_297#_c_548_n N_A_27_47#_c_885_n 0.00711741f $X=2.36 $Y=0.73 $X2=0
+ $Y2=0
cc_460 N_A_193_297#_M1020_s N_A_27_47#_c_886_n 0.00304656f $X=2.225 $Y=0.235
+ $X2=0 $Y2=0
cc_461 N_A_193_297#_c_548_n N_A_27_47#_c_886_n 0.0162134f $X=2.36 $Y=0.73 $X2=0
+ $Y2=0
cc_462 N_A_193_297#_c_519_n N_A_27_47#_c_886_n 0.00345006f $X=2.36 $Y=1.96 $X2=0
+ $Y2=0
cc_463 N_A_193_297#_c_513_n N_VGND_c_949_n 0.0015308f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_464 N_A_193_297#_c_524_n N_VGND_c_949_n 0.00388941f $X=5.165 $Y=1.53 $X2=0
+ $Y2=0
cc_465 N_A_193_297#_c_513_n N_VGND_c_950_n 0.00542163f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_466 N_A_193_297#_c_514_n N_VGND_c_950_n 0.00424138f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_467 N_A_193_297#_c_514_n N_VGND_c_951_n 0.00146448f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_468 N_A_193_297#_c_515_n N_VGND_c_951_n 0.00146448f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_469 N_A_193_297#_c_516_n N_VGND_c_952_n 0.00316354f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_470 N_A_193_297#_c_515_n N_VGND_c_961_n 0.00424138f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_471 N_A_193_297#_c_516_n N_VGND_c_961_n 0.00424138f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_193_297#_M1020_s N_VGND_c_964_n 0.00216833f $X=2.225 $Y=0.235 $X2=0
+ $Y2=0
cc_473 N_A_193_297#_c_513_n N_VGND_c_964_n 0.00952972f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_193_297#_c_514_n N_VGND_c_964_n 0.00571728f $X=5.61 $Y=0.995 $X2=0
+ $Y2=0
cc_475 N_A_193_297#_c_515_n N_VGND_c_964_n 0.00571728f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_A_193_297#_c_516_n N_VGND_c_964_n 0.00704335f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_477 N_A_193_297#_c_524_n N_A_717_47#_c_1064_n 0.00145512f $X=5.165 $Y=1.53
+ $X2=0 $Y2=0
cc_478 N_VPWR_c_670_n N_A_109_297#_M1019_d 0.00246446f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_479 N_VPWR_c_670_n N_A_109_297#_M1003_d 0.00219968f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_679_n N_A_109_297#_c_793_n 0.0330174f $X=1.815 $Y=2.72 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_670_n N_A_109_297#_c_793_n 0.0204667f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_679_n N_A_109_297#_c_804_n 0.0143053f $X=1.815 $Y=2.72 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_670_n N_A_109_297#_c_804_n 0.00962794f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_679_n N_A_109_297#_c_799_n 0.0137033f $X=1.815 $Y=2.72 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_670_n N_A_109_297#_c_799_n 0.00938745f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_670_n N_X_M1000_d 0.00254126f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_487 N_VPWR_c_670_n N_X_M1005_d 0.00254126f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_488 N_VPWR_c_676_n N_X_c_856_n 0.0142343f $X=5.695 $Y=2.72 $X2=0 $Y2=0
cc_489 N_VPWR_c_670_n N_X_c_856_n 0.00955092f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_490 N_VPWR_M1002_s N_X_c_820_n 0.00441488f $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_491 N_VPWR_c_677_n N_X_c_820_n 0.0102703f $X=5.82 $Y=2.33 $X2=0 $Y2=0
cc_492 N_VPWR_c_670_n N_X_c_820_n 0.0110135f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_493 N_VPWR_c_685_n N_X_c_861_n 0.0142343f $X=6.535 $Y=2.72 $X2=0 $Y2=0
cc_494 N_VPWR_c_670_n N_X_c_861_n 0.00955092f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_495 N_VPWR_M1026_s X 0.00298019f $X=6.525 $Y=1.485 $X2=0 $Y2=0
cc_496 N_VPWR_c_678_n X 0.0180643f $X=6.66 $Y=1.99 $X2=0 $Y2=0
cc_497 N_X_c_808_n N_VGND_M1010_s 0.00162089f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_498 N_X_c_810_n N_VGND_M1017_s 0.00324398f $X=6.605 $Y=0.815 $X2=0 $Y2=0
cc_499 N_X_c_809_n N_VGND_c_949_n 0.00750114f $X=5.565 $Y=0.815 $X2=0 $Y2=0
cc_500 N_X_c_817_n N_VGND_c_950_n 0.0167046f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_501 N_X_c_808_n N_VGND_c_950_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_502 N_X_c_808_n N_VGND_c_951_n 0.0122559f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_503 N_X_c_810_n N_VGND_c_952_n 0.0137936f $X=6.605 $Y=0.815 $X2=0 $Y2=0
cc_504 N_X_c_808_n N_VGND_c_961_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_505 N_X_c_838_n N_VGND_c_961_n 0.0167046f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_506 N_X_c_810_n N_VGND_c_961_n 0.00198695f $X=6.605 $Y=0.815 $X2=0 $Y2=0
cc_507 N_X_c_810_n N_VGND_c_963_n 0.00276263f $X=6.605 $Y=0.815 $X2=0 $Y2=0
cc_508 N_X_M1006_d N_VGND_c_964_n 0.00216035f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_509 N_X_M1011_d N_VGND_c_964_n 0.00216035f $X=6.105 $Y=0.235 $X2=0 $Y2=0
cc_510 N_X_c_817_n N_VGND_c_964_n 0.0120721f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_511 N_X_c_808_n N_VGND_c_964_n 0.00835832f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_512 N_X_c_838_n N_VGND_c_964_n 0.0120721f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_513 N_X_c_810_n N_VGND_c_964_n 0.00925667f $X=6.605 $Y=0.815 $X2=0 $Y2=0
cc_514 N_A_27_47#_c_883_n N_VGND_M1016_s 0.00162089f $X=0.935 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_515 N_A_27_47#_c_885_n N_VGND_M1018_s 0.00165819f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_c_883_n N_VGND_c_946_n 0.0122559f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_885_n N_VGND_c_947_n 0.0116528f $X=1.775 $Y=0.82 $X2=0 $Y2=0
cc_518 N_A_27_47#_c_886_n N_VGND_c_948_n 0.0130084f $X=2.78 $Y=0.39 $X2=0 $Y2=0
cc_519 N_A_27_47#_c_882_n N_VGND_c_953_n 0.0209752f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_520 N_A_27_47#_c_883_n N_VGND_c_953_n 0.00198695f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_c_883_n N_VGND_c_955_n 0.00198695f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_895_n N_VGND_c_955_n 0.0188551f $X=1.1 $Y=0.39 $X2=0 $Y2=0
cc_523 N_A_27_47#_c_885_n N_VGND_c_955_n 0.00193763f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_524 N_A_27_47#_c_885_n N_VGND_c_957_n 0.00193763f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_525 N_A_27_47#_c_901_n N_VGND_c_957_n 0.0152108f $X=1.9 $Y=0.475 $X2=0 $Y2=0
cc_526 N_A_27_47#_c_886_n N_VGND_c_957_n 0.0522924f $X=2.78 $Y=0.39 $X2=0 $Y2=0
cc_527 N_A_27_47#_M1016_d N_VGND_c_964_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_528 N_A_27_47#_M1013_d N_VGND_c_964_n 0.00215201f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_529 N_A_27_47#_M1027_d N_VGND_c_964_n 0.00215206f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_530 N_A_27_47#_M1024_d N_VGND_c_964_n 0.00209344f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_531 N_A_27_47#_c_882_n N_VGND_c_964_n 0.0124119f $X=0.26 $Y=0.39 $X2=0 $Y2=0
cc_532 N_A_27_47#_c_883_n N_VGND_c_964_n 0.00835832f $X=0.935 $Y=0.815 $X2=0
+ $Y2=0
cc_533 N_A_27_47#_c_895_n N_VGND_c_964_n 0.0122069f $X=1.1 $Y=0.39 $X2=0 $Y2=0
cc_534 N_A_27_47#_c_885_n N_VGND_c_964_n 0.00827287f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_535 N_A_27_47#_c_901_n N_VGND_c_964_n 0.00940698f $X=1.9 $Y=0.475 $X2=0 $Y2=0
cc_536 N_A_27_47#_c_886_n N_VGND_c_964_n 0.0329455f $X=2.78 $Y=0.39 $X2=0 $Y2=0
cc_537 N_VGND_c_964_n N_A_717_47#_M1008_d 0.00218617f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_538 N_VGND_c_964_n N_A_717_47#_M1014_s 0.00218529f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_c_959_n N_A_717_47#_c_1066_n 0.0378883f $X=4.895 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_c_964_n N_A_717_47#_c_1066_n 0.031469f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_959_n N_A_717_47#_c_1071_n 0.0114667f $X=4.895 $Y=0 $X2=0 $Y2=0
cc_542 N_VGND_c_964_n N_A_717_47#_c_1071_n 0.00913547f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_949_n N_A_717_47#_c_1064_n 0.0154056f $X=4.98 $Y=0.39 $X2=0
+ $Y2=0

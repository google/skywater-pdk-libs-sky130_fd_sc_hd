* File: sky130_fd_sc_hd__dfbbn_2.spice.pex
* Created: Thu Aug 27 14:14:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFBBN_2%CLK_N 4 5 7 8 10 13 17 19 20 24 26
c45 13 0 2.71124e-20 $X=0.47 $Y=0.805
r46 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r47 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r48 19 20 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.262 $Y=1.19
+ $X2=0.262 $Y2=1.53
r49 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r50 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r51 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r52 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r53 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r54 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r55 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r56 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r57 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r58 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r59 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_27_47# 1 2 9 13 17 19 20 23 26 27 29 32 36
+ 40 41 42 46 47 49 51 52 55 58 59 61 62 63 66 70 71 74 81 84
c261 61 0 9.18873e-20 $X=3.032 $Y=1.12
c262 49 0 1.20913e-19 $X=6.652 $Y=1.305
c263 47 0 1.7288e-19 $X=6.335 $Y=0.87
c264 17 0 4.43992e-20 $X=2.305 $Y=2.275
r265 84 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=0.93
+ $X2=2.905 $Y2=1.095
r266 84 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=0.93
+ $X2=2.905 $Y2=0.765
r267 78 81 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r268 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r269 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.225 $Y=1.19
+ $X2=6.225 $Y2=1.19
r270 71 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=0.93 $X2=2.905 $Y2=0.93
r271 70 72 0.0716299 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=2.985 $Y=0.85
+ $X2=2.985 $Y2=0.965
r272 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.985 $Y=0.85
+ $X2=2.985 $Y2=0.85
r273 66 79 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.725 $Y=0.85
+ $X2=0.725 $Y2=1.235
r274 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=0.85
+ $X2=0.695 $Y2=0.85
r275 62 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=1.19
+ $X2=6.225 $Y2=1.19
r276 62 63 3.65098 $w=1.4e-07 $l=2.95e-06 $layer=MET1_cond $X=6.08 $Y=1.19
+ $X2=3.13 $Y2=1.19
r277 61 63 0.0723178 $w=1.4e-07 $l=1.28312e-07 $layer=MET1_cond $X=3.032 $Y=1.12
+ $X2=3.13 $Y2=1.19
r278 61 72 0.12202 $w=1.95e-07 $l=1.55e-07 $layer=MET1_cond $X=3.032 $Y=1.12
+ $X2=3.032 $Y2=0.965
r279 59 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=0.85
+ $X2=0.695 $Y2=0.85
r280 58 70 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.84 $Y=0.85
+ $X2=2.985 $Y2=0.85
r281 58 59 2.47524 $w=1.4e-07 $l=2e-06 $layer=MET1_cond $X=2.84 $Y=0.85 $X2=0.84
+ $Y2=0.85
r282 57 79 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r283 56 66 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=0.85
r284 52 94 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.67 $Y=1.74
+ $X2=6.67 $Y2=1.875
r285 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.67
+ $Y=1.74 $X2=6.67 $Y2=1.74
r286 49 75 26.3101 $w=1.78e-07 $l=4.27e-07 $layer=LI1_cond $X=6.652 $Y=1.215
+ $X2=6.225 $Y2=1.215
r287 49 51 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=6.652 $Y=1.305
+ $X2=6.652 $Y2=1.74
r288 47 88 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.335 $Y=0.87
+ $X2=6.21 $Y2=0.87
r289 46 75 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=6.277 $Y=0.87
+ $X2=6.277 $Y2=1.125
r290 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.335
+ $Y=0.87 $X2=6.335 $Y2=0.87
r291 43 55 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r292 42 57 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.795
r293 42 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r294 40 56 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r295 40 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r296 34 41 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r297 34 36 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r298 32 94 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.64 $Y=2.275
+ $X2=6.64 $Y2=1.875
r299 27 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=0.705
+ $X2=6.21 $Y2=0.87
r300 27 29 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.21 $Y=0.705
+ $X2=6.21 $Y2=0.415
r301 26 87 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.845 $Y=1.245
+ $X2=2.845 $Y2=1.095
r302 23 86 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.845 $Y=0.415
+ $X2=2.845 $Y2=0.765
r303 19 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.77 $Y=1.32
+ $X2=2.845 $Y2=1.245
r304 19 20 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.77 $Y=1.32
+ $X2=2.38 $Y2=1.32
r305 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.305 $Y=1.395
+ $X2=2.38 $Y2=1.32
r306 15 17 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.305 $Y=1.395
+ $X2=2.305 $Y2=2.275
r307 11 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r308 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r309 7 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r310 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r311 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r312 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%D 3 7 9 10 14 15
c41 7 0 1.779e-19 $X=1.83 $Y=2.275
r42 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.17
+ $X2=1.845 $Y2=1.335
r43 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.17
+ $X2=1.845 $Y2=1.005
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.17 $X2=1.845 $Y2=1.17
r45 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.965 $Y=1.19
+ $X2=1.965 $Y2=1.53
r46 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.965 $Y=1.19
+ $X2=1.965 $Y2=1.17
r47 7 17 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.83 $Y=2.275 $X2=1.83
+ $Y2=1.335
r48 3 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.83 $Y=0.445
+ $X2=1.83 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_193_47# 1 2 7 9 12 18 20 21 24 28 29 31 32
+ 33 34 43 51 52 56 57 58 61
c202 56 0 2.05666e-19 $X=6.16 $Y=1.74
c203 33 0 1.55301e-20 $X=6.08 $Y=1.87
c204 29 0 9.18873e-20 $X=2.425 $Y=0.87
c205 28 0 1.779e-19 $X=2.425 $Y=0.87
c206 18 0 3.84972e-20 $X=6.22 $Y=2.275
r207 56 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.74
+ $X2=6.16 $Y2=1.905
r208 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.74
+ $X2=6.16 $Y2=1.575
r209 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.16
+ $Y=1.74 $X2=6.16 $Y2=1.74
r210 51 54 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.755 $Y=1.74
+ $X2=2.755 $Y2=1.875
r211 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.755
+ $Y=1.74 $X2=2.755 $Y2=1.74
r212 43 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.225 $Y=1.87
+ $X2=6.225 $Y2=1.87
r213 41 52 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=2.545 $Y=1.765
+ $X2=2.755 $Y2=1.765
r214 41 69 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.545 $Y=1.765
+ $X2=2.45 $Y2=1.765
r215 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.545 $Y=1.87
+ $X2=2.545 $Y2=1.87
r216 37 61 69.6588 $w=2.23e-07 $l=1.36e-06 $layer=LI1_cond $X=1.127 $Y=1.87
+ $X2=1.127 $Y2=0.51
r217 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r218 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.69 $Y=1.87
+ $X2=2.545 $Y2=1.87
r219 33 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.08 $Y=1.87
+ $X2=6.225 $Y2=1.87
r220 33 34 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=6.08 $Y=1.87
+ $X2=2.69 $Y2=1.87
r221 32 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r222 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.4 $Y=1.87
+ $X2=2.545 $Y2=1.87
r223 31 32 1.36138 $w=1.4e-07 $l=1.1e-06 $layer=MET1_cond $X=2.4 $Y=1.87 $X2=1.3
+ $Y2=1.87
r224 29 46 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.425 $Y=0.87
+ $X2=2.305 $Y2=0.87
r225 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.425
+ $Y=0.87 $X2=2.425 $Y2=0.87
r226 26 69 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.45 $Y=1.575
+ $X2=2.45 $Y2=1.765
r227 26 28 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.45 $Y=1.575
+ $X2=2.45 $Y2=0.87
r228 22 24 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=6.755 $Y=1.245
+ $X2=6.755 $Y2=0.415
r229 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.68 $Y=1.32
+ $X2=6.755 $Y2=1.245
r230 20 21 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.68 $Y=1.32
+ $X2=6.295 $Y2=1.32
r231 18 59 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.22 $Y=2.275
+ $X2=6.22 $Y2=1.905
r232 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.22 $Y=1.395
+ $X2=6.295 $Y2=1.32
r233 14 58 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.22 $Y=1.395
+ $X2=6.22 $Y2=1.575
r234 12 54 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.725 $Y=2.275
+ $X2=2.725 $Y2=1.875
r235 7 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r236 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r237 2 37 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r238 1 61 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_650_21# 1 2 9 13 17 19 21 22 26 28 30 31
+ 32 35 36 41 45 49
c145 9 0 7.56837e-20 $X=3.325 $Y=0.445
r146 49 56 10.4783 $w=2.76e-07 $l=6e-08 $layer=POLY_cond $X=5.675 $Y=1.15
+ $X2=5.735 $Y2=1.15
r147 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.675
+ $Y=1.15 $X2=5.675 $Y2=1.15
r148 45 48 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.675 $Y=0.98
+ $X2=5.675 $Y2=1.15
r149 43 44 14.1313 $w=2.59e-07 $l=3e-07 $layer=LI1_cond $X=4.585 $Y=0.68
+ $X2=4.585 $Y2=0.98
r150 36 53 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.74
+ $X2=3.41 $Y2=1.905
r151 36 52 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.74
+ $X2=3.41 $Y2=1.575
r152 35 38 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.475 $Y=1.74
+ $X2=3.475 $Y2=1.91
r153 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.435
+ $Y=1.74 $X2=3.435 $Y2=1.74
r154 33 44 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=0.98
+ $X2=4.585 $Y2=0.98
r155 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=0.98
+ $X2=5.675 $Y2=0.98
r156 32 33 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.51 $Y=0.98
+ $X2=4.75 $Y2=0.98
r157 30 44 5.44435 $w=2.59e-07 $l=9.88686e-08 $layer=LI1_cond $X=4.615 $Y=1.065
+ $X2=4.585 $Y2=0.98
r158 30 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.615 $Y=1.065
+ $X2=4.615 $Y2=1.785
r159 29 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=1.91
+ $X2=4.185 $Y2=1.91
r160 28 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.53 $Y=1.91
+ $X2=4.615 $Y2=1.785
r161 28 29 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=4.53 $Y=1.91
+ $X2=4.27 $Y2=1.91
r162 24 41 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=2.035
+ $X2=4.185 $Y2=1.91
r163 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.185 $Y=2.035
+ $X2=4.185 $Y2=2.21
r164 23 38 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=1.91
+ $X2=3.475 $Y2=1.91
r165 22 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=1.91
+ $X2=4.185 $Y2=1.91
r166 22 23 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=4.1 $Y=1.91 $X2=3.6
+ $Y2=1.91
r167 19 56 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=0.985
+ $X2=5.735 $Y2=1.15
r168 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.735 $Y=0.985
+ $X2=5.735 $Y2=0.555
r169 15 49 30.5616 $w=2.76e-07 $l=2.43926e-07 $layer=POLY_cond $X=5.5 $Y=1.315
+ $X2=5.675 $Y2=1.15
r170 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.5 $Y=1.315
+ $X2=5.5 $Y2=2.065
r171 13 53 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.325 $Y=2.275
+ $X2=3.325 $Y2=1.905
r172 9 52 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.325 $Y=0.445
+ $X2=3.325 $Y2=1.575
r173 2 41 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=2.065 $X2=4.185 $Y2=1.87
r174 2 26 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=2.065 $X2=4.185 $Y2=2.21
r175 1 43 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.235 $X2=4.585 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%SET_B 1 3 7 11 15 17 19 20 26 27 33
c131 33 0 1.0279e-19 $X=7.65 $Y=0.98
c132 19 0 1.0411e-19 $X=7.46 $Y=0.85
c133 15 0 1.0852e-19 $X=7.77 $Y=2.275
r134 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.68 $Y=0.98
+ $X2=7.68 $Y2=1.145
r135 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.68 $Y=0.98
+ $X2=7.68 $Y2=0.815
r136 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.65
+ $Y=0.98 $X2=7.65 $Y2=0.98
r137 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.605 $Y=0.85
+ $X2=7.605 $Y2=0.85
r138 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.07 $Y=0.85
+ $X2=3.925 $Y2=0.85
r139 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.46 $Y=0.85
+ $X2=7.605 $Y2=0.85
r140 19 20 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=7.46 $Y=0.85
+ $X2=4.07 $Y2=0.85
r141 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.765
+ $Y=0.98 $X2=3.765 $Y2=0.98
r142 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.925 $Y=0.85
+ $X2=3.925 $Y2=0.85
r143 15 36 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.77 $Y=2.275
+ $X2=7.77 $Y2=1.145
r144 11 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.66 $Y=0.445
+ $X2=7.66 $Y2=0.815
r145 5 30 38.532 $w=3.09e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.875 $Y=0.815
+ $X2=3.79 $Y2=0.98
r146 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.875 $Y=0.815
+ $X2=3.875 $Y2=0.445
r147 1 30 38.532 $w=3.09e-07 $l=1.94808e-07 $layer=POLY_cond $X=3.855 $Y=1.145
+ $X2=3.79 $Y2=0.98
r148 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.855 $Y=1.145
+ $X2=3.855 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_476_47# 1 2 9 13 15 19 24 26 27 32 35
c105 35 0 1.0411e-19 $X=4.275 $Y=1.32
c106 32 0 4.43992e-20 $X=3.41 $Y=1.3
r107 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.32
+ $X2=4.305 $Y2=1.485
r108 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.32
+ $X2=4.305 $Y2=1.155
r109 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.275
+ $Y=1.32 $X2=4.275 $Y2=1.32
r110 31 32 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=1.3
+ $X2=3.41 $Y2=1.3
r111 29 31 12.1472 $w=2.08e-07 $l=2.3e-07 $layer=LI1_cond $X=3.095 $Y=1.3
+ $X2=3.325 $Y2=1.3
r112 27 34 8.9562 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.11 $Y=1.32
+ $X2=4.275 $Y2=1.32
r113 27 32 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.11 $Y=1.32 $X2=3.41
+ $Y2=1.32
r114 26 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.325 $Y=1.195
+ $X2=3.325 $Y2=1.3
r115 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.325 $Y=0.465
+ $X2=3.325 $Y2=1.195
r116 23 29 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=1.405
+ $X2=3.095 $Y2=1.3
r117 23 24 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.095 $Y=1.405
+ $X2=3.095 $Y2=2.25
r118 19 25 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.24 $Y=0.365
+ $X2=3.325 $Y2=0.465
r119 19 21 36.6 $w=1.98e-07 $l=6.6e-07 $layer=LI1_cond $X=3.24 $Y=0.365 $X2=2.58
+ $Y2=0.365
r120 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.01 $Y=2.335
+ $X2=3.095 $Y2=2.25
r121 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.01 $Y=2.335
+ $X2=2.515 $Y2=2.335
r122 13 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.395 $Y=2.065
+ $X2=4.395 $Y2=1.485
r123 9 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.375 $Y=0.555
+ $X2=4.375 $Y2=1.155
r124 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=2.065 $X2=2.515 $Y2=2.335
r125 1 21 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.58 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_944_21# 1 2 9 13 17 21 23 24 25 27 31 34
+ 35 42 43 46 49 57 60
c158 57 0 1.89563e-19 $X=8.67 $Y=1.32
c159 42 0 2.58372e-20 $X=8.84 $Y=1.53
c160 35 0 1.55301e-20 $X=5.035 $Y=1.32
c161 27 0 1.48493e-19 $X=9.405 $Y=1.66
r162 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.88
+ $Y=1.32 $X2=8.88 $Y2=1.32
r163 57 59 32.9707 $w=3.07e-07 $l=2.1e-07 $layer=POLY_cond $X=8.67 $Y=1.32
+ $X2=8.88 $Y2=1.32
r164 56 57 9.4202 $w=3.07e-07 $l=6e-08 $layer=POLY_cond $X=8.61 $Y=1.32 $X2=8.67
+ $Y2=1.32
r165 50 60 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=8.932 $Y=1.53
+ $X2=8.932 $Y2=1.32
r166 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.985 $Y=1.53
+ $X2=8.985 $Y2=1.53
r167 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.765 $Y=1.53
+ $X2=5.765 $Y2=1.53
r168 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.91 $Y=1.53
+ $X2=5.765 $Y2=1.53
r169 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.84 $Y=1.53
+ $X2=8.985 $Y2=1.53
r170 42 43 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=8.84 $Y=1.53
+ $X2=5.91 $Y2=1.53
r171 41 50 1.88582 $w=2.73e-07 $l=4.5e-08 $layer=LI1_cond $X=8.932 $Y=1.575
+ $X2=8.932 $Y2=1.53
r172 40 60 16.5533 $w=2.73e-07 $l=3.95e-07 $layer=LI1_cond $X=8.932 $Y=0.925
+ $X2=8.932 $Y2=1.32
r173 38 46 27.1304 $w=2.38e-07 $l=5.65e-07 $layer=LI1_cond $X=5.2 $Y=1.535
+ $X2=5.765 $Y2=1.535
r174 37 38 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=1.535
+ $X2=5.2 $Y2=1.535
r175 35 52 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=5.035 $Y=1.32
+ $X2=4.795 $Y2=1.32
r176 34 37 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.035 $Y=1.32
+ $X2=5.035 $Y2=1.535
r177 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.035
+ $Y=1.32 $X2=5.035 $Y2=1.32
r178 29 31 17.0247 $w=2.18e-07 $l=3.25e-07 $layer=LI1_cond $X=9.39 $Y=0.755
+ $X2=9.39 $Y2=0.43
r179 25 41 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=9.07 $Y=1.66
+ $X2=8.932 $Y2=1.575
r180 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.07 $Y=1.66
+ $X2=9.405 $Y2=1.66
r181 24 40 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=9.07 $Y=0.84
+ $X2=8.932 $Y2=0.925
r182 23 29 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=9.28 $Y=0.84
+ $X2=9.39 $Y2=0.755
r183 23 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.28 $Y=0.84
+ $X2=9.07 $Y2=0.84
r184 19 57 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=1.155
+ $X2=8.67 $Y2=1.32
r185 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.67 $Y=1.155 $X2=8.67
+ $Y2=0.555
r186 15 56 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.485
+ $X2=8.61 $Y2=1.32
r187 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.61 $Y=1.485
+ $X2=8.61 $Y2=2.065
r188 11 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.795 $Y=1.485
+ $X2=4.795 $Y2=1.32
r189 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.795 $Y=1.485
+ $X2=4.795 $Y2=2.065
r190 7 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.795 $Y=1.155
+ $X2=4.795 $Y2=1.32
r191 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.795 $Y=1.155 $X2=4.795
+ $Y2=0.555
r192 2 27 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=9.28
+ $Y=1.505 $X2=9.405 $Y2=1.66
r193 1 31 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=9.29
+ $Y=0.235 $X2=9.415 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_1431_21# 1 2 9 13 15 17 20 24 28 30 31 33
+ 35 36 38 39 41 44 46 49 53 54 56 57 60 62 65 66 69 70 74 76 78
c196 78 0 1.15981e-19 $X=10.055 $Y=1.16
c197 74 0 1.22108e-19 $X=8.535 $Y=0.687
c198 20 0 1.48493e-19 $X=10.115 $Y=1.985
c199 9 0 8.81272e-20 $X=7.23 $Y=0.445
r200 79 86 9.87031 $w=2.93e-07 $l=6e-08 $layer=POLY_cond $X=10.055 $Y=1.16
+ $X2=10.115 $Y2=1.16
r201 78 81 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=10.02 $Y=1.16
+ $X2=10.02 $Y2=1.325
r202 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.055
+ $Y=1.16 $X2=10.055 $Y2=1.16
r203 72 74 4.49631 $w=1.83e-07 $l=7.5e-08 $layer=LI1_cond $X=8.46 $Y=0.687
+ $X2=8.535 $Y2=0.687
r204 69 81 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.985 $Y=1.915
+ $X2=9.985 $Y2=1.325
r205 67 76 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.625 $Y=2 $X2=8.535
+ $Y2=2
r206 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.9 $Y=2
+ $X2=9.985 $Y2=1.915
r207 66 67 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=9.9 $Y=2
+ $X2=8.625 $Y2=2
r208 65 76 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.535 $Y=1.915
+ $X2=8.535 $Y2=2
r209 64 74 0.88302 $w=1.8e-07 $l=9.3e-08 $layer=LI1_cond $X=8.535 $Y=0.78
+ $X2=8.535 $Y2=0.687
r210 64 65 69.9343 $w=1.78e-07 $l=1.135e-06 $layer=LI1_cond $X=8.535 $Y=0.78
+ $X2=8.535 $Y2=1.915
r211 63 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.125 $Y=2 $X2=8.04
+ $Y2=2
r212 62 76 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=8.445 $Y=2 $X2=8.535
+ $Y2=2
r213 62 63 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.445 $Y=2 $X2=8.125
+ $Y2=2
r214 58 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=2.085
+ $X2=8.04 $Y2=2
r215 58 60 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.04 $Y=2.085
+ $X2=8.04 $Y2=2.21
r216 56 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=2 $X2=8.04
+ $Y2=2
r217 56 57 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.955 $Y=2
+ $X2=7.515 $Y2=2
r218 54 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.32 $Y=1.74
+ $X2=7.32 $Y2=1.905
r219 54 83 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.32 $Y=1.74
+ $X2=7.32 $Y2=1.575
r220 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.35
+ $Y=1.74 $X2=7.35 $Y2=1.74
r221 51 57 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.39 $Y=1.915
+ $X2=7.515 $Y2=2
r222 51 53 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=7.39 $Y=1.915
+ $X2=7.39 $Y2=1.74
r223 47 49 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=11.385 $Y=1.61
+ $X2=11.515 $Y2=1.61
r224 42 44 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=11.385 $Y=0.805
+ $X2=11.515 $Y2=0.805
r225 39 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.515 $Y=1.685
+ $X2=11.515 $Y2=1.61
r226 39 41 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=11.515 $Y=1.685
+ $X2=11.515 $Y2=2.085
r227 36 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.515 $Y=0.73
+ $X2=11.515 $Y2=0.805
r228 36 38 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.515 $Y=0.73
+ $X2=11.515 $Y2=0.445
r229 35 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.385 $Y=1.535
+ $X2=11.385 $Y2=1.61
r230 34 46 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.385 $Y=1.295
+ $X2=11.385 $Y2=1.16
r231 34 35 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.385 $Y=1.295
+ $X2=11.385 $Y2=1.535
r232 33 46 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.385 $Y=1.025
+ $X2=11.385 $Y2=1.16
r233 32 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.385 $Y=0.88
+ $X2=11.385 $Y2=0.805
r234 32 33 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=11.385 $Y=0.88
+ $X2=11.385 $Y2=1.025
r235 30 46 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=11.31 $Y=1.16
+ $X2=11.385 $Y2=1.16
r236 30 31 155.522 $w=2.7e-07 $l=7e-07 $layer=POLY_cond $X=11.31 $Y=1.16
+ $X2=10.61 $Y2=1.16
r237 22 31 12.7172 $w=2.93e-07 $l=7.5e-08 $layer=POLY_cond $X=10.535 $Y=1.16
+ $X2=10.61 $Y2=1.16
r238 22 86 69.0921 $w=2.93e-07 $l=4.2e-07 $layer=POLY_cond $X=10.535 $Y=1.16
+ $X2=10.115 $Y2=1.16
r239 22 28 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.535 $Y=1.295
+ $X2=10.535 $Y2=1.985
r240 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.535 $Y=1.025
+ $X2=10.535 $Y2=0.56
r241 18 86 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.115 $Y=1.325
+ $X2=10.115 $Y2=1.16
r242 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.115 $Y=1.325
+ $X2=10.115 $Y2=1.985
r243 15 86 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.115 $Y=0.995
+ $X2=10.115 $Y2=1.16
r244 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.115 $Y=0.995
+ $X2=10.115 $Y2=0.56
r245 13 84 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.23 $Y=2.275
+ $X2=7.23 $Y2=1.905
r246 9 83 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.23 $Y=0.445
+ $X2=7.23 $Y2=1.575
r247 2 60 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=7.845
+ $Y=2.065 $X2=8.04 $Y2=2.21
r248 1 72 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.235 $X2=8.46 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_1257_47# 1 2 9 13 15 19 24 26 27 29 31 32
c99 32 0 2.58372e-20 $X=8.19 $Y=1.24
c100 31 0 1.75976e-19 $X=8.19 $Y=1.24
c101 26 0 3.84972e-20 $X=7.01 $Y=2.25
r102 32 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.19 $Y=1.24
+ $X2=8.19 $Y2=1.405
r103 32 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.19 $Y=1.24
+ $X2=8.19 $Y2=1.075
r104 31 34 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=8.165 $Y=1.24
+ $X2=8.165 $Y2=1.32
r105 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.19
+ $Y=1.24 $X2=8.19 $Y2=1.24
r106 28 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=1.32
+ $X2=7.01 $Y2=1.32
r107 27 34 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=8.055 $Y=1.32
+ $X2=8.165 $Y2=1.32
r108 27 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.055 $Y=1.32
+ $X2=7.095 $Y2=1.32
r109 25 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=1.405
+ $X2=7.01 $Y2=1.32
r110 25 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=7.01 $Y=1.405
+ $X2=7.01 $Y2=2.25
r111 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=1.235
+ $X2=7.01 $Y2=1.32
r112 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.01 $Y=0.465
+ $X2=7.01 $Y2=1.235
r113 19 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.925 $Y=0.365
+ $X2=7.01 $Y2=0.465
r114 19 21 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=6.925 $Y=0.365
+ $X2=6.495 $Y2=0.365
r115 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.925 $Y=2.335
+ $X2=7.01 $Y2=2.25
r116 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.925 $Y=2.335
+ $X2=6.43 $Y2=2.335
r117 13 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.25 $Y=2.065
+ $X2=8.25 $Y2=1.405
r118 9 37 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.25 $Y=0.555
+ $X2=8.25 $Y2=1.075
r119 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=2.065 $X2=6.43 $Y2=2.335
r120 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.495 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%RESET_B 3 7 9 15
r36 12 15 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=9.415 $Y=1.18
+ $X2=9.63 $Y2=1.18
r37 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.415
+ $Y=1.18 $X2=9.415 $Y2=1.18
r38 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=1.345
+ $X2=9.63 $Y2=1.18
r39 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.63 $Y=1.345 $X2=9.63
+ $Y2=1.825
r40 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=1.015
+ $X2=9.63 $Y2=1.18
r41 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=9.63 $Y=1.015 $X2=9.63
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_2236_47# 1 2 7 9 12 14 16 19 23 27 31 34
+ 38
c72 38 0 3.03687e-19 $X=12.41 $Y=1.16
r73 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=11.99 $Y=1.16
+ $X2=12.41 $Y2=1.16
r74 32 37 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=11.905 $Y=1.16
+ $X2=11.99 $Y2=1.16
r75 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.905
+ $Y=1.16 $X2=11.905 $Y2=1.16
r76 29 34 0.432806 $w=3.3e-07 $l=1.28e-07 $layer=LI1_cond $X=11.47 $Y=1.16
+ $X2=11.342 $Y2=1.16
r77 29 31 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=11.47 $Y=1.16
+ $X2=11.905 $Y2=1.16
r78 25 34 6.36606 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=11.342 $Y=1.325
+ $X2=11.342 $Y2=1.16
r79 25 27 26.4384 $w=2.53e-07 $l=5.85e-07 $layer=LI1_cond $X=11.342 $Y=1.325
+ $X2=11.342 $Y2=1.91
r80 21 34 6.36606 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=11.342 $Y=0.995
+ $X2=11.342 $Y2=1.16
r81 21 23 21.919 $w=2.53e-07 $l=4.85e-07 $layer=LI1_cond $X=11.342 $Y=0.995
+ $X2=11.342 $Y2=0.51
r82 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.41 $Y=1.325
+ $X2=12.41 $Y2=1.16
r83 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.41 $Y=1.325
+ $X2=12.41 $Y2=1.985
r84 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.41 $Y2=1.16
r85 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.41 $Y2=0.56
r86 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.99 $Y=1.325
+ $X2=11.99 $Y2=1.16
r87 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.99 $Y=1.325
+ $X2=11.99 $Y2=1.985
r88 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.99 $Y=0.995
+ $X2=11.99 $Y2=1.16
r89 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.99 $Y=0.995
+ $X2=11.99 $Y2=0.56
r90 2 27 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.18
+ $Y=1.765 $X2=11.305 $Y2=1.91
r91 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=11.18
+ $Y=0.235 $X2=11.305 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 59 61 66 67 68 72 73 75 77 83 88 100 111 115 120 126 129 132 135 146 148
+ 151 155 158
r201 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r202 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r203 149 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r204 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r205 145 146 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.905 $Y=2.53
+ $X2=10.07 $Y2=2.53
r206 142 145 0.326203 $w=5.48e-07 $l=1.5e-08 $layer=LI1_cond $X=9.89 $Y=2.53
+ $X2=9.905 $Y2=2.53
r207 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r208 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r209 135 138 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=7.525 $Y=2.34
+ $X2=7.525 $Y2=2.72
r210 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r211 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r212 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r213 124 155 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=12.65 $Y2=2.72
r214 124 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r215 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r216 121 151 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=11.945 $Y=2.72
+ $X2=11.797 $Y2=2.72
r217 121 123 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.945 $Y=2.72
+ $X2=12.19 $Y2=2.72
r218 120 154 4.33505 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=12.515 $Y=2.72
+ $X2=12.697 $Y2=2.72
r219 120 123 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.515 $Y=2.72
+ $X2=12.19 $Y2=2.72
r220 119 149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r221 119 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.89 $Y2=2.72
r222 118 146 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.35 $Y=2.72
+ $X2=10.07 $Y2=2.72
r223 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r224 115 148 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=10.68 $Y=2.72
+ $X2=10.795 $Y2=2.72
r225 115 118 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.68 $Y=2.72
+ $X2=10.35 $Y2=2.72
r226 114 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r227 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r228 111 142 2.06595 $w=5.48e-07 $l=9.5e-08 $layer=LI1_cond $X=9.795 $Y=2.53
+ $X2=9.89 $Y2=2.53
r229 111 113 17.9412 $w=5.48e-07 $l=8.25e-07 $layer=LI1_cond $X=9.795 $Y=2.53
+ $X2=8.97 $Y2=2.53
r230 110 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r231 110 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=7.59 $Y2=2.72
r232 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r233 107 138 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.715 $Y=2.72
+ $X2=7.525 $Y2=2.72
r234 107 109 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=7.715 $Y=2.72
+ $X2=8.51 $Y2=2.72
r235 106 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r236 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r237 103 106 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r238 102 105 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r239 102 103 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r240 100 138 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.525 $Y2=2.72
r241 100 105 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.13 $Y2=2.72
r242 99 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r243 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r244 96 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r245 96 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r246 95 98 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r247 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r248 93 132 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.8 $Y=2.72
+ $X2=3.61 $Y2=2.72
r249 93 95 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.8 $Y=2.72
+ $X2=3.91 $Y2=2.72
r250 92 133 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r251 92 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r252 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r253 89 129 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.615 $Y2=2.72
r254 89 91 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r255 88 132 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.42 $Y=2.72
+ $X2=3.61 $Y2=2.72
r256 88 91 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.42 $Y=2.72
+ $X2=2.07 $Y2=2.72
r257 87 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r258 87 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r259 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r260 84 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r261 84 86 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r262 83 129 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.615 $Y2=2.72
r263 83 86 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=2.72
+ $X2=1.15 $Y2=2.72
r264 77 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r265 75 127 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r266 75 158 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r267 73 77 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r268 73 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r269 72 109 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.655 $Y=2.72
+ $X2=8.51 $Y2=2.72
r270 71 72 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.82 $Y=2.53
+ $X2=8.655 $Y2=2.53
r271 68 113 0.869875 $w=5.48e-07 $l=4e-08 $layer=LI1_cond $X=8.93 $Y=2.53
+ $X2=8.97 $Y2=2.53
r272 68 71 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=8.93 $Y=2.53
+ $X2=8.82 $Y2=2.53
r273 66 98 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.89 $Y=2.72 $X2=4.83
+ $Y2=2.72
r274 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.89 $Y=2.72
+ $X2=5.055 $Y2=2.72
r275 65 102 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.22 $Y=2.72
+ $X2=5.29 $Y2=2.72
r276 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.22 $Y=2.72
+ $X2=5.055 $Y2=2.72
r277 61 64 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=12.655 $Y=1.63
+ $X2=12.655 $Y2=2.31
r278 59 154 3.02501 $w=2.8e-07 $l=1.03899e-07 $layer=LI1_cond $X=12.655 $Y=2.635
+ $X2=12.697 $Y2=2.72
r279 59 64 13.3766 $w=2.78e-07 $l=3.25e-07 $layer=LI1_cond $X=12.655 $Y=2.635
+ $X2=12.655 $Y2=2.31
r280 55 151 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=11.797 $Y=2.635
+ $X2=11.797 $Y2=2.72
r281 55 57 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=11.797 $Y=2.635
+ $X2=11.797 $Y2=1.94
r282 54 148 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=10.91 $Y=2.72
+ $X2=10.795 $Y2=2.72
r283 53 151 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=11.65 $Y=2.72
+ $X2=11.797 $Y2=2.72
r284 53 54 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.65 $Y=2.72
+ $X2=10.91 $Y2=2.72
r285 49 52 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.795 $Y=1.63
+ $X2=10.795 $Y2=2.31
r286 47 148 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.795 $Y=2.635
+ $X2=10.795 $Y2=2.72
r287 47 52 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=10.795 $Y=2.635
+ $X2=10.795 $Y2=2.31
r288 43 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=2.635
+ $X2=5.055 $Y2=2.72
r289 43 45 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.055 $Y=2.635
+ $X2=5.055 $Y2=2
r290 39 132 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=2.635
+ $X2=3.61 $Y2=2.72
r291 39 41 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=3.61 $Y=2.635
+ $X2=3.61 $Y2=2.29
r292 35 129 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=2.635
+ $X2=1.615 $Y2=2.72
r293 35 37 14.0666 $w=3.38e-07 $l=4.15e-07 $layer=LI1_cond $X=1.615 $Y=2.635
+ $X2=1.615 $Y2=2.22
r294 31 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r295 31 33 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r296 10 64 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.62 $Y2=2.31
r297 10 61 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.62 $Y2=1.63
r298 9 57 300 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=2 $X=11.59
+ $Y=1.765 $X2=11.78 $Y2=1.94
r299 8 52 400 $w=1.7e-07 $l=9.08295e-07 $layer=licon1_PDIFF $count=1 $X=10.61
+ $Y=1.485 $X2=10.785 $Y2=2.31
r300 8 49 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.61
+ $Y=1.485 $X2=10.785 $Y2=1.63
r301 7 145 600 $w=1.7e-07 $l=9.29637e-07 $layer=licon1_PDIFF $count=1 $X=9.705
+ $Y=1.505 $X2=9.905 $Y2=2.34
r302 6 71 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=8.685
+ $Y=1.645 $X2=8.82 $Y2=2.34
r303 5 135 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=7.305
+ $Y=2.065 $X2=7.5 $Y2=2.34
r304 4 45 300 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_PDIFF $count=2 $X=4.87
+ $Y=1.645 $X2=5.055 $Y2=2
r305 3 41 600 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=2.065 $X2=3.585 $Y2=2.29
r306 2 37 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.065 $X2=1.62 $Y2=2.22
r307 1 33 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_381_47# 1 2 8 9 10 11 12 15 19
r58 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=1.965
+ $X2=2.04 $Y2=2.3
r59 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r60 11 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.965
r61 11 12 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.59 $Y2=1.88
r62 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r63 9 10 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=1.59 $Y2=0.73
r64 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=1.795
+ $X2=1.59 $Y2=1.88
r65 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.505 $Y=0.825
+ $X2=1.59 $Y2=0.73
r66 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.505 $Y=0.825
+ $X2=1.505 $Y2=1.795
r67 2 19 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.065 $X2=2.04 $Y2=2.3
r68 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%Q_N 1 2 9 10 11 12 13 18 21
r23 18 21 3.51923 $w=2.6e-07 $l=7.5e-08 $layer=LI1_cond $X=10.37 $Y=0.585
+ $X2=10.37 $Y2=0.51
r24 12 13 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=10.37 $Y=1.815
+ $X2=10.37 $Y2=2.21
r25 11 30 6.64242 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=10.37 $Y=0.59
+ $X2=10.37 $Y2=0.715
r26 11 18 0.221624 $w=2.58e-07 $l=5e-09 $layer=LI1_cond $X=10.37 $Y=0.59
+ $X2=10.37 $Y2=0.585
r27 11 21 0.234615 $w=2.6e-07 $l=5e-09 $layer=LI1_cond $X=10.37 $Y=0.505
+ $X2=10.37 $Y2=0.51
r28 10 30 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=10.41 $Y=1.63
+ $X2=10.41 $Y2=0.715
r29 9 12 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=10.37 $Y=1.76
+ $X2=10.37 $Y2=1.815
r30 9 10 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=10.37 $Y=1.76
+ $X2=10.37 $Y2=1.63
r31 2 12 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=10.19
+ $Y=1.485 $X2=10.325 $Y2=1.815
r32 1 21 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=10.19
+ $Y=0.235 $X2=10.325 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%Q 1 2 10 11 12 13 14 15
c22 11 0 1.58152e-19 $X=12.23 $Y=1.56
c23 10 0 1.45535e-19 $X=12.23 $Y=0.825
r24 14 15 19.5414 $w=2.28e-07 $l=3.9e-07 $layer=LI1_cond $X=12.23 $Y=1.82
+ $X2=12.23 $Y2=2.21
r25 11 14 13.0276 $w=2.28e-07 $l=2.6e-07 $layer=LI1_cond $X=12.23 $Y=1.56
+ $X2=12.23 $Y2=1.82
r26 11 12 6.23684 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=12.23 $Y=1.56
+ $X2=12.23 $Y2=1.445
r27 10 12 37.1695 $w=1.83e-07 $l=6.2e-07 $layer=LI1_cond $X=12.252 $Y=0.825
+ $X2=12.252 $Y2=1.445
r28 9 13 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=12.23 $Y=0.71 $X2=12.23
+ $Y2=0.51
r29 9 10 6.23684 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=12.23 $Y=0.71
+ $X2=12.23 $Y2=0.825
r30 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=12.065
+ $Y=1.485 $X2=12.2 $Y2=1.82
r31 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=12.065
+ $Y=0.235 $X2=12.2 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 56 60 62 64 67 68 70 71 73 74 75 77 79 85 86 110 117 122 128 131 134 137 140
+ 144 147
c207 144 0 2.71124e-20 $X=12.65 $Y=0
c208 46 0 1.0279e-19 $X=7.45 $Y=0.36
r209 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r210 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r211 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r212 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r213 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r214 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r215 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r216 126 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=12.65 $Y2=0
r217 126 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r218 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r219 123 140 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=11.945 $Y=0
+ $X2=11.797 $Y2=0
r220 123 125 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.945 $Y=0
+ $X2=12.19 $Y2=0
r221 122 143 4.33505 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.697 $Y2=0
r222 122 125 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.19 $Y2=0
r223 121 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r224 121 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=9.89 $Y2=0
r225 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r226 118 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.07 $Y=0
+ $X2=9.905 $Y2=0
r227 118 120 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.07 $Y=0
+ $X2=10.35 $Y2=0
r228 117 137 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=10.68 $Y=0
+ $X2=10.795 $Y2=0
r229 117 120 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.68 $Y=0
+ $X2=10.35 $Y2=0
r230 116 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r231 115 116 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r232 113 116 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r233 112 115 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r234 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r235 110 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.74 $Y=0
+ $X2=9.905 $Y2=0
r236 110 115 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.74 $Y=0
+ $X2=9.43 $Y2=0
r237 109 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r238 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r239 106 109 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=7.13 $Y2=0
r240 105 108 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=7.13 $Y2=0
r241 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r242 103 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r243 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r244 100 103 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r245 99 102 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r246 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r247 97 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r248 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r249 94 97 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r250 94 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r251 93 96 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r252 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r253 91 131 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.615 $Y2=0
r254 91 93 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r255 90 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r256 90 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r257 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r258 87 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r259 87 89 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r260 86 131 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.445 $Y=0
+ $X2=1.615 $Y2=0
r261 86 89 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.15
+ $Y2=0
r262 79 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r263 79 85 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.245
+ $Y2=0
r264 77 129 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r265 77 147 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r266 75 85 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.245
+ $Y2=0
r267 75 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r268 73 108 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.13 $Y2=0
r269 73 74 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.275 $Y=0 $X2=7.405
+ $Y2=0
r270 72 112 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.535 $Y=0
+ $X2=7.59 $Y2=0
r271 72 74 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.405
+ $Y2=0
r272 70 102 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.29
+ $Y2=0
r273 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.525
+ $Y2=0
r274 69 105 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.69 $Y=0 $X2=5.75
+ $Y2=0
r275 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.69 $Y=0 $X2=5.525
+ $Y2=0
r276 67 96 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.45
+ $Y2=0
r277 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.665
+ $Y2=0
r278 66 99 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.91
+ $Y2=0
r279 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.665
+ $Y2=0
r280 62 143 3.02501 $w=2.8e-07 $l=1.03899e-07 $layer=LI1_cond $X=12.655 $Y=0.085
+ $X2=12.697 $Y2=0
r281 62 64 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=12.655 $Y=0.085
+ $X2=12.655 $Y2=0.38
r282 58 140 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=11.797 $Y=0.085
+ $X2=11.797 $Y2=0
r283 58 60 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=11.797 $Y=0.085
+ $X2=11.797 $Y2=0.38
r284 57 137 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=10.91 $Y=0
+ $X2=10.795 $Y2=0
r285 56 140 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=11.797 $Y2=0
r286 56 57 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=10.91 $Y2=0
r287 52 137 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.795 $Y=0.085
+ $X2=10.795 $Y2=0
r288 52 54 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.795 $Y=0.085
+ $X2=10.795 $Y2=0.38
r289 48 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.905 $Y=0.085
+ $X2=9.905 $Y2=0
r290 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.905 $Y=0.085
+ $X2=9.905 $Y2=0.38
r291 44 74 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=0.085
+ $X2=7.405 $Y2=0
r292 44 46 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=7.405 $Y=0.085
+ $X2=7.405 $Y2=0.36
r293 40 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.525 $Y=0.085
+ $X2=5.525 $Y2=0
r294 40 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.525 $Y=0.085
+ $X2=5.525 $Y2=0.38
r295 36 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=0.085
+ $X2=3.665 $Y2=0
r296 36 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.665 $Y=0.085
+ $X2=3.665 $Y2=0.36
r297 32 131 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0
r298 32 34 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.38
r299 28 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r300 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r301 9 64 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.485
+ $Y=0.235 $X2=12.62 $Y2=0.38
r302 8 60 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=11.59
+ $Y=0.235 $X2=11.78 $Y2=0.38
r303 7 54 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=10.61
+ $Y=0.235 $X2=10.785 $Y2=0.38
r304 6 50 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=9.705
+ $Y=0.235 $X2=9.905 $Y2=0.38
r305 5 46 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.305
+ $Y=0.235 $X2=7.45 $Y2=0.36
r306 4 42 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.235 $X2=5.525 $Y2=0.38
r307 3 38 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.235 $X2=3.665 $Y2=0.36
r308 2 34 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r309 1 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_790_47# 1 2 7 11 13
c28 13 0 7.56837e-20 $X=4.085 $Y=0.34
r29 13 16 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.085 $Y=0.34
+ $X2=4.085 $Y2=0.46
r30 9 11 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.045 $Y=0.425
+ $X2=5.045 $Y2=0.55
r31 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.25 $Y=0.34
+ $X2=4.085 $Y2=0.34
r32 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.92 $Y=0.34
+ $X2=5.045 $Y2=0.425
r33 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.92 $Y=0.34 $X2=4.25
+ $Y2=0.34
r34 2 11 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=5.005 $Y2=0.55
r35 1 16 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.235 $X2=4.085 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_2%A_1547_47# 1 2 7 9 16
r22 9 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.96 $Y=0.34 $X2=7.96
+ $Y2=0.46
r23 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=0.34 $X2=7.96
+ $Y2=0.34
r24 7 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.795 $Y=0.34
+ $X2=8.88 $Y2=0.34
r25 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.795 $Y=0.34
+ $X2=8.125 $Y2=0.34
r26 2 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.745
+ $Y=0.235 $X2=8.88 $Y2=0.42
r27 1 12 182 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=1 $X=7.735
+ $Y=0.235 $X2=7.96 $Y2=0.46
.ends


* File: sky130_fd_sc_hd__sdfsbp_2.pxi.spice
* Created: Tue Sep  1 19:30:37 2020
* 
x_PM_SKY130_FD_SC_HD__SDFSBP_2%SCD N_SCD_c_295_n N_SCD_c_299_n N_SCD_c_296_n
+ N_SCD_M1041_g N_SCD_c_300_n N_SCD_M1025_g N_SCD_c_301_n SCD SCD
+ PM_SKY130_FD_SC_HD__SDFSBP_2%SCD
x_PM_SKY130_FD_SC_HD__SDFSBP_2%SCE N_SCE_M1016_g N_SCE_c_328_n N_SCE_M1001_g
+ N_SCE_M1024_g N_SCE_M1029_g SCE N_SCE_c_331_n N_SCE_c_352_n N_SCE_c_332_n
+ N_SCE_c_333_n N_SCE_c_334_n PM_SKY130_FD_SC_HD__SDFSBP_2%SCE
x_PM_SKY130_FD_SC_HD__SDFSBP_2%D N_D_c_433_n N_D_M1027_g N_D_M1004_g D D
+ N_D_c_436_n PM_SKY130_FD_SC_HD__SDFSBP_2%D
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_328_21# N_A_328_21#_M1024_s N_A_328_21#_M1029_s
+ N_A_328_21#_M1036_g N_A_328_21#_M1032_g N_A_328_21#_c_477_n
+ N_A_328_21#_c_478_n N_A_328_21#_c_479_n N_A_328_21#_c_480_n
+ N_A_328_21#_c_484_n N_A_328_21#_c_485_n PM_SKY130_FD_SC_HD__SDFSBP_2%A_328_21#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%CLK N_CLK_c_561_n N_CLK_c_555_n N_CLK_M1003_g
+ N_CLK_c_562_n N_CLK_M1010_g N_CLK_c_556_n N_CLK_c_563_n CLK CLK CLK CLK
+ N_CLK_c_559_n N_CLK_c_560_n PM_SKY130_FD_SC_HD__SDFSBP_2%CLK
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_652_47# N_A_652_47#_M1003_s N_A_652_47#_M1010_s
+ N_A_652_47#_c_633_n N_A_652_47#_c_634_n N_A_652_47#_M1045_g
+ N_A_652_47#_c_635_n N_A_652_47#_M1031_g N_A_652_47#_c_636_n
+ N_A_652_47#_c_637_n N_A_652_47#_M1030_g N_A_652_47#_M1034_g
+ N_A_652_47#_M1021_g N_A_652_47#_M1018_g N_A_652_47#_c_639_n
+ N_A_652_47#_c_640_n N_A_652_47#_c_665_n N_A_652_47#_c_641_n
+ N_A_652_47#_c_642_n N_A_652_47#_c_654_n N_A_652_47#_c_655_n
+ N_A_652_47#_c_729_p N_A_652_47#_c_643_n N_A_652_47#_c_644_n
+ N_A_652_47#_c_645_n N_A_652_47#_c_646_n N_A_652_47#_c_647_n
+ N_A_652_47#_c_648_n N_A_652_47#_c_649_n N_A_652_47#_c_714_p
+ N_A_652_47#_c_659_n N_A_652_47#_c_731_p N_A_652_47#_c_660_n
+ N_A_652_47#_c_661_n N_A_652_47#_c_775_p N_A_652_47#_c_662_n
+ N_A_652_47#_c_663_n PM_SKY130_FD_SC_HD__SDFSBP_2%A_652_47#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_818_47# N_A_818_47#_M1045_d N_A_818_47#_M1031_d
+ N_A_818_47#_c_933_n N_A_818_47#_c_921_n N_A_818_47#_c_934_n
+ N_A_818_47#_M1007_g N_A_818_47#_c_922_n N_A_818_47#_M1019_g
+ N_A_818_47#_M1043_g N_A_818_47#_c_936_n N_A_818_47#_M1039_g
+ N_A_818_47#_c_938_n N_A_818_47#_c_924_n N_A_818_47#_c_925_n
+ N_A_818_47#_c_973_n N_A_818_47#_c_939_n N_A_818_47#_c_940_n
+ N_A_818_47#_c_926_n N_A_818_47#_c_927_n N_A_818_47#_c_928_n
+ N_A_818_47#_c_929_n N_A_818_47#_c_930_n N_A_818_47#_c_931_n
+ N_A_818_47#_c_932_n PM_SKY130_FD_SC_HD__SDFSBP_2%A_818_47#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_1132_21# N_A_1132_21#_M1002_s
+ N_A_1132_21#_M1008_d N_A_1132_21#_M1022_g N_A_1132_21#_c_1115_n
+ N_A_1132_21#_M1044_g N_A_1132_21#_c_1123_n N_A_1132_21#_c_1124_n
+ N_A_1132_21#_c_1116_n N_A_1132_21#_c_1125_n N_A_1132_21#_c_1126_n
+ N_A_1132_21#_c_1117_n N_A_1132_21#_c_1194_p N_A_1132_21#_c_1118_n
+ N_A_1132_21#_c_1119_n N_A_1132_21#_c_1120_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%A_1132_21#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_1006_47# N_A_1006_47#_M1030_d
+ N_A_1006_47#_M1007_d N_A_1006_47#_M1008_g N_A_1006_47#_c_1216_n
+ N_A_1006_47#_M1002_g N_A_1006_47#_M1023_g N_A_1006_47#_M1015_g
+ N_A_1006_47#_c_1217_n N_A_1006_47#_c_1218_n N_A_1006_47#_c_1245_n
+ N_A_1006_47#_c_1219_n N_A_1006_47#_c_1220_n N_A_1006_47#_c_1234_n
+ N_A_1006_47#_c_1221_n N_A_1006_47#_c_1222_n N_A_1006_47#_c_1223_n
+ N_A_1006_47#_c_1224_n N_A_1006_47#_c_1225_n N_A_1006_47#_c_1226_n
+ N_A_1006_47#_c_1227_n N_A_1006_47#_c_1228_n N_A_1006_47#_c_1229_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%A_1006_47#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%SET_B N_SET_B_M1033_g N_SET_B_M1037_g
+ N_SET_B_c_1378_n N_SET_B_M1013_g N_SET_B_M1014_g N_SET_B_c_1376_n
+ N_SET_B_c_1381_n N_SET_B_c_1382_n N_SET_B_c_1383_n N_SET_B_c_1384_n SET_B
+ N_SET_B_c_1385_n N_SET_B_c_1386_n N_SET_B_c_1387_n N_SET_B_c_1388_n
+ N_SET_B_c_1389_n N_SET_B_c_1390_n N_SET_B_c_1391_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%SET_B
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_1781_295# N_A_1781_295#_M1000_d
+ N_A_1781_295#_M1026_d N_A_1781_295#_M1009_g N_A_1781_295#_c_1518_n
+ N_A_1781_295#_c_1519_n N_A_1781_295#_M1020_g N_A_1781_295#_c_1511_n
+ N_A_1781_295#_c_1512_n N_A_1781_295#_c_1513_n N_A_1781_295#_c_1514_n
+ N_A_1781_295#_c_1522_n N_A_1781_295#_c_1523_n N_A_1781_295#_c_1515_n
+ N_A_1781_295#_c_1516_n N_A_1781_295#_c_1524_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%A_1781_295#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_1597_329# N_A_1597_329#_M1043_d
+ N_A_1597_329#_M1021_d N_A_1597_329#_M1013_d N_A_1597_329#_c_1613_n
+ N_A_1597_329#_M1000_g N_A_1597_329#_c_1614_n N_A_1597_329#_M1026_g
+ N_A_1597_329#_c_1615_n N_A_1597_329#_c_1616_n N_A_1597_329#_M1035_g
+ N_A_1597_329#_M1012_g N_A_1597_329#_c_1617_n N_A_1597_329#_M1038_g
+ N_A_1597_329#_M1028_g N_A_1597_329#_c_1618_n N_A_1597_329#_c_1619_n
+ N_A_1597_329#_M1011_g N_A_1597_329#_M1005_g N_A_1597_329#_c_1621_n
+ N_A_1597_329#_c_1644_n N_A_1597_329#_c_1645_n N_A_1597_329#_c_1634_n
+ N_A_1597_329#_c_1635_n N_A_1597_329#_c_1622_n N_A_1597_329#_c_1623_n
+ N_A_1597_329#_c_1624_n N_A_1597_329#_c_1636_n N_A_1597_329#_c_1637_n
+ N_A_1597_329#_c_1638_n N_A_1597_329#_c_1639_n N_A_1597_329#_c_1679_n
+ N_A_1597_329#_c_1640_n PM_SKY130_FD_SC_HD__SDFSBP_2%A_1597_329#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_2501_47# N_A_2501_47#_M1011_s
+ N_A_2501_47#_M1005_s N_A_2501_47#_c_1793_n N_A_2501_47#_M1040_g
+ N_A_2501_47#_M1006_g N_A_2501_47#_c_1794_n N_A_2501_47#_M1042_g
+ N_A_2501_47#_M1017_g N_A_2501_47#_c_1795_n N_A_2501_47#_c_1800_n
+ N_A_2501_47#_c_1796_n N_A_2501_47#_c_1811_n N_A_2501_47#_c_1797_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%A_2501_47#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_27_369# N_A_27_369#_M1025_s N_A_27_369#_M1032_d
+ N_A_27_369#_c_1853_n N_A_27_369#_c_1867_n N_A_27_369#_c_1868_n
+ N_A_27_369#_c_1854_n N_A_27_369#_c_1855_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%A_27_369#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%VPWR N_VPWR_M1025_d N_VPWR_M1029_d N_VPWR_M1010_d
+ N_VPWR_M1044_d N_VPWR_M1033_d N_VPWR_M1009_d N_VPWR_M1026_s N_VPWR_M1012_d
+ N_VPWR_M1028_d N_VPWR_M1005_d N_VPWR_M1017_d N_VPWR_c_1895_n N_VPWR_c_1896_n
+ N_VPWR_c_1897_n N_VPWR_c_1898_n N_VPWR_c_1899_n N_VPWR_c_1900_n
+ N_VPWR_c_1901_n N_VPWR_c_1902_n N_VPWR_c_1903_n N_VPWR_c_1904_n
+ N_VPWR_c_1905_n N_VPWR_c_1906_n N_VPWR_c_1907_n N_VPWR_c_1908_n
+ N_VPWR_c_1909_n N_VPWR_c_1910_n N_VPWR_c_1911_n VPWR N_VPWR_c_1912_n
+ N_VPWR_c_1913_n N_VPWR_c_1914_n N_VPWR_c_1915_n N_VPWR_c_1916_n
+ N_VPWR_c_1917_n N_VPWR_c_1918_n N_VPWR_c_1919_n N_VPWR_c_1920_n
+ N_VPWR_c_1921_n N_VPWR_c_1922_n N_VPWR_c_1923_n N_VPWR_c_1924_n
+ N_VPWR_c_1925_n N_VPWR_c_1926_n N_VPWR_c_1894_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%VPWR
x_PM_SKY130_FD_SC_HD__SDFSBP_2%A_181_47# N_A_181_47#_M1016_d N_A_181_47#_M1030_s
+ N_A_181_47#_M1004_d N_A_181_47#_M1007_s N_A_181_47#_c_2116_n
+ N_A_181_47#_c_2117_n N_A_181_47#_c_2121_n N_A_181_47#_c_2122_n
+ N_A_181_47#_c_2118_n N_A_181_47#_c_2132_n N_A_181_47#_c_2119_n
+ N_A_181_47#_c_2124_n N_A_181_47#_c_2125_n N_A_181_47#_c_2120_n
+ N_A_181_47#_c_2127_n PM_SKY130_FD_SC_HD__SDFSBP_2%A_181_47#
x_PM_SKY130_FD_SC_HD__SDFSBP_2%Q_N N_Q_N_M1035_s N_Q_N_M1012_s Q_N Q_N Q_N Q_N
+ Q_N Q_N N_Q_N_c_2249_n PM_SKY130_FD_SC_HD__SDFSBP_2%Q_N
x_PM_SKY130_FD_SC_HD__SDFSBP_2%Q N_Q_M1040_s N_Q_M1006_s Q Q Q Q Q Q
+ N_Q_c_2273_n Q Q PM_SKY130_FD_SC_HD__SDFSBP_2%Q
x_PM_SKY130_FD_SC_HD__SDFSBP_2%VGND N_VGND_M1041_s N_VGND_M1036_d N_VGND_M1024_d
+ N_VGND_M1003_d N_VGND_M1022_d N_VGND_M1037_d N_VGND_M1014_d N_VGND_M1035_d
+ N_VGND_M1038_d N_VGND_M1011_d N_VGND_M1042_d N_VGND_c_2290_n N_VGND_c_2291_n
+ N_VGND_c_2292_n N_VGND_c_2293_n N_VGND_c_2294_n N_VGND_c_2295_n
+ N_VGND_c_2296_n N_VGND_c_2297_n N_VGND_c_2298_n N_VGND_c_2299_n
+ N_VGND_c_2300_n N_VGND_c_2301_n N_VGND_c_2302_n N_VGND_c_2303_n
+ N_VGND_c_2304_n VGND N_VGND_c_2305_n N_VGND_c_2306_n N_VGND_c_2307_n
+ N_VGND_c_2308_n N_VGND_c_2309_n N_VGND_c_2310_n N_VGND_c_2311_n
+ N_VGND_c_2312_n N_VGND_c_2313_n N_VGND_c_2314_n N_VGND_c_2315_n
+ N_VGND_c_2316_n N_VGND_c_2317_n N_VGND_c_2318_n N_VGND_c_2319_n
+ PM_SKY130_FD_SC_HD__SDFSBP_2%VGND
cc_1 VNB N_SCD_c_295_n 0.0592907f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.325
cc_2 VNB N_SCD_c_296_n 0.017218f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB SCD 0.0208496f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_SCE_M1016_g 0.030725f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_5 VNB N_SCE_c_328_n 0.0195372f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_6 VNB N_SCE_M1024_g 0.0378941f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.695
cc_7 VNB SCE 0.00509679f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_8 VNB N_SCE_c_331_n 0.00914897f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_9 VNB N_SCE_c_332_n 0.00100889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_333_n 0.00258872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_SCE_c_334_n 0.0261434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_D_c_433_n 0.0167893f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.325
cc_13 VNB N_D_M1004_g 0.00900213f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.77
cc_14 VNB D 0.00525725f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_15 VNB N_D_c_436_n 0.0258198f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_16 VNB N_A_328_21#_M1036_g 0.0312417f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_17 VNB N_A_328_21#_c_477_n 0.00409066f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_18 VNB N_A_328_21#_c_478_n 0.039298f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_19 VNB N_A_328_21#_c_479_n 0.0124639f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_20 VNB N_A_328_21#_c_480_n 0.00706038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_CLK_c_555_n 0.0170609f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_22 VNB N_CLK_c_556_n 0.0152719f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_23 VNB CLK 0.0102177f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_24 VNB CLK 0.0134917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_CLK_c_559_n 0.0163974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_CLK_c_560_n 0.0133326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_652_47#_c_633_n 0.0110155f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_28 VNB N_A_652_47#_c_634_n 0.0173626f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_29 VNB N_A_652_47#_c_635_n 0.0160921f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_652_47#_c_636_n 0.0510371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_652_47#_c_637_n 0.0179438f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_32 VNB N_A_652_47#_M1018_g 0.0241734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_652_47#_c_639_n 0.00632952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_652_47#_c_640_n 0.00133693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_652_47#_c_641_n 0.00586117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_652_47#_c_642_n 0.00227297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_652_47#_c_643_n 0.00316033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_652_47#_c_644_n 0.00199626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_652_47#_c_645_n 0.0263197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_652_47#_c_646_n 0.00960826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_652_47#_c_647_n 2.52613e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_652_47#_c_648_n 0.00451712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_652_47#_c_649_n 0.0280058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_818_47#_c_921_n 0.0383145f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_45 VNB N_A_818_47#_c_922_n 0.0129031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_818_47#_M1043_g 0.036405f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_818_47#_c_924_n 0.0136171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_818_47#_c_925_n 0.00923607f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_818_47#_c_926_n 0.0188967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_818_47#_c_927_n 0.0027097f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_818_47#_c_928_n 0.00326418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_818_47#_c_929_n 0.00365861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_818_47#_c_930_n 0.00174312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_818_47#_c_931_n 0.0191844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_818_47#_c_932_n 0.0048019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1132_21#_c_1115_n 0.0107737f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.695
cc_57 VNB N_A_1132_21#_c_1116_n 0.00766843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1132_21#_c_1117_n 0.00385507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1132_21#_c_1118_n 0.0057123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1132_21#_c_1119_n 0.0297274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1132_21#_c_1120_n 0.0171303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1006_47#_c_1216_n 0.0162044f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_63 VNB N_A_1006_47#_c_1217_n 0.0213622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1006_47#_c_1218_n 0.00675227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1006_47#_c_1219_n 0.00237615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1006_47#_c_1220_n 0.00215563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1006_47#_c_1221_n 6.99033e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1006_47#_c_1222_n 0.0188701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1006_47#_c_1223_n 0.00170342f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1006_47#_c_1224_n 0.00230045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1006_47#_c_1225_n 0.00355589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1006_47#_c_1226_n 0.0209471f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1006_47#_c_1227_n 0.0113035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1006_47#_c_1228_n 0.012284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1006_47#_c_1229_n 0.0192224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_SET_B_M1037_g 0.0360613f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_77 VNB N_SET_B_M1014_g 0.0433163f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_SET_B_c_1376_n 0.00656881f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_79 VNB N_A_1781_295#_M1020_g 0.0213855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1781_295#_c_1511_n 0.00630515f $X=-0.19 $Y=-0.24 $X2=0.255
+ $Y2=1.16
cc_81 VNB N_A_1781_295#_c_1512_n 0.00102967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1781_295#_c_1513_n 0.0287182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1781_295#_c_1514_n 0.00638132f $X=-0.19 $Y=-0.24 $X2=0.212
+ $Y2=1.53
cc_84 VNB N_A_1781_295#_c_1515_n 0.00904914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1781_295#_c_1516_n 0.00793305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1597_329#_c_1613_n 0.0201172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1597_329#_c_1614_n 0.0360377f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=0.765
cc_88 VNB N_A_1597_329#_c_1615_n 0.0480885f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_89 VNB N_A_1597_329#_c_1616_n 0.0193019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1597_329#_c_1617_n 0.0197007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1597_329#_c_1618_n 0.0513144f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_1597_329#_c_1619_n 0.021326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_1597_329#_M1011_g 0.0319861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_1597_329#_c_1621_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_1597_329#_c_1622_n 0.00189779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_1597_329#_c_1623_n 0.00171166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_1597_329#_c_1624_n 0.00888098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_2501_47#_c_1793_n 0.0167001f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_99 VNB N_A_2501_47#_c_1794_n 0.0215032f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_100 VNB N_A_2501_47#_c_1795_n 0.00685394f $X=-0.19 $Y=-0.24 $X2=0.212
+ $Y2=1.16
cc_101 VNB N_A_2501_47#_c_1796_n 0.00194757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_A_2501_47#_c_1797_n 0.0478635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VPWR_c_1894_n 0.592346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_A_181_47#_c_2116_n 7.98501e-19 $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=0.765
cc_105 VNB N_A_181_47#_c_2117_n 0.00536944f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_106 VNB N_A_181_47#_c_2118_n 0.00335328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_A_181_47#_c_2119_n 0.00147615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_A_181_47#_c_2120_n 0.00327965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB Q 0.00106334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2290_n 0.00752609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2291_n 0.00701999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2292_n 0.0025484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2293_n 0.00240024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2294_n 0.00645503f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2295_n 0.0143512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2296_n 0.00303296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2297_n 0.0100096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2298_n 0.0337748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2299_n 0.0281049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2300_n 0.00477715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2301_n 0.0588928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2302_n 0.00356769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2303_n 0.0212793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2304_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2305_n 0.015123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2306_n 0.0135577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2307_n 0.0437877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2308_n 0.0193843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2309_n 0.0153065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2310_n 0.0182896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2311_n 0.0338415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2312_n 0.00642278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2313_n 0.00449945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2314_n 0.0134872f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2315_n 0.013792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2316_n 0.0173854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2317_n 0.00557475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2318_n 0.00558559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2319_n 0.668909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VPB N_SCD_c_295_n 0.00536633f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.325
cc_141 VPB N_SCD_c_299_n 0.019303f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.62
cc_142 VPB N_SCD_c_300_n 0.0190089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.77
cc_143 VPB N_SCD_c_301_n 0.0259455f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_144 VPB SCD 0.0148037f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_145 VPB N_SCE_c_328_n 0.0133475f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_146 VPB N_SCE_M1001_g 0.0314422f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_147 VPB N_SCE_M1029_g 0.0499623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB SCE 0.00452509f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_149 VPB N_SCE_c_333_n 0.00426864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_SCE_c_334_n 0.00558169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_D_M1004_g 0.0348977f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.77
cc_152 VPB D 0.00582207f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_153 VPB N_A_328_21#_M1032_g 0.0429677f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_154 VPB N_A_328_21#_c_477_n 0.00918755f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_155 VPB N_A_328_21#_c_478_n 0.0147307f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_156 VPB N_A_328_21#_c_484_n 0.00509652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_328_21#_c_485_n 0.0114079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_CLK_c_561_n 0.0106726f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_159 VPB N_CLK_c_562_n 0.0174348f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_160 VPB N_CLK_c_563_n 0.0183991f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_161 VPB CLK 0.00879878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB CLK 0.0143572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_CLK_c_559_n 0.0103664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_652_47#_c_635_n 0.0272914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_652_47#_M1031_g 0.021706f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_166 VPB N_A_652_47#_M1034_g 0.0194363f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_167 VPB N_A_652_47#_M1021_g 0.0245732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_652_47#_c_654_n 9.44198e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_652_47#_c_655_n 0.00140884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_652_47#_c_643_n 0.00351449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_652_47#_c_644_n 0.0023723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_652_47#_c_645_n 0.00502468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_652_47#_c_659_n 0.00655951f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_652_47#_c_660_n 0.00699976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_652_47#_c_661_n 0.00163014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_652_47#_c_662_n 0.0309552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_652_47#_c_663_n 0.00480233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_818_47#_c_933_n 0.0245892f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_179 VPB N_A_818_47#_c_934_n 0.0183942f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_180 VPB N_A_818_47#_M1043_g 0.0159101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_818_47#_c_936_n 0.0362831f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_182 VPB N_A_818_47#_M1039_g 0.0213627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_818_47#_c_938_n 0.0280669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_818_47#_c_939_n 0.00416446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_818_47#_c_940_n 0.00953737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_818_47#_c_928_n 0.00121793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_818_47#_c_929_n 3.90977e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_818_47#_c_930_n 0.0046846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_818_47#_c_931_n 0.0195903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1132_21#_c_1115_n 0.0163932f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_191 VPB N_A_1132_21#_M1044_g 0.0207249f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_192 VPB N_A_1132_21#_c_1123_n 0.00186016f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_193 VPB N_A_1132_21#_c_1124_n 0.0378508f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_194 VPB N_A_1132_21#_c_1125_n 0.00527575f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.16
cc_195 VPB N_A_1132_21#_c_1126_n 7.27868e-19 $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.53
cc_196 VPB N_A_1006_47#_M1008_g 0.0474078f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_197 VPB N_A_1006_47#_M1015_g 0.0264674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1006_47#_c_1219_n 0.00213496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1006_47#_c_1220_n 0.00336726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1006_47#_c_1234_n 0.0124408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1006_47#_c_1222_n 0.00929565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_1006_47#_c_1223_n 0.00278293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1006_47#_c_1224_n 0.00131078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1006_47#_c_1225_n 9.00638e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1006_47#_c_1226_n 0.00612855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_SET_B_M1033_g 0.0241763f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_207 VPB N_SET_B_c_1378_n 0.0185321f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_208 VPB N_SET_B_M1014_g 0.00935824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_SET_B_c_1376_n 0.00612012f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_210 VPB N_SET_B_c_1381_n 0.0275591f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_211 VPB N_SET_B_c_1382_n 0.0119113f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_SET_B_c_1383_n 0.00718944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_SET_B_c_1384_n 0.0148843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_SET_B_c_1385_n 0.0175592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_SET_B_c_1386_n 0.00490784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_SET_B_c_1387_n 0.00625323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_SET_B_c_1388_n 0.0278775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_SET_B_c_1389_n 0.00931593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_SET_B_c_1390_n 0.00833156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_SET_B_c_1391_n 0.00385115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1781_295#_M1009_g 0.0341907f $X=-0.19 $Y=1.305 $X2=0.315
+ $Y2=1.695
cc_222 VPB N_A_1781_295#_c_1518_n 0.0265033f $X=-0.19 $Y=1.305 $X2=0.47
+ $Y2=1.695
cc_223 VPB N_A_1781_295#_c_1519_n 0.00628592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1781_295#_c_1511_n 0.0109338f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_225 VPB N_A_1781_295#_c_1514_n 0.00703029f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.53
cc_226 VPB N_A_1781_295#_c_1522_n 7.16388e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1781_295#_c_1523_n 0.0195654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1781_295#_c_1524_n 0.00297807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_1597_329#_c_1614_n 9.23577e-19 $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=0.765
cc_230 VPB N_A_1597_329#_M1026_g 0.0293397f $X=-0.19 $Y=1.305 $X2=0.325 $Y2=1.16
cc_231 VPB N_A_1597_329#_c_1615_n 0.0221781f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_232 VPB N_A_1597_329#_M1012_g 0.0222507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_1597_329#_M1028_g 0.022668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_1597_329#_c_1618_n 0.0252244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_1597_329#_c_1619_n 0.00378286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_1597_329#_M1005_g 0.0423423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_A_1597_329#_c_1621_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_1597_329#_c_1634_n 0.00734199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_A_1597_329#_c_1635_n 0.00462018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_1597_329#_c_1636_n 0.00531894f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_A_1597_329#_c_1637_n 0.00442575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_A_1597_329#_c_1638_n 0.0321498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_A_1597_329#_c_1639_n 0.00235934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_A_1597_329#_c_1640_n 0.0169018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_A_2501_47#_M1006_g 0.0193854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_A_2501_47#_M1017_g 0.0252966f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_247 VPB N_A_2501_47#_c_1800_n 0.0121614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_A_2501_47#_c_1796_n 0.00246016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_A_2501_47#_c_1797_n 0.00816398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_A_27_369#_c_1853_n 0.00117506f $X=-0.19 $Y=1.305 $X2=0.315
+ $Y2=1.695
cc_251 VPB N_A_27_369#_c_1854_n 0.00247045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_A_27_369#_c_1855_n 0.0266682f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_253 VPB N_VPWR_c_1895_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1896_n 0.00752066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1897_n 4.01796e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1898_n 0.0056301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1899_n 0.0026976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1900_n 0.00472716f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1901_n 0.00661141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1902_n 0.0180927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1903_n 0.00321952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1904_n 0.00998368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1905_n 0.0471703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1906_n 0.0271668f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1907_n 0.00507122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1908_n 0.0143691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1909_n 0.00507288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1910_n 0.0172878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1911_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1912_n 0.0143088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1913_n 0.0425618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1914_n 0.0141341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1915_n 0.0510056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1916_n 0.0193843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1917_n 0.0153065f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1918_n 0.0182605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1919_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1920_n 0.00632819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1921_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1922_n 0.00631318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1923_n 0.0199409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1924_n 0.0192332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1925_n 0.00554886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1926_n 0.0055597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1894_n 0.0825425f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_286 VPB N_A_181_47#_c_2121_n 0.00378515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_287 VPB N_A_181_47#_c_2122_n 0.0022281f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_288 VPB N_A_181_47#_c_2118_n 0.00201708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_289 VPB N_A_181_47#_c_2124_n 0.0273128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_290 VPB N_A_181_47#_c_2125_n 0.00231687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_291 VPB N_A_181_47#_c_2120_n 0.00329791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_292 VPB N_A_181_47#_c_2127_n 0.0042939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_293 VPB Q 0.00116001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_294 N_SCD_c_295_n N_SCE_M1016_g 0.00583208f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_295 N_SCD_c_296_n N_SCE_M1016_g 0.0484084f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_296 SCD N_SCE_M1016_g 2.56735e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_297 N_SCD_c_295_n N_SCE_c_328_n 0.0200842f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_298 SCD N_SCE_c_328_n 3.421e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_299 N_SCD_c_299_n N_SCE_M1001_g 0.00453523f $X=0.315 $Y=1.62 $X2=0 $Y2=0
cc_300 N_SCD_c_301_n N_SCE_M1001_g 0.0326857f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_301 SCD N_SCE_M1001_g 2.04234e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_302 N_SCD_c_295_n SCE 0.00799654f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_303 N_SCD_c_301_n SCE 0.00146655f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_304 SCD SCE 0.0593537f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_305 SCD N_SCE_c_352_n 0.00158165f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_306 N_SCD_c_300_n N_A_27_369#_c_1853_n 0.0154938f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_307 N_SCD_c_295_n N_A_27_369#_c_1855_n 5.05332e-19 $X=0.315 $Y=1.325 $X2=0
+ $Y2=0
cc_308 N_SCD_c_301_n N_A_27_369#_c_1855_n 0.00316572f $X=0.47 $Y=1.695 $X2=0
+ $Y2=0
cc_309 SCD N_A_27_369#_c_1855_n 0.0226954f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_310 N_SCD_c_300_n N_VPWR_c_1895_n 0.00808197f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_311 N_SCD_c_300_n N_VPWR_c_1912_n 0.00340533f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_312 N_SCD_c_300_n N_VPWR_c_1894_n 0.00499747f $X=0.47 $Y=1.77 $X2=0 $Y2=0
cc_313 N_SCD_c_296_n N_A_181_47#_c_2116_n 2.6495e-19 $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_314 N_SCD_c_295_n N_VGND_c_2311_n 0.00480402f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_315 N_SCD_c_296_n N_VGND_c_2311_n 0.0218413f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_316 SCD N_VGND_c_2311_n 0.0221354f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_317 SCD N_VGND_c_2319_n 9.88088e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_318 N_SCE_M1016_g N_D_c_433_n 0.0148828f $X=0.83 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_319 N_SCE_c_328_n N_D_M1004_g 0.0912898f $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_320 SCE N_D_M1004_g 6.11571e-19 $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_321 N_SCE_M1016_g D 0.00302957f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_322 N_SCE_c_328_n D 0.00293745f $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_323 SCE D 0.0531526f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_324 N_SCE_c_331_n D 0.0225619f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_325 N_SCE_c_352_n D 0.00219522f $X=0.835 $Y=1.19 $X2=0 $Y2=0
cc_326 N_SCE_M1016_g N_D_c_436_n 0.0194304f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_327 SCE N_D_c_436_n 3.39482e-19 $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_328 N_SCE_c_331_n N_D_c_436_n 0.00134139f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_329 N_SCE_M1024_g N_A_328_21#_c_477_n 0.00176491f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_330 N_SCE_M1029_g N_A_328_21#_c_477_n 0.00449189f $X=2.66 $Y=2.165 $X2=0
+ $Y2=0
cc_331 N_SCE_c_331_n N_A_328_21#_c_477_n 0.014286f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_332 N_SCE_c_332_n N_A_328_21#_c_477_n 0.00266192f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_333 N_SCE_c_333_n N_A_328_21#_c_477_n 0.0382385f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_334 N_SCE_c_334_n N_A_328_21#_c_477_n 0.0015262f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_335 N_SCE_c_331_n N_A_328_21#_c_478_n 0.0100047f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_336 N_SCE_c_333_n N_A_328_21#_c_478_n 6.13531e-19 $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_337 N_SCE_c_334_n N_A_328_21#_c_478_n 0.0184786f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_338 N_SCE_M1024_g N_A_328_21#_c_479_n 0.00518112f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_339 N_SCE_c_331_n N_A_328_21#_c_479_n 0.0076772f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_340 N_SCE_c_332_n N_A_328_21#_c_479_n 0.00404451f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_341 N_SCE_c_333_n N_A_328_21#_c_479_n 0.00808528f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_342 N_SCE_c_334_n N_A_328_21#_c_479_n 0.00234786f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_343 N_SCE_M1024_g N_A_328_21#_c_480_n 0.00283811f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_344 N_SCE_M1029_g N_A_328_21#_c_485_n 0.00222738f $X=2.66 $Y=2.165 $X2=0
+ $Y2=0
cc_345 N_SCE_c_333_n N_A_328_21#_c_485_n 0.00910591f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_346 N_SCE_c_334_n N_A_328_21#_c_485_n 4.11404e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_347 N_SCE_M1029_g N_CLK_c_561_n 0.0035615f $X=2.66 $Y=2.165 $X2=0 $Y2=0
cc_348 N_SCE_M1024_g N_CLK_c_556_n 0.00249428f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_349 N_SCE_M1024_g CLK 0.00341058f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_350 N_SCE_c_334_n CLK 9.32708e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_351 N_SCE_M1029_g CLK 0.0064941f $X=2.66 $Y=2.165 $X2=0 $Y2=0
cc_352 N_SCE_M1029_g CLK 3.68886e-19 $X=2.66 $Y=2.165 $X2=0 $Y2=0
cc_353 N_SCE_c_332_n CLK 0.00161909f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_354 N_SCE_c_333_n CLK 0.039758f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_355 N_SCE_c_334_n CLK 0.0027156f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_356 N_SCE_c_333_n N_CLK_c_559_n 2.49383e-19 $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_357 N_SCE_c_334_n N_CLK_c_559_n 0.00515768f $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_358 N_SCE_c_334_n N_CLK_c_560_n 9.62133e-19 $X=2.57 $Y=1.16 $X2=0 $Y2=0
cc_359 N_SCE_M1024_g N_A_652_47#_c_640_n 0.00355226f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_360 N_SCE_M1029_g N_A_652_47#_c_665_n 0.00356206f $X=2.66 $Y=2.165 $X2=0
+ $Y2=0
cc_361 N_SCE_M1024_g N_A_652_47#_c_642_n 5.26825e-19 $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_362 N_SCE_M1029_g N_A_652_47#_c_655_n 0.00106055f $X=2.66 $Y=2.165 $X2=0
+ $Y2=0
cc_363 N_SCE_c_328_n N_A_27_369#_c_1853_n 7.77528e-19 $X=0.89 $Y=1.415 $X2=0
+ $Y2=0
cc_364 N_SCE_M1001_g N_A_27_369#_c_1853_n 0.0145203f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_365 SCE N_A_27_369#_c_1853_n 0.0188059f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_366 N_SCE_c_331_n N_A_27_369#_c_1853_n 0.00676074f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_367 N_SCE_c_352_n N_A_27_369#_c_1853_n 0.00144701f $X=0.835 $Y=1.19 $X2=0
+ $Y2=0
cc_368 N_SCE_M1001_g N_VPWR_c_1895_n 0.00755808f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_369 N_SCE_M1029_g N_VPWR_c_1896_n 0.0113293f $X=2.66 $Y=2.165 $X2=0 $Y2=0
cc_370 N_SCE_c_333_n N_VPWR_c_1896_n 4.57941e-19 $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_371 N_SCE_M1001_g N_VPWR_c_1913_n 0.00340533f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_372 N_SCE_M1029_g N_VPWR_c_1913_n 0.0046653f $X=2.66 $Y=2.165 $X2=0 $Y2=0
cc_373 N_SCE_M1001_g N_VPWR_c_1894_n 0.00387201f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_374 N_SCE_M1029_g N_VPWR_c_1894_n 0.00934473f $X=2.66 $Y=2.165 $X2=0 $Y2=0
cc_375 N_SCE_M1016_g N_A_181_47#_c_2116_n 0.00473765f $X=0.83 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_SCE_c_328_n N_A_181_47#_c_2116_n 9.02625e-19 $X=0.89 $Y=1.415 $X2=0
+ $Y2=0
cc_377 N_SCE_c_331_n N_A_181_47#_c_2116_n 0.0130638f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_378 N_SCE_c_331_n N_A_181_47#_c_2132_n 0.00354885f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_379 N_SCE_M1029_g N_A_181_47#_c_2124_n 0.00717814f $X=2.66 $Y=2.165 $X2=0
+ $Y2=0
cc_380 N_SCE_c_331_n N_A_181_47#_c_2124_n 0.0498114f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_381 N_SCE_c_332_n N_A_181_47#_c_2124_n 0.0251568f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_382 N_SCE_c_333_n N_A_181_47#_c_2124_n 0.0167673f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_383 N_SCE_c_331_n N_A_181_47#_c_2125_n 0.0258668f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_384 N_SCE_c_331_n N_A_181_47#_c_2120_n 0.0188281f $X=2.385 $Y=1.19 $X2=0
+ $Y2=0
cc_385 N_SCE_M1024_g N_VGND_c_2290_n 0.00187853f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_386 N_SCE_c_331_n N_VGND_c_2290_n 0.00450255f $X=2.385 $Y=1.19 $X2=0 $Y2=0
cc_387 N_SCE_M1024_g N_VGND_c_2291_n 0.00959953f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_388 N_SCE_c_333_n N_VGND_c_2291_n 0.00101546f $X=2.53 $Y=1.19 $X2=0 $Y2=0
cc_389 N_SCE_M1016_g N_VGND_c_2299_n 0.005323f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_390 N_SCE_M1024_g N_VGND_c_2305_n 0.0046653f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_391 N_SCE_M1016_g N_VGND_c_2311_n 0.00412734f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_392 N_SCE_c_328_n N_VGND_c_2311_n 3.91104e-19 $X=0.89 $Y=1.415 $X2=0 $Y2=0
cc_393 SCE N_VGND_c_2311_n 0.0111408f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_394 N_SCE_c_352_n N_VGND_c_2311_n 6.88562e-19 $X=0.835 $Y=1.19 $X2=0 $Y2=0
cc_395 N_SCE_M1016_g N_VGND_c_2319_n 0.00728858f $X=0.83 $Y=0.445 $X2=0 $Y2=0
cc_396 N_SCE_M1024_g N_VGND_c_2319_n 0.00934473f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_397 SCE N_VGND_c_2319_n 0.00510613f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_398 N_D_c_433_n N_A_328_21#_M1036_g 0.025603f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_399 D N_A_328_21#_M1036_g 3.06083e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_400 N_D_c_436_n N_A_328_21#_M1036_g 0.0156608f $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_401 N_D_M1004_g N_A_328_21#_M1032_g 0.0356733f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_402 D N_A_328_21#_M1032_g 8.81974e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_403 N_D_M1004_g N_A_328_21#_c_478_n 0.00893563f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_404 D N_A_328_21#_c_478_n 5.01903e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_405 N_D_M1004_g N_A_27_369#_c_1853_n 0.00432785f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_406 D N_A_27_369#_c_1853_n 0.00945908f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_407 N_D_M1004_g N_A_27_369#_c_1867_n 0.00396011f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_408 N_D_M1004_g N_A_27_369#_c_1868_n 0.00152167f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_409 N_D_M1004_g N_A_27_369#_c_1854_n 0.0104505f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_410 D N_A_27_369#_c_1854_n 0.00408716f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_411 N_D_M1004_g N_VPWR_c_1895_n 0.00137466f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_412 N_D_M1004_g N_VPWR_c_1913_n 0.00357863f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_413 N_D_M1004_g N_VPWR_c_1894_n 0.00530374f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_414 N_D_c_433_n N_A_181_47#_c_2116_n 0.0151453f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_415 D N_A_181_47#_c_2116_n 0.0192545f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_416 N_D_c_436_n N_A_181_47#_c_2116_n 0.0013923f $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_417 D N_A_181_47#_c_2125_n 0.00763475f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_418 N_D_c_433_n N_A_181_47#_c_2120_n 9.34382e-19 $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_419 N_D_M1004_g N_A_181_47#_c_2120_n 0.0053499f $X=1.25 $Y=2.165 $X2=0 $Y2=0
cc_420 D N_A_181_47#_c_2120_n 0.0669028f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_421 N_D_c_436_n N_A_181_47#_c_2120_n 0.00210142f $X=1.25 $Y=0.93 $X2=0 $Y2=0
cc_422 N_D_c_433_n N_VGND_c_2299_n 0.00357877f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_423 N_D_c_433_n N_VGND_c_2319_n 0.0053916f $X=1.25 $Y=0.765 $X2=0 $Y2=0
cc_424 N_A_328_21#_c_477_n CLK 0.00445597f $X=2.065 $Y=1.16 $X2=0 $Y2=0
cc_425 N_A_328_21#_c_479_n CLK 0.00862596f $X=2.395 $Y=0.715 $X2=0 $Y2=0
cc_426 N_A_328_21#_c_477_n CLK 0.00431415f $X=2.065 $Y=1.16 $X2=0 $Y2=0
cc_427 N_A_328_21#_c_485_n CLK 0.00668113f $X=2.45 $Y=1.99 $X2=0 $Y2=0
cc_428 N_A_328_21#_c_477_n CLK 0.00126367f $X=2.065 $Y=1.16 $X2=0 $Y2=0
cc_429 N_A_328_21#_c_485_n N_A_27_369#_M1032_d 0.00431967f $X=2.45 $Y=1.99 $X2=0
+ $Y2=0
cc_430 N_A_328_21#_M1032_g N_A_27_369#_c_1867_n 6.173e-19 $X=1.73 $Y=2.165 $X2=0
+ $Y2=0
cc_431 N_A_328_21#_M1032_g N_A_27_369#_c_1854_n 0.0112284f $X=1.73 $Y=2.165
+ $X2=0 $Y2=0
cc_432 N_A_328_21#_c_484_n N_A_27_369#_c_1854_n 0.0180913f $X=2.405 $Y=1.922
+ $X2=0 $Y2=0
cc_433 N_A_328_21#_c_485_n N_A_27_369#_c_1854_n 0.00930147f $X=2.45 $Y=1.99
+ $X2=0 $Y2=0
cc_434 N_A_328_21#_M1032_g N_VPWR_c_1913_n 0.00357877f $X=1.73 $Y=2.165 $X2=0
+ $Y2=0
cc_435 N_A_328_21#_c_484_n N_VPWR_c_1913_n 0.0172798f $X=2.405 $Y=1.922 $X2=0
+ $Y2=0
cc_436 N_A_328_21#_c_485_n N_VPWR_c_1913_n 0.00328493f $X=2.45 $Y=1.99 $X2=0
+ $Y2=0
cc_437 N_A_328_21#_M1029_s N_VPWR_c_1894_n 0.00374699f $X=2.325 $Y=1.845 $X2=0
+ $Y2=0
cc_438 N_A_328_21#_M1032_g N_VPWR_c_1894_n 0.00672549f $X=1.73 $Y=2.165 $X2=0
+ $Y2=0
cc_439 N_A_328_21#_c_484_n N_VPWR_c_1894_n 0.00979174f $X=2.405 $Y=1.922 $X2=0
+ $Y2=0
cc_440 N_A_328_21#_c_485_n N_VPWR_c_1894_n 0.00528232f $X=2.45 $Y=1.99 $X2=0
+ $Y2=0
cc_441 N_A_328_21#_M1036_g N_A_181_47#_c_2116_n 0.0133544f $X=1.715 $Y=0.445
+ $X2=0 $Y2=0
cc_442 N_A_328_21#_c_480_n N_A_181_47#_c_2116_n 0.00519792f $X=2.445 $Y=0.44
+ $X2=0 $Y2=0
cc_443 N_A_328_21#_M1032_g N_A_181_47#_c_2132_n 0.004135f $X=1.73 $Y=2.165 $X2=0
+ $Y2=0
cc_444 N_A_328_21#_c_485_n N_A_181_47#_c_2132_n 0.0130658f $X=2.45 $Y=1.99 $X2=0
+ $Y2=0
cc_445 N_A_328_21#_M1032_g N_A_181_47#_c_2124_n 0.0048301f $X=1.73 $Y=2.165
+ $X2=0 $Y2=0
cc_446 N_A_328_21#_c_477_n N_A_181_47#_c_2124_n 0.01438f $X=2.065 $Y=1.16 $X2=0
+ $Y2=0
cc_447 N_A_328_21#_c_478_n N_A_181_47#_c_2124_n 0.0027371f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_448 N_A_328_21#_c_485_n N_A_181_47#_c_2124_n 0.0130547f $X=2.45 $Y=1.99 $X2=0
+ $Y2=0
cc_449 N_A_328_21#_M1032_g N_A_181_47#_c_2125_n 0.00229183f $X=1.73 $Y=2.165
+ $X2=0 $Y2=0
cc_450 N_A_328_21#_c_477_n N_A_181_47#_c_2125_n 0.00225271f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_451 N_A_328_21#_M1036_g N_A_181_47#_c_2120_n 0.00610463f $X=1.715 $Y=0.445
+ $X2=0 $Y2=0
cc_452 N_A_328_21#_M1032_g N_A_181_47#_c_2120_n 0.011049f $X=1.73 $Y=2.165 $X2=0
+ $Y2=0
cc_453 N_A_328_21#_c_477_n N_A_181_47#_c_2120_n 0.0376443f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_454 N_A_328_21#_c_478_n N_A_181_47#_c_2120_n 0.00961581f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_455 N_A_328_21#_c_479_n N_A_181_47#_c_2120_n 0.00997646f $X=2.395 $Y=0.715
+ $X2=0 $Y2=0
cc_456 N_A_328_21#_c_485_n N_A_181_47#_c_2120_n 0.00456819f $X=2.45 $Y=1.99
+ $X2=0 $Y2=0
cc_457 N_A_328_21#_M1036_g N_VGND_c_2290_n 0.0044954f $X=1.715 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_328_21#_c_478_n N_VGND_c_2290_n 0.00443575f $X=2.065 $Y=1.16 $X2=0
+ $Y2=0
cc_459 N_A_328_21#_c_479_n N_VGND_c_2290_n 0.00851697f $X=2.395 $Y=0.715 $X2=0
+ $Y2=0
cc_460 N_A_328_21#_c_480_n N_VGND_c_2290_n 0.0232895f $X=2.445 $Y=0.44 $X2=0
+ $Y2=0
cc_461 N_A_328_21#_M1036_g N_VGND_c_2299_n 0.00513347f $X=1.715 $Y=0.445 $X2=0
+ $Y2=0
cc_462 N_A_328_21#_c_479_n N_VGND_c_2305_n 0.00268684f $X=2.395 $Y=0.715 $X2=0
+ $Y2=0
cc_463 N_A_328_21#_c_480_n N_VGND_c_2305_n 0.0181977f $X=2.445 $Y=0.44 $X2=0
+ $Y2=0
cc_464 N_A_328_21#_M1024_s N_VGND_c_2319_n 0.00382897f $X=2.32 $Y=0.235 $X2=0
+ $Y2=0
cc_465 N_A_328_21#_M1036_g N_VGND_c_2319_n 0.0101499f $X=1.715 $Y=0.445 $X2=0
+ $Y2=0
cc_466 N_A_328_21#_c_479_n N_VGND_c_2319_n 0.00506824f $X=2.395 $Y=0.715 $X2=0
+ $Y2=0
cc_467 N_A_328_21#_c_480_n N_VGND_c_2319_n 0.0102186f $X=2.445 $Y=0.44 $X2=0
+ $Y2=0
cc_468 N_CLK_c_560_n N_A_652_47#_c_633_n 0.0064798f $X=3.43 $Y=1.09 $X2=0 $Y2=0
cc_469 N_CLK_c_555_n N_A_652_47#_c_634_n 0.0141259f $X=3.595 $Y=0.73 $X2=0 $Y2=0
cc_470 N_CLK_c_561_n N_A_652_47#_c_635_n 0.00752524f $X=3.49 $Y=1.62 $X2=0 $Y2=0
cc_471 N_CLK_c_563_n N_A_652_47#_c_635_n 0.00363391f $X=3.6 $Y=1.695 $X2=0 $Y2=0
cc_472 CLK N_A_652_47#_c_635_n 6.44849e-19 $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_473 N_CLK_c_559_n N_A_652_47#_c_635_n 0.0213743f $X=3.43 $Y=1.255 $X2=0 $Y2=0
cc_474 N_CLK_c_563_n N_A_652_47#_M1031_g 0.0277592f $X=3.6 $Y=1.695 $X2=0 $Y2=0
cc_475 N_CLK_c_556_n N_A_652_47#_c_639_n 0.00827288f $X=3.595 $Y=0.805 $X2=0
+ $Y2=0
cc_476 N_CLK_c_555_n N_A_652_47#_c_640_n 0.00273103f $X=3.595 $Y=0.73 $X2=0
+ $Y2=0
cc_477 N_CLK_c_555_n N_A_652_47#_c_641_n 0.00390827f $X=3.595 $Y=0.73 $X2=0
+ $Y2=0
cc_478 N_CLK_c_556_n N_A_652_47#_c_641_n 0.00649316f $X=3.595 $Y=0.805 $X2=0
+ $Y2=0
cc_479 CLK N_A_652_47#_c_641_n 0.00687961f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_480 N_CLK_c_560_n N_A_652_47#_c_641_n 0.00130904f $X=3.43 $Y=1.09 $X2=0 $Y2=0
cc_481 N_CLK_c_556_n N_A_652_47#_c_642_n 0.00404447f $X=3.595 $Y=0.805 $X2=0
+ $Y2=0
cc_482 CLK N_A_652_47#_c_642_n 0.0136403f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_483 CLK N_A_652_47#_c_642_n 0.0173161f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_484 N_CLK_c_559_n N_A_652_47#_c_642_n 8.54762e-19 $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_485 N_CLK_c_560_n N_A_652_47#_c_642_n 7.77662e-19 $X=3.43 $Y=1.09 $X2=0 $Y2=0
cc_486 N_CLK_c_562_n N_A_652_47#_c_654_n 0.0125884f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_487 N_CLK_c_563_n N_A_652_47#_c_654_n 0.00152901f $X=3.6 $Y=1.695 $X2=0 $Y2=0
cc_488 CLK N_A_652_47#_c_654_n 0.00507511f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_489 N_CLK_c_563_n N_A_652_47#_c_655_n 0.0018976f $X=3.6 $Y=1.695 $X2=0 $Y2=0
cc_490 CLK N_A_652_47#_c_655_n 0.0117145f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_491 CLK N_A_652_47#_c_655_n 0.013475f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_492 N_CLK_c_559_n N_A_652_47#_c_655_n 5.89316e-19 $X=3.43 $Y=1.255 $X2=0
+ $Y2=0
cc_493 N_CLK_c_563_n N_A_652_47#_c_643_n 0.0028039f $X=3.6 $Y=1.695 $X2=0 $Y2=0
cc_494 CLK N_A_652_47#_c_643_n 0.0052596f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_495 CLK N_A_652_47#_c_643_n 0.00664496f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_496 CLK N_A_652_47#_c_643_n 0.0439523f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_497 N_CLK_c_560_n N_A_652_47#_c_643_n 0.00373637f $X=3.43 $Y=1.09 $X2=0 $Y2=0
cc_498 CLK N_VPWR_M1029_d 0.00300367f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_499 N_CLK_c_562_n N_VPWR_c_1896_n 0.00418408f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_500 CLK N_VPWR_c_1896_n 0.0158561f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_501 N_CLK_c_562_n N_VPWR_c_1897_n 0.00802611f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_502 N_CLK_c_562_n N_VPWR_c_1914_n 0.00348948f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_503 N_CLK_c_562_n N_VPWR_c_1894_n 0.00553267f $X=3.6 $Y=1.77 $X2=0 $Y2=0
cc_504 CLK N_VPWR_c_1894_n 7.52808e-19 $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_505 N_CLK_c_561_n N_A_181_47#_c_2124_n 9.84938e-19 $X=3.49 $Y=1.62 $X2=0
+ $Y2=0
cc_506 N_CLK_c_563_n N_A_181_47#_c_2124_n 0.0033491f $X=3.6 $Y=1.695 $X2=0 $Y2=0
cc_507 CLK N_A_181_47#_c_2124_n 5.20642e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_508 CLK N_A_181_47#_c_2124_n 0.00419839f $X=2.905 $Y=1.785 $X2=0 $Y2=0
cc_509 CLK N_A_181_47#_c_2124_n 0.0426481f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_510 N_CLK_c_555_n N_VGND_c_2291_n 0.00218807f $X=3.595 $Y=0.73 $X2=0 $Y2=0
cc_511 CLK N_VGND_c_2291_n 0.0163337f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_512 N_CLK_c_555_n N_VGND_c_2292_n 0.00750008f $X=3.595 $Y=0.73 $X2=0 $Y2=0
cc_513 N_CLK_c_555_n N_VGND_c_2306_n 0.00348405f $X=3.595 $Y=0.73 $X2=0 $Y2=0
cc_514 N_CLK_c_556_n N_VGND_c_2306_n 3.16884e-19 $X=3.595 $Y=0.805 $X2=0 $Y2=0
cc_515 N_CLK_c_555_n N_VGND_c_2319_n 0.00552264f $X=3.595 $Y=0.73 $X2=0 $Y2=0
cc_516 CLK N_VGND_c_2319_n 7.78553e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_517 N_A_652_47#_c_659_n N_A_818_47#_M1031_d 8.60715e-19 $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_518 N_A_652_47#_c_635_n N_A_818_47#_c_933_n 0.00693195f $X=4.02 $Y=1.68 $X2=0
+ $Y2=0
cc_519 N_A_652_47#_c_659_n N_A_818_47#_c_933_n 0.00109756f $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_520 N_A_652_47#_c_662_n N_A_818_47#_c_933_n 0.00337278f $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_521 N_A_652_47#_c_663_n N_A_818_47#_c_933_n 5.29703e-19 $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_522 N_A_652_47#_c_662_n N_A_818_47#_c_921_n 0.00558999f $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_523 N_A_652_47#_c_663_n N_A_818_47#_c_921_n 3.53e-19 $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_524 N_A_652_47#_M1021_g N_A_818_47#_M1043_g 0.0143433f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_525 N_A_652_47#_M1018_g N_A_818_47#_M1043_g 0.0179266f $X=8.99 $Y=0.445 $X2=0
+ $Y2=0
cc_526 N_A_652_47#_c_644_n N_A_818_47#_M1043_g 0.00684887f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_527 N_A_652_47#_c_645_n N_A_818_47#_M1043_g 0.0212722f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_528 N_A_652_47#_c_646_n N_A_818_47#_M1043_g 0.0164384f $X=8.83 $Y=0.795 $X2=0
+ $Y2=0
cc_529 N_A_652_47#_c_648_n N_A_818_47#_M1043_g 0.00171168f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_530 N_A_652_47#_c_649_n N_A_818_47#_M1043_g 0.0119544f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_531 N_A_652_47#_M1021_g N_A_818_47#_c_936_n 0.00430564f $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_532 N_A_652_47#_c_646_n N_A_818_47#_c_936_n 0.00125328f $X=8.83 $Y=0.795
+ $X2=0 $Y2=0
cc_533 N_A_652_47#_c_714_p N_A_818_47#_c_936_n 0.00105592f $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_534 N_A_652_47#_M1021_g N_A_818_47#_M1039_g 0.0125874f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_535 N_A_652_47#_c_714_p N_A_818_47#_M1039_g 0.00109295f $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_536 N_A_652_47#_M1031_g N_A_818_47#_c_938_n 0.00434334f $X=4.02 $Y=2.165
+ $X2=0 $Y2=0
cc_537 N_A_652_47#_M1034_g N_A_818_47#_c_938_n 0.0129984f $X=5.435 $Y=2.275
+ $X2=0 $Y2=0
cc_538 N_A_652_47#_c_659_n N_A_818_47#_c_938_n 0.00543369f $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_539 N_A_652_47#_c_661_n N_A_818_47#_c_938_n 7.44986e-19 $X=5.49 $Y=1.87 $X2=0
+ $Y2=0
cc_540 N_A_652_47#_c_662_n N_A_818_47#_c_938_n 0.00442966f $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_541 N_A_652_47#_c_663_n N_A_818_47#_c_938_n 7.11308e-19 $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_542 N_A_652_47#_c_637_n N_A_818_47#_c_924_n 0.0115863f $X=4.955 $Y=0.73 $X2=0
+ $Y2=0
cc_543 N_A_652_47#_c_636_n N_A_818_47#_c_925_n 0.00974012f $X=4.88 $Y=0.805
+ $X2=0 $Y2=0
cc_544 N_A_652_47#_c_662_n N_A_818_47#_c_925_n 4.68998e-19 $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_545 N_A_652_47#_c_637_n N_A_818_47#_c_973_n 7.9339e-19 $X=4.955 $Y=0.73 $X2=0
+ $Y2=0
cc_546 N_A_652_47#_c_659_n N_A_818_47#_c_939_n 6.29265e-19 $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_547 N_A_652_47#_c_635_n N_A_818_47#_c_940_n 0.00908669f $X=4.02 $Y=1.68 $X2=0
+ $Y2=0
cc_548 N_A_652_47#_c_729_p N_A_818_47#_c_940_n 0.0116011f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_549 N_A_652_47#_c_659_n N_A_818_47#_c_940_n 0.0194461f $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_550 N_A_652_47#_c_731_p N_A_818_47#_c_940_n 0.00243106f $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_551 N_A_652_47#_c_636_n N_A_818_47#_c_926_n 8.56524e-19 $X=4.88 $Y=0.805
+ $X2=0 $Y2=0
cc_552 N_A_652_47#_c_644_n N_A_818_47#_c_926_n 0.0171369f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_553 N_A_652_47#_c_645_n N_A_818_47#_c_926_n 0.00425451f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_554 N_A_652_47#_c_646_n N_A_818_47#_c_926_n 0.0149498f $X=8.83 $Y=0.795 $X2=0
+ $Y2=0
cc_555 N_A_652_47#_c_659_n N_A_818_47#_c_926_n 0.00752192f $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_556 N_A_652_47#_c_660_n N_A_818_47#_c_926_n 0.0448163f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_557 N_A_652_47#_c_661_n N_A_818_47#_c_926_n 0.0123623f $X=5.49 $Y=1.87 $X2=0
+ $Y2=0
cc_558 N_A_652_47#_c_663_n N_A_818_47#_c_926_n 8.48602e-19 $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_559 N_A_652_47#_c_636_n N_A_818_47#_c_927_n 0.00234075f $X=4.88 $Y=0.805
+ $X2=0 $Y2=0
cc_560 N_A_652_47#_c_643_n N_A_818_47#_c_927_n 0.00138833f $X=3.91 $Y=1.255
+ $X2=0 $Y2=0
cc_561 N_A_652_47#_c_635_n N_A_818_47#_c_928_n 0.00372602f $X=4.02 $Y=1.68 $X2=0
+ $Y2=0
cc_562 N_A_652_47#_c_636_n N_A_818_47#_c_928_n 0.00183262f $X=4.88 $Y=0.805
+ $X2=0 $Y2=0
cc_563 N_A_652_47#_c_644_n N_A_818_47#_c_929_n 0.001872f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_564 N_A_652_47#_c_645_n N_A_818_47#_c_929_n 4.40906e-19 $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_565 N_A_652_47#_c_646_n N_A_818_47#_c_929_n 0.00465383f $X=8.83 $Y=0.795
+ $X2=0 $Y2=0
cc_566 N_A_652_47#_c_648_n N_A_818_47#_c_929_n 0.00641513f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_567 N_A_652_47#_c_649_n N_A_818_47#_c_929_n 0.00388112f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_568 N_A_652_47#_M1021_g N_A_818_47#_c_930_n 0.0011294f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_569 N_A_652_47#_c_644_n N_A_818_47#_c_930_n 0.0205397f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_570 N_A_652_47#_c_645_n N_A_818_47#_c_930_n 8.3813e-19 $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_571 N_A_652_47#_c_646_n N_A_818_47#_c_930_n 0.0144401f $X=8.83 $Y=0.795 $X2=0
+ $Y2=0
cc_572 N_A_652_47#_c_648_n N_A_818_47#_c_930_n 0.0114642f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_573 N_A_652_47#_c_649_n N_A_818_47#_c_930_n 0.00126492f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_574 N_A_652_47#_c_714_p N_A_818_47#_c_930_n 0.00966933f $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_575 N_A_652_47#_c_635_n N_A_818_47#_c_931_n 0.0203168f $X=4.02 $Y=1.68 $X2=0
+ $Y2=0
cc_576 N_A_652_47#_c_636_n N_A_818_47#_c_931_n 0.0494337f $X=4.88 $Y=0.805 $X2=0
+ $Y2=0
cc_577 N_A_652_47#_c_643_n N_A_818_47#_c_931_n 3.0071e-19 $X=3.91 $Y=1.255 $X2=0
+ $Y2=0
cc_578 N_A_652_47#_c_633_n N_A_818_47#_c_932_n 0.00372602f $X=3.985 $Y=1.09
+ $X2=0 $Y2=0
cc_579 N_A_652_47#_c_634_n N_A_818_47#_c_932_n 0.00465654f $X=4.015 $Y=0.73
+ $X2=0 $Y2=0
cc_580 N_A_652_47#_c_636_n N_A_818_47#_c_932_n 0.012902f $X=4.88 $Y=0.805 $X2=0
+ $Y2=0
cc_581 N_A_652_47#_c_641_n N_A_818_47#_c_932_n 0.0129402f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_582 N_A_652_47#_c_643_n N_A_818_47#_c_932_n 0.0686518f $X=3.91 $Y=1.255 $X2=0
+ $Y2=0
cc_583 N_A_652_47#_M1034_g N_A_1132_21#_M1044_g 0.026736f $X=5.435 $Y=2.275
+ $X2=0 $Y2=0
cc_584 N_A_652_47#_c_660_n N_A_1132_21#_M1044_g 0.00300937f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_585 N_A_652_47#_c_660_n N_A_1132_21#_c_1123_n 0.0108654f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_586 N_A_652_47#_c_660_n N_A_1132_21#_c_1124_n 0.00397683f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_587 N_A_652_47#_c_662_n N_A_1132_21#_c_1124_n 0.0133445f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_588 N_A_652_47#_c_714_p N_A_1132_21#_c_1125_n 6.25817e-19 $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_589 N_A_652_47#_c_660_n N_A_1132_21#_c_1125_n 0.023552f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_590 N_A_652_47#_c_660_n N_A_1132_21#_c_1126_n 0.00323561f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_591 N_A_652_47#_c_660_n N_A_1006_47#_M1008_g 0.00367443f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_592 N_A_652_47#_M1021_g N_A_1006_47#_M1015_g 0.052059f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_593 N_A_652_47#_c_714_p N_A_1006_47#_M1015_g 0.0121762f $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_594 N_A_652_47#_c_775_p N_A_1006_47#_M1015_g 0.00166615f $X=7.645 $Y=1.87
+ $X2=0 $Y2=0
cc_595 N_A_652_47#_c_637_n N_A_1006_47#_c_1218_n 0.00204386f $X=4.955 $Y=0.73
+ $X2=0 $Y2=0
cc_596 N_A_652_47#_M1034_g N_A_1006_47#_c_1245_n 0.0115873f $X=5.435 $Y=2.275
+ $X2=0 $Y2=0
cc_597 N_A_652_47#_c_659_n N_A_1006_47#_c_1245_n 0.00461962f $X=5.2 $Y=1.87
+ $X2=0 $Y2=0
cc_598 N_A_652_47#_c_660_n N_A_1006_47#_c_1245_n 0.00465741f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_599 N_A_652_47#_c_661_n N_A_1006_47#_c_1245_n 0.00385089f $X=5.49 $Y=1.87
+ $X2=0 $Y2=0
cc_600 N_A_652_47#_c_662_n N_A_1006_47#_c_1245_n 6.03921e-19 $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_601 N_A_652_47#_c_663_n N_A_1006_47#_c_1245_n 0.0143644f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_602 N_A_652_47#_c_660_n N_A_1006_47#_c_1219_n 0.00337041f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_603 N_A_652_47#_c_661_n N_A_1006_47#_c_1219_n 6.59679e-19 $X=5.49 $Y=1.87
+ $X2=0 $Y2=0
cc_604 N_A_652_47#_c_662_n N_A_1006_47#_c_1219_n 0.00216854f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_605 N_A_652_47#_c_663_n N_A_1006_47#_c_1219_n 8.5205e-19 $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_606 N_A_652_47#_c_659_n N_A_1006_47#_c_1220_n 0.00396196f $X=5.2 $Y=1.87
+ $X2=0 $Y2=0
cc_607 N_A_652_47#_c_661_n N_A_1006_47#_c_1220_n 0.00107185f $X=5.49 $Y=1.87
+ $X2=0 $Y2=0
cc_608 N_A_652_47#_c_662_n N_A_1006_47#_c_1220_n 9.08724e-19 $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_609 N_A_652_47#_c_663_n N_A_1006_47#_c_1220_n 0.0174492f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_610 N_A_652_47#_M1034_g N_A_1006_47#_c_1234_n 0.00422822f $X=5.435 $Y=2.275
+ $X2=0 $Y2=0
cc_611 N_A_652_47#_c_660_n N_A_1006_47#_c_1234_n 0.0149262f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_612 N_A_652_47#_c_661_n N_A_1006_47#_c_1234_n 0.00291663f $X=5.49 $Y=1.87
+ $X2=0 $Y2=0
cc_613 N_A_652_47#_c_662_n N_A_1006_47#_c_1234_n 0.00210597f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_614 N_A_652_47#_c_663_n N_A_1006_47#_c_1234_n 0.0264226f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_615 N_A_652_47#_c_660_n N_A_1006_47#_c_1223_n 0.0072615f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_616 N_A_652_47#_c_644_n N_A_1006_47#_c_1225_n 0.0251285f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_617 N_A_652_47#_c_645_n N_A_1006_47#_c_1225_n 0.00191818f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_618 N_A_652_47#_c_714_p N_A_1006_47#_c_1225_n 0.00546057f $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_619 N_A_652_47#_c_644_n N_A_1006_47#_c_1226_n 0.00313024f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_620 N_A_652_47#_c_645_n N_A_1006_47#_c_1226_n 0.052059f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_621 N_A_652_47#_c_714_p N_A_1006_47#_c_1226_n 0.00169347f $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_622 N_A_652_47#_c_660_n N_A_1006_47#_c_1227_n 0.00149088f $X=7.5 $Y=1.87
+ $X2=0 $Y2=0
cc_623 N_A_652_47#_c_644_n N_A_1006_47#_c_1229_n 0.00249477f $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_624 N_A_652_47#_c_647_n N_A_1006_47#_c_1229_n 0.00390485f $X=8.055 $Y=0.795
+ $X2=0 $Y2=0
cc_625 N_A_652_47#_c_660_n N_SET_B_M1033_g 0.00452095f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_626 N_A_652_47#_M1021_g N_SET_B_c_1385_n 0.00162178f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_627 N_A_652_47#_c_644_n N_SET_B_c_1385_n 0.0156963f $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_628 N_A_652_47#_c_645_n N_SET_B_c_1385_n 7.93137e-19 $X=7.97 $Y=1.16 $X2=0
+ $Y2=0
cc_629 N_A_652_47#_c_646_n N_SET_B_c_1385_n 0.00445119f $X=8.83 $Y=0.795 $X2=0
+ $Y2=0
cc_630 N_A_652_47#_c_648_n N_SET_B_c_1385_n 0.0015071f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_631 N_A_652_47#_c_649_n N_SET_B_c_1385_n 8.56178e-19 $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_632 N_A_652_47#_c_714_p N_SET_B_c_1385_n 0.0100297f $X=7.885 $Y=1.83 $X2=0
+ $Y2=0
cc_633 N_A_652_47#_c_660_n N_SET_B_c_1385_n 0.0506964f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_634 N_A_652_47#_c_775_p N_SET_B_c_1385_n 0.0261745f $X=7.645 $Y=1.87 $X2=0
+ $Y2=0
cc_635 N_A_652_47#_c_660_n N_SET_B_c_1386_n 0.0265307f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_636 N_A_652_47#_c_648_n N_SET_B_c_1387_n 0.00580626f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_637 N_A_652_47#_c_714_p N_SET_B_c_1388_n 0.00326884f $X=7.885 $Y=1.83 $X2=0
+ $Y2=0
cc_638 N_A_652_47#_c_660_n N_SET_B_c_1388_n 0.00390363f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_639 N_A_652_47#_c_714_p N_SET_B_c_1389_n 0.00318955f $X=7.885 $Y=1.83 $X2=0
+ $Y2=0
cc_640 N_A_652_47#_c_660_n N_SET_B_c_1389_n 0.00855439f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_641 N_A_652_47#_c_648_n N_SET_B_c_1391_n 0.0141629f $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_642 N_A_652_47#_c_649_n N_SET_B_c_1391_n 5.77505e-19 $X=8.93 $Y=1.1 $X2=0
+ $Y2=0
cc_643 N_A_652_47#_c_649_n N_A_1781_295#_c_1519_n 0.0104254f $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_644 N_A_652_47#_M1018_g N_A_1781_295#_M1020_g 0.0365671f $X=8.99 $Y=0.445
+ $X2=0 $Y2=0
cc_645 N_A_652_47#_c_646_n N_A_1781_295#_M1020_g 0.00205168f $X=8.83 $Y=0.795
+ $X2=0 $Y2=0
cc_646 N_A_652_47#_M1018_g N_A_1781_295#_c_1512_n 3.97377e-19 $X=8.99 $Y=0.445
+ $X2=0 $Y2=0
cc_647 N_A_652_47#_c_646_n N_A_1781_295#_c_1512_n 0.00291473f $X=8.83 $Y=0.795
+ $X2=0 $Y2=0
cc_648 N_A_652_47#_c_648_n N_A_1781_295#_c_1512_n 0.0190455f $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_649 N_A_652_47#_c_648_n N_A_1781_295#_c_1513_n 0.00201993f $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_650 N_A_652_47#_c_649_n N_A_1781_295#_c_1513_n 0.0365671f $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_651 N_A_652_47#_c_648_n N_A_1781_295#_c_1522_n 0.00554642f $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_652 N_A_652_47#_c_646_n N_A_1597_329#_M1043_d 0.00232367f $X=8.83 $Y=0.795
+ $X2=-0.19 $Y2=-0.24
cc_653 N_A_652_47#_c_644_n N_A_1597_329#_M1021_d 7.02761e-19 $X=7.97 $Y=1.16
+ $X2=0 $Y2=0
cc_654 N_A_652_47#_c_714_p N_A_1597_329#_M1021_d 0.0036765f $X=7.885 $Y=1.83
+ $X2=0 $Y2=0
cc_655 N_A_652_47#_M1021_g N_A_1597_329#_c_1644_n 0.00138656f $X=7.91 $Y=2.065
+ $X2=0 $Y2=0
cc_656 N_A_652_47#_M1018_g N_A_1597_329#_c_1645_n 0.012991f $X=8.99 $Y=0.445
+ $X2=0 $Y2=0
cc_657 N_A_652_47#_c_646_n N_A_1597_329#_c_1645_n 0.0365254f $X=8.83 $Y=0.795
+ $X2=0 $Y2=0
cc_658 N_A_652_47#_c_649_n N_A_1597_329#_c_1645_n 3.3555e-19 $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_659 N_A_652_47#_c_646_n N_A_1597_329#_c_1622_n 0.00518737f $X=8.83 $Y=0.795
+ $X2=0 $Y2=0
cc_660 N_A_652_47#_c_646_n N_A_1597_329#_c_1623_n 3.83724e-19 $X=8.83 $Y=0.795
+ $X2=0 $Y2=0
cc_661 N_A_652_47#_c_648_n N_A_1597_329#_c_1639_n 6.22675e-19 $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_662 N_A_652_47#_c_649_n N_A_1597_329#_c_1639_n 5.91567e-19 $X=8.93 $Y=1.1
+ $X2=0 $Y2=0
cc_663 N_A_652_47#_c_729_p N_VPWR_M1010_d 0.00204119f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_664 N_A_652_47#_c_714_p N_VPWR_M1033_d 0.00457308f $X=7.885 $Y=1.83 $X2=0
+ $Y2=0
cc_665 N_A_652_47#_c_660_n N_VPWR_M1033_d 0.00245698f $X=7.5 $Y=1.87 $X2=0 $Y2=0
cc_666 N_A_652_47#_c_665_n N_VPWR_c_1896_n 0.0148242f $X=3.39 $Y=2.16 $X2=0
+ $Y2=0
cc_667 N_A_652_47#_M1031_g N_VPWR_c_1897_n 0.00819473f $X=4.02 $Y=2.165 $X2=0
+ $Y2=0
cc_668 N_A_652_47#_c_654_n N_VPWR_c_1897_n 0.00139915f $X=3.735 $Y=1.915 $X2=0
+ $Y2=0
cc_669 N_A_652_47#_c_729_p N_VPWR_c_1897_n 0.00862024f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_670 N_A_652_47#_c_731_p N_VPWR_c_1897_n 0.00112064f $X=4.055 $Y=1.87 $X2=0
+ $Y2=0
cc_671 N_A_652_47#_c_660_n N_VPWR_c_1898_n 0.00119074f $X=7.5 $Y=1.87 $X2=0
+ $Y2=0
cc_672 N_A_652_47#_c_665_n N_VPWR_c_1914_n 0.00719182f $X=3.39 $Y=2.16 $X2=0
+ $Y2=0
cc_673 N_A_652_47#_c_654_n N_VPWR_c_1914_n 0.0020032f $X=3.735 $Y=1.915 $X2=0
+ $Y2=0
cc_674 N_A_652_47#_M1031_g N_VPWR_c_1915_n 0.00447739f $X=4.02 $Y=2.165 $X2=0
+ $Y2=0
cc_675 N_A_652_47#_M1034_g N_VPWR_c_1915_n 0.00357877f $X=5.435 $Y=2.275 $X2=0
+ $Y2=0
cc_676 N_A_652_47#_c_729_p N_VPWR_c_1915_n 2.83312e-19 $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_677 N_A_652_47#_M1021_g N_VPWR_c_1924_n 0.0199583f $X=7.91 $Y=2.065 $X2=0
+ $Y2=0
cc_678 N_A_652_47#_c_714_p N_VPWR_c_1924_n 0.0317948f $X=7.885 $Y=1.83 $X2=0
+ $Y2=0
cc_679 N_A_652_47#_c_660_n N_VPWR_c_1924_n 0.0126308f $X=7.5 $Y=1.87 $X2=0 $Y2=0
cc_680 N_A_652_47#_c_775_p N_VPWR_c_1924_n 0.00338024f $X=7.645 $Y=1.87 $X2=0
+ $Y2=0
cc_681 N_A_652_47#_M1010_s N_VPWR_c_1894_n 0.0026885f $X=3.265 $Y=1.845 $X2=0
+ $Y2=0
cc_682 N_A_652_47#_M1031_g N_VPWR_c_1894_n 0.00555929f $X=4.02 $Y=2.165 $X2=0
+ $Y2=0
cc_683 N_A_652_47#_M1034_g N_VPWR_c_1894_n 0.00539092f $X=5.435 $Y=2.275 $X2=0
+ $Y2=0
cc_684 N_A_652_47#_c_665_n N_VPWR_c_1894_n 0.00714172f $X=3.39 $Y=2.16 $X2=0
+ $Y2=0
cc_685 N_A_652_47#_c_654_n N_VPWR_c_1894_n 0.00432974f $X=3.735 $Y=1.915 $X2=0
+ $Y2=0
cc_686 N_A_652_47#_c_729_p N_VPWR_c_1894_n 0.00121239f $X=3.865 $Y=1.83 $X2=0
+ $Y2=0
cc_687 N_A_652_47#_c_714_p N_VPWR_c_1894_n 0.00298002f $X=7.885 $Y=1.83 $X2=0
+ $Y2=0
cc_688 N_A_652_47#_c_659_n N_VPWR_c_1894_n 0.0557464f $X=5.2 $Y=1.87 $X2=0 $Y2=0
cc_689 N_A_652_47#_c_731_p N_VPWR_c_1894_n 0.0137798f $X=4.055 $Y=1.87 $X2=0
+ $Y2=0
cc_690 N_A_652_47#_c_660_n N_VPWR_c_1894_n 0.0920009f $X=7.5 $Y=1.87 $X2=0 $Y2=0
cc_691 N_A_652_47#_c_661_n N_VPWR_c_1894_n 0.0156836f $X=5.49 $Y=1.87 $X2=0
+ $Y2=0
cc_692 N_A_652_47#_c_775_p N_VPWR_c_1894_n 0.0143849f $X=7.645 $Y=1.87 $X2=0
+ $Y2=0
cc_693 N_A_652_47#_c_637_n N_A_181_47#_c_2117_n 0.00655099f $X=4.955 $Y=0.73
+ $X2=0 $Y2=0
cc_694 N_A_652_47#_c_659_n N_A_181_47#_c_2121_n 5.67924e-19 $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_695 N_A_652_47#_c_663_n N_A_181_47#_c_2121_n 0.00195457f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_696 N_A_652_47#_M1034_g N_A_181_47#_c_2122_n 8.05795e-19 $X=5.435 $Y=2.275
+ $X2=0 $Y2=0
cc_697 N_A_652_47#_c_659_n N_A_181_47#_c_2122_n 0.0168696f $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_698 N_A_652_47#_c_661_n N_A_181_47#_c_2122_n 0.002781f $X=5.49 $Y=1.87 $X2=0
+ $Y2=0
cc_699 N_A_652_47#_c_662_n N_A_181_47#_c_2122_n 0.00107694f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_700 N_A_652_47#_c_663_n N_A_181_47#_c_2122_n 0.0139595f $X=5.38 $Y=1.74 $X2=0
+ $Y2=0
cc_701 N_A_652_47#_c_636_n N_A_181_47#_c_2119_n 0.017038f $X=4.88 $Y=0.805 $X2=0
+ $Y2=0
cc_702 N_A_652_47#_c_635_n N_A_181_47#_c_2124_n 0.00523679f $X=4.02 $Y=1.68
+ $X2=0 $Y2=0
cc_703 N_A_652_47#_c_639_n N_A_181_47#_c_2124_n 0.00199031f $X=4 $Y=0.805 $X2=0
+ $Y2=0
cc_704 N_A_652_47#_c_641_n N_A_181_47#_c_2124_n 0.00554925f $X=3.735 $Y=0.8
+ $X2=0 $Y2=0
cc_705 N_A_652_47#_c_642_n N_A_181_47#_c_2124_n 7.61163e-19 $X=3.47 $Y=0.8 $X2=0
+ $Y2=0
cc_706 N_A_652_47#_c_654_n N_A_181_47#_c_2124_n 0.00747114f $X=3.735 $Y=1.915
+ $X2=0 $Y2=0
cc_707 N_A_652_47#_c_655_n N_A_181_47#_c_2124_n 0.00164507f $X=3.475 $Y=1.915
+ $X2=0 $Y2=0
cc_708 N_A_652_47#_c_643_n N_A_181_47#_c_2124_n 0.022041f $X=3.91 $Y=1.255 $X2=0
+ $Y2=0
cc_709 N_A_652_47#_c_659_n N_A_181_47#_c_2124_n 0.0535603f $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_710 N_A_652_47#_c_731_p N_A_181_47#_c_2124_n 0.0254302f $X=4.055 $Y=1.87
+ $X2=0 $Y2=0
cc_711 N_A_652_47#_c_659_n N_A_181_47#_c_2127_n 0.026422f $X=5.2 $Y=1.87 $X2=0
+ $Y2=0
cc_712 N_A_652_47#_c_663_n N_A_181_47#_c_2127_n 0.00223839f $X=5.38 $Y=1.74
+ $X2=0 $Y2=0
cc_713 N_A_652_47#_c_714_p A_1525_329# 0.00170472f $X=7.885 $Y=1.83 $X2=-0.19
+ $Y2=-0.24
cc_714 N_A_652_47#_c_775_p A_1525_329# 0.00159132f $X=7.645 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_715 N_A_652_47#_c_640_n N_VGND_c_2291_n 0.0240223f $X=3.385 $Y=0.44 $X2=0
+ $Y2=0
cc_716 N_A_652_47#_c_634_n N_VGND_c_2292_n 0.00309854f $X=4.015 $Y=0.73 $X2=0
+ $Y2=0
cc_717 N_A_652_47#_c_635_n N_VGND_c_2292_n 4.44358e-19 $X=4.02 $Y=1.68 $X2=0
+ $Y2=0
cc_718 N_A_652_47#_c_641_n N_VGND_c_2292_n 0.0201015f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_719 N_A_652_47#_M1018_g N_VGND_c_2301_n 0.00362032f $X=8.99 $Y=0.445 $X2=0
+ $Y2=0
cc_720 N_A_652_47#_c_646_n N_VGND_c_2301_n 0.00579644f $X=8.83 $Y=0.795 $X2=0
+ $Y2=0
cc_721 N_A_652_47#_c_647_n N_VGND_c_2301_n 0.00289816f $X=8.055 $Y=0.795 $X2=0
+ $Y2=0
cc_722 N_A_652_47#_c_640_n N_VGND_c_2306_n 0.0136391f $X=3.385 $Y=0.44 $X2=0
+ $Y2=0
cc_723 N_A_652_47#_c_641_n N_VGND_c_2306_n 0.00240298f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_724 N_A_652_47#_c_634_n N_VGND_c_2307_n 0.00529955f $X=4.015 $Y=0.73 $X2=0
+ $Y2=0
cc_725 N_A_652_47#_c_636_n N_VGND_c_2307_n 0.00382472f $X=4.88 $Y=0.805 $X2=0
+ $Y2=0
cc_726 N_A_652_47#_c_637_n N_VGND_c_2307_n 0.00579312f $X=4.955 $Y=0.73 $X2=0
+ $Y2=0
cc_727 N_A_652_47#_c_641_n N_VGND_c_2307_n 8.20832e-19 $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_728 N_A_652_47#_c_647_n N_VGND_c_2316_n 0.00941377f $X=8.055 $Y=0.795 $X2=0
+ $Y2=0
cc_729 N_A_652_47#_M1003_s N_VGND_c_2319_n 0.00271619f $X=3.26 $Y=0.235 $X2=0
+ $Y2=0
cc_730 N_A_652_47#_c_634_n N_VGND_c_2319_n 0.0100522f $X=4.015 $Y=0.73 $X2=0
+ $Y2=0
cc_731 N_A_652_47#_c_636_n N_VGND_c_2319_n 0.00371212f $X=4.88 $Y=0.805 $X2=0
+ $Y2=0
cc_732 N_A_652_47#_c_637_n N_VGND_c_2319_n 0.011875f $X=4.955 $Y=0.73 $X2=0
+ $Y2=0
cc_733 N_A_652_47#_M1018_g N_VGND_c_2319_n 0.00555751f $X=8.99 $Y=0.445 $X2=0
+ $Y2=0
cc_734 N_A_652_47#_c_640_n N_VGND_c_2319_n 0.00761007f $X=3.385 $Y=0.44 $X2=0
+ $Y2=0
cc_735 N_A_652_47#_c_641_n N_VGND_c_2319_n 0.00648481f $X=3.735 $Y=0.8 $X2=0
+ $Y2=0
cc_736 N_A_652_47#_c_646_n N_VGND_c_2319_n 0.0110862f $X=8.83 $Y=0.795 $X2=0
+ $Y2=0
cc_737 N_A_652_47#_c_647_n N_VGND_c_2319_n 0.00489372f $X=8.055 $Y=0.795 $X2=0
+ $Y2=0
cc_738 N_A_652_47#_c_646_n A_1517_47# 0.00430463f $X=8.83 $Y=0.795 $X2=-0.19
+ $Y2=-0.24
cc_739 N_A_652_47#_c_647_n A_1517_47# 0.00654797f $X=8.055 $Y=0.795 $X2=-0.19
+ $Y2=-0.24
cc_740 N_A_818_47#_c_921_n N_A_1132_21#_c_1115_n 0.00415828f $X=5.24 $Y=1.165
+ $X2=0 $Y2=0
cc_741 N_A_818_47#_c_926_n N_A_1132_21#_c_1115_n 0.00268968f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_742 N_A_818_47#_c_926_n N_A_1132_21#_c_1123_n 5.84337e-19 $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_743 N_A_818_47#_c_926_n N_A_1132_21#_c_1116_n 0.00817983f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_744 N_A_818_47#_c_922_n N_A_1132_21#_c_1118_n 4.89802e-19 $X=5.32 $Y=1.09
+ $X2=0 $Y2=0
cc_745 N_A_818_47#_c_924_n N_A_1132_21#_c_1118_n 0.0011462f $X=5.345 $Y=0.73
+ $X2=0 $Y2=0
cc_746 N_A_818_47#_c_926_n N_A_1132_21#_c_1118_n 0.0104686f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_747 N_A_818_47#_c_922_n N_A_1132_21#_c_1119_n 0.0114272f $X=5.32 $Y=1.09
+ $X2=0 $Y2=0
cc_748 N_A_818_47#_c_925_n N_A_1132_21#_c_1119_n 0.0226044f $X=5.345 $Y=0.86
+ $X2=0 $Y2=0
cc_749 N_A_818_47#_c_926_n N_A_1132_21#_c_1119_n 0.0045534f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_750 N_A_818_47#_c_924_n N_A_1132_21#_c_1120_n 0.0226044f $X=5.345 $Y=0.73
+ $X2=0 $Y2=0
cc_751 N_A_818_47#_c_921_n N_A_1006_47#_c_1218_n 0.0108945f $X=5.24 $Y=1.165
+ $X2=0 $Y2=0
cc_752 N_A_818_47#_c_922_n N_A_1006_47#_c_1218_n 0.00826036f $X=5.32 $Y=1.09
+ $X2=0 $Y2=0
cc_753 N_A_818_47#_c_924_n N_A_1006_47#_c_1218_n 0.0126947f $X=5.345 $Y=0.73
+ $X2=0 $Y2=0
cc_754 N_A_818_47#_c_925_n N_A_1006_47#_c_1218_n 0.00625103f $X=5.345 $Y=0.86
+ $X2=0 $Y2=0
cc_755 N_A_818_47#_c_926_n N_A_1006_47#_c_1218_n 0.0288745f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_756 N_A_818_47#_c_926_n N_A_1006_47#_c_1219_n 0.00841601f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_757 N_A_818_47#_c_921_n N_A_1006_47#_c_1220_n 0.00525632f $X=5.24 $Y=1.165
+ $X2=0 $Y2=0
cc_758 N_A_818_47#_c_926_n N_A_1006_47#_c_1220_n 0.00857227f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_759 N_A_818_47#_c_931_n N_A_1006_47#_c_1220_n 3.67371e-19 $X=4.745 $Y=1.255
+ $X2=0 $Y2=0
cc_760 N_A_818_47#_c_926_n N_A_1006_47#_c_1221_n 0.00653615f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_761 N_A_818_47#_c_926_n N_A_1006_47#_c_1222_n 0.00137673f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_762 N_A_818_47#_c_926_n N_A_1006_47#_c_1223_n 0.0157171f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_763 N_A_818_47#_c_926_n N_A_1006_47#_c_1224_n 0.0111406f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_764 N_A_818_47#_c_926_n N_A_1006_47#_c_1225_n 0.0144608f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_765 N_A_818_47#_c_926_n N_A_1006_47#_c_1227_n 0.0332696f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_766 N_A_818_47#_M1043_g N_SET_B_c_1385_n 0.00169335f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_767 N_A_818_47#_c_936_n N_SET_B_c_1385_n 0.00258644f $X=8.54 $Y=1.905 $X2=0
+ $Y2=0
cc_768 N_A_818_47#_c_926_n N_SET_B_c_1385_n 0.12203f $X=8.42 $Y=1.19 $X2=0 $Y2=0
cc_769 N_A_818_47#_c_929_n N_SET_B_c_1385_n 0.0255536f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_770 N_A_818_47#_c_930_n N_SET_B_c_1385_n 0.0148271f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_771 N_A_818_47#_c_926_n N_SET_B_c_1386_n 0.0264445f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_772 N_A_818_47#_c_930_n N_SET_B_c_1387_n 0.00148131f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_773 N_A_818_47#_c_926_n N_SET_B_c_1389_n 9.31754e-19 $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_774 N_A_818_47#_M1043_g N_SET_B_c_1391_n 3.56571e-19 $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_775 N_A_818_47#_c_936_n N_SET_B_c_1391_n 9.30315e-19 $X=8.54 $Y=1.905 $X2=0
+ $Y2=0
cc_776 N_A_818_47#_c_930_n N_SET_B_c_1391_n 0.0159952f $X=8.565 $Y=1.19 $X2=0
+ $Y2=0
cc_777 N_A_818_47#_M1039_g N_A_1781_295#_M1009_g 0.0304162f $X=8.54 $Y=2.275
+ $X2=0 $Y2=0
cc_778 N_A_818_47#_c_930_n N_A_1781_295#_M1009_g 0.0010368f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_779 N_A_818_47#_M1043_g N_A_1781_295#_c_1519_n 0.00238821f $X=8.39 $Y=0.555
+ $X2=0 $Y2=0
cc_780 N_A_818_47#_c_936_n N_A_1781_295#_c_1519_n 0.0209749f $X=8.54 $Y=1.905
+ $X2=0 $Y2=0
cc_781 N_A_818_47#_c_930_n N_A_1781_295#_c_1519_n 4.7495e-19 $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_782 N_A_818_47#_c_929_n N_A_1781_295#_c_1511_n 7.56349e-19 $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_783 N_A_818_47#_c_930_n N_A_1781_295#_c_1511_n 0.00303247f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_784 N_A_818_47#_c_929_n N_A_1781_295#_c_1522_n 0.00104583f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_785 N_A_818_47#_c_930_n N_A_1781_295#_c_1522_n 0.00211352f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_786 N_A_818_47#_c_936_n N_A_1597_329#_c_1644_n 0.00480909f $X=8.54 $Y=1.905
+ $X2=0 $Y2=0
cc_787 N_A_818_47#_M1039_g N_A_1597_329#_c_1644_n 0.0113397f $X=8.54 $Y=2.275
+ $X2=0 $Y2=0
cc_788 N_A_818_47#_c_930_n N_A_1597_329#_c_1644_n 0.0110537f $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_789 N_A_818_47#_M1039_g N_A_1597_329#_c_1639_n 0.00469548f $X=8.54 $Y=2.275
+ $X2=0 $Y2=0
cc_790 N_A_818_47#_c_930_n N_A_1597_329#_c_1639_n 7.3132e-19 $X=8.565 $Y=1.19
+ $X2=0 $Y2=0
cc_791 N_A_818_47#_M1039_g N_VPWR_c_1906_n 0.00358923f $X=8.54 $Y=2.275 $X2=0
+ $Y2=0
cc_792 N_A_818_47#_c_934_n N_VPWR_c_1915_n 0.00579312f $X=4.96 $Y=1.99 $X2=0
+ $Y2=0
cc_793 N_A_818_47#_c_938_n N_VPWR_c_1915_n 0.00197896f $X=4.96 $Y=1.915 $X2=0
+ $Y2=0
cc_794 N_A_818_47#_c_939_n N_VPWR_c_1915_n 0.0204643f $X=4.23 $Y=2.3 $X2=0 $Y2=0
cc_795 N_A_818_47#_M1039_g N_VPWR_c_1924_n 0.00159206f $X=8.54 $Y=2.275 $X2=0
+ $Y2=0
cc_796 N_A_818_47#_M1031_d N_VPWR_c_1894_n 0.0021132f $X=4.095 $Y=1.845 $X2=0
+ $Y2=0
cc_797 N_A_818_47#_c_934_n N_VPWR_c_1894_n 0.00777633f $X=4.96 $Y=1.99 $X2=0
+ $Y2=0
cc_798 N_A_818_47#_M1039_g N_VPWR_c_1894_n 0.0057638f $X=8.54 $Y=2.275 $X2=0
+ $Y2=0
cc_799 N_A_818_47#_c_938_n N_VPWR_c_1894_n 0.00127223f $X=4.96 $Y=1.915 $X2=0
+ $Y2=0
cc_800 N_A_818_47#_c_939_n N_VPWR_c_1894_n 0.00536207f $X=4.23 $Y=2.3 $X2=0
+ $Y2=0
cc_801 N_A_818_47#_c_973_n N_A_181_47#_c_2117_n 0.0260149f $X=4.225 $Y=0.42
+ $X2=0 $Y2=0
cc_802 N_A_818_47#_c_933_n N_A_181_47#_c_2121_n 0.00565936f $X=4.67 $Y=1.84
+ $X2=0 $Y2=0
cc_803 N_A_818_47#_c_921_n N_A_181_47#_c_2121_n 0.0015014f $X=5.24 $Y=1.165
+ $X2=0 $Y2=0
cc_804 N_A_818_47#_c_938_n N_A_181_47#_c_2121_n 0.00142271f $X=4.96 $Y=1.915
+ $X2=0 $Y2=0
cc_805 N_A_818_47#_c_940_n N_A_181_47#_c_2121_n 0.00740664f $X=4.292 $Y=2.135
+ $X2=0 $Y2=0
cc_806 N_A_818_47#_c_926_n N_A_181_47#_c_2121_n 9.25945e-19 $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_807 N_A_818_47#_c_933_n N_A_181_47#_c_2122_n 0.00481946f $X=4.67 $Y=1.84
+ $X2=0 $Y2=0
cc_808 N_A_818_47#_c_934_n N_A_181_47#_c_2122_n 0.00744813f $X=4.96 $Y=1.99
+ $X2=0 $Y2=0
cc_809 N_A_818_47#_c_938_n N_A_181_47#_c_2122_n 0.0128233f $X=4.96 $Y=1.915
+ $X2=0 $Y2=0
cc_810 N_A_818_47#_c_940_n N_A_181_47#_c_2122_n 0.0517431f $X=4.292 $Y=2.135
+ $X2=0 $Y2=0
cc_811 N_A_818_47#_c_933_n N_A_181_47#_c_2118_n 7.0296e-19 $X=4.67 $Y=1.84 $X2=0
+ $Y2=0
cc_812 N_A_818_47#_c_921_n N_A_181_47#_c_2118_n 0.00723713f $X=5.24 $Y=1.165
+ $X2=0 $Y2=0
cc_813 N_A_818_47#_c_940_n N_A_181_47#_c_2118_n 0.00102314f $X=4.292 $Y=2.135
+ $X2=0 $Y2=0
cc_814 N_A_818_47#_c_926_n N_A_181_47#_c_2118_n 0.0123859f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_815 N_A_818_47#_c_927_n N_A_181_47#_c_2118_n 0.00226234f $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_816 N_A_818_47#_c_928_n N_A_181_47#_c_2118_n 0.0164614f $X=4.37 $Y=1.19 $X2=0
+ $Y2=0
cc_817 N_A_818_47#_c_931_n N_A_181_47#_c_2118_n 0.00697892f $X=4.745 $Y=1.255
+ $X2=0 $Y2=0
cc_818 N_A_818_47#_c_932_n N_A_181_47#_c_2118_n 0.00706773f $X=4.327 $Y=1.09
+ $X2=0 $Y2=0
cc_819 N_A_818_47#_c_922_n N_A_181_47#_c_2119_n 9.74224e-19 $X=5.32 $Y=1.09
+ $X2=0 $Y2=0
cc_820 N_A_818_47#_c_926_n N_A_181_47#_c_2119_n 0.00856991f $X=8.42 $Y=1.19
+ $X2=0 $Y2=0
cc_821 N_A_818_47#_c_927_n N_A_181_47#_c_2119_n 5.00901e-19 $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_822 N_A_818_47#_c_931_n N_A_181_47#_c_2119_n 0.00497404f $X=4.745 $Y=1.255
+ $X2=0 $Y2=0
cc_823 N_A_818_47#_c_932_n N_A_181_47#_c_2119_n 0.0260149f $X=4.327 $Y=1.09
+ $X2=0 $Y2=0
cc_824 N_A_818_47#_c_933_n N_A_181_47#_c_2124_n 0.00307322f $X=4.67 $Y=1.84
+ $X2=0 $Y2=0
cc_825 N_A_818_47#_c_940_n N_A_181_47#_c_2124_n 0.0166962f $X=4.292 $Y=2.135
+ $X2=0 $Y2=0
cc_826 N_A_818_47#_c_926_n N_A_181_47#_c_2124_n 0.0181259f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_827 N_A_818_47#_c_927_n N_A_181_47#_c_2124_n 0.0254082f $X=4.515 $Y=1.19
+ $X2=0 $Y2=0
cc_828 N_A_818_47#_c_928_n N_A_181_47#_c_2124_n 0.0014472f $X=4.37 $Y=1.19 $X2=0
+ $Y2=0
cc_829 N_A_818_47#_c_931_n N_A_181_47#_c_2124_n 0.00175281f $X=4.745 $Y=1.255
+ $X2=0 $Y2=0
cc_830 N_A_818_47#_c_921_n N_A_181_47#_c_2127_n 4.09059e-19 $X=5.24 $Y=1.165
+ $X2=0 $Y2=0
cc_831 N_A_818_47#_c_938_n N_A_181_47#_c_2127_n 3.99374e-19 $X=4.96 $Y=1.915
+ $X2=0 $Y2=0
cc_832 N_A_818_47#_c_940_n N_A_181_47#_c_2127_n 5.63414e-19 $X=4.292 $Y=2.135
+ $X2=0 $Y2=0
cc_833 N_A_818_47#_c_926_n N_A_181_47#_c_2127_n 0.0264737f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_834 N_A_818_47#_M1043_g N_VGND_c_2301_n 0.00433717f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_835 N_A_818_47#_c_924_n N_VGND_c_2307_n 0.00359186f $X=5.345 $Y=0.73 $X2=0
+ $Y2=0
cc_836 N_A_818_47#_c_973_n N_VGND_c_2307_n 0.0143635f $X=4.225 $Y=0.42 $X2=0
+ $Y2=0
cc_837 N_A_818_47#_c_924_n N_VGND_c_2314_n 0.0022254f $X=5.345 $Y=0.73 $X2=0
+ $Y2=0
cc_838 N_A_818_47#_M1043_g N_VGND_c_2316_n 0.0140829f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_839 N_A_818_47#_c_926_n N_VGND_c_2316_n 0.00591877f $X=8.42 $Y=1.19 $X2=0
+ $Y2=0
cc_840 N_A_818_47#_M1045_d N_VGND_c_2319_n 0.0029715f $X=4.09 $Y=0.235 $X2=0
+ $Y2=0
cc_841 N_A_818_47#_M1043_g N_VGND_c_2319_n 0.00776391f $X=8.39 $Y=0.555 $X2=0
+ $Y2=0
cc_842 N_A_818_47#_c_924_n N_VGND_c_2319_n 0.00510857f $X=5.345 $Y=0.73 $X2=0
+ $Y2=0
cc_843 N_A_818_47#_c_973_n N_VGND_c_2319_n 0.0085511f $X=4.225 $Y=0.42 $X2=0
+ $Y2=0
cc_844 N_A_1132_21#_c_1115_n N_A_1006_47#_M1008_g 0.00519515f $X=5.885 $Y=1.575
+ $X2=0 $Y2=0
cc_845 N_A_1132_21#_M1044_g N_A_1006_47#_M1008_g 0.0159634f $X=5.885 $Y=2.275
+ $X2=0 $Y2=0
cc_846 N_A_1132_21#_c_1123_n N_A_1006_47#_M1008_g 0.00225299f $X=6.06 $Y=1.74
+ $X2=0 $Y2=0
cc_847 N_A_1132_21#_c_1124_n N_A_1006_47#_M1008_g 0.0213433f $X=6.06 $Y=1.74
+ $X2=0 $Y2=0
cc_848 N_A_1132_21#_c_1125_n N_A_1006_47#_M1008_g 0.0128904f $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_849 N_A_1132_21#_c_1116_n N_A_1006_47#_c_1216_n 0.00169518f $X=6.335 $Y=0.72
+ $X2=0 $Y2=0
cc_850 N_A_1132_21#_c_1116_n N_A_1006_47#_c_1217_n 0.00843421f $X=6.335 $Y=0.72
+ $X2=0 $Y2=0
cc_851 N_A_1132_21#_c_1118_n N_A_1006_47#_c_1217_n 0.0035496f $X=5.817 $Y=0.72
+ $X2=0 $Y2=0
cc_852 N_A_1132_21#_c_1119_n N_A_1006_47#_c_1217_n 0.00757926f $X=5.795 $Y=0.93
+ $X2=0 $Y2=0
cc_853 N_A_1132_21#_c_1120_n N_A_1006_47#_c_1217_n 4.77792e-19 $X=5.81 $Y=0.765
+ $X2=0 $Y2=0
cc_854 N_A_1132_21#_c_1115_n N_A_1006_47#_c_1218_n 0.00187677f $X=5.885 $Y=1.575
+ $X2=0 $Y2=0
cc_855 N_A_1132_21#_c_1118_n N_A_1006_47#_c_1218_n 0.0306216f $X=5.817 $Y=0.72
+ $X2=0 $Y2=0
cc_856 N_A_1132_21#_c_1119_n N_A_1006_47#_c_1218_n 0.00238433f $X=5.795 $Y=0.93
+ $X2=0 $Y2=0
cc_857 N_A_1132_21#_c_1120_n N_A_1006_47#_c_1218_n 0.00202497f $X=5.81 $Y=0.765
+ $X2=0 $Y2=0
cc_858 N_A_1132_21#_c_1118_n N_A_1006_47#_c_1219_n 7.44766e-19 $X=5.817 $Y=0.72
+ $X2=0 $Y2=0
cc_859 N_A_1132_21#_c_1115_n N_A_1006_47#_c_1234_n 0.0117953f $X=5.885 $Y=1.575
+ $X2=0 $Y2=0
cc_860 N_A_1132_21#_c_1123_n N_A_1006_47#_c_1234_n 0.0251678f $X=6.06 $Y=1.74
+ $X2=0 $Y2=0
cc_861 N_A_1132_21#_c_1126_n N_A_1006_47#_c_1234_n 0.0106732f $X=6.145 $Y=2.02
+ $X2=0 $Y2=0
cc_862 N_A_1132_21#_c_1118_n N_A_1006_47#_c_1221_n 0.00921157f $X=5.817 $Y=0.72
+ $X2=0 $Y2=0
cc_863 N_A_1132_21#_c_1119_n N_A_1006_47#_c_1221_n 0.00406544f $X=5.795 $Y=0.93
+ $X2=0 $Y2=0
cc_864 N_A_1132_21#_c_1115_n N_A_1006_47#_c_1222_n 0.0137286f $X=5.885 $Y=1.575
+ $X2=0 $Y2=0
cc_865 N_A_1132_21#_c_1116_n N_A_1006_47#_c_1222_n 0.00223241f $X=6.335 $Y=0.72
+ $X2=0 $Y2=0
cc_866 N_A_1132_21#_c_1125_n N_A_1006_47#_c_1222_n 6.97279e-19 $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_867 N_A_1132_21#_c_1115_n N_A_1006_47#_c_1223_n 0.0126813f $X=5.885 $Y=1.575
+ $X2=0 $Y2=0
cc_868 N_A_1132_21#_c_1123_n N_A_1006_47#_c_1223_n 0.0109804f $X=6.06 $Y=1.74
+ $X2=0 $Y2=0
cc_869 N_A_1132_21#_c_1124_n N_A_1006_47#_c_1223_n 0.00309725f $X=6.06 $Y=1.74
+ $X2=0 $Y2=0
cc_870 N_A_1132_21#_c_1116_n N_A_1006_47#_c_1223_n 0.00704107f $X=6.335 $Y=0.72
+ $X2=0 $Y2=0
cc_871 N_A_1132_21#_c_1125_n N_A_1006_47#_c_1223_n 0.00602228f $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_872 N_A_1132_21#_c_1118_n N_A_1006_47#_c_1223_n 0.0105929f $X=5.817 $Y=0.72
+ $X2=0 $Y2=0
cc_873 N_A_1132_21#_c_1115_n N_A_1006_47#_c_1224_n 0.00108886f $X=5.885 $Y=1.575
+ $X2=0 $Y2=0
cc_874 N_A_1132_21#_c_1116_n N_A_1006_47#_c_1224_n 0.0186643f $X=6.335 $Y=0.72
+ $X2=0 $Y2=0
cc_875 N_A_1132_21#_c_1118_n N_A_1006_47#_c_1224_n 0.00240735f $X=5.817 $Y=0.72
+ $X2=0 $Y2=0
cc_876 N_A_1132_21#_c_1119_n N_A_1006_47#_c_1224_n 0.0021169f $X=5.795 $Y=0.93
+ $X2=0 $Y2=0
cc_877 N_A_1132_21#_c_1125_n N_A_1006_47#_c_1227_n 0.00198283f $X=6.605 $Y=2.02
+ $X2=0 $Y2=0
cc_878 N_A_1132_21#_c_1125_n N_SET_B_M1033_g 0.00497375f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_879 N_A_1132_21#_c_1123_n N_SET_B_c_1386_n 0.00174961f $X=6.06 $Y=1.74 $X2=0
+ $Y2=0
cc_880 N_A_1132_21#_c_1125_n N_SET_B_c_1386_n 3.32046e-19 $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_881 N_A_1132_21#_c_1125_n N_SET_B_c_1388_n 0.00107555f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_882 N_A_1132_21#_c_1123_n N_SET_B_c_1389_n 0.00551177f $X=6.06 $Y=1.74 $X2=0
+ $Y2=0
cc_883 N_A_1132_21#_c_1125_n N_SET_B_c_1389_n 0.0122653f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_884 N_A_1132_21#_c_1125_n N_VPWR_M1044_d 0.00225394f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_885 N_A_1132_21#_c_1126_n N_VPWR_M1044_d 0.0014782f $X=6.145 $Y=2.02 $X2=0
+ $Y2=0
cc_886 N_A_1132_21#_M1044_g N_VPWR_c_1898_n 0.00453186f $X=5.885 $Y=2.275 $X2=0
+ $Y2=0
cc_887 N_A_1132_21#_c_1124_n N_VPWR_c_1898_n 7.72184e-19 $X=6.06 $Y=1.74 $X2=0
+ $Y2=0
cc_888 N_A_1132_21#_c_1125_n N_VPWR_c_1898_n 0.0129414f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_889 N_A_1132_21#_c_1126_n N_VPWR_c_1898_n 0.00985859f $X=6.145 $Y=2.02 $X2=0
+ $Y2=0
cc_890 N_A_1132_21#_M1044_g N_VPWR_c_1915_n 0.00585385f $X=5.885 $Y=2.275 $X2=0
+ $Y2=0
cc_891 N_A_1132_21#_c_1125_n N_VPWR_c_1923_n 0.00398868f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_892 N_A_1132_21#_c_1194_p N_VPWR_c_1923_n 0.0132089f $X=6.715 $Y=2.285 $X2=0
+ $Y2=0
cc_893 N_A_1132_21#_M1008_d N_VPWR_c_1894_n 0.00275725f $X=6.555 $Y=2.065 $X2=0
+ $Y2=0
cc_894 N_A_1132_21#_M1044_g N_VPWR_c_1894_n 0.00680616f $X=5.885 $Y=2.275 $X2=0
+ $Y2=0
cc_895 N_A_1132_21#_c_1125_n N_VPWR_c_1894_n 0.00360571f $X=6.605 $Y=2.02 $X2=0
+ $Y2=0
cc_896 N_A_1132_21#_c_1126_n N_VPWR_c_1894_n 8.36043e-19 $X=6.145 $Y=2.02 $X2=0
+ $Y2=0
cc_897 N_A_1132_21#_c_1194_p N_VPWR_c_1894_n 0.00381852f $X=6.715 $Y=2.285 $X2=0
+ $Y2=0
cc_898 N_A_1132_21#_c_1116_n N_VGND_M1022_d 6.08904e-19 $X=6.335 $Y=0.72 $X2=0
+ $Y2=0
cc_899 N_A_1132_21#_c_1118_n N_VGND_M1022_d 0.00158965f $X=5.817 $Y=0.72 $X2=0
+ $Y2=0
cc_900 N_A_1132_21#_c_1118_n N_VGND_c_2307_n 4.68982e-19 $X=5.817 $Y=0.72 $X2=0
+ $Y2=0
cc_901 N_A_1132_21#_c_1116_n N_VGND_c_2314_n 0.0116402f $X=6.335 $Y=0.72 $X2=0
+ $Y2=0
cc_902 N_A_1132_21#_c_1117_n N_VGND_c_2314_n 0.0175033f $X=6.465 $Y=0.51 $X2=0
+ $Y2=0
cc_903 N_A_1132_21#_c_1118_n N_VGND_c_2314_n 0.0227777f $X=5.817 $Y=0.72 $X2=0
+ $Y2=0
cc_904 N_A_1132_21#_c_1119_n N_VGND_c_2314_n 7.06418e-19 $X=5.795 $Y=0.93 $X2=0
+ $Y2=0
cc_905 N_A_1132_21#_c_1120_n N_VGND_c_2314_n 0.0158202f $X=5.81 $Y=0.765 $X2=0
+ $Y2=0
cc_906 N_A_1132_21#_c_1116_n N_VGND_c_2315_n 0.00309842f $X=6.335 $Y=0.72 $X2=0
+ $Y2=0
cc_907 N_A_1132_21#_c_1117_n N_VGND_c_2315_n 0.0145511f $X=6.465 $Y=0.51 $X2=0
+ $Y2=0
cc_908 N_A_1132_21#_c_1116_n N_VGND_c_2316_n 0.0134722f $X=6.335 $Y=0.72 $X2=0
+ $Y2=0
cc_909 N_A_1132_21#_M1002_s N_VGND_c_2319_n 0.00268769f $X=6.34 $Y=0.235 $X2=0
+ $Y2=0
cc_910 N_A_1132_21#_c_1116_n N_VGND_c_2319_n 0.00551338f $X=6.335 $Y=0.72 $X2=0
+ $Y2=0
cc_911 N_A_1132_21#_c_1117_n N_VGND_c_2319_n 0.008158f $X=6.465 $Y=0.51 $X2=0
+ $Y2=0
cc_912 N_A_1132_21#_c_1118_n N_VGND_c_2319_n 0.00290347f $X=5.817 $Y=0.72 $X2=0
+ $Y2=0
cc_913 N_A_1132_21#_c_1120_n N_VGND_c_2319_n 8.07363e-19 $X=5.81 $Y=0.765 $X2=0
+ $Y2=0
cc_914 N_A_1006_47#_M1008_g N_SET_B_M1033_g 0.0138848f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_915 N_A_1006_47#_c_1216_n N_SET_B_M1037_g 0.0503265f $X=6.675 $Y=0.73 $X2=0
+ $Y2=0
cc_916 N_A_1006_47#_c_1226_n N_SET_B_M1037_g 0.0213561f $X=7.455 $Y=1.16 $X2=0
+ $Y2=0
cc_917 N_A_1006_47#_c_1227_n N_SET_B_M1037_g 0.0113502f $X=7.355 $Y=1.15 $X2=0
+ $Y2=0
cc_918 N_A_1006_47#_c_1228_n N_SET_B_M1037_g 0.00994643f $X=6.39 $Y=1.095 $X2=0
+ $Y2=0
cc_919 N_A_1006_47#_c_1229_n N_SET_B_M1037_g 0.0223839f $X=7.472 $Y=0.995 $X2=0
+ $Y2=0
cc_920 N_A_1006_47#_M1015_g N_SET_B_c_1376_n 0.00162366f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_921 N_A_1006_47#_c_1222_n N_SET_B_c_1376_n 0.00546402f $X=6.39 $Y=1.23 $X2=0
+ $Y2=0
cc_922 N_A_1006_47#_c_1224_n N_SET_B_c_1376_n 6.21737e-19 $X=6.475 $Y=1.185
+ $X2=0 $Y2=0
cc_923 N_A_1006_47#_c_1225_n N_SET_B_c_1376_n 3.0927e-19 $X=7.455 $Y=1.16 $X2=0
+ $Y2=0
cc_924 N_A_1006_47#_c_1227_n N_SET_B_c_1376_n 0.00659956f $X=7.355 $Y=1.15 $X2=0
+ $Y2=0
cc_925 N_A_1006_47#_M1015_g N_SET_B_c_1385_n 0.00455115f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_926 N_A_1006_47#_c_1225_n N_SET_B_c_1385_n 0.00394848f $X=7.455 $Y=1.16 $X2=0
+ $Y2=0
cc_927 N_A_1006_47#_c_1226_n N_SET_B_c_1385_n 0.00256245f $X=7.455 $Y=1.16 $X2=0
+ $Y2=0
cc_928 N_A_1006_47#_c_1227_n N_SET_B_c_1385_n 0.00862879f $X=7.355 $Y=1.15 $X2=0
+ $Y2=0
cc_929 N_A_1006_47#_M1008_g N_SET_B_c_1386_n 0.00451637f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_930 N_A_1006_47#_c_1227_n N_SET_B_c_1386_n 0.00232629f $X=7.355 $Y=1.15 $X2=0
+ $Y2=0
cc_931 N_A_1006_47#_M1008_g N_SET_B_c_1388_n 0.0201171f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_932 N_A_1006_47#_c_1227_n N_SET_B_c_1388_n 7.95701e-19 $X=7.355 $Y=1.15 $X2=0
+ $Y2=0
cc_933 N_A_1006_47#_M1008_g N_SET_B_c_1389_n 0.00478519f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_934 N_A_1006_47#_M1015_g N_SET_B_c_1389_n 0.00429264f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_935 N_A_1006_47#_c_1227_n N_SET_B_c_1389_n 0.0278918f $X=7.355 $Y=1.15 $X2=0
+ $Y2=0
cc_936 N_A_1006_47#_M1008_g N_SET_B_c_1390_n 0.00546402f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_937 N_A_1006_47#_M1015_g N_SET_B_c_1390_n 0.0293548f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_938 N_A_1006_47#_M1008_g N_VPWR_c_1898_n 0.00579022f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_939 N_A_1006_47#_c_1245_n N_VPWR_c_1915_n 0.0433516f $X=5.635 $Y=2.3 $X2=0
+ $Y2=0
cc_940 N_A_1006_47#_M1008_g N_VPWR_c_1923_n 0.00422112f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_941 N_A_1006_47#_M1015_g N_VPWR_c_1924_n 0.0234385f $X=7.55 $Y=2.065 $X2=0
+ $Y2=0
cc_942 N_A_1006_47#_M1007_d N_VPWR_c_1894_n 0.00228352f $X=5.035 $Y=2.065 $X2=0
+ $Y2=0
cc_943 N_A_1006_47#_M1008_g N_VPWR_c_1894_n 0.00611683f $X=6.48 $Y=2.275 $X2=0
+ $Y2=0
cc_944 N_A_1006_47#_c_1245_n N_VPWR_c_1894_n 0.0126591f $X=5.635 $Y=2.3 $X2=0
+ $Y2=0
cc_945 N_A_1006_47#_c_1218_n N_A_181_47#_c_2117_n 0.0594178f $X=5.165 $Y=0.42
+ $X2=0 $Y2=0
cc_946 N_A_1006_47#_c_1234_n N_A_181_47#_c_2121_n 0.0019891f $X=5.72 $Y=2.135
+ $X2=0 $Y2=0
cc_947 N_A_1006_47#_c_1220_n N_A_181_47#_c_2118_n 0.0112919f $X=5.45 $Y=1.31
+ $X2=0 $Y2=0
cc_948 N_A_1006_47#_c_1234_n N_A_181_47#_c_2127_n 0.00425696f $X=5.72 $Y=2.135
+ $X2=0 $Y2=0
cc_949 N_A_1006_47#_c_1245_n A_1102_413# 0.00390174f $X=5.635 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_950 N_A_1006_47#_c_1234_n A_1102_413# 0.00101971f $X=5.72 $Y=2.135 $X2=-0.19
+ $Y2=-0.24
cc_951 N_A_1006_47#_c_1218_n N_VGND_c_2307_n 0.0242185f $X=5.165 $Y=0.42 $X2=0
+ $Y2=0
cc_952 N_A_1006_47#_c_1216_n N_VGND_c_2314_n 0.00215107f $X=6.675 $Y=0.73 $X2=0
+ $Y2=0
cc_953 N_A_1006_47#_c_1218_n N_VGND_c_2314_n 0.0136716f $X=5.165 $Y=0.42 $X2=0
+ $Y2=0
cc_954 N_A_1006_47#_c_1216_n N_VGND_c_2315_n 0.0046653f $X=6.675 $Y=0.73 $X2=0
+ $Y2=0
cc_955 N_A_1006_47#_c_1217_n N_VGND_c_2315_n 0.00117078f $X=6.675 $Y=0.805 $X2=0
+ $Y2=0
cc_956 N_A_1006_47#_c_1216_n N_VGND_c_2316_n 0.0135898f $X=6.675 $Y=0.73 $X2=0
+ $Y2=0
cc_957 N_A_1006_47#_c_1217_n N_VGND_c_2316_n 0.00215986f $X=6.675 $Y=0.805 $X2=0
+ $Y2=0
cc_958 N_A_1006_47#_c_1226_n N_VGND_c_2316_n 7.09791e-19 $X=7.455 $Y=1.16 $X2=0
+ $Y2=0
cc_959 N_A_1006_47#_c_1227_n N_VGND_c_2316_n 0.072947f $X=7.355 $Y=1.15 $X2=0
+ $Y2=0
cc_960 N_A_1006_47#_c_1229_n N_VGND_c_2316_n 0.0313595f $X=7.472 $Y=0.995 $X2=0
+ $Y2=0
cc_961 N_A_1006_47#_M1030_d N_VGND_c_2319_n 0.0030199f $X=5.03 $Y=0.235 $X2=0
+ $Y2=0
cc_962 N_A_1006_47#_c_1216_n N_VGND_c_2319_n 0.00929621f $X=6.675 $Y=0.73 $X2=0
+ $Y2=0
cc_963 N_A_1006_47#_c_1217_n N_VGND_c_2319_n 0.00111946f $X=6.675 $Y=0.805 $X2=0
+ $Y2=0
cc_964 N_A_1006_47#_c_1218_n N_VGND_c_2319_n 0.0143813f $X=5.165 $Y=0.42 $X2=0
+ $Y2=0
cc_965 N_SET_B_c_1381_n N_A_1781_295#_M1009_g 0.0170808f $X=9.78 $Y=1.835 $X2=0
+ $Y2=0
cc_966 N_SET_B_c_1384_n N_A_1781_295#_M1009_g 0.00446321f $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_967 N_SET_B_c_1391_n N_A_1781_295#_M1009_g 0.00552373f $X=9.115 $Y=1.58 $X2=0
+ $Y2=0
cc_968 N_SET_B_c_1382_n N_A_1781_295#_c_1518_n 0.0101264f $X=9.78 $Y=1.62 $X2=0
+ $Y2=0
cc_969 N_SET_B_c_1383_n N_A_1781_295#_c_1518_n 0.0160423f $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_970 N_SET_B_c_1387_n N_A_1781_295#_c_1518_n 0.00146845f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_971 N_SET_B_c_1391_n N_A_1781_295#_c_1518_n 0.00363216f $X=9.115 $Y=1.58
+ $X2=0 $Y2=0
cc_972 N_SET_B_c_1391_n N_A_1781_295#_c_1519_n 0.00327833f $X=9.115 $Y=1.58
+ $X2=0 $Y2=0
cc_973 N_SET_B_M1014_g N_A_1781_295#_M1020_g 0.0250034f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_974 N_SET_B_M1014_g N_A_1781_295#_c_1511_n 0.0104404f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_975 N_SET_B_c_1387_n N_A_1781_295#_c_1511_n 0.00154091f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_976 N_SET_B_c_1391_n N_A_1781_295#_c_1511_n 0.00121518f $X=9.115 $Y=1.58
+ $X2=0 $Y2=0
cc_977 N_SET_B_M1014_g N_A_1781_295#_c_1512_n 0.00116147f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_978 N_SET_B_M1014_g N_A_1781_295#_c_1513_n 0.020675f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_979 N_SET_B_c_1381_n N_A_1781_295#_c_1513_n 0.00119817f $X=9.78 $Y=1.835
+ $X2=0 $Y2=0
cc_980 N_SET_B_c_1383_n N_A_1781_295#_c_1513_n 3.13661e-19 $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_981 N_SET_B_M1014_g N_A_1781_295#_c_1514_n 0.0110789f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_982 N_SET_B_c_1382_n N_A_1781_295#_c_1514_n 0.00364149f $X=9.78 $Y=1.62 $X2=0
+ $Y2=0
cc_983 N_SET_B_c_1383_n N_A_1781_295#_c_1514_n 0.0303022f $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_984 N_SET_B_c_1383_n N_A_1781_295#_c_1522_n 0.0180161f $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_985 N_SET_B_M1014_g N_A_1597_329#_c_1613_n 0.0223093f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_986 N_SET_B_c_1382_n N_A_1597_329#_c_1614_n 0.0223093f $X=9.78 $Y=1.62 $X2=0
+ $Y2=0
cc_987 N_SET_B_c_1384_n N_A_1597_329#_M1026_g 0.0032976f $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_988 N_SET_B_c_1385_n N_A_1597_329#_c_1644_n 0.0145657f $X=8.88 $Y=1.53 $X2=0
+ $Y2=0
cc_989 N_SET_B_M1014_g N_A_1597_329#_c_1645_n 0.00751876f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_990 N_SET_B_c_1378_n N_A_1597_329#_c_1634_n 0.00739124f $X=9.535 $Y=1.985
+ $X2=0 $Y2=0
cc_991 N_SET_B_c_1381_n N_A_1597_329#_c_1634_n 0.00533673f $X=9.78 $Y=1.835
+ $X2=0 $Y2=0
cc_992 N_SET_B_c_1387_n N_A_1597_329#_c_1634_n 0.00108108f $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_993 N_SET_B_c_1391_n N_A_1597_329#_c_1634_n 0.0488989f $X=9.115 $Y=1.58 $X2=0
+ $Y2=0
cc_994 N_SET_B_M1014_g N_A_1597_329#_c_1622_n 0.00943202f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_995 N_SET_B_M1014_g N_A_1597_329#_c_1623_n 0.00316304f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_996 N_SET_B_M1014_g N_A_1597_329#_c_1624_n 0.00597361f $X=9.85 $Y=0.445 $X2=0
+ $Y2=0
cc_997 N_SET_B_c_1383_n N_A_1597_329#_c_1636_n 3.43563e-19 $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_998 N_SET_B_c_1382_n N_A_1597_329#_c_1637_n 6.42775e-19 $X=9.78 $Y=1.62 $X2=0
+ $Y2=0
cc_999 N_SET_B_c_1383_n N_A_1597_329#_c_1637_n 0.0174901f $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_1000 N_SET_B_c_1384_n N_A_1597_329#_c_1637_n 0.00413664f $X=9.77 $Y=1.64
+ $X2=0 $Y2=0
cc_1001 N_SET_B_c_1382_n N_A_1597_329#_c_1638_n 0.0172113f $X=9.78 $Y=1.62 $X2=0
+ $Y2=0
cc_1002 N_SET_B_c_1383_n N_A_1597_329#_c_1638_n 5.95759e-19 $X=9.77 $Y=1.64
+ $X2=0 $Y2=0
cc_1003 N_SET_B_c_1378_n N_A_1597_329#_c_1639_n 4.13646e-19 $X=9.535 $Y=1.985
+ $X2=0 $Y2=0
cc_1004 N_SET_B_c_1385_n N_A_1597_329#_c_1639_n 0.00185617f $X=8.88 $Y=1.53
+ $X2=0 $Y2=0
cc_1005 N_SET_B_c_1387_n N_A_1597_329#_c_1639_n 7.07036e-19 $X=9.025 $Y=1.53
+ $X2=0 $Y2=0
cc_1006 N_SET_B_c_1391_n N_A_1597_329#_c_1639_n 0.00798957f $X=9.115 $Y=1.58
+ $X2=0 $Y2=0
cc_1007 N_SET_B_c_1381_n N_A_1597_329#_c_1679_n 0.0134625f $X=9.78 $Y=1.835
+ $X2=0 $Y2=0
cc_1008 N_SET_B_c_1383_n N_A_1597_329#_c_1679_n 0.0204978f $X=9.77 $Y=1.64 $X2=0
+ $Y2=0
cc_1009 N_SET_B_c_1378_n N_VPWR_c_1899_n 0.00758954f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1010 N_SET_B_c_1378_n N_VPWR_c_1900_n 0.00181984f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1011 N_SET_B_c_1378_n N_VPWR_c_1908_n 0.00341689f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1012 N_SET_B_c_1381_n N_VPWR_c_1908_n 7.95779e-19 $X=9.78 $Y=1.835 $X2=0
+ $Y2=0
cc_1013 N_SET_B_M1033_g N_VPWR_c_1923_n 0.00585385f $X=6.97 $Y=2.275 $X2=0 $Y2=0
cc_1014 N_SET_B_M1033_g N_VPWR_c_1924_n 0.00385005f $X=6.97 $Y=2.275 $X2=0 $Y2=0
cc_1015 N_SET_B_c_1385_n N_VPWR_c_1924_n 0.00126181f $X=8.88 $Y=1.53 $X2=0 $Y2=0
cc_1016 N_SET_B_M1033_g N_VPWR_c_1894_n 0.00672875f $X=6.97 $Y=2.275 $X2=0 $Y2=0
cc_1017 N_SET_B_c_1378_n N_VPWR_c_1894_n 0.00538978f $X=9.535 $Y=1.985 $X2=0
+ $Y2=0
cc_1018 N_SET_B_c_1388_n N_VPWR_c_1894_n 4.0446e-19 $X=6.9 $Y=1.68 $X2=0 $Y2=0
cc_1019 N_SET_B_M1014_g N_VGND_c_2293_n 0.00409726f $X=9.85 $Y=0.445 $X2=0 $Y2=0
cc_1020 N_SET_B_M1014_g N_VGND_c_2301_n 0.00466154f $X=9.85 $Y=0.445 $X2=0 $Y2=0
cc_1021 N_SET_B_M1037_g N_VGND_c_2316_n 0.0259455f $X=7.035 $Y=0.445 $X2=0 $Y2=0
cc_1022 N_SET_B_c_1376_n N_VGND_c_2316_n 2.97882e-19 $X=7.002 $Y=1.365 $X2=0
+ $Y2=0
cc_1023 N_SET_B_M1014_g N_VGND_c_2319_n 0.00614767f $X=9.85 $Y=0.445 $X2=0 $Y2=0
cc_1024 N_A_1781_295#_c_1515_n N_A_1597_329#_c_1613_n 0.00484049f $X=10.82
+ $Y=1.185 $X2=0 $Y2=0
cc_1025 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1614_n 0.00968539f $X=10.6
+ $Y=1.27 $X2=0 $Y2=0
cc_1026 N_A_1781_295#_c_1515_n N_A_1597_329#_c_1614_n 0.00386519f $X=10.82
+ $Y=1.185 $X2=0 $Y2=0
cc_1027 N_A_1781_295#_c_1516_n N_A_1597_329#_c_1614_n 0.00178633f $X=10.82
+ $Y=0.42 $X2=0 $Y2=0
cc_1028 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1615_n 0.00179299f $X=10.6
+ $Y=1.27 $X2=0 $Y2=0
cc_1029 N_A_1781_295#_c_1515_n N_A_1597_329#_c_1615_n 0.0193219f $X=10.82
+ $Y=1.185 $X2=0 $Y2=0
cc_1030 N_A_1781_295#_c_1516_n N_A_1597_329#_c_1615_n 0.00284737f $X=10.82
+ $Y=0.42 $X2=0 $Y2=0
cc_1031 N_A_1781_295#_c_1524_n N_A_1597_329#_c_1615_n 0.0167159f $X=10.755
+ $Y=1.27 $X2=0 $Y2=0
cc_1032 N_A_1781_295#_c_1515_n N_A_1597_329#_c_1616_n 0.00232817f $X=10.82
+ $Y=1.185 $X2=0 $Y2=0
cc_1033 N_A_1781_295#_c_1523_n N_A_1597_329#_M1012_g 0.00382912f $X=10.685
+ $Y=2.285 $X2=0 $Y2=0
cc_1034 N_A_1781_295#_c_1524_n N_A_1597_329#_M1012_g 5.3403e-19 $X=10.755
+ $Y=1.27 $X2=0 $Y2=0
cc_1035 N_A_1781_295#_M1009_g N_A_1597_329#_c_1644_n 5.40489e-19 $X=8.98
+ $Y=2.275 $X2=0 $Y2=0
cc_1036 N_A_1781_295#_M1020_g N_A_1597_329#_c_1645_n 0.0135566f $X=9.35 $Y=0.445
+ $X2=0 $Y2=0
cc_1037 N_A_1781_295#_c_1512_n N_A_1597_329#_c_1645_n 0.00772659f $X=9.43
+ $Y=1.02 $X2=0 $Y2=0
cc_1038 N_A_1781_295#_c_1513_n N_A_1597_329#_c_1645_n 0.00154099f $X=9.43
+ $Y=1.02 $X2=0 $Y2=0
cc_1039 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1645_n 0.00472301f $X=10.6
+ $Y=1.27 $X2=0 $Y2=0
cc_1040 N_A_1781_295#_M1009_g N_A_1597_329#_c_1634_n 0.00649005f $X=8.98
+ $Y=2.275 $X2=0 $Y2=0
cc_1041 N_A_1781_295#_c_1518_n N_A_1597_329#_c_1634_n 0.00202703f $X=9.275
+ $Y=1.55 $X2=0 $Y2=0
cc_1042 N_A_1781_295#_M1020_g N_A_1597_329#_c_1622_n 0.00477677f $X=9.35
+ $Y=0.445 $X2=0 $Y2=0
cc_1043 N_A_1781_295#_c_1512_n N_A_1597_329#_c_1623_n 0.0131676f $X=9.43 $Y=1.02
+ $X2=0 $Y2=0
cc_1044 N_A_1781_295#_c_1513_n N_A_1597_329#_c_1623_n 0.00106925f $X=9.43
+ $Y=1.02 $X2=0 $Y2=0
cc_1045 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1623_n 0.0136954f $X=10.6 $Y=1.27
+ $X2=0 $Y2=0
cc_1046 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1624_n 0.0502028f $X=10.6 $Y=1.27
+ $X2=0 $Y2=0
cc_1047 N_A_1781_295#_c_1515_n N_A_1597_329#_c_1624_n 0.0140849f $X=10.82
+ $Y=1.185 $X2=0 $Y2=0
cc_1048 N_A_1781_295#_c_1516_n N_A_1597_329#_c_1624_n 0.00480877f $X=10.82
+ $Y=0.42 $X2=0 $Y2=0
cc_1049 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1636_n 0.00572977f $X=10.6
+ $Y=1.27 $X2=0 $Y2=0
cc_1050 N_A_1781_295#_c_1523_n N_A_1597_329#_c_1636_n 0.0139105f $X=10.685
+ $Y=2.285 $X2=0 $Y2=0
cc_1051 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1637_n 0.0253887f $X=10.6 $Y=1.27
+ $X2=0 $Y2=0
cc_1052 N_A_1781_295#_c_1523_n N_A_1597_329#_c_1637_n 0.0284538f $X=10.685
+ $Y=2.285 $X2=0 $Y2=0
cc_1053 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1638_n 8.12073e-19 $X=10.6
+ $Y=1.27 $X2=0 $Y2=0
cc_1054 N_A_1781_295#_M1009_g N_A_1597_329#_c_1639_n 0.014405f $X=8.98 $Y=2.275
+ $X2=0 $Y2=0
cc_1055 N_A_1781_295#_c_1514_n N_A_1597_329#_c_1640_n 0.00939164f $X=10.6
+ $Y=1.27 $X2=0 $Y2=0
cc_1056 N_A_1781_295#_c_1523_n N_A_1597_329#_c_1640_n 0.0213766f $X=10.685
+ $Y=2.285 $X2=0 $Y2=0
cc_1057 N_A_1781_295#_M1009_g N_VPWR_c_1899_n 0.00520032f $X=8.98 $Y=2.275 $X2=0
+ $Y2=0
cc_1058 N_A_1781_295#_c_1523_n N_VPWR_c_1901_n 0.0600397f $X=10.685 $Y=2.285
+ $X2=0 $Y2=0
cc_1059 N_A_1781_295#_M1009_g N_VPWR_c_1906_n 0.00390259f $X=8.98 $Y=2.275 $X2=0
+ $Y2=0
cc_1060 N_A_1781_295#_c_1523_n N_VPWR_c_1910_n 0.0169256f $X=10.685 $Y=2.285
+ $X2=0 $Y2=0
cc_1061 N_A_1781_295#_M1026_d N_VPWR_c_1894_n 0.00382897f $X=10.55 $Y=2.065
+ $X2=0 $Y2=0
cc_1062 N_A_1781_295#_M1009_g N_VPWR_c_1894_n 0.00595646f $X=8.98 $Y=2.275 $X2=0
+ $Y2=0
cc_1063 N_A_1781_295#_c_1523_n N_VPWR_c_1894_n 0.00935836f $X=10.685 $Y=2.285
+ $X2=0 $Y2=0
cc_1064 N_A_1781_295#_c_1523_n N_Q_N_c_2249_n 0.00382073f $X=10.685 $Y=2.285
+ $X2=0 $Y2=0
cc_1065 N_A_1781_295#_c_1515_n N_Q_N_c_2249_n 0.00870919f $X=10.82 $Y=1.185
+ $X2=0 $Y2=0
cc_1066 N_A_1781_295#_c_1524_n N_Q_N_c_2249_n 0.00534895f $X=10.755 $Y=1.27
+ $X2=0 $Y2=0
cc_1067 N_A_1781_295#_c_1515_n N_VGND_c_2294_n 0.0191429f $X=10.82 $Y=1.185
+ $X2=0 $Y2=0
cc_1068 N_A_1781_295#_c_1516_n N_VGND_c_2294_n 0.0225931f $X=10.82 $Y=0.42 $X2=0
+ $Y2=0
cc_1069 N_A_1781_295#_M1020_g N_VGND_c_2301_n 0.00362032f $X=9.35 $Y=0.445 $X2=0
+ $Y2=0
cc_1070 N_A_1781_295#_c_1516_n N_VGND_c_2303_n 0.0297315f $X=10.82 $Y=0.42 $X2=0
+ $Y2=0
cc_1071 N_A_1781_295#_M1000_d N_VGND_c_2319_n 0.0024997f $X=10.41 $Y=0.235 $X2=0
+ $Y2=0
cc_1072 N_A_1781_295#_M1020_g N_VGND_c_2319_n 0.00535444f $X=9.35 $Y=0.445 $X2=0
+ $Y2=0
cc_1073 N_A_1781_295#_c_1516_n N_VGND_c_2319_n 0.0168122f $X=10.82 $Y=0.42 $X2=0
+ $Y2=0
cc_1074 N_A_1597_329#_M1011_g N_A_2501_47#_c_1793_n 0.0202173f $X=12.84 $Y=0.445
+ $X2=0 $Y2=0
cc_1075 N_A_1597_329#_M1005_g N_A_2501_47#_M1006_g 0.0219329f $X=12.84 $Y=2.1
+ $X2=0 $Y2=0
cc_1076 N_A_1597_329#_c_1617_n N_A_2501_47#_c_1795_n 0.00231059f $X=11.835
+ $Y=0.995 $X2=0 $Y2=0
cc_1077 N_A_1597_329#_M1011_g N_A_2501_47#_c_1795_n 0.0108047f $X=12.84 $Y=0.445
+ $X2=0 $Y2=0
cc_1078 N_A_1597_329#_M1028_g N_A_2501_47#_c_1800_n 0.00344615f $X=11.835
+ $Y=1.985 $X2=0 $Y2=0
cc_1079 N_A_1597_329#_M1005_g N_A_2501_47#_c_1800_n 0.0163772f $X=12.84 $Y=2.1
+ $X2=0 $Y2=0
cc_1080 N_A_1597_329#_c_1618_n N_A_2501_47#_c_1796_n 0.00606691f $X=12.765
+ $Y=1.16 $X2=0 $Y2=0
cc_1081 N_A_1597_329#_c_1621_n N_A_2501_47#_c_1796_n 0.0201727f $X=12.84 $Y=1.16
+ $X2=0 $Y2=0
cc_1082 N_A_1597_329#_c_1618_n N_A_2501_47#_c_1811_n 0.0230864f $X=12.765
+ $Y=1.16 $X2=0 $Y2=0
cc_1083 N_A_1597_329#_c_1621_n N_A_2501_47#_c_1797_n 0.0216153f $X=12.84 $Y=1.16
+ $X2=0 $Y2=0
cc_1084 N_A_1597_329#_c_1636_n N_VPWR_M1026_s 0.00275838f $X=10.105 $Y=1.98
+ $X2=0 $Y2=0
cc_1085 N_A_1597_329#_c_1634_n N_VPWR_c_1899_n 0.022845f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1086 N_A_1597_329#_c_1639_n N_VPWR_c_1899_n 0.0166484f $X=8.905 $Y=1.98 $X2=0
+ $Y2=0
cc_1087 N_A_1597_329#_M1026_g N_VPWR_c_1900_n 0.00843927f $X=10.475 $Y=2.275
+ $X2=0 $Y2=0
cc_1088 N_A_1597_329#_c_1635_n N_VPWR_c_1900_n 0.0176349f $X=9.745 $Y=2.285
+ $X2=0 $Y2=0
cc_1089 N_A_1597_329#_c_1636_n N_VPWR_c_1900_n 0.0244506f $X=10.105 $Y=1.98
+ $X2=0 $Y2=0
cc_1090 N_A_1597_329#_c_1638_n N_VPWR_c_1900_n 0.00108855f $X=10.3 $Y=1.69 $X2=0
+ $Y2=0
cc_1091 N_A_1597_329#_M1026_g N_VPWR_c_1901_n 0.0029163f $X=10.475 $Y=2.275
+ $X2=0 $Y2=0
cc_1092 N_A_1597_329#_c_1615_n N_VPWR_c_1901_n 0.00563428f $X=11.34 $Y=1.16
+ $X2=0 $Y2=0
cc_1093 N_A_1597_329#_M1012_g N_VPWR_c_1901_n 0.00444548f $X=11.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1094 N_A_1597_329#_M1028_g N_VPWR_c_1902_n 0.0250461f $X=11.835 $Y=1.985
+ $X2=0 $Y2=0
cc_1095 N_A_1597_329#_c_1618_n N_VPWR_c_1902_n 0.00856698f $X=12.765 $Y=1.16
+ $X2=0 $Y2=0
cc_1096 N_A_1597_329#_M1005_g N_VPWR_c_1902_n 0.0035148f $X=12.84 $Y=2.1 $X2=0
+ $Y2=0
cc_1097 N_A_1597_329#_M1005_g N_VPWR_c_1903_n 0.0164475f $X=12.84 $Y=2.1 $X2=0
+ $Y2=0
cc_1098 N_A_1597_329#_c_1644_n N_VPWR_c_1906_n 0.0371085f $X=8.82 $Y=2.292 $X2=0
+ $Y2=0
cc_1099 N_A_1597_329#_c_1634_n N_VPWR_c_1906_n 0.00284657f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1100 N_A_1597_329#_c_1639_n N_VPWR_c_1906_n 0.00925064f $X=8.905 $Y=1.98
+ $X2=0 $Y2=0
cc_1101 N_A_1597_329#_c_1634_n N_VPWR_c_1908_n 0.00273399f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1102 N_A_1597_329#_c_1635_n N_VPWR_c_1908_n 0.0168316f $X=9.745 $Y=2.285
+ $X2=0 $Y2=0
cc_1103 N_A_1597_329#_c_1636_n N_VPWR_c_1908_n 0.00296166f $X=10.105 $Y=1.98
+ $X2=0 $Y2=0
cc_1104 N_A_1597_329#_M1026_g N_VPWR_c_1910_n 0.0046653f $X=10.475 $Y=2.275
+ $X2=0 $Y2=0
cc_1105 N_A_1597_329#_M1012_g N_VPWR_c_1916_n 0.00541359f $X=11.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1106 N_A_1597_329#_M1028_g N_VPWR_c_1916_n 0.00442682f $X=11.835 $Y=1.985
+ $X2=0 $Y2=0
cc_1107 N_A_1597_329#_M1005_g N_VPWR_c_1917_n 0.0046653f $X=12.84 $Y=2.1 $X2=0
+ $Y2=0
cc_1108 N_A_1597_329#_M1021_d N_VPWR_c_1894_n 0.00832535f $X=7.985 $Y=1.645
+ $X2=0 $Y2=0
cc_1109 N_A_1597_329#_M1013_d N_VPWR_c_1894_n 0.00228252f $X=9.61 $Y=2.065 $X2=0
+ $Y2=0
cc_1110 N_A_1597_329#_M1026_g N_VPWR_c_1894_n 0.00929867f $X=10.475 $Y=2.275
+ $X2=0 $Y2=0
cc_1111 N_A_1597_329#_M1012_g N_VPWR_c_1894_n 0.0108276f $X=11.415 $Y=1.985
+ $X2=0 $Y2=0
cc_1112 N_A_1597_329#_M1028_g N_VPWR_c_1894_n 0.00867323f $X=11.835 $Y=1.985
+ $X2=0 $Y2=0
cc_1113 N_A_1597_329#_M1005_g N_VPWR_c_1894_n 0.00934473f $X=12.84 $Y=2.1 $X2=0
+ $Y2=0
cc_1114 N_A_1597_329#_c_1644_n N_VPWR_c_1894_n 0.0231897f $X=8.82 $Y=2.292 $X2=0
+ $Y2=0
cc_1115 N_A_1597_329#_c_1634_n N_VPWR_c_1894_n 0.00998273f $X=9.66 $Y=1.98 $X2=0
+ $Y2=0
cc_1116 N_A_1597_329#_c_1635_n N_VPWR_c_1894_n 0.0101906f $X=9.745 $Y=2.285
+ $X2=0 $Y2=0
cc_1117 N_A_1597_329#_c_1636_n N_VPWR_c_1894_n 0.00630672f $X=10.105 $Y=1.98
+ $X2=0 $Y2=0
cc_1118 N_A_1597_329#_c_1639_n N_VPWR_c_1894_n 0.00603799f $X=8.905 $Y=1.98
+ $X2=0 $Y2=0
cc_1119 N_A_1597_329#_c_1644_n A_1723_413# 0.00493444f $X=8.82 $Y=2.292
+ $X2=-0.19 $Y2=-0.24
cc_1120 N_A_1597_329#_c_1639_n A_1723_413# 0.00180472f $X=8.905 $Y=1.98
+ $X2=-0.19 $Y2=-0.24
cc_1121 N_A_1597_329#_c_1616_n N_Q_N_c_2249_n 0.0106186f $X=11.415 $Y=0.995
+ $X2=0 $Y2=0
cc_1122 N_A_1597_329#_M1012_g N_Q_N_c_2249_n 0.016255f $X=11.415 $Y=1.985 $X2=0
+ $Y2=0
cc_1123 N_A_1597_329#_c_1617_n N_Q_N_c_2249_n 0.0146644f $X=11.835 $Y=0.995
+ $X2=0 $Y2=0
cc_1124 N_A_1597_329#_M1028_g N_Q_N_c_2249_n 0.0219643f $X=11.835 $Y=1.985 $X2=0
+ $Y2=0
cc_1125 N_A_1597_329#_c_1619_n N_Q_N_c_2249_n 0.0355255f $X=11.91 $Y=1.16 $X2=0
+ $Y2=0
cc_1126 N_A_1597_329#_c_1613_n N_VGND_c_2293_n 0.00894049f $X=10.335 $Y=0.765
+ $X2=0 $Y2=0
cc_1127 N_A_1597_329#_c_1645_n N_VGND_c_2293_n 0.0185403f $X=9.685 $Y=0.395
+ $X2=0 $Y2=0
cc_1128 N_A_1597_329#_c_1622_n N_VGND_c_2293_n 0.00204496f $X=9.77 $Y=0.845
+ $X2=0 $Y2=0
cc_1129 N_A_1597_329#_c_1624_n N_VGND_c_2293_n 0.0106024f $X=10.395 $Y=0.93
+ $X2=0 $Y2=0
cc_1130 N_A_1597_329#_c_1615_n N_VGND_c_2294_n 0.00410222f $X=11.34 $Y=1.16
+ $X2=0 $Y2=0
cc_1131 N_A_1597_329#_c_1616_n N_VGND_c_2294_n 0.00438629f $X=11.415 $Y=0.995
+ $X2=0 $Y2=0
cc_1132 N_A_1597_329#_c_1617_n N_VGND_c_2295_n 0.0177979f $X=11.835 $Y=0.995
+ $X2=0 $Y2=0
cc_1133 N_A_1597_329#_c_1618_n N_VGND_c_2295_n 0.00915844f $X=12.765 $Y=1.16
+ $X2=0 $Y2=0
cc_1134 N_A_1597_329#_M1011_g N_VGND_c_2295_n 0.00274822f $X=12.84 $Y=0.445
+ $X2=0 $Y2=0
cc_1135 N_A_1597_329#_M1011_g N_VGND_c_2296_n 0.0141499f $X=12.84 $Y=0.445 $X2=0
+ $Y2=0
cc_1136 N_A_1597_329#_c_1645_n N_VGND_c_2301_n 0.0709356f $X=9.685 $Y=0.395
+ $X2=0 $Y2=0
cc_1137 N_A_1597_329#_c_1613_n N_VGND_c_2303_n 0.00486043f $X=10.335 $Y=0.765
+ $X2=0 $Y2=0
cc_1138 N_A_1597_329#_c_1614_n N_VGND_c_2303_n 0.00112301f $X=10.405 $Y=1.325
+ $X2=0 $Y2=0
cc_1139 N_A_1597_329#_c_1616_n N_VGND_c_2308_n 0.00541359f $X=11.415 $Y=0.995
+ $X2=0 $Y2=0
cc_1140 N_A_1597_329#_c_1617_n N_VGND_c_2308_n 0.00442682f $X=11.835 $Y=0.995
+ $X2=0 $Y2=0
cc_1141 N_A_1597_329#_M1011_g N_VGND_c_2309_n 0.0046653f $X=12.84 $Y=0.445 $X2=0
+ $Y2=0
cc_1142 N_A_1597_329#_M1043_d N_VGND_c_2319_n 0.0036355f $X=8.465 $Y=0.235 $X2=0
+ $Y2=0
cc_1143 N_A_1597_329#_c_1613_n N_VGND_c_2319_n 0.0058467f $X=10.335 $Y=0.765
+ $X2=0 $Y2=0
cc_1144 N_A_1597_329#_c_1614_n N_VGND_c_2319_n 0.00144869f $X=10.405 $Y=1.325
+ $X2=0 $Y2=0
cc_1145 N_A_1597_329#_c_1616_n N_VGND_c_2319_n 0.0108276f $X=11.415 $Y=0.995
+ $X2=0 $Y2=0
cc_1146 N_A_1597_329#_c_1617_n N_VGND_c_2319_n 0.00867323f $X=11.835 $Y=0.995
+ $X2=0 $Y2=0
cc_1147 N_A_1597_329#_M1011_g N_VGND_c_2319_n 0.00934473f $X=12.84 $Y=0.445
+ $X2=0 $Y2=0
cc_1148 N_A_1597_329#_c_1645_n N_VGND_c_2319_n 0.0499447f $X=9.685 $Y=0.395
+ $X2=0 $Y2=0
cc_1149 N_A_1597_329#_c_1624_n N_VGND_c_2319_n 0.0118873f $X=10.395 $Y=0.93
+ $X2=0 $Y2=0
cc_1150 N_A_1597_329#_c_1645_n A_1813_47# 0.004771f $X=9.685 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_1151 N_A_1597_329#_c_1645_n A_1885_47# 0.00608206f $X=9.685 $Y=0.395
+ $X2=-0.19 $Y2=-0.24
cc_1152 N_A_1597_329#_c_1622_n A_1885_47# 0.00172677f $X=9.77 $Y=0.845 $X2=-0.19
+ $Y2=-0.24
cc_1153 N_A_2501_47#_c_1800_n N_VPWR_c_1902_n 0.0647312f $X=12.63 $Y=1.935 $X2=0
+ $Y2=0
cc_1154 N_A_2501_47#_M1006_g N_VPWR_c_1903_n 0.00251482f $X=13.315 $Y=1.985
+ $X2=0 $Y2=0
cc_1155 N_A_2501_47#_c_1800_n N_VPWR_c_1903_n 0.0386585f $X=12.63 $Y=1.935 $X2=0
+ $Y2=0
cc_1156 N_A_2501_47#_c_1796_n N_VPWR_c_1903_n 0.0177211f $X=13.26 $Y=1.16 $X2=0
+ $Y2=0
cc_1157 N_A_2501_47#_c_1797_n N_VPWR_c_1903_n 0.00222195f $X=13.735 $Y=1.16
+ $X2=0 $Y2=0
cc_1158 N_A_2501_47#_M1017_g N_VPWR_c_1905_n 0.00590436f $X=13.735 $Y=1.985
+ $X2=0 $Y2=0
cc_1159 N_A_2501_47#_c_1800_n N_VPWR_c_1917_n 0.0131202f $X=12.63 $Y=1.935 $X2=0
+ $Y2=0
cc_1160 N_A_2501_47#_M1006_g N_VPWR_c_1918_n 0.00583607f $X=13.315 $Y=1.985
+ $X2=0 $Y2=0
cc_1161 N_A_2501_47#_M1017_g N_VPWR_c_1918_n 0.004671f $X=13.735 $Y=1.985 $X2=0
+ $Y2=0
cc_1162 N_A_2501_47#_M1006_g N_VPWR_c_1894_n 0.0106798f $X=13.315 $Y=1.985 $X2=0
+ $Y2=0
cc_1163 N_A_2501_47#_M1017_g N_VPWR_c_1894_n 0.00880968f $X=13.735 $Y=1.985
+ $X2=0 $Y2=0
cc_1164 N_A_2501_47#_c_1800_n N_VPWR_c_1894_n 0.00704765f $X=12.63 $Y=1.935
+ $X2=0 $Y2=0
cc_1165 N_A_2501_47#_c_1795_n N_Q_N_c_2249_n 0.00291039f $X=12.63 $Y=0.44 $X2=0
+ $Y2=0
cc_1166 N_A_2501_47#_c_1800_n N_Q_N_c_2249_n 0.00424543f $X=12.63 $Y=1.935 $X2=0
+ $Y2=0
cc_1167 N_A_2501_47#_c_1811_n N_Q_N_c_2249_n 0.00839287f $X=12.622 $Y=1.16 $X2=0
+ $Y2=0
cc_1168 N_A_2501_47#_c_1794_n Q 0.00391291f $X=13.735 $Y=0.995 $X2=0 $Y2=0
cc_1169 N_A_2501_47#_c_1797_n Q 0.00103509f $X=13.735 $Y=1.16 $X2=0 $Y2=0
cc_1170 N_A_2501_47#_M1017_g Q 0.0128627f $X=13.735 $Y=1.985 $X2=0 $Y2=0
cc_1171 N_A_2501_47#_c_1794_n N_Q_c_2273_n 0.00646675f $X=13.735 $Y=0.995 $X2=0
+ $Y2=0
cc_1172 N_A_2501_47#_c_1793_n Q 0.00275116f $X=13.315 $Y=0.995 $X2=0 $Y2=0
cc_1173 N_A_2501_47#_M1006_g Q 0.00275116f $X=13.315 $Y=1.985 $X2=0 $Y2=0
cc_1174 N_A_2501_47#_c_1794_n Q 0.00727939f $X=13.735 $Y=0.995 $X2=0 $Y2=0
cc_1175 N_A_2501_47#_M1017_g Q 0.00907839f $X=13.735 $Y=1.985 $X2=0 $Y2=0
cc_1176 N_A_2501_47#_c_1796_n Q 0.0254774f $X=13.26 $Y=1.16 $X2=0 $Y2=0
cc_1177 N_A_2501_47#_c_1797_n Q 0.0267269f $X=13.735 $Y=1.16 $X2=0 $Y2=0
cc_1178 N_A_2501_47#_M1017_g Q 0.00391291f $X=13.735 $Y=1.985 $X2=0 $Y2=0
cc_1179 N_A_2501_47#_c_1797_n Q 0.00105578f $X=13.735 $Y=1.16 $X2=0 $Y2=0
cc_1180 N_A_2501_47#_c_1795_n N_VGND_c_2295_n 0.0416294f $X=12.63 $Y=0.44 $X2=0
+ $Y2=0
cc_1181 N_A_2501_47#_c_1793_n N_VGND_c_2296_n 0.00330487f $X=13.315 $Y=0.995
+ $X2=0 $Y2=0
cc_1182 N_A_2501_47#_c_1795_n N_VGND_c_2296_n 0.0280689f $X=12.63 $Y=0.44 $X2=0
+ $Y2=0
cc_1183 N_A_2501_47#_c_1796_n N_VGND_c_2296_n 0.0275537f $X=13.26 $Y=1.16 $X2=0
+ $Y2=0
cc_1184 N_A_2501_47#_c_1797_n N_VGND_c_2296_n 0.00248507f $X=13.735 $Y=1.16
+ $X2=0 $Y2=0
cc_1185 N_A_2501_47#_c_1794_n N_VGND_c_2298_n 0.00495486f $X=13.735 $Y=0.995
+ $X2=0 $Y2=0
cc_1186 N_A_2501_47#_c_1795_n N_VGND_c_2309_n 0.0126596f $X=12.63 $Y=0.44 $X2=0
+ $Y2=0
cc_1187 N_A_2501_47#_c_1793_n N_VGND_c_2310_n 0.00583607f $X=13.315 $Y=0.995
+ $X2=0 $Y2=0
cc_1188 N_A_2501_47#_c_1794_n N_VGND_c_2310_n 0.00467644f $X=13.735 $Y=0.995
+ $X2=0 $Y2=0
cc_1189 N_A_2501_47#_M1011_s N_VGND_c_2319_n 0.00477433f $X=12.505 $Y=0.235
+ $X2=0 $Y2=0
cc_1190 N_A_2501_47#_c_1793_n N_VGND_c_2319_n 0.0106371f $X=13.315 $Y=0.995
+ $X2=0 $Y2=0
cc_1191 N_A_2501_47#_c_1794_n N_VGND_c_2319_n 0.00881968f $X=13.735 $Y=0.995
+ $X2=0 $Y2=0
cc_1192 N_A_2501_47#_c_1795_n N_VGND_c_2319_n 0.00704765f $X=12.63 $Y=0.44 $X2=0
+ $Y2=0
cc_1193 N_A_27_369#_c_1853_n N_VPWR_M1025_d 0.00315122f $X=1.015 $Y=1.96
+ $X2=-0.19 $Y2=1.305
cc_1194 N_A_27_369#_c_1853_n N_VPWR_c_1895_n 0.0140834f $X=1.015 $Y=1.96 $X2=0
+ $Y2=0
cc_1195 N_A_27_369#_c_1853_n N_VPWR_c_1912_n 0.00241588f $X=1.015 $Y=1.96 $X2=0
+ $Y2=0
cc_1196 N_A_27_369#_c_1855_n N_VPWR_c_1912_n 0.0178803f $X=0.26 $Y=2.07 $X2=0
+ $Y2=0
cc_1197 N_A_27_369#_c_1853_n N_VPWR_c_1913_n 0.00242264f $X=1.015 $Y=1.96 $X2=0
+ $Y2=0
cc_1198 N_A_27_369#_c_1868_n N_VPWR_c_1913_n 0.00965331f $X=1.185 $Y=2.36 $X2=0
+ $Y2=0
cc_1199 N_A_27_369#_c_1854_n N_VPWR_c_1913_n 0.0536236f $X=1.94 $Y=2.34 $X2=0
+ $Y2=0
cc_1200 N_A_27_369#_M1025_s N_VPWR_c_1894_n 0.00228283f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_1201 N_A_27_369#_M1032_d N_VPWR_c_1894_n 0.00209344f $X=1.805 $Y=1.845 $X2=0
+ $Y2=0
cc_1202 N_A_27_369#_c_1853_n N_VPWR_c_1894_n 0.0100664f $X=1.015 $Y=1.96 $X2=0
+ $Y2=0
cc_1203 N_A_27_369#_c_1868_n N_VPWR_c_1894_n 0.00648546f $X=1.185 $Y=2.36 $X2=0
+ $Y2=0
cc_1204 N_A_27_369#_c_1854_n N_VPWR_c_1894_n 0.0330273f $X=1.94 $Y=2.34 $X2=0
+ $Y2=0
cc_1205 N_A_27_369#_c_1855_n N_VPWR_c_1894_n 0.00991202f $X=0.26 $Y=2.07 $X2=0
+ $Y2=0
cc_1206 N_A_27_369#_c_1853_n A_193_369# 0.00140409f $X=1.015 $Y=1.96 $X2=-0.19
+ $Y2=1.305
cc_1207 N_A_27_369#_c_1868_n A_193_369# 9.36188e-19 $X=1.185 $Y=2.36 $X2=-0.19
+ $Y2=1.305
cc_1208 N_A_27_369#_c_1854_n N_A_181_47#_M1004_d 0.00434085f $X=1.94 $Y=2.34
+ $X2=0 $Y2=0
cc_1209 N_A_27_369#_c_1854_n N_A_181_47#_c_2132_n 0.0178345f $X=1.94 $Y=2.34
+ $X2=0 $Y2=0
cc_1210 N_A_27_369#_c_1854_n N_A_181_47#_c_2125_n 0.00152909f $X=1.94 $Y=2.34
+ $X2=0 $Y2=0
cc_1211 N_VPWR_c_1894_n A_193_369# 0.00187591f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1212 N_VPWR_c_1894_n N_A_181_47#_M1004_d 0.00265018f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1213 N_VPWR_c_1894_n N_A_181_47#_M1007_s 0.00194602f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1214 N_VPWR_c_1915_n N_A_181_47#_c_2122_n 0.0136544f $X=6 $Y=2.72 $X2=0 $Y2=0
cc_1215 N_VPWR_c_1894_n N_A_181_47#_c_2122_n 0.00404777f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1216 N_VPWR_c_1896_n N_A_181_47#_c_2124_n 0.00717133f $X=2.87 $Y=2.34 $X2=0
+ $Y2=0
cc_1217 N_VPWR_c_1894_n A_1102_413# 0.00202059f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1218 N_VPWR_c_1924_n A_1525_329# 9.61034e-19 $X=8.015 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1219 N_VPWR_c_1894_n A_1723_413# 0.00232248f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1220 N_VPWR_c_1894_n N_Q_N_M1012_s 0.00215201f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1221 N_VPWR_c_1902_n N_Q_N_c_2249_n 0.0763475f $X=12.11 $Y=1.66 $X2=0 $Y2=0
cc_1222 N_VPWR_c_1916_n N_Q_N_c_2249_n 0.0233356f $X=12.025 $Y=2.72 $X2=0 $Y2=0
cc_1223 N_VPWR_c_1894_n N_Q_N_c_2249_n 0.0144277f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1224 N_VPWR_c_1894_n N_Q_M1006_s 0.00285153f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1225 N_VPWR_c_1918_n Q 0.0179105f $X=13.91 $Y=2.72 $X2=0 $Y2=0
cc_1226 N_VPWR_c_1894_n Q 0.0121049f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1227 N_VPWR_c_1905_n Q 0.0736255f $X=13.995 $Y=1.66 $X2=0 $Y2=0
cc_1228 N_VPWR_c_1901_n N_VGND_c_2294_n 0.00562283f $X=11.205 $Y=1.66 $X2=0
+ $Y2=0
cc_1229 N_VPWR_c_1902_n N_VGND_c_2295_n 0.0102631f $X=12.11 $Y=1.66 $X2=0 $Y2=0
cc_1230 N_VPWR_c_1905_n N_VGND_c_2298_n 0.00938925f $X=13.995 $Y=1.66 $X2=0
+ $Y2=0
cc_1231 N_A_181_47#_c_2116_n N_VGND_c_2299_n 0.0464212f $X=1.495 $Y=0.425 $X2=0
+ $Y2=0
cc_1232 N_A_181_47#_c_2117_n N_VGND_c_2307_n 0.024686f $X=4.745 $Y=0.42 $X2=0
+ $Y2=0
cc_1233 N_A_181_47#_M1016_d N_VGND_c_2319_n 0.00215227f $X=0.905 $Y=0.235 $X2=0
+ $Y2=0
cc_1234 N_A_181_47#_M1030_s N_VGND_c_2319_n 0.00209319f $X=4.62 $Y=0.235 $X2=0
+ $Y2=0
cc_1235 N_A_181_47#_c_2116_n N_VGND_c_2319_n 0.0298675f $X=1.495 $Y=0.425 $X2=0
+ $Y2=0
cc_1236 N_A_181_47#_c_2117_n N_VGND_c_2319_n 0.014462f $X=4.745 $Y=0.42 $X2=0
+ $Y2=0
cc_1237 N_A_181_47#_c_2116_n A_265_47# 0.00487325f $X=1.495 $Y=0.425 $X2=-0.19
+ $Y2=-0.24
cc_1238 N_Q_N_c_2249_n N_VGND_c_2295_n 0.0490806f $X=11.625 $Y=0.38 $X2=0 $Y2=0
cc_1239 N_Q_N_c_2249_n N_VGND_c_2308_n 0.0233356f $X=11.625 $Y=0.38 $X2=0 $Y2=0
cc_1240 N_Q_N_M1035_s N_VGND_c_2319_n 0.00215201f $X=11.49 $Y=0.235 $X2=0 $Y2=0
cc_1241 N_Q_N_c_2249_n N_VGND_c_2319_n 0.0144277f $X=11.625 $Y=0.38 $X2=0 $Y2=0
cc_1242 N_Q_c_2273_n N_VGND_c_2298_n 0.0466822f $X=13.525 $Y=0.44 $X2=0 $Y2=0
cc_1243 N_Q_c_2273_n N_VGND_c_2310_n 0.0173391f $X=13.525 $Y=0.44 $X2=0 $Y2=0
cc_1244 N_Q_M1040_s N_VGND_c_2319_n 0.00290484f $X=13.39 $Y=0.235 $X2=0 $Y2=0
cc_1245 N_Q_c_2273_n N_VGND_c_2319_n 0.0121108f $X=13.525 $Y=0.44 $X2=0 $Y2=0
cc_1246 N_VGND_c_2311_n A_109_47# 9.17637e-19 $X=0.23 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1247 N_VGND_c_2319_n A_109_47# 7.33531e-19 $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1248 N_VGND_c_2319_n A_265_47# 0.00252958f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1249 N_VGND_c_2319_n A_1090_47# 0.00776438f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1250 N_VGND_c_2316_n A_1517_47# 0.0109537f $X=7.705 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1251 N_VGND_c_2319_n A_1517_47# 0.0131461f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1252 N_VGND_c_2319_n A_1813_47# 0.00169327f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1253 N_VGND_c_2319_n A_1885_47# 0.00282192f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__and2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.765000 0.450000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.645000 2.200000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.580000 2.680000 2.365000 ;
        RECT 2.445000 0.255000 2.680000 0.775000 ;
        RECT 2.505000 0.775000 2.680000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.590000 ;
        RECT 1.875000  0.085000 2.275000 0.580000 ;
        RECT 2.865000  0.085000 3.135000 0.720000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 0.515000 2.185000 0.845000 2.635000 ;
        RECT 1.510000 2.165000 2.195000 2.635000 ;
        RECT 2.865000 1.680000 3.135000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 1.785000 0.855000 2.015000 ;
      RECT 0.175000 2.015000 0.345000 2.445000 ;
      RECT 0.595000 0.280000 0.835000 0.655000 ;
      RECT 0.620000 0.655000 0.835000 0.805000 ;
      RECT 0.620000 0.805000 1.175000 1.135000 ;
      RECT 0.620000 1.135000 0.855000 1.785000 ;
      RECT 1.045000 1.305000 2.335000 1.325000 ;
      RECT 1.045000 1.325000 1.905000 1.475000 ;
      RECT 1.045000 1.475000 1.330000 2.420000 ;
      RECT 1.115000 0.270000 1.285000 0.415000 ;
      RECT 1.115000 0.415000 1.515000 0.610000 ;
      RECT 1.345000 0.610000 1.515000 0.945000 ;
      RECT 1.345000 0.945000 2.335000 1.305000 ;
  END
END sky130_fd_sc_hd__and2b_2
END LIBRARY

* File: sky130_fd_sc_hd__lpflow_decapkapwr_12.pex.spice
* Created: Tue Sep  1 19:11:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%VGND 1 9 10 11 12 14 22 34 37
r28 36 37 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r29 34 36 0.448529 $w=8.16e-07 $l=3e-08 $layer=LI1_cond $X=5.26 $Y=0.385
+ $X2=5.29 $Y2=0.385
r30 31 37 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=5.29
+ $Y2=0
r31 30 31 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r32 24 27 0.25811 $w=1.418e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.645
+ $X2=0.26 $Y2=0.645
r33 21 30 15.4006 $w=1.418e-06 $l=1.79e-06 $layer=LI1_cond $X=2.48 $Y=0.645
+ $X2=0.69 $Y2=0.645
r34 20 22 8.47369 $w=1.49e-06 $l=1.65e-07 $layer=POLY_cond $X=2.48 $Y=1.87
+ $X2=2.645 $Y2=1.87
r35 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.48
+ $Y=1.29 $X2=2.48 $Y2=1.29
r36 17 30 1.11848 $w=1.418e-06 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=0.645
+ $X2=0.69 $Y2=0.645
r37 17 27 2.5811 $w=1.418e-06 $l=3e-07 $layer=LI1_cond $X=0.56 $Y=0.645 $X2=0.26
+ $Y2=0.645
r38 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.56
+ $Y=1.29 $X2=0.56 $Y2=1.29
r39 14 20 19.2327 $w=1.49e-06 $l=5.8e-07 $layer=POLY_cond $X=1.9 $Y=1.87
+ $X2=2.48 $Y2=1.87
r40 14 16 44.4343 $w=1.49e-06 $l=1.34e-06 $layer=POLY_cond $X=1.9 $Y=1.87
+ $X2=0.56 $Y2=1.87
r41 12 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r42 12 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r43 11 21 2.97997 $w=1.418e-06 $l=3.40147e-07 $layer=LI1_cond $X=2.665 $Y=0.385
+ $X2=2.48 $Y2=0.645
r44 10 34 4.13877 $w=9.4e-07 $l=3e-07 $layer=LI1_cond $X=4.96 $Y=0.385 $X2=5.26
+ $Y2=0.385
r45 10 11 29.7862 $w=9.38e-07 $l=2.295e-06 $layer=LI1_cond $X=4.96 $Y=0.385
+ $X2=2.665 $Y2=0.385
r46 9 22 4.90531 $w=1.13e-06 $l=1.15e-07 $layer=POLY_cond $X=2.76 $Y=2.05
+ $X2=2.645 $Y2=2.05
r47 1 34 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=5.125 $Y=0.235
+ $X2=5.26 $Y2=0.475
r48 1 27 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%KAPWR 1 9 10 15 18 22 24 37 38
+ 40 42
c30 38 0 1.06778e-19 $X=5.29 $Y=2.21
r31 40 42 0.0085136 $w=2.6e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=2.21
+ $X2=0.23 $Y2=2.21
r32 37 38 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=5.29 $Y=2.21
+ $X2=5.29 $Y2=2.21
r33 35 37 0.254167 $w=1.438e-06 $l=3e-08 $layer=LI1_cond $X=5.26 $Y=1.745
+ $X2=5.29 $Y2=1.745
r34 28 32 0.397826 $w=9.18e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=2.005
+ $X2=0.26 $Y2=2.005
r35 28 42 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.23 $Y=2.21
+ $X2=0.23 $Y2=2.21
r36 25 35 2.71111 $w=1.438e-06 $l=3.2e-07 $layer=LI1_cond $X=4.94 $Y=1.745
+ $X2=5.26 $Y2=1.745
r37 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.94
+ $Y=1.11 $X2=4.94 $Y2=1.11
r38 18 40 0.0120192 $w=2.6e-07 $l=2.5e-08 $layer=MET1_cond $X=0.19 $Y=2.21
+ $X2=0.215 $Y2=2.21
r39 18 38 2.84524 $w=2.6e-07 $l=5.013e-06 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=5.29 $Y2=2.21
r40 18 42 0.0266759 $w=2.6e-07 $l=4.7e-08 $layer=MET1_cond $X=0.277 $Y=2.21
+ $X2=0.23 $Y2=2.21
r41 15 32 34.1467 $w=9.18e-07 $l=2.575e-06 $layer=LI1_cond $X=2.835 $Y=2.005
+ $X2=0.26 $Y2=2.005
r42 14 24 84.3769 $w=1.17e-06 $l=1.92e-06 $layer=POLY_cond $X=3.02 $Y=0.69
+ $X2=4.94 $Y2=0.69
r43 14 22 12.167 $w=1.17e-06 $l=1.65e-07 $layer=POLY_cond $X=3.02 $Y=0.69
+ $X2=2.855 $Y2=0.69
r44 13 15 3.1528 $w=1.438e-06 $l=1.85e-07 $layer=LI1_cond $X=3.02 $Y=1.745
+ $X2=2.835 $Y2=1.745
r45 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.02
+ $Y=1.11 $X2=3.02 $Y2=1.11
r46 10 25 11.734 $w=1.438e-06 $l=1.385e-06 $layer=LI1_cond $X=3.555 $Y=1.745
+ $X2=4.94 $Y2=1.745
r47 10 13 4.53264 $w=1.438e-06 $l=5.35e-07 $layer=LI1_cond $X=3.555 $Y=1.745
+ $X2=3.02 $Y2=1.745
r48 9 22 5.65309 $w=8.1e-07 $l=9.5e-08 $layer=POLY_cond $X=2.76 $Y=0.51
+ $X2=2.855 $Y2=0.51
r49 1 35 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.615 $X2=5.26 $Y2=1.83
r50 1 32 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_DECAPKAPWR_12%VPWR 1 8 9
c11 8 0 1.06778e-19 $X=5.29 $Y=2.72
r12 8 9 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r13 4 8 330.118 $w=1.68e-07 $l=5.06e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=5.29
+ $Y2=2.72
r14 1 9 1.43978 $w=4.8e-07 $l=5.06e-06 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=5.29
+ $Y2=2.72
r15 1 4 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
.ends


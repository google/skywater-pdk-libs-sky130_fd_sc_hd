* File: sky130_fd_sc_hd__a41o_4.spice.pex
* Created: Thu Aug 27 14:06:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A41O_4%A_79_21# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 38 47 49 50 51 52 53 56 60 66 67 69 76
r125 73 74 61.7195 $w=3.28e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r126 63 69 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=1.955
+ $X2=2.88 $Y2=2.04
r127 63 65 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.88 $Y=1.955
+ $X2=2.88 $Y2=1.7
r128 62 65 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.88 $Y=1.625
+ $X2=2.88 $Y2=1.7
r129 58 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.73
+ $X2=2.38 $Y2=0.73
r130 58 60 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=2.465 $Y=0.73
+ $X2=3.74 $Y2=0.73
r131 54 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=0.645
+ $X2=2.38 $Y2=0.73
r132 54 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.38 $Y=0.645
+ $X2=2.38 $Y2=0.42
r133 52 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.795 $Y=1.54
+ $X2=2.88 $Y2=1.625
r134 52 53 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.795 $Y=1.54
+ $X2=1.945 $Y2=1.54
r135 50 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=0.73
+ $X2=2.38 $Y2=0.73
r136 50 51 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.295 $Y=0.73
+ $X2=1.945 $Y2=0.73
r137 49 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.86 $Y=1.455
+ $X2=1.945 $Y2=1.54
r138 48 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=1.245
+ $X2=1.86 $Y2=1.16
r139 48 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.86 $Y=1.245
+ $X2=1.86 $Y2=1.455
r140 47 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=1.075
+ $X2=1.86 $Y2=1.16
r141 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.86 $Y=0.815
+ $X2=1.945 $Y2=0.73
r142 46 47 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.86 $Y=0.815
+ $X2=1.86 $Y2=1.075
r143 45 76 8.08232 $w=3.28e-07 $l=5.5e-08 $layer=POLY_cond $X=1.675 $Y=1.16
+ $X2=1.73 $Y2=1.16
r144 45 74 53.6372 $w=3.28e-07 $l=3.65e-07 $layer=POLY_cond $X=1.675 $Y=1.16
+ $X2=1.31 $Y2=1.16
r145 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r146 41 73 34.5335 $w=3.28e-07 $l=2.35e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.89 $Y2=1.16
r147 41 71 27.186 $w=3.28e-07 $l=1.85e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.47 $Y2=1.16
r148 40 44 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.655 $Y=1.16
+ $X2=1.675 $Y2=1.16
r149 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.655
+ $Y=1.16 $X2=0.655 $Y2=1.16
r150 38 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=1.16
+ $X2=1.86 $Y2=1.16
r151 38 44 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.775 $Y=1.16
+ $X2=1.675 $Y2=1.16
r152 34 76 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r153 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r154 31 76 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r155 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r156 27 74 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r157 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r158 24 74 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r159 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r160 20 73 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r161 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r162 17 73 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r163 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r164 13 71 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r165 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r166 10 71 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r167 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r168 3 69 600 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2.04
r169 3 65 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.7
r170 2 60 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.235 $X2=3.74 $Y2=0.73
r171 1 56 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%B1 1 3 4 6 9 13 15 16 29
r52 27 29 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.98 $Y=1.16
+ $X2=3.09 $Y2=1.16
r53 25 27 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=2.67 $Y=1.16 $X2=2.98
+ $Y2=1.16
r54 24 25 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.59 $Y=1.16 $X2=2.67
+ $Y2=1.16
r55 22 24 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=2.3 $Y=1.16 $X2=2.59
+ $Y2=1.16
r56 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=1.16 $X2=2.3 $Y2=1.16
r57 19 22 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.17 $Y=1.16 $X2=2.3
+ $Y2=1.16
r58 16 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=1.16 $X2=2.98 $Y2=1.16
r59 15 16 22.9933 $w=2.03e-07 $l=4.25e-07 $layer=LI1_cond $X=2.555 $Y=1.177
+ $X2=2.98 $Y2=1.177
r60 15 23 13.796 $w=2.03e-07 $l=2.55e-07 $layer=LI1_cond $X=2.555 $Y=1.177
+ $X2=2.3 $Y2=1.177
r61 11 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.325
+ $X2=3.09 $Y2=1.16
r62 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.09 $Y=1.325
+ $X2=3.09 $Y2=1.985
r63 7 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.325
+ $X2=2.67 $Y2=1.16
r64 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.67 $Y=1.325 $X2=2.67
+ $Y2=1.985
r65 4 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.16
r66 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995 $X2=2.59
+ $Y2=0.56
r67 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r68 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995 $X2=2.17
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A1 1 3 6 8 10 13 15 16 23
c42 23 0 1.90366e-19 $X=3.95 $Y=1.16
c43 8 0 1.21078e-19 $X=3.95 $Y=0.995
r44 21 23 7.50779 $w=3.21e-07 $l=5e-08 $layer=POLY_cond $X=3.9 $Y=1.16 $X2=3.95
+ $Y2=1.16
r45 19 21 55.5576 $w=3.21e-07 $l=3.7e-07 $layer=POLY_cond $X=3.53 $Y=1.16
+ $X2=3.9 $Y2=1.16
r46 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.9 $Y=1.16
+ $X2=3.9 $Y2=1.16
r47 15 16 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=3.495 $Y=1.185
+ $X2=3.9 $Y2=1.185
r48 11 23 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.325
+ $X2=3.95 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.95 $Y=1.325
+ $X2=3.95 $Y2=1.985
r50 8 23 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.95 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.95 $Y2=0.56
r52 4 19 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.53 $Y=1.325 $X2=3.53
+ $Y2=1.985
r54 1 19 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.53 $Y=0.995 $X2=3.53
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A2 3 7 11 15 17 18 26
r43 24 26 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=4.78 $Y=1.16 $X2=4.79
+ $Y2=1.16
r44 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.78
+ $Y=1.16 $X2=4.78 $Y2=1.16
r45 21 24 91.0912 $w=2.7e-07 $l=4.1e-07 $layer=POLY_cond $X=4.37 $Y=1.16
+ $X2=4.78 $Y2=1.16
r46 18 25 5.01732 $w=2.08e-07 $l=9.5e-08 $layer=LI1_cond $X=4.875 $Y=1.18
+ $X2=4.78 $Y2=1.18
r47 17 25 19.2771 $w=2.08e-07 $l=3.65e-07 $layer=LI1_cond $X=4.415 $Y=1.18
+ $X2=4.78 $Y2=1.18
r48 13 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.79 $Y=1.295
+ $X2=4.79 $Y2=1.16
r49 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.79 $Y=1.295
+ $X2=4.79 $Y2=1.985
r50 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.79 $Y=1.025
+ $X2=4.79 $Y2=1.16
r51 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.79 $Y=1.025
+ $X2=4.79 $Y2=0.56
r52 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.37 $Y=1.295
+ $X2=4.37 $Y2=1.16
r53 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.37 $Y=1.295 $X2=4.37
+ $Y2=1.985
r54 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.37 $Y=1.025
+ $X2=4.37 $Y2=1.16
r55 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.37 $Y=1.025
+ $X2=4.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A3 3 7 11 15 17 18 19 22 29 30
r49 28 30 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=6.02 $Y=1.16
+ $X2=6.15 $Y2=1.16
r50 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.02
+ $Y=1.16 $X2=6.02 $Y2=1.16
r51 26 28 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=5.73 $Y=1.16
+ $X2=6.02 $Y2=1.16
r52 22 26 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.655 $Y=1.16
+ $X2=5.73 $Y2=1.16
r53 22 24 74.4282 $w=2.7e-07 $l=3.35e-07 $layer=POLY_cond $X=5.655 $Y=1.16
+ $X2=5.32 $Y2=1.16
r54 19 29 10.7387 $w=2.18e-07 $l=2.05e-07 $layer=LI1_cond $X=5.815 $Y=1.185
+ $X2=6.02 $Y2=1.185
r55 18 19 25.93 $w=2.18e-07 $l=4.95e-07 $layer=LI1_cond $X=5.32 $Y=1.185
+ $X2=5.815 $Y2=1.185
r56 18 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.32
+ $Y=1.16 $X2=5.32 $Y2=1.16
r57 17 24 3.33261 $w=2.7e-07 $l=1.5e-08 $layer=POLY_cond $X=5.305 $Y=1.16
+ $X2=5.32 $Y2=1.16
r58 13 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.15 $Y=1.295
+ $X2=6.15 $Y2=1.16
r59 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.15 $Y=1.295
+ $X2=6.15 $Y2=1.985
r60 9 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.15 $Y=1.025
+ $X2=6.15 $Y2=1.16
r61 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.15 $Y=1.025
+ $X2=6.15 $Y2=0.56
r62 5 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.73 $Y=1.025
+ $X2=5.73 $Y2=1.16
r63 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.73 $Y=1.025
+ $X2=5.73 $Y2=0.56
r64 1 17 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=5.23 $Y=1.295
+ $X2=5.305 $Y2=1.16
r65 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.23 $Y=1.295 $X2=5.23
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A4 3 7 11 15 17 18 21 23 24
r38 29 31 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=6.66 $Y=1.16
+ $X2=6.99 $Y2=1.16
r39 26 29 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.57 $Y=1.16 $X2=6.66
+ $Y2=1.16
r40 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.16 $X2=7.34 $Y2=1.16
r41 21 31 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=7.065 $Y=1.16
+ $X2=6.99 $Y2=1.16
r42 21 23 61.0978 $w=2.7e-07 $l=2.75e-07 $layer=POLY_cond $X=7.065 $Y=1.16
+ $X2=7.34 $Y2=1.16
r43 18 24 7.59565 $w=2.18e-07 $l=1.45e-07 $layer=LI1_cond $X=7.195 $Y=1.185
+ $X2=7.34 $Y2=1.185
r44 17 18 28.0253 $w=2.18e-07 $l=5.35e-07 $layer=LI1_cond $X=6.66 $Y=1.185
+ $X2=7.195 $Y2=1.185
r45 17 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.16 $X2=6.66 $Y2=1.16
r46 13 31 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.99 $Y=1.295
+ $X2=6.99 $Y2=1.16
r47 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.99 $Y=1.295
+ $X2=6.99 $Y2=1.985
r48 9 31 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.99 $Y=1.025
+ $X2=6.99 $Y2=1.16
r49 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.99 $Y=1.025
+ $X2=6.99 $Y2=0.56
r50 5 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.57 $Y=1.295
+ $X2=6.57 $Y2=1.16
r51 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.57 $Y=1.295 $X2=6.57
+ $Y2=1.985
r52 1 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.57 $Y=1.025
+ $X2=6.57 $Y2=1.16
r53 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.57 $Y=1.025
+ $X2=6.57 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46 50
+ 53 54 56 57 58 60 65 77 83 84 90 93 96 99
r120 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r121 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r122 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r123 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r125 84 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r126 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r127 81 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=6.78 $Y2=2.72
r128 81 83 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.945 $Y=2.72
+ $X2=7.59 $Y2=2.72
r129 80 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r130 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r131 77 96 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.69 $Y2=2.72
r132 77 79 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r133 76 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r135 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r136 73 94 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r137 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r138 70 93 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=1.95 $Y2=2.72
r139 70 72 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=3.45 $Y2=2.72
r140 69 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 69 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r142 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r143 66 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.1 $Y2=2.72
r144 66 68 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.61 $Y2=2.72
r145 65 93 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.95 $Y2=2.72
r146 65 68 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.61 $Y2=2.72
r147 64 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r149 61 87 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r150 61 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 60 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.1 $Y2=2.72
r152 60 63 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r153 58 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 58 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 56 75 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.415 $Y=2.72
+ $X2=4.37 $Y2=2.72
r156 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=2.72
+ $X2=4.58 $Y2=2.72
r157 55 79 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.745 $Y=2.72
+ $X2=5.29 $Y2=2.72
r158 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=2.72
+ $X2=4.58 $Y2=2.72
r159 53 72 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=2.72
+ $X2=3.45 $Y2=2.72
r160 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=2.72
+ $X2=3.74 $Y2=2.72
r161 52 75 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.905 $Y=2.72
+ $X2=4.37 $Y2=2.72
r162 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=2.72
+ $X2=3.74 $Y2=2.72
r163 48 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.78 $Y=2.635
+ $X2=6.78 $Y2=2.72
r164 48 50 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.78 $Y=2.635
+ $X2=6.78 $Y2=2
r165 47 96 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=6.035 $Y=2.72
+ $X2=5.69 $Y2=2.72
r166 46 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.615 $Y=2.72
+ $X2=6.78 $Y2=2.72
r167 46 47 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.615 $Y=2.72
+ $X2=6.035 $Y2=2.72
r168 42 96 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.69 $Y=2.635
+ $X2=5.69 $Y2=2.72
r169 42 44 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=5.69 $Y=2.635
+ $X2=5.69 $Y2=2
r170 38 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=2.635
+ $X2=4.58 $Y2=2.72
r171 38 40 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.58 $Y=2.635
+ $X2=4.58 $Y2=2
r172 34 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=2.635
+ $X2=3.74 $Y2=2.72
r173 34 36 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.74 $Y=2.635
+ $X2=3.74 $Y2=2
r174 30 93 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=2.635
+ $X2=1.95 $Y2=2.72
r175 30 32 20.9086 $w=3.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.95 $Y=2.635
+ $X2=1.95 $Y2=2
r176 26 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r177 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r178 22 87 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r179 22 24 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2
r180 7 50 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.645
+ $Y=1.485 $X2=6.78 $Y2=2
r181 6 44 150 $w=1.7e-07 $l=7.81153e-07 $layer=licon1_PDIFF $count=4 $X=5.305
+ $Y=1.485 $X2=5.87 $Y2=2
r182 5 40 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.445
+ $Y=1.485 $X2=4.58 $Y2=2
r183 4 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.605
+ $Y=1.485 $X2=3.74 $Y2=2
r184 3 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r185 2 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r186 1 24 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%X 1 2 3 4 15 19 21 23 27 31 33 34 35 36 37 38
+ 39 47 48 50 56
r52 48 56 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.235 $Y=1.575
+ $X2=0.235 $Y2=1.53
r53 47 50 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.235 $Y=0.805
+ $X2=0.235 $Y2=0.85
r54 39 48 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=1.66
+ $X2=0.235 $Y2=1.575
r55 39 56 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.235 $Y=1.51
+ $X2=0.235 $Y2=1.53
r56 38 39 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.235 $Y=1.19
+ $X2=0.235 $Y2=1.51
r57 37 47 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=0.72
+ $X2=0.235 $Y2=0.805
r58 37 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.235 $Y=0.87
+ $X2=0.235 $Y2=1.19
r59 37 50 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.235 $Y=0.87
+ $X2=0.235 $Y2=0.85
r60 35 39 14.9587 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=0.595 $Y=1.66
+ $X2=0.32 $Y2=1.66
r61 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=1.66
+ $X2=0.68 $Y2=1.66
r62 33 37 14.9587 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=0.595 $Y=0.72
+ $X2=0.32 $Y2=0.72
r63 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0.72
+ $X2=0.68 $Y2=0.72
r64 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.52 $Y=1.745
+ $X2=1.52 $Y2=1.96
r65 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.52 $Y=0.635
+ $X2=1.52 $Y2=0.42
r66 24 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.66
+ $X2=0.68 $Y2=1.66
r67 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=1.52 $Y2=1.745
r68 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=0.765 $Y2=1.66
r69 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.72
+ $X2=0.68 $Y2=0.72
r70 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=1.52 $Y2=0.635
r71 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=0.72
+ $X2=0.765 $Y2=0.72
r72 17 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=1.745
+ $X2=0.68 $Y2=1.66
r73 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=1.745
+ $X2=0.68 $Y2=1.96
r74 13 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.68 $Y2=0.72
r75 13 15 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=0.635
+ $X2=0.68 $Y2=0.42
r76 4 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r77 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
r78 2 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.42
r79 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A_467_297# 1 2 3 4 5 6 21 23 24 28 29 30 33
+ 35 39 41 45 47 51 54
c62 30 0 1.90366e-19 $X=3.405 $Y=1.62
r63 49 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.2 $Y=1.705
+ $X2=7.2 $Y2=1.96
r64 48 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.445 $Y=1.62
+ $X2=6.36 $Y2=1.62
r65 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.115 $Y=1.62
+ $X2=7.2 $Y2=1.705
r66 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.115 $Y=1.62
+ $X2=6.445 $Y2=1.62
r67 43 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.36 $Y=1.705
+ $X2=6.36 $Y2=1.62
r68 43 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.36 $Y=1.705
+ $X2=6.36 $Y2=1.96
r69 42 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=1.62
+ $X2=5.02 $Y2=1.62
r70 41 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.275 $Y=1.62
+ $X2=6.36 $Y2=1.62
r71 41 42 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=6.275 $Y=1.62
+ $X2=5.105 $Y2=1.62
r72 37 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.02 $Y=1.705
+ $X2=5.02 $Y2=1.62
r73 37 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.02 $Y=1.705
+ $X2=5.02 $Y2=1.96
r74 36 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=1.62
+ $X2=4.16 $Y2=1.62
r75 35 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=1.62
+ $X2=5.02 $Y2=1.62
r76 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.935 $Y=1.62
+ $X2=4.245 $Y2=1.62
r77 31 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.705
+ $X2=4.16 $Y2=1.62
r78 31 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.16 $Y=1.705
+ $X2=4.16 $Y2=1.96
r79 29 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=1.62
+ $X2=4.16 $Y2=1.62
r80 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.075 $Y=1.62
+ $X2=3.405 $Y2=1.62
r81 26 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.32 $Y=2.295
+ $X2=3.32 $Y2=1.96
r82 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.32 $Y=1.705
+ $X2=3.405 $Y2=1.62
r83 25 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.32 $Y=1.705
+ $X2=3.32 $Y2=1.96
r84 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.235 $Y=2.38
+ $X2=3.32 $Y2=2.295
r85 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.235 $Y=2.38
+ $X2=2.545 $Y2=2.38
r86 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=2.295
+ $X2=2.545 $Y2=2.38
r87 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.46 $Y=2.295
+ $X2=2.46 $Y2=1.96
r88 6 51 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.065
+ $Y=1.485 $X2=7.2 $Y2=1.96
r89 5 45 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.225
+ $Y=1.485 $X2=6.36 $Y2=1.96
r90 4 39 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5.02 $Y2=1.96
r91 3 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.025
+ $Y=1.485 $X2=4.16 $Y2=1.96
r92 2 28 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.485 $X2=3.32 $Y2=1.96
r93 1 21 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 42 44 56 62 63 69 72
r119 72 73 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r120 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r121 63 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=6.67
+ $Y2=0
r122 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r123 60 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.945 $Y=0 $X2=6.78
+ $Y2=0
r124 60 62 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=7.59 $Y2=0
r125 59 73 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=6.67
+ $Y2=0
r126 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r127 56 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.615 $Y=0 $X2=6.78
+ $Y2=0
r128 56 58 236.497 $w=1.68e-07 $l=3.625e-06 $layer=LI1_cond $X=6.615 $Y=0
+ $X2=2.99 $Y2=0
r129 55 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r130 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r131 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r132 52 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r133 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r134 49 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r135 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r136 48 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r137 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r138 45 66 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r139 45 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r140 44 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r141 44 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r142 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r143 42 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r144 40 54 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=0
+ $X2=2.53 $Y2=0
r145 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.8
+ $Y2=0
r146 39 58 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.99
+ $Y2=0
r147 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.8
+ $Y2=0
r148 37 51 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.61 $Y2=0
r149 37 38 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.95
+ $Y2=0
r150 36 54 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=0
+ $X2=2.53 $Y2=0
r151 36 38 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.95
+ $Y2=0
r152 32 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.78 $Y=0.085
+ $X2=6.78 $Y2=0
r153 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.78 $Y=0.085
+ $X2=6.78 $Y2=0.38
r154 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r155 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.38
r156 24 38 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0
r157 24 26 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0.38
r158 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r159 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.38
r160 16 66 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r161 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r162 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.645
+ $Y=0.235 $X2=6.78 $Y2=0.38
r163 4 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.38
r164 3 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r165 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r166 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A_639_47# 1 2 3 10 18
r26 16 21 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.73
+ $X2=4.16 $Y2=0.73
r27 16 18 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.245 $Y=0.73 $X2=5
+ $Y2=0.73
r28 15 21 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=0.645
+ $X2=4.16 $Y2=0.73
r29 14 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.16 $Y=0.465
+ $X2=4.16 $Y2=0.645
r30 10 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.075 $Y=0.38
+ $X2=4.16 $Y2=0.465
r31 10 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.075 $Y=0.38
+ $X2=3.32 $Y2=0.38
r32 3 18 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5 $Y2=0.73
r33 2 21 182 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.235 $X2=4.16 $Y2=0.65
r34 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.235 $X2=3.32 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A_889_47# 1 2 11
c19 11 0 1.21078e-19 $X=5.94 $Y=0.38
r20 8 11 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.58 $Y=0.38
+ $X2=5.94 $Y2=0.38
r21 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.805
+ $Y=0.235 $X2=5.94 $Y2=0.38
r22 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.58 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41O_4%A_1079_47# 1 2 3 10 18
r25 16 18 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.2 $Y=0.645
+ $X2=7.2 $Y2=0.42
r26 12 15 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.52 $Y=0.73
+ $X2=6.36 $Y2=0.73
r27 10 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.115 $Y=0.73
+ $X2=7.2 $Y2=0.645
r28 10 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.115 $Y=0.73
+ $X2=6.36 $Y2=0.73
r29 3 18 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=7.065
+ $Y=0.235 $X2=7.2 $Y2=0.42
r30 2 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=6.225
+ $Y=0.235 $X2=6.36 $Y2=0.73
r31 1 12 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.52 $Y2=0.73
.ends


* File: sky130_fd_sc_hd__nand3b_4.spice
* Created: Thu Aug 27 14:29:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand3b_4.pex.spice"
.subckt sky130_fd_sc_hd__nand3b_4  VNB VPB A_N B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_A_N_M1023_g N_A_27_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_215_47#_M1004_d N_A_27_47#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1006 N_A_215_47#_M1006_d N_A_27_47#_M1006_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1008 N_A_215_47#_M1006_d N_A_27_47#_M1008_g N_Y_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1014 N_A_215_47#_M1014_d N_A_27_47#_M1014_g N_Y_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1007 N_A_633_47#_M1007_d N_B_M1007_g N_A_215_47#_M1014_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.9 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1009 N_A_633_47#_M1007_d N_B_M1009_g N_A_215_47#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.3 SB=75001 A=0.0975 P=1.6 MULT=1
MM1012 N_A_633_47#_M1012_d N_B_M1012_g N_A_215_47#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75002.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1013 N_A_633_47#_M1012_d N_B_M1013_g N_A_215_47#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_C_M1000_g N_A_633_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_C_M1003_g N_A_633_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1003_d N_C_M1005_g N_A_633_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1025_d N_C_M1025_g N_A_633_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.234 AS=0.08775 PD=2.02 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1018 N_VPWR_M1018_d N_A_N_M1018_g N_A_27_47#_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A_27_47#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1001_d N_A_27_47#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1019 N_Y_M1019_d N_A_27_47#_M1019_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1020 N_Y_M1019_d N_A_27_47#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1010_d N_B_M1010_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1011 N_Y_M1010_d N_B_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1016 N_Y_M1016_d N_B_M1016_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1021 N_Y_M1016_d N_B_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1 SB=75000.2 A=0.15
+ P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_C_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_C_M1017_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1017_d N_C_M1022_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.7 A=0.15
+ P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_C_M1024_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1 AD=0.36
+ AS=0.135 PD=2.72 PS=1.27 NRD=14.775 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75000.3
+ A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=12.4227 P=18.69
*
.include "sky130_fd_sc_hd__nand3b_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a221oi_1.pxi.spice
* Created: Thu Aug 27 14:01:59 2020
* 
x_PM_SKY130_FD_SC_HD__A221OI_1%C1 N_C1_c_57_n N_C1_M1008_g N_C1_M1005_g C1
+ N_C1_c_59_n PM_SKY130_FD_SC_HD__A221OI_1%C1
x_PM_SKY130_FD_SC_HD__A221OI_1%B2 N_B2_M1002_g N_B2_M1009_g B2 N_B2_c_84_n
+ N_B2_c_85_n N_B2_c_86_n PM_SKY130_FD_SC_HD__A221OI_1%B2
x_PM_SKY130_FD_SC_HD__A221OI_1%B1 N_B1_M1004_g N_B1_M1000_g B1 B1 N_B1_c_115_n
+ N_B1_c_116_n PM_SKY130_FD_SC_HD__A221OI_1%B1
x_PM_SKY130_FD_SC_HD__A221OI_1%A1 N_A1_M1003_g N_A1_M1006_g A1 A1 N_A1_c_157_n
+ N_A1_c_158_n PM_SKY130_FD_SC_HD__A221OI_1%A1
x_PM_SKY130_FD_SC_HD__A221OI_1%A2 N_A2_M1001_g N_A2_M1007_g A2 N_A2_c_194_n
+ N_A2_c_195_n N_A2_c_196_n PM_SKY130_FD_SC_HD__A221OI_1%A2
x_PM_SKY130_FD_SC_HD__A221OI_1%Y N_Y_M1008_s N_Y_M1004_d N_Y_M1003_s N_Y_M1005_s
+ N_Y_c_309_p N_Y_c_298_p N_Y_c_226_n N_Y_c_227_n N_Y_c_231_n N_Y_c_228_n
+ N_Y_c_259_n N_Y_c_268_n N_Y_c_275_n N_Y_c_277_n N_Y_c_232_n N_Y_c_271_n Y Y Y
+ N_Y_c_229_n N_Y_c_233_n Y PM_SKY130_FD_SC_HD__A221OI_1%Y
x_PM_SKY130_FD_SC_HD__A221OI_1%A_109_297# N_A_109_297#_M1005_d
+ N_A_109_297#_M1000_d N_A_109_297#_c_328_n N_A_109_297#_c_329_n
+ N_A_109_297#_c_327_n N_A_109_297#_c_330_n
+ PM_SKY130_FD_SC_HD__A221OI_1%A_109_297#
x_PM_SKY130_FD_SC_HD__A221OI_1%A_193_297# N_A_193_297#_M1002_d
+ N_A_193_297#_M1006_d N_A_193_297#_c_349_n N_A_193_297#_c_353_n
+ N_A_193_297#_c_359_n N_A_193_297#_c_371_p N_A_193_297#_c_352_n
+ N_A_193_297#_c_350_n PM_SKY130_FD_SC_HD__A221OI_1%A_193_297#
x_PM_SKY130_FD_SC_HD__A221OI_1%VPWR N_VPWR_M1006_s N_VPWR_M1007_d N_VPWR_c_378_n
+ N_VPWR_c_379_n N_VPWR_c_380_n VPWR N_VPWR_c_381_n N_VPWR_c_382_n
+ N_VPWR_c_383_n N_VPWR_c_377_n PM_SKY130_FD_SC_HD__A221OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A221OI_1%VGND N_VGND_M1008_d N_VGND_M1001_d N_VGND_c_425_n
+ N_VGND_c_426_n N_VGND_c_427_n VGND N_VGND_c_428_n N_VGND_c_429_n
+ N_VGND_c_430_n N_VGND_c_431_n PM_SKY130_FD_SC_HD__A221OI_1%VGND
cc_1 VNB N_C1_c_57_n 0.0219373f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB C1 0.00922438f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_C1_c_59_n 0.0394737f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B2_c_84_n 0.0193929f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_5 VNB N_B2_c_85_n 0.00565245f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_6 VNB N_B2_c_86_n 0.0161745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB B1 0.00529535f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_8 VNB B1 0.00498335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_115_n 0.0236812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_c_116_n 0.0187209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A1 0.00154951f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_12 VNB A1 0.00190929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A1_c_157_n 0.0282713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_158_n 0.020504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_194_n 0.0220842f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_16 VNB N_A2_c_195_n 0.00266591f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_17 VNB N_A2_c_196_n 0.0189107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_226_n 0.00585349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_227_n 0.0018364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_228_n 0.0127894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_229_n 0.00791786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB Y 0.0228665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_377_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_425_n 0.00280434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_426_n 0.0115039f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_26 VNB N_VGND_c_427_n 0.00281836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_428_n 0.0152294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_429_n 0.0434593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_430_n 0.00507731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_431_n 0.184413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_C1_M1005_g 0.0255531f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_32 VPB N_C1_c_59_n 0.0111003f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_33 VPB N_B2_M1002_g 0.0187873f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_34 VPB N_B2_c_84_n 0.00418691f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_35 VPB N_B1_M1000_g 0.0255531f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_36 VPB N_B1_c_115_n 0.0048989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A1_M1006_g 0.0252293f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_38 VPB N_A1_c_157_n 0.00630163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A2_M1007_g 0.0227111f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_40 VPB N_A2_c_194_n 0.00412822f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_41 VPB N_A2_c_195_n 7.95285e-19 $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_42 VPB N_Y_c_231_n 0.00227642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_Y_c_232_n 0.0223637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_Y_c_233_n 0.00803945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB Y 0.00947859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_109_297#_c_327_n 0.00255716f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_47 VPB N_A_193_297#_c_349_n 0.00782532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_193_297#_c_350_n 4.02524e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_378_n 0.00589481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_379_n 0.0115529f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_51 VPB N_VPWR_c_380_n 0.0288934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_381_n 0.0480855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_382_n 0.0146253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_383_n 0.00507404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_377_n 0.0475114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 N_C1_M1005_g N_B2_M1002_g 0.0283323f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_57 N_C1_c_59_n N_B2_c_84_n 0.0222415f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_58 C1 N_B2_c_85_n 0.0162774f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_59 N_C1_c_59_n N_B2_c_85_n 0.00157241f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_60 N_C1_c_57_n N_B2_c_86_n 0.019333f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_61 N_C1_c_57_n N_Y_c_226_n 0.0141809f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_62 C1 N_Y_c_226_n 0.00631464f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_63 N_C1_c_59_n N_Y_c_226_n 0.0012291f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_64 C1 N_Y_c_227_n 0.0143329f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_65 N_C1_c_59_n N_Y_c_227_n 0.00447564f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_66 C1 N_Y_c_231_n 0.0139774f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_67 N_C1_c_59_n N_Y_c_231_n 0.00415326f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_68 N_C1_M1005_g N_Y_c_232_n 0.0138373f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 C1 N_Y_c_232_n 0.00631482f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_70 N_C1_c_59_n N_Y_c_232_n 0.00117204f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_71 N_C1_M1005_g N_A_109_297#_c_328_n 0.00589212f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_72 N_C1_M1005_g N_A_109_297#_c_329_n 0.00211624f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_73 N_C1_M1005_g N_VPWR_c_381_n 0.00539841f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_74 N_C1_M1005_g N_VPWR_c_377_n 0.0105687f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_75 N_C1_c_57_n N_VGND_c_425_n 0.00955426f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_76 N_C1_c_57_n N_VGND_c_428_n 0.00350562f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_77 N_C1_c_57_n N_VGND_c_431_n 0.00517665f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B2_M1002_g N_B1_M1000_g 0.0445512f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_79 N_B2_c_84_n B1 3.80321e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B2_c_84_n B1 6.76372e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B2_c_85_n B1 0.0183385f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B2_c_84_n N_B1_c_115_n 0.0219687f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B2_c_85_n N_B1_c_115_n 7.0101e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B2_c_86_n N_B1_c_116_n 0.0516652f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B2_c_84_n N_Y_c_226_n 0.00319406f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B2_c_85_n N_Y_c_226_n 0.0320614f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B2_c_86_n N_Y_c_226_n 0.0120179f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B2_M1002_g N_Y_c_232_n 0.0125579f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_89 N_B2_c_84_n N_Y_c_232_n 0.00304642f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B2_c_85_n N_Y_c_232_n 0.0320618f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B2_M1002_g N_A_109_297#_c_330_n 0.00984328f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B2_M1002_g N_VPWR_c_381_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 N_B2_M1002_g N_VPWR_c_377_n 0.00528062f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_94 N_B2_c_86_n N_VGND_c_425_n 0.00315422f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B2_c_86_n N_VGND_c_429_n 0.00439206f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B2_c_86_n N_VGND_c_431_n 0.00597996f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_97 B1 A1 0.0242987f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_98 N_B1_c_115_n A1 2.24093e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_99 B1 A1 0.0136402f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_100 N_B1_c_115_n A1 6.14088e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_101 B1 N_A1_c_157_n 3.07641e-19 $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_102 B1 N_A1_c_157_n 8.63992e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B1_c_115_n N_A1_c_157_n 0.00835431f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_104 B1 N_A1_c_158_n 0.00140229f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_105 B1 N_Y_M1004_d 0.0036585f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_106 B1 N_Y_c_226_n 0.00758187f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_107 B1 N_Y_c_226_n 8.53788e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B1_c_116_n N_Y_c_226_n 0.00141492f $X=1.382 $Y=0.995 $X2=0 $Y2=0
cc_109 B1 N_Y_c_228_n 0.0194133f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_110 B1 N_Y_c_228_n 0.00433948f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B1_c_115_n N_Y_c_228_n 3.80467e-19 $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B1_c_116_n N_Y_c_228_n 0.0087337f $X=1.382 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B1_c_116_n N_Y_c_259_n 0.00155357f $X=1.382 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B1_M1000_g N_Y_c_232_n 0.0124265f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_115 B1 N_Y_c_232_n 0.0342605f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B1_c_115_n N_Y_c_232_n 0.00340764f $X=1.39 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B1_M1000_g N_A_109_297#_c_327_n 0.00188941f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_B1_M1000_g N_A_109_297#_c_330_n 0.00679304f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_B1_M1000_g N_A_193_297#_c_349_n 0.0137052f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B1_M1000_g N_A_193_297#_c_352_n 0.00325589f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_B1_M1000_g N_VPWR_c_378_n 0.00236436f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_M1000_g N_VPWR_c_381_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_M1000_g N_VPWR_c_377_n 0.00657948f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_c_116_n N_VGND_c_429_n 0.00357877f $X=1.382 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B1_c_116_n N_VGND_c_431_n 0.00643093f $X=1.382 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A1_M1006_g N_A2_M1007_g 0.024119f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_127 A1 N_A2_c_194_n 2.14944e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_128 N_A1_c_157_n N_A2_c_194_n 0.0206359f $X=2.11 $Y=1.16 $X2=0 $Y2=0
cc_129 A1 N_A2_c_195_n 0.00428688f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_130 A1 N_A2_c_195_n 0.0148854f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_131 N_A1_c_157_n N_A2_c_195_n 0.00279312f $X=2.11 $Y=1.16 $X2=0 $Y2=0
cc_132 A1 N_A2_c_196_n 9.30735e-19 $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_133 N_A1_c_158_n N_A2_c_196_n 0.0328126f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_134 A1 N_Y_M1003_s 0.00463034f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_135 A1 N_Y_c_228_n 0.0153116f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_136 A1 N_Y_c_228_n 0.00194388f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A1_c_157_n N_Y_c_228_n 6.52469e-19 $X=2.11 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A1_c_158_n N_Y_c_228_n 0.0119735f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_M1006_g N_Y_c_268_n 0.00387315f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_140 A1 N_Y_c_232_n 0.0253905f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A1_c_157_n N_Y_c_232_n 0.00469821f $X=2.11 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A1_M1006_g N_Y_c_271_n 0.0118949f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A1_M1006_g N_A_193_297#_c_353_n 0.0132419f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A1_M1006_g N_A_193_297#_c_350_n 0.0016383f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A1_M1006_g N_VPWR_c_378_n 0.00836739f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A1_M1006_g N_VPWR_c_382_n 0.00343969f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A1_M1006_g N_VPWR_c_377_n 0.00413318f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A1_c_158_n N_VGND_c_427_n 0.00126016f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A1_c_158_n N_VGND_c_429_n 0.00357877f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A1_c_158_n N_VGND_c_431_n 0.00666658f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A2_M1007_g N_Y_c_268_n 0.0170474f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A2_c_194_n N_Y_c_268_n 0.0020049f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A2_c_195_n N_Y_c_268_n 0.018938f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A2_c_195_n N_Y_c_275_n 0.0108027f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A2_c_196_n N_Y_c_275_n 0.0131626f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_c_194_n N_Y_c_277_n 0.00102097f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_195_n N_Y_c_277_n 0.00891746f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A2_M1007_g Y 0.00566597f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A2_c_194_n Y 0.00760128f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A2_c_195_n Y 0.0249027f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A2_c_196_n Y 0.00609508f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_M1007_g N_VPWR_c_378_n 5.27646e-19 $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A2_M1007_g N_VPWR_c_380_n 0.00338373f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A2_M1007_g N_VPWR_c_382_n 0.00585385f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A2_M1007_g N_VPWR_c_377_n 0.0115551f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A2_c_196_n N_VGND_c_427_n 0.0091689f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_c_196_n N_VGND_c_429_n 0.00341689f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_c_196_n N_VGND_c_431_n 0.00414154f $X=2.67 $Y=0.995 $X2=0 $Y2=0
cc_169 N_Y_c_232_n N_A_109_297#_M1005_d 0.00165831f $X=2.15 $Y=1.56 $X2=-0.19
+ $Y2=-0.24
cc_170 N_Y_c_232_n N_A_109_297#_M1000_d 0.00277869f $X=2.15 $Y=1.56 $X2=0 $Y2=0
cc_171 N_Y_c_232_n N_A_109_297#_c_328_n 0.0148409f $X=2.15 $Y=1.56 $X2=0 $Y2=0
cc_172 N_Y_c_232_n N_A_109_297#_c_330_n 0.00321995f $X=2.15 $Y=1.56 $X2=0 $Y2=0
cc_173 N_Y_c_232_n N_A_193_297#_M1002_d 0.00166235f $X=2.15 $Y=1.56 $X2=-0.19
+ $Y2=-0.24
cc_174 N_Y_c_268_n N_A_193_297#_M1006_d 0.00480277f $X=2.925 $Y=1.58 $X2=0 $Y2=0
cc_175 N_Y_c_232_n N_A_193_297#_c_353_n 0.00583797f $X=2.15 $Y=1.56 $X2=0 $Y2=0
cc_176 N_Y_c_271_n N_A_193_297#_c_353_n 0.010406f $X=2.3 $Y=1.56 $X2=0 $Y2=0
cc_177 N_Y_c_268_n N_A_193_297#_c_359_n 0.0154429f $X=2.925 $Y=1.58 $X2=0 $Y2=0
cc_178 N_Y_c_232_n N_A_193_297#_c_352_n 0.0666481f $X=2.15 $Y=1.56 $X2=0 $Y2=0
cc_179 N_Y_c_232_n N_VPWR_M1006_s 0.00287335f $X=2.15 $Y=1.56 $X2=-0.19
+ $Y2=-0.24
cc_180 N_Y_c_268_n N_VPWR_M1007_d 0.00275678f $X=2.925 $Y=1.58 $X2=0 $Y2=0
cc_181 N_Y_c_233_n N_VPWR_M1007_d 0.00310605f $X=3.03 $Y=1.495 $X2=0 $Y2=0
cc_182 N_Y_c_268_n N_VPWR_c_380_n 0.00608658f $X=2.925 $Y=1.58 $X2=0 $Y2=0
cc_183 N_Y_c_233_n N_VPWR_c_380_n 0.0154232f $X=3.03 $Y=1.495 $X2=0 $Y2=0
cc_184 N_Y_c_298_p N_VPWR_c_381_n 0.0116048f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_185 N_Y_M1005_s N_VPWR_c_377_n 0.00525232f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_186 N_Y_c_298_p N_VPWR_c_377_n 0.00646998f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_187 N_Y_c_226_n N_VGND_M1008_d 0.00219123f $X=1.065 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_188 N_Y_c_275_n N_VGND_M1001_d 0.00263626f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_189 N_Y_c_229_n N_VGND_M1001_d 0.00291499f $X=3.03 $Y=0.825 $X2=0 $Y2=0
cc_190 Y N_VGND_M1001_d 0.00109932f $X=3.015 $Y=0.85 $X2=0 $Y2=0
cc_191 N_Y_c_226_n N_VGND_c_425_n 0.0186461f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_192 N_Y_c_229_n N_VGND_c_426_n 0.00107004f $X=3.03 $Y=0.825 $X2=0 $Y2=0
cc_193 N_Y_c_275_n N_VGND_c_427_n 0.00876529f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_194 N_Y_c_229_n N_VGND_c_427_n 0.0130592f $X=3.03 $Y=0.825 $X2=0 $Y2=0
cc_195 N_Y_c_309_p N_VGND_c_428_n 0.0119176f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_196 N_Y_c_226_n N_VGND_c_428_n 0.00193763f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_197 N_Y_c_226_n N_VGND_c_429_n 0.00248756f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_198 N_Y_c_228_n N_VGND_c_429_n 0.082677f $X=2.38 $Y=0.38 $X2=0 $Y2=0
cc_199 N_Y_c_259_n N_VGND_c_429_n 0.00952712f $X=1.235 $Y=0.38 $X2=0 $Y2=0
cc_200 N_Y_c_275_n N_VGND_c_429_n 0.0023303f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_201 N_Y_M1008_s N_VGND_c_431_n 0.00359898f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_202 N_Y_M1004_d N_VGND_c_431_n 0.00209344f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_203 N_Y_M1003_s N_VGND_c_431_n 0.00209344f $X=1.915 $Y=0.235 $X2=0 $Y2=0
cc_204 N_Y_c_309_p N_VGND_c_431_n 0.00665463f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_205 N_Y_c_226_n N_VGND_c_431_n 0.0101058f $X=1.065 $Y=0.82 $X2=0 $Y2=0
cc_206 N_Y_c_228_n N_VGND_c_431_n 0.0491463f $X=2.38 $Y=0.38 $X2=0 $Y2=0
cc_207 N_Y_c_259_n N_VGND_c_431_n 0.00653924f $X=1.235 $Y=0.38 $X2=0 $Y2=0
cc_208 N_Y_c_275_n N_VGND_c_431_n 0.0049037f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_209 N_Y_c_229_n N_VGND_c_431_n 0.00242556f $X=3.03 $Y=0.825 $X2=0 $Y2=0
cc_210 N_Y_c_259_n A_204_47# 9.86369e-19 $X=1.235 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_211 N_Y_c_228_n A_465_47# 0.00266519f $X=2.38 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_212 N_Y_c_277_n A_465_47# 0.00330503f $X=2.58 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_213 N_A_109_297#_c_330_n N_A_193_297#_M1002_d 0.00312752f $X=1.355 $Y=2.36
+ $X2=-0.19 $Y2=1.305
cc_214 N_A_109_297#_M1000_d N_A_193_297#_c_349_n 0.00548815f $X=1.385 $Y=1.485
+ $X2=0 $Y2=0
cc_215 N_A_109_297#_c_327_n N_A_193_297#_c_349_n 0.0164139f $X=1.52 $Y=2.34
+ $X2=0 $Y2=0
cc_216 N_A_109_297#_c_330_n N_A_193_297#_c_349_n 0.00527315f $X=1.355 $Y=2.36
+ $X2=0 $Y2=0
cc_217 N_A_109_297#_c_330_n N_A_193_297#_c_352_n 0.0114974f $X=1.355 $Y=2.36
+ $X2=0 $Y2=0
cc_218 N_A_109_297#_c_327_n N_VPWR_c_378_n 0.0168338f $X=1.52 $Y=2.34 $X2=0
+ $Y2=0
cc_219 N_A_109_297#_c_329_n N_VPWR_c_381_n 0.0152068f $X=0.765 $Y=2.38 $X2=0
+ $Y2=0
cc_220 N_A_109_297#_c_330_n N_VPWR_c_381_n 0.0517525f $X=1.355 $Y=2.36 $X2=0
+ $Y2=0
cc_221 N_A_109_297#_M1005_d N_VPWR_c_377_n 0.00215206f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_222 N_A_109_297#_M1000_d N_VPWR_c_377_n 0.00209344f $X=1.385 $Y=1.485 $X2=0
+ $Y2=0
cc_223 N_A_109_297#_c_329_n N_VPWR_c_377_n 0.00940996f $X=0.765 $Y=2.38 $X2=0
+ $Y2=0
cc_224 N_A_109_297#_c_330_n N_VPWR_c_377_n 0.0328097f $X=1.355 $Y=2.36 $X2=0
+ $Y2=0
cc_225 N_A_193_297#_c_353_n N_VPWR_M1006_s 0.00191164f $X=2.375 $Y=1.94
+ $X2=-0.19 $Y2=1.305
cc_226 N_A_193_297#_c_350_n N_VPWR_M1006_s 0.00389374f $X=2.025 $Y=1.92
+ $X2=-0.19 $Y2=1.305
cc_227 N_A_193_297#_c_349_n N_VPWR_c_378_n 0.0212138f $X=1.9 $Y=1.92 $X2=0 $Y2=0
cc_228 N_A_193_297#_c_349_n N_VPWR_c_381_n 0.00327883f $X=1.9 $Y=1.92 $X2=0
+ $Y2=0
cc_229 N_A_193_297#_c_353_n N_VPWR_c_382_n 0.00224243f $X=2.375 $Y=1.94 $X2=0
+ $Y2=0
cc_230 N_A_193_297#_c_371_p N_VPWR_c_382_n 0.0153787f $X=2.46 $Y=2.3 $X2=0 $Y2=0
cc_231 N_A_193_297#_M1002_d N_VPWR_c_377_n 0.00216833f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_193_297#_M1006_d N_VPWR_c_377_n 0.00280591f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_A_193_297#_c_349_n N_VPWR_c_377_n 0.00775536f $X=1.9 $Y=1.92 $X2=0
+ $Y2=0
cc_234 N_A_193_297#_c_353_n N_VPWR_c_377_n 0.00408444f $X=2.375 $Y=1.94 $X2=0
+ $Y2=0
cc_235 N_A_193_297#_c_371_p N_VPWR_c_377_n 0.0095318f $X=2.46 $Y=2.3 $X2=0 $Y2=0
cc_236 N_VGND_c_431_n A_204_47# 0.00195685f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_237 N_VGND_c_431_n A_465_47# 0.00264607f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

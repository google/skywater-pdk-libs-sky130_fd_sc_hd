* File: sky130_fd_sc_hd__dfbbn_1.spice.pex
* Created: Thu Aug 27 14:13:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFBBN_1%CLK_N 4 5 7 8 10 13 17 19 20 24 26
c45 13 0 2.71124e-20 $X=0.47 $Y=0.805
r46 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r47 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r48 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r49 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r50 15 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=1.665
+ $X2=0.47 $Y2=1.665
r51 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.47 $Y2=0.805
r52 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r53 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r54 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r55 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r56 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r57 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r58 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r59 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_27_47# 1 2 9 13 17 19 20 23 26 27 29 32 36
+ 40 41 42 46 47 51 52 55 58 59 61 62 63 66 70 74 81 84 85 99
c262 99 0 8.91099e-20 $X=6.295 $Y=1.182
c263 61 0 9.6376e-20 $X=3.027 $Y=1.12
c264 47 0 1.06217e-19 $X=6.32 $Y=0.87
c265 46 0 1.43345e-19 $X=6.32 $Y=0.87
c266 17 0 4.43992e-20 $X=2.29 $Y=2.275
r267 99 100 19.6811 $w=2.12e-07 $l=3.42e-07 $layer=LI1_cond $X=6.295 $Y=1.182
+ $X2=6.637 $Y2=1.182
r268 84 87 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=0.93
+ $X2=2.89 $Y2=1.095
r269 84 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=0.93
+ $X2=2.89 $Y2=0.765
r270 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.89
+ $Y=0.93 $X2=2.89 $Y2=0.93
r271 78 81 31.1043 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=0.75 $Y=1.235
+ $X2=0.89 $Y2=1.235
r272 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.235 $X2=0.75 $Y2=1.235
r273 75 99 4.89151 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=1.182
+ $X2=6.295 $Y2=1.182
r274 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=1.19
+ $X2=6.21 $Y2=1.19
r275 70 72 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.965
r276 70 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.85
r277 66 79 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.725 $Y=0.85
+ $X2=0.725 $Y2=1.235
r278 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=0.85
+ $X2=0.695 $Y2=0.85
r279 62 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.065 $Y=1.19
+ $X2=6.21 $Y2=1.19
r280 62 63 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=6.065 $Y=1.19
+ $X2=3.135 $Y2=1.19
r281 61 63 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.135 $Y2=1.19
r282 61 72 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.027 $Y2=0.965
r283 59 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=0.85
+ $X2=0.695 $Y2=0.85
r284 58 70 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=2.99 $Y2=0.85
r285 58 59 2.48143 $w=1.4e-07 $l=2.005e-06 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=0.84 $Y2=0.85
r286 57 79 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r287 56 66 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=0.85
r288 52 92 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.655 $Y=1.74
+ $X2=6.655 $Y2=1.875
r289 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.655
+ $Y=1.74 $X2=6.655 $Y2=1.74
r290 49 100 0.949179 $w=2.05e-07 $l=1.23e-07 $layer=LI1_cond $X=6.637 $Y=1.305
+ $X2=6.637 $Y2=1.182
r291 49 51 23.5344 $w=2.03e-07 $l=4.35e-07 $layer=LI1_cond $X=6.637 $Y=1.305
+ $X2=6.637 $Y2=1.74
r292 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.32
+ $Y=0.87 $X2=6.32 $Y2=0.87
r293 44 99 0.489344 $w=2.2e-07 $l=1.22e-07 $layer=LI1_cond $X=6.295 $Y=1.06
+ $X2=6.295 $Y2=1.182
r294 44 46 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=6.295 $Y=1.06
+ $X2=6.295 $Y2=0.87
r295 43 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r296 42 57 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.795
r297 42 43 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r298 40 56 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r299 40 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r300 34 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r301 34 36 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r302 32 92 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.625 $Y=2.275
+ $X2=6.625 $Y2=1.875
r303 27 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.32 $Y=0.705
+ $X2=6.32 $Y2=0.87
r304 27 29 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.32 $Y=0.705
+ $X2=6.32 $Y2=0.415
r305 26 87 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.83 $Y=1.245
+ $X2=2.83 $Y2=1.095
r306 23 86 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.83 $Y=0.415
+ $X2=2.83 $Y2=0.765
r307 19 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.755 $Y=1.32
+ $X2=2.83 $Y2=1.245
r308 19 20 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.755 $Y=1.32
+ $X2=2.365 $Y2=1.32
r309 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.29 $Y=1.395
+ $X2=2.365 $Y2=1.32
r310 15 17 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.29 $Y=1.395
+ $X2=2.29 $Y2=2.275
r311 11 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r312 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r313 7 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r314 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r315 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r316 1 36 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%D 3 7 9 10 14 15
c41 7 0 1.80024e-19 $X=1.83 $Y=2.275
r42 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.17 $X2=1.83 $Y2=1.17
r43 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.95 $Y=1.19 $X2=1.95
+ $Y2=1.53
r44 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.95 $Y=1.19 $X2=1.95
+ $Y2=1.17
r45 5 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.335
+ $X2=1.83 $Y2=1.17
r46 5 7 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.83 $Y=1.335 $X2=1.83
+ $Y2=2.275
r47 1 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.005
+ $X2=1.83 $Y2=1.17
r48 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.83 $Y=1.005 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_193_47# 1 2 7 9 12 18 20 21 24 28 29 31 32
+ 33 34 43 51 52 56 57 58 61
c202 57 0 9.11072e-20 $X=6.145 $Y=1.74
c203 29 0 2.53399e-19 $X=2.41 $Y=0.87
c204 28 0 1.80024e-19 $X=2.41 $Y=0.87
c205 18 0 3.84972e-20 $X=6.205 $Y=2.275
r206 56 59 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.145 $Y=1.74
+ $X2=6.145 $Y2=1.905
r207 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.145 $Y=1.74
+ $X2=6.145 $Y2=1.575
r208 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.145
+ $Y=1.74 $X2=6.145 $Y2=1.74
r209 51 54 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.74 $Y=1.74
+ $X2=2.74 $Y2=1.875
r210 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.74 $X2=2.74 $Y2=1.74
r211 43 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=1.87
+ $X2=6.21 $Y2=1.87
r212 41 52 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.74 $Y2=1.765
r213 41 69 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.435 $Y2=1.765
r214 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=1.87
r215 37 61 71.2419 $w=2.18e-07 $l=1.36e-06 $layer=LI1_cond $X=1.125 $Y=1.87
+ $X2=1.125 $Y2=0.51
r216 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.87
+ $X2=1.15 $Y2=1.87
r217 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.87
+ $X2=2.53 $Y2=1.87
r218 33 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.065 $Y=1.87
+ $X2=6.21 $Y2=1.87
r219 33 34 4.19554 $w=1.4e-07 $l=3.39e-06 $layer=MET1_cond $X=6.065 $Y=1.87
+ $X2=2.675 $Y2=1.87
r220 32 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.87
+ $X2=1.15 $Y2=1.87
r221 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=2.53 $Y2=1.87
r222 31 32 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=1.295 $Y2=1.87
r223 29 46 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=2.41 $Y=0.87
+ $X2=2.305 $Y2=0.87
r224 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=0.87 $X2=2.41 $Y2=0.87
r225 26 69 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.435 $Y=1.575
+ $X2=2.435 $Y2=1.765
r226 26 28 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.435 $Y=1.575
+ $X2=2.435 $Y2=0.87
r227 22 24 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=6.74 $Y=1.245
+ $X2=6.74 $Y2=0.415
r228 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.665 $Y=1.32
+ $X2=6.74 $Y2=1.245
r229 20 21 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.665 $Y=1.32
+ $X2=6.28 $Y2=1.32
r230 18 59 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.205 $Y=2.275
+ $X2=6.205 $Y2=1.905
r231 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.205 $Y=1.395
+ $X2=6.28 $Y2=1.32
r232 14 58 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.205 $Y=1.395
+ $X2=6.205 $Y2=1.575
r233 12 54 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.71 $Y=2.275
+ $X2=2.71 $Y2=1.875
r234 7 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r235 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r236 2 37 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r237 1 61 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_647_21# 1 2 9 13 17 19 21 22 26 28 30 31
+ 32 35 36 41 45 49
c147 49 0 1.43345e-19 $X=5.66 $Y=1.15
r148 49 56 10.4783 $w=2.76e-07 $l=6e-08 $layer=POLY_cond $X=5.66 $Y=1.15
+ $X2=5.72 $Y2=1.15
r149 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.66
+ $Y=1.15 $X2=5.66 $Y2=1.15
r150 45 48 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.66 $Y=0.98
+ $X2=5.66 $Y2=1.15
r151 43 44 14.1313 $w=2.59e-07 $l=3e-07 $layer=LI1_cond $X=4.57 $Y=0.68 $X2=4.57
+ $Y2=0.98
r152 36 53 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.74
+ $X2=3.395 $Y2=1.905
r153 36 52 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.74
+ $X2=3.395 $Y2=1.575
r154 35 38 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.46 $Y=1.74
+ $X2=3.46 $Y2=1.91
r155 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.74 $X2=3.42 $Y2=1.74
r156 33 44 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=0.98
+ $X2=4.57 $Y2=0.98
r157 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=0.98
+ $X2=5.66 $Y2=0.98
r158 32 33 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.495 $Y=0.98
+ $X2=4.735 $Y2=0.98
r159 30 44 5.44435 $w=2.59e-07 $l=9.88686e-08 $layer=LI1_cond $X=4.6 $Y=1.065
+ $X2=4.57 $Y2=0.98
r160 30 31 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.6 $Y=1.065
+ $X2=4.6 $Y2=1.785
r161 29 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=1.91
+ $X2=4.17 $Y2=1.91
r162 28 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.515 $Y=1.91
+ $X2=4.6 $Y2=1.785
r163 28 29 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=4.515 $Y=1.91
+ $X2=4.255 $Y2=1.91
r164 24 41 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.17 $Y=2.035
+ $X2=4.17 $Y2=1.91
r165 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.17 $Y=2.035
+ $X2=4.17 $Y2=2.21
r166 23 38 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.585 $Y=1.91
+ $X2=3.46 $Y2=1.91
r167 22 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=1.91
+ $X2=4.17 $Y2=1.91
r168 22 23 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=4.085 $Y=1.91
+ $X2=3.585 $Y2=1.91
r169 19 56 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.72 $Y=0.985
+ $X2=5.72 $Y2=1.15
r170 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.72 $Y=0.985
+ $X2=5.72 $Y2=0.555
r171 15 49 30.5616 $w=2.76e-07 $l=2.43926e-07 $layer=POLY_cond $X=5.485 $Y=1.315
+ $X2=5.66 $Y2=1.15
r172 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.485 $Y=1.315
+ $X2=5.485 $Y2=2.065
r173 13 53 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.31 $Y=2.275
+ $X2=3.31 $Y2=1.905
r174 9 52 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.31 $Y=0.445
+ $X2=3.31 $Y2=1.575
r175 2 41 600 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=2.065 $X2=4.17 $Y2=1.87
r176 2 26 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=2.065 $X2=4.17 $Y2=2.21
r177 1 43 182 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_NDIFF $count=1 $X=4.435
+ $Y=0.235 $X2=4.57 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%SET_B 1 3 7 11 13 15 17 19 20 26 27
c132 19 0 1.0411e-19 $X=7.515 $Y=0.85
c133 15 0 1.0852e-19 $X=7.755 $Y=2.275
c134 11 0 9.90542e-21 $X=7.7 $Y=0.445
r135 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.64
+ $Y=0.98 $X2=7.64 $Y2=0.98
r136 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.66 $Y=0.85
+ $X2=7.66 $Y2=0.85
r137 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=0.85
+ $X2=3.91 $Y2=0.85
r138 19 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.515 $Y=0.85
+ $X2=7.66 $Y2=0.85
r139 19 20 4.28217 $w=1.4e-07 $l=3.46e-06 $layer=MET1_cond $X=7.515 $Y=0.85
+ $X2=4.055 $Y2=0.85
r140 17 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.75
+ $Y=0.98 $X2=3.75 $Y2=0.98
r141 17 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0.85
+ $X2=3.91 $Y2=0.85
r142 13 33 44.3765 $w=2.92e-07 $l=2.4e-07 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.667 $Y2=0.98
r143 13 15 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.755 $Y2=2.275
r144 9 33 38.5991 $w=2.92e-07 $l=1.80748e-07 $layer=POLY_cond $X=7.7 $Y=0.815
+ $X2=7.667 $Y2=0.98
r145 9 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.7 $Y=0.815 $X2=7.7
+ $Y2=0.445
r146 5 30 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.88 $Y=0.815
+ $X2=3.785 $Y2=0.98
r147 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.88 $Y=0.815
+ $X2=3.88 $Y2=0.445
r148 1 30 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.84 $Y=1.145
+ $X2=3.785 $Y2=0.98
r149 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.84 $Y=1.145
+ $X2=3.84 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_473_413# 1 2 9 13 15 19 24 26 27 32 35
c105 35 0 1.0411e-19 $X=4.26 $Y=1.32
c106 32 0 4.43992e-20 $X=3.415 $Y=1.3
r107 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.29 $Y=1.32
+ $X2=4.29 $Y2=1.485
r108 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.29 $Y=1.32
+ $X2=4.29 $Y2=1.155
r109 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.26
+ $Y=1.32 $X2=4.26 $Y2=1.32
r110 31 32 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=1.3
+ $X2=3.415 $Y2=1.3
r111 29 31 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=3.08 $Y=1.3
+ $X2=3.33 $Y2=1.3
r112 27 34 8.9562 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=1.32
+ $X2=4.26 $Y2=1.32
r113 27 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.095 $Y=1.32
+ $X2=3.415 $Y2=1.32
r114 26 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.33 $Y=1.195
+ $X2=3.33 $Y2=1.3
r115 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.33 $Y=0.465
+ $X2=3.33 $Y2=1.195
r116 23 29 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.08 $Y=1.405
+ $X2=3.08 $Y2=1.3
r117 23 24 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.08 $Y=1.405
+ $X2=3.08 $Y2=2.25
r118 19 25 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.245 $Y=0.365
+ $X2=3.33 $Y2=0.465
r119 19 21 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.245 $Y=0.365
+ $X2=2.565 $Y2=0.365
r120 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=2.335
+ $X2=3.08 $Y2=2.25
r121 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.995 $Y=2.335
+ $X2=2.5 $Y2=2.335
r122 13 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.38 $Y=2.065
+ $X2=4.38 $Y2=1.485
r123 9 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.36 $Y=0.555 $X2=4.36
+ $Y2=1.155
r124 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=2.065 $X2=2.5 $Y2=2.335
r125 1 21 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.565 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_941_21# 1 2 9 13 17 21 25 26 27 29 33 36
+ 37 42 43 45 46 49 52 64 65
c168 45 0 2.58372e-20 $X=8.795 $Y=1.53
c169 29 0 1.52865e-19 $X=9.375 $Y=1.66
c170 21 0 6.55176e-20 $X=8.66 $Y=0.555
r171 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.855
+ $Y=1.32 $X2=8.855 $Y2=1.32
r172 62 64 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=8.66 $Y=1.32
+ $X2=8.855 $Y2=1.32
r173 60 62 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.645 $Y=1.32
+ $X2=8.66 $Y2=1.32
r174 55 57 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.78 $Y=1.32 $X2=4.8
+ $Y2=1.32
r175 53 65 8.49168 $w=2.83e-07 $l=2.1e-07 $layer=LI1_cond $X=8.912 $Y=1.53
+ $X2=8.912 $Y2=1.32
r176 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.94 $Y=1.53
+ $X2=8.94 $Y2=1.53
r177 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=1.53
+ $X2=5.75 $Y2=1.53
r178 46 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.895 $Y=1.53
+ $X2=5.75 $Y2=1.53
r179 45 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.795 $Y=1.53
+ $X2=8.94 $Y2=1.53
r180 45 46 3.5891 $w=1.4e-07 $l=2.9e-06 $layer=MET1_cond $X=8.795 $Y=1.53
+ $X2=5.895 $Y2=1.53
r181 44 53 1.81965 $w=2.83e-07 $l=4.5e-08 $layer=LI1_cond $X=8.912 $Y=1.575
+ $X2=8.912 $Y2=1.53
r182 42 65 2.74969 $w=2.83e-07 $l=6.8e-08 $layer=LI1_cond $X=8.912 $Y=1.252
+ $X2=8.912 $Y2=1.32
r183 42 43 6.37134 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=8.912 $Y=1.252
+ $X2=8.912 $Y2=1.11
r184 40 49 27.1304 $w=2.38e-07 $l=5.65e-07 $layer=LI1_cond $X=5.185 $Y=1.535
+ $X2=5.75 $Y2=1.535
r185 39 40 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.02 $Y=1.535
+ $X2=5.185 $Y2=1.535
r186 37 57 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.02 $Y=1.32
+ $X2=4.8 $Y2=1.32
r187 36 39 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.02 $Y=1.32
+ $X2=5.02 $Y2=1.535
r188 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.02
+ $Y=1.32 $X2=5.02 $Y2=1.32
r189 31 33 17.1645 $w=2.08e-07 $l=3.25e-07 $layer=LI1_cond $X=9.37 $Y=0.755
+ $X2=9.37 $Y2=0.43
r190 27 44 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=9.055 $Y=1.66
+ $X2=8.912 $Y2=1.575
r191 27 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.055 $Y=1.66
+ $X2=9.375 $Y2=1.66
r192 25 31 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.265 $Y=0.84
+ $X2=9.37 $Y2=0.755
r193 25 26 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.265 $Y=0.84
+ $X2=9.055 $Y2=0.84
r194 23 26 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=8.945 $Y=0.925
+ $X2=9.055 $Y2=0.84
r195 23 43 9.691 $w=2.18e-07 $l=1.85e-07 $layer=LI1_cond $X=8.945 $Y=0.925
+ $X2=8.945 $Y2=1.11
r196 19 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.66 $Y=1.155
+ $X2=8.66 $Y2=1.32
r197 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.66 $Y=1.155 $X2=8.66
+ $Y2=0.555
r198 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.485
+ $X2=8.645 $Y2=1.32
r199 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.645 $Y=1.485
+ $X2=8.645 $Y2=2.065
r200 11 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.8 $Y=1.485
+ $X2=4.8 $Y2=1.32
r201 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.8 $Y=1.485
+ $X2=4.8 $Y2=2.065
r202 7 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.78 $Y=1.155
+ $X2=4.78 $Y2=1.32
r203 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.78 $Y=1.155 $X2=4.78
+ $Y2=0.555
r204 2 29 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=9.25
+ $Y=1.505 $X2=9.375 $Y2=1.66
r205 1 33 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=9.265
+ $Y=0.235 $X2=9.39 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_1415_315# 1 2 9 13 15 17 20 22 23 25 27 28
+ 30 31 33 36 38 41 45 46 48 49 52 54 57 58 61 62 64 66 70
c195 20 0 1.52865e-19 $X=10.075 $Y=1.985
c196 13 0 8.91099e-20 $X=7.215 $Y=0.445
r197 73 75 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.15 $Y=1.74
+ $X2=7.215 $Y2=1.74
r198 71 79 5.15902 $w=3.27e-07 $l=3.5e-08 $layer=POLY_cond $X=10.04 $Y=1.16
+ $X2=10.075 $Y2=1.16
r199 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.04
+ $Y=1.16 $X2=10.04 $Y2=1.16
r200 67 70 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=9.945 $Y=1.16
+ $X2=10.04 $Y2=1.16
r201 64 65 4.61047 $w=1.72e-07 $l=6.5e-08 $layer=LI1_cond $X=8.45 $Y=0.752
+ $X2=8.515 $Y2=0.752
r202 60 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.945 $Y=1.325
+ $X2=9.945 $Y2=1.16
r203 60 61 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.945 $Y=1.325
+ $X2=9.945 $Y2=1.915
r204 59 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.6 $Y=2 $X2=8.515
+ $Y2=2
r205 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.86 $Y=2
+ $X2=9.945 $Y2=1.915
r206 58 59 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=9.86 $Y=2 $X2=8.6
+ $Y2=2
r207 57 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.515 $Y=1.915
+ $X2=8.515 $Y2=2
r208 56 65 0.787725 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=8.515 $Y=0.84
+ $X2=8.515 $Y2=0.752
r209 56 57 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=8.515 $Y=0.84
+ $X2=8.515 $Y2=1.915
r210 55 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=2 $X2=8.025
+ $Y2=2
r211 54 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=2 $X2=8.515
+ $Y2=2
r212 54 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.43 $Y=2 $X2=8.11
+ $Y2=2
r213 50 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=2.085
+ $X2=8.025 $Y2=2
r214 50 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=2.085
+ $X2=8.025 $Y2=2.21
r215 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=2 $X2=8.025
+ $Y2=2
r216 48 49 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.94 $Y=2 $X2=7.5
+ $Y2=2
r217 46 75 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=7.335 $Y=1.74
+ $X2=7.215 $Y2=1.74
r218 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.335
+ $Y=1.74 $X2=7.335 $Y2=1.74
r219 43 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.375 $Y=1.915
+ $X2=7.5 $Y2=2
r220 43 45 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=7.375 $Y=1.915
+ $X2=7.375 $Y2=1.74
r221 39 41 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=10.89 $Y=1.61
+ $X2=11.015 $Y2=1.61
r222 34 36 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=10.89 $Y=0.805
+ $X2=11.015 $Y2=0.805
r223 31 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=1.685
+ $X2=11.015 $Y2=1.61
r224 31 33 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=11.015 $Y=1.685
+ $X2=11.015 $Y2=2.085
r225 28 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=0.73
+ $X2=11.015 $Y2=0.805
r226 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.015 $Y=0.73
+ $X2=11.015 $Y2=0.445
r227 27 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.89 $Y=1.535
+ $X2=10.89 $Y2=1.61
r228 26 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.89 $Y=1.295
+ $X2=10.89 $Y2=1.16
r229 26 27 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.89 $Y=1.295
+ $X2=10.89 $Y2=1.535
r230 25 38 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.89 $Y=1.025
+ $X2=10.89 $Y2=1.16
r231 24 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.89 $Y=0.88
+ $X2=10.89 $Y2=0.805
r232 24 25 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=10.89 $Y=0.88
+ $X2=10.89 $Y2=1.025
r233 23 79 16.3472 $w=3.27e-07 $l=1e-07 $layer=POLY_cond $X=10.175 $Y=1.16
+ $X2=10.075 $Y2=1.16
r234 22 38 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=10.815 $Y=1.16
+ $X2=10.89 $Y2=1.16
r235 22 23 142.191 $w=2.7e-07 $l=6.4e-07 $layer=POLY_cond $X=10.815 $Y=1.16
+ $X2=10.175 $Y2=1.16
r236 18 79 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.075 $Y=1.325
+ $X2=10.075 $Y2=1.16
r237 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.075 $Y=1.325
+ $X2=10.075 $Y2=1.985
r238 15 79 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.075 $Y=0.995
+ $X2=10.075 $Y2=1.16
r239 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.075 $Y=0.995
+ $X2=10.075 $Y2=0.56
r240 11 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.215 $Y=1.575
+ $X2=7.215 $Y2=1.74
r241 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.215 $Y=1.575
+ $X2=7.215 $Y2=0.445
r242 7 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.15 $Y=1.905
+ $X2=7.15 $Y2=1.74
r243 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.15 $Y=1.905
+ $X2=7.15 $Y2=2.275
r244 2 52 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=7.83
+ $Y=2.065 $X2=8.025 $Y2=2.21
r245 1 64 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=8.315
+ $Y=0.235 $X2=8.45 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_1256_413# 1 2 9 13 15 19 24 26 27 29 31 32
c112 32 0 2.15595e-19 $X=8.175 $Y=1.24
c113 31 0 1.74038e-19 $X=8.175 $Y=1.24
c114 26 0 3.84972e-20 $X=6.995 $Y=2.25
r115 32 38 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.2 $Y=1.24
+ $X2=8.2 $Y2=1.405
r116 32 37 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.2 $Y=1.24
+ $X2=8.2 $Y2=1.075
r117 31 34 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=8.15 $Y=1.24 $X2=8.15
+ $Y2=1.32
r118 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.175
+ $Y=1.24 $X2=8.175 $Y2=1.24
r119 28 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=1.32
+ $X2=6.995 $Y2=1.32
r120 27 34 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=8.04 $Y=1.32 $X2=8.15
+ $Y2=1.32
r121 27 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.04 $Y=1.32
+ $X2=7.08 $Y2=1.32
r122 25 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=1.405
+ $X2=6.995 $Y2=1.32
r123 25 26 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=6.995 $Y=1.405
+ $X2=6.995 $Y2=2.25
r124 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=1.235
+ $X2=6.995 $Y2=1.32
r125 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.995 $Y=0.465
+ $X2=6.995 $Y2=1.235
r126 19 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.91 $Y=0.365
+ $X2=6.995 $Y2=0.465
r127 19 21 21.0727 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=6.91 $Y=0.365
+ $X2=6.53 $Y2=0.365
r128 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.91 $Y=2.335
+ $X2=6.995 $Y2=2.25
r129 15 17 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.91 $Y=2.335
+ $X2=6.415 $Y2=2.335
r130 13 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.285 $Y=2.065
+ $X2=8.285 $Y2=1.405
r131 9 37 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.24 $Y=0.555
+ $X2=8.24 $Y2=1.075
r132 2 17 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=2.065 $X2=6.415 $Y2=2.335
r133 1 21 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.395
+ $Y=0.235 $X2=6.53 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%RESET_B 3 7 9 16
r39 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=9.59 $Y=1.18 $X2=9.6
+ $Y2=1.18
r40 12 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=9.4 $Y=1.18 $X2=9.59
+ $Y2=1.18
r41 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.4 $Y=1.18
+ $X2=9.4 $Y2=1.18
r42 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.6 $Y=1.015 $X2=9.6
+ $Y2=1.18
r43 5 7 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=9.6 $Y=1.015 $X2=9.6
+ $Y2=0.445
r44 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.59 $Y=1.345
+ $X2=9.59 $Y2=1.18
r45 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.59 $Y=1.345 $X2=9.59
+ $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_2136_47# 1 2 9 12 16 20 24 25 27 29
c54 27 0 1.39343e-19 $X=10.817 $Y=1.16
r55 25 30 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.422 $Y=1.16
+ $X2=11.422 $Y2=1.325
r56 25 29 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.422 $Y=1.16
+ $X2=11.422 $Y2=0.995
r57 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.41
+ $Y=1.16 $X2=11.41 $Y2=1.16
r58 22 27 1.17559 $w=3.3e-07 $l=1.58e-07 $layer=LI1_cond $X=10.975 $Y=1.16
+ $X2=10.817 $Y2=1.16
r59 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=10.975 $Y=1.16
+ $X2=11.41 $Y2=1.16
r60 18 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=10.817 $Y=1.325
+ $X2=10.817 $Y2=1.16
r61 18 20 21.4025 $w=3.13e-07 $l=5.85e-07 $layer=LI1_cond $X=10.817 $Y=1.325
+ $X2=10.817 $Y2=1.91
r62 14 27 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=10.817 $Y=0.995
+ $X2=10.817 $Y2=1.16
r63 14 16 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=10.817 $Y=0.995
+ $X2=10.817 $Y2=0.51
r64 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.49 $Y=1.985
+ $X2=11.49 $Y2=1.325
r65 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.49 $Y=0.56
+ $X2=11.49 $Y2=0.995
r66 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.68
+ $Y=1.765 $X2=10.805 $Y2=1.91
r67 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=10.68
+ $Y=0.235 $X2=10.805 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 46 47 48
+ 52 53 55 57 63 68 80 91 95 102 103 106 109 112 115 126 128
r184 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r185 124 126 9.28831 $w=5.48e-07 $l=1.4e-07 $layer=LI1_cond $X=9.89 $Y=2.53
+ $X2=10.03 $Y2=2.53
r186 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r187 122 124 0.543672 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=9.865 $Y=2.53
+ $X2=9.89 $Y2=2.53
r188 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r189 115 118 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=7.51 $Y=2.34
+ $X2=7.51 $Y2=2.72
r190 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r191 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r192 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r193 103 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r194 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r195 100 128 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.445 $Y=2.72
+ $X2=11.3 $Y2=2.72
r196 100 102 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.445 $Y=2.72
+ $X2=11.73 $Y2=2.72
r197 99 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r198 99 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=9.89 $Y2=2.72
r199 98 126 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=10.03 $Y2=2.72
r200 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r201 95 128 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.155 $Y=2.72
+ $X2=11.3 $Y2=2.72
r202 95 98 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.155 $Y=2.72
+ $X2=10.81 $Y2=2.72
r203 94 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r204 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r205 91 122 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=9.755 $Y=2.53
+ $X2=9.865 $Y2=2.53
r206 91 93 17.0713 $w=5.48e-07 $l=7.85e-07 $layer=LI1_cond $X=9.755 $Y=2.53
+ $X2=8.97 $Y2=2.53
r207 90 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r208 90 119 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=7.59 $Y2=2.72
r209 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r210 87 118 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.7 $Y=2.72
+ $X2=7.51 $Y2=2.72
r211 87 89 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=7.7 $Y=2.72
+ $X2=8.51 $Y2=2.72
r212 86 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r213 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r214 83 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r215 82 85 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=7.13 $Y2=2.72
r216 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r217 80 118 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.32 $Y=2.72
+ $X2=7.51 $Y2=2.72
r218 80 85 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.32 $Y=2.72
+ $X2=7.13 $Y2=2.72
r219 79 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r220 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r221 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r222 76 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r223 75 78 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r224 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r225 73 112 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.595 $Y2=2.72
r226 73 75 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.91 $Y2=2.72
r227 72 113 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r228 72 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r229 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r230 69 109 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.607 $Y2=2.72
r231 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r232 68 112 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.405 $Y=2.72
+ $X2=3.595 $Y2=2.72
r233 68 71 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=3.405 $Y=2.72
+ $X2=2.07 $Y2=2.72
r234 67 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r235 67 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r236 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r237 64 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r238 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r239 63 109 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.607 $Y2=2.72
r240 63 66 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.15 $Y2=2.72
r241 57 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r242 55 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r243 53 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r244 53 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r245 52 89 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=8.64 $Y=2.72
+ $X2=8.51 $Y2=2.72
r246 51 52 10.9193 $w=5.48e-07 $l=2.15e-07 $layer=LI1_cond $X=8.855 $Y=2.53
+ $X2=8.64 $Y2=2.53
r247 48 93 1.19608 $w=5.48e-07 $l=5.5e-08 $layer=LI1_cond $X=8.915 $Y=2.53
+ $X2=8.97 $Y2=2.53
r248 48 51 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=8.915 $Y=2.53
+ $X2=8.855 $Y2=2.53
r249 46 78 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=4.83 $Y2=2.72
r250 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=5.04 $Y2=2.72
r251 45 82 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=2.72
+ $X2=5.29 $Y2=2.72
r252 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=2.72
+ $X2=5.04 $Y2=2.72
r253 41 128 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.3 $Y=2.635
+ $X2=11.3 $Y2=2.72
r254 41 43 27.6189 $w=2.88e-07 $l=6.95e-07 $layer=LI1_cond $X=11.3 $Y=2.635
+ $X2=11.3 $Y2=1.94
r255 37 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=2.635
+ $X2=5.04 $Y2=2.72
r256 37 39 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.04 $Y=2.635
+ $X2=5.04 $Y2=2
r257 33 112 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=2.635
+ $X2=3.595 $Y2=2.72
r258 33 35 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=3.595 $Y=2.635
+ $X2=3.595 $Y2=2.29
r259 29 109 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.72
r260 29 31 13.4722 $w=3.53e-07 $l=4.15e-07 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.22
r261 25 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r262 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r263 8 43 300 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=2 $X=11.09
+ $Y=1.765 $X2=11.28 $Y2=1.94
r264 7 122 600 $w=1.7e-07 $l=9.29637e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.505 $X2=9.865 $Y2=2.34
r265 6 51 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.645 $X2=8.855 $Y2=2.34
r266 5 115 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=2.065 $X2=7.485 $Y2=2.34
r267 4 39 300 $w=1.7e-07 $l=4.29651e-07 $layer=licon1_PDIFF $count=2 $X=4.875
+ $Y=1.645 $X2=5.04 $Y2=2
r268 3 35 600 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=2.065 $X2=3.57 $Y2=2.29
r269 2 31 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.065 $X2=1.62 $Y2=2.22
r270 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_381_47# 1 2 8 9 10 11 12 15 19
r58 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.04 $Y=1.965
+ $X2=2.04 $Y2=2.3
r59 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r60 11 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.965
r61 11 12 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.575 $Y2=1.88
r62 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r63 9 10 22.1818 $w=1.88e-07 $l=3.8e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=1.575 $Y2=0.73
r64 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.49 $Y=1.795
+ $X2=1.575 $Y2=1.88
r65 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.49 $Y=0.825
+ $X2=1.575 $Y2=0.73
r66 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.49 $Y=0.825 $X2=1.49
+ $Y2=1.795
r67 2 19 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=2.065 $X2=2.04 $Y2=2.3
r68 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%Q_N 1 2 9 10 11 12 13 18 21
r31 18 21 2.69684 $w=2.85e-07 $l=6.3e-08 $layer=LI1_cond $X=10.342 $Y=0.573
+ $X2=10.342 $Y2=0.51
r32 12 13 15.9725 $w=2.83e-07 $l=3.95e-07 $layer=LI1_cond $X=10.342 $Y=1.815
+ $X2=10.342 $Y2=2.21
r33 11 30 6.85431 $w=2.83e-07 $l=1.31e-07 $layer=LI1_cond $X=10.342 $Y=0.584
+ $X2=10.342 $Y2=0.715
r34 11 18 0.444803 $w=2.83e-07 $l=1.1e-08 $layer=LI1_cond $X=10.342 $Y=0.584
+ $X2=10.342 $Y2=0.573
r35 11 21 0.470877 $w=2.85e-07 $l=1.1e-08 $layer=LI1_cond $X=10.342 $Y=0.499
+ $X2=10.342 $Y2=0.51
r36 10 30 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=10.395 $Y=1.63
+ $X2=10.395 $Y2=0.715
r37 9 12 1.73877 $w=2.83e-07 $l=4.3e-08 $layer=LI1_cond $X=10.342 $Y=1.772
+ $X2=10.342 $Y2=1.815
r38 9 10 7.29911 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=10.342 $Y=1.772
+ $X2=10.342 $Y2=1.63
r39 2 12 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=10.15
+ $Y=1.485 $X2=10.285 $Y2=1.815
r40 1 21 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=10.15
+ $Y=0.235 $X2=10.285 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%Q 1 2 10 11 12 13 14 15
r18 14 15 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=11.745 $Y=1.82
+ $X2=11.745 $Y2=2.21
r19 11 14 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=11.745 $Y=1.585
+ $X2=11.745 $Y2=1.82
r20 11 12 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=11.745 $Y=1.585
+ $X2=11.745 $Y2=1.455
r21 10 12 33.2727 $w=2.08e-07 $l=6.3e-07 $layer=LI1_cond $X=11.77 $Y=0.825
+ $X2=11.77 $Y2=1.455
r22 9 13 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=11.745 $Y=0.695
+ $X2=11.745 $Y2=0.51
r23 9 10 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=11.745 $Y=0.695
+ $X2=11.745 $Y2=0.825
r24 2 14 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=11.565
+ $Y=1.485 $X2=11.7 $Y2=1.82
r25 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=11.565
+ $Y=0.235 $X2=11.7 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 48 51
+ 52 54 55 57 58 59 61 63 69 93 100 107 108 111 114 117 120
c187 108 0 4.22219e-20 $X=11.73 $Y=0
c188 51 0 1.57023e-19 $X=3.585 $Y=0
r189 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r190 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r191 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r192 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r193 108 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r194 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r195 105 120 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=11.445 $Y=0
+ $X2=11.297 $Y2=0
r196 105 107 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.445 $Y=0
+ $X2=11.73 $Y2=0
r197 104 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r198 104 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=9.89 $Y2=0
r199 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r200 101 117 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=10.03 $Y=0
+ $X2=9.877 $Y2=0
r201 101 103 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=10.03 $Y=0
+ $X2=10.81 $Y2=0
r202 100 120 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=11.297 $Y2=0
r203 100 103 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=10.81 $Y2=0
r204 99 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r205 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r206 96 99 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r207 95 98 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=0 $X2=9.43
+ $Y2=0
r208 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r209 93 117 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=9.725 $Y=0
+ $X2=9.877 $Y2=0
r210 93 98 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.725 $Y=0 $X2=9.43
+ $Y2=0
r211 92 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r212 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r213 89 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=7.13 $Y2=0
r214 88 91 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=7.13
+ $Y2=0
r215 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r216 86 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r217 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r218 83 86 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r219 82 85 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r220 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r221 80 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r222 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r223 77 80 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r224 77 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r225 76 79 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r226 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r227 74 114 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.607 $Y2=0
r228 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r229 73 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r230 73 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r231 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r232 70 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r233 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r234 69 114 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.43 $Y=0
+ $X2=1.607 $Y2=0
r235 69 72 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.43 $Y=0 $X2=1.15
+ $Y2=0
r236 63 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r237 61 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r238 59 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r239 59 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r240 57 91 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.25 $Y=0 $X2=7.13
+ $Y2=0
r241 57 58 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=7.25 $Y=0 $X2=7.412
+ $Y2=0
r242 56 95 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.575 $Y=0 $X2=7.59
+ $Y2=0
r243 56 58 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=7.575 $Y=0 $X2=7.412
+ $Y2=0
r244 54 85 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.29
+ $Y2=0
r245 54 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.5
+ $Y2=0
r246 53 88 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.675 $Y=0 $X2=5.75
+ $Y2=0
r247 53 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.675 $Y=0 $X2=5.5
+ $Y2=0
r248 51 79 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.585 $Y=0
+ $X2=3.45 $Y2=0
r249 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.67
+ $Y2=0
r250 50 82 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.755 $Y=0
+ $X2=3.91 $Y2=0
r251 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.67
+ $Y2=0
r252 46 120 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=11.297 $Y=0.085
+ $X2=11.297 $Y2=0
r253 46 48 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=11.297 $Y=0.085
+ $X2=11.297 $Y2=0.38
r254 42 117 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.877 $Y=0.085
+ $X2=9.877 $Y2=0
r255 42 44 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=9.877 $Y=0.085
+ $X2=9.877 $Y2=0.38
r256 38 58 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.412 $Y=0.085
+ $X2=7.412 $Y2=0
r257 38 40 9.75144 $w=3.23e-07 $l=2.75e-07 $layer=LI1_cond $X=7.412 $Y=0.085
+ $X2=7.412 $Y2=0.36
r258 34 55 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r259 34 36 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.38
r260 30 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0.085
+ $X2=3.67 $Y2=0
r261 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.67 $Y=0.085
+ $X2=3.67 $Y2=0.36
r262 26 114 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.607 $Y=0.085
+ $X2=1.607 $Y2=0
r263 26 28 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.607 $Y=0.085
+ $X2=1.607 $Y2=0.38
r264 22 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r265 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r266 7 48 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=11.09
+ $Y=0.235 $X2=11.28 $Y2=0.38
r267 6 44 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=9.675
+ $Y=0.235 $X2=9.865 $Y2=0.38
r268 5 40 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=7.29
+ $Y=0.235 $X2=7.49 $Y2=0.36
r269 4 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.235 $X2=5.51 $Y2=0.38
r270 3 32 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=3.385
+ $Y=0.235 $X2=3.67 $Y2=0.36
r271 2 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r272 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_791_47# 1 2 7 11 16
r26 14 16 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0.38
+ $X2=4.255 $Y2=0.38
r27 9 11 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.99 $Y=0.425
+ $X2=4.99 $Y2=0.55
r28 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.905 $Y=0.34
+ $X2=4.99 $Y2=0.425
r29 7 16 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.905 $Y=0.34
+ $X2=4.255 $Y2=0.34
r30 2 11 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.235 $X2=4.99 $Y2=0.55
r31 1 14 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.235 $X2=4.09 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFBBN_1%A_1555_47# 1 2 7 9 16
c26 9 0 1.89757e-19 $X=7.91 $Y=0.34
c27 7 0 9.90542e-21 $X=8.785 $Y=0.34
r28 9 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.91 $Y=0.34 $X2=7.91
+ $Y2=0.46
r29 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0.34 $X2=7.91
+ $Y2=0.34
r30 7 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.34
+ $X2=8.87 $Y2=0.34
r31 7 8 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.785 $Y=0.34
+ $X2=8.075 $Y2=0.34
r32 2 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.235 $X2=8.87 $Y2=0.42
r33 1 12 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=7.775
+ $Y=0.235 $X2=7.91 $Y2=0.46
.ends


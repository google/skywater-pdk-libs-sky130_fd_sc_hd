* File: sky130_fd_sc_hd__a2bb2o_2.spice.pex
* Created: Thu Aug 27 14:03:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%A_82_21# 1 2 7 9 12 14 16 19 22 23 24 26 27
+ 28 30 33 36 37 41 45
c114 45 0 7.18975e-20 $X=2.945 $Y=0.785
c115 41 0 1.71567e-19 $X=2.585 $Y=2.275
c116 36 0 1.32536e-19 $X=0.95 $Y=1.16
r117 47 49 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.485 $Y=1.16
+ $X2=0.905 $Y2=1.16
r118 43 45 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.765 $Y=0.785
+ $X2=2.945 $Y2=0.785
r119 41 42 0.446886 $w=2.73e-07 $l=1e-08 $layer=LI1_cond $X=2.645 $Y=2.275
+ $X2=2.645 $Y2=2.285
r120 37 49 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=0.905 $Y2=1.16
r121 36 39 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.992 $Y=1.16
+ $X2=0.992 $Y2=1.325
r122 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.16 $X2=0.95 $Y2=1.16
r123 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.7
+ $X2=2.945 $Y2=0.785
r124 31 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.945 $Y=0.7
+ $X2=2.945 $Y2=0.445
r125 30 41 18.7084 $w=2.73e-07 $l=4.3589e-07 $layer=LI1_cond $X=2.765 $Y=1.895
+ $X2=2.645 $Y2=2.275
r126 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=0.87
+ $X2=2.765 $Y2=0.785
r127 29 30 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.765 $Y=0.87
+ $X2=2.765 $Y2=1.895
r128 27 42 3.50848 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.44 $Y=2.285
+ $X2=2.645 $Y2=2.285
r129 27 28 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.44 $Y=2.285
+ $X2=1.71 $Y2=2.285
r130 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.625 $Y=2.2
+ $X2=1.71 $Y2=2.285
r131 25 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.625 $Y=1.975
+ $X2=1.625 $Y2=2.2
r132 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.54 $Y=1.89
+ $X2=1.625 $Y2=1.975
r133 23 24 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.54 $Y=1.89
+ $X2=1.12 $Y2=1.89
r134 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=1.805
+ $X2=1.12 $Y2=1.89
r135 22 39 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.035 $Y=1.805
+ $X2=1.035 $Y2=1.325
r136 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r137 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r138 14 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r139 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r140 10 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.16
r141 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.985
r142 7 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.16
r143 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
r144 2 41 600 $w=1.7e-07 $l=4.88518e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.845 $X2=2.585 $Y2=2.275
r145 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.235 $X2=2.945 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%A1_N 3 7 9 10 14 15
c37 7 0 1.85041e-19 $X=1.49 $Y=1.805
r38 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.43 $Y2=1.325
r39 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.43 $Y2=0.995
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.16 $X2=1.43 $Y2=1.16
r41 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.51 $Y=1.19 $X2=1.51
+ $Y2=1.53
r42 9 15 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.51 $Y=1.19 $X2=1.51
+ $Y2=1.16
r43 7 17 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.49 $Y=1.805
+ $X2=1.49 $Y2=1.325
r44 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.49 $Y=0.445
+ $X2=1.49 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%A2_N 1 3 6 8
c31 6 0 7.18975e-20 $X=1.91 $Y=0.445
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.16 $X2=1.93 $Y2=1.16
r33 8 12 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=2.05 $Y=1.185
+ $X2=1.93 $Y2=1.185
r34 4 11 38.945 $w=2.68e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.91 $Y=0.995
+ $X2=1.92 $Y2=1.16
r35 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.91 $Y=0.995 $X2=1.91
+ $Y2=0.445
r36 1 11 47.9375 $w=2.68e-07 $l=2.47538e-07 $layer=POLY_cond $X=1.85 $Y=1.375
+ $X2=1.92 $Y2=1.16
r37 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.85 $Y=1.375 $X2=1.85
+ $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%A_313_47# 1 2 7 9 10 12 16 18 19 20 25 29
c61 25 0 1.04517e-19 $X=2.425 $Y=1.155
c62 10 0 1.46486e-19 $X=2.795 $Y=1.435
r63 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.425
+ $Y=1.155 $X2=2.425 $Y2=1.155
r64 23 25 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.425 $Y=1.545
+ $X2=2.425 $Y2=1.155
r65 22 25 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.425 $Y=0.825
+ $X2=2.425 $Y2=1.155
r66 21 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=1.63
+ $X2=2.06 $Y2=1.63
r67 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.34 $Y=1.63
+ $X2=2.425 $Y2=1.545
r68 20 21 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.34 $Y=1.63
+ $X2=2.145 $Y2=1.63
r69 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.34 $Y=0.74
+ $X2=2.425 $Y2=0.825
r70 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.34 $Y=0.74
+ $X2=1.785 $Y2=0.74
r71 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.7 $Y=0.655
+ $X2=1.785 $Y2=0.74
r72 14 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.7 $Y=0.655 $X2=1.7
+ $Y2=0.445
r73 10 26 53.3539 $w=5.54e-07 $l=3.7229e-07 $layer=POLY_cond $X=2.795 $Y=1.435
+ $X2=2.58 $Y2=1.155
r74 10 12 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.795 $Y=1.435
+ $X2=2.795 $Y2=2.165
r75 7 26 62.9243 $w=5.54e-07 $l=4.61031e-07 $layer=POLY_cond $X=2.735 $Y=0.765
+ $X2=2.58 $Y2=1.155
r76 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.735 $Y=0.765
+ $X2=2.735 $Y2=0.445
r77 2 29 600 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=1.485 $X2=2.06 $Y2=1.71
r78 1 16 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.7 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%B2 3 7 11 14 20
c45 20 0 1.46486e-19 $X=3.4 $Y=1.505
c46 14 0 1.64941e-19 $X=3.215 $Y=1.47
c47 11 0 1.22353e-19 $X=3.445 $Y=1.53
c48 7 0 1.85736e-19 $X=3.25 $Y=2.165
c49 3 0 1.04517e-19 $X=3.155 $Y=0.445
r50 15 20 7.10673 $w=2.98e-07 $l=1.85e-07 $layer=LI1_cond $X=3.215 $Y=1.505
+ $X2=3.4 $Y2=1.505
r51 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.47
+ $X2=3.215 $Y2=1.635
r52 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.47
+ $X2=3.215 $Y2=1.305
r53 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=1.47 $X2=3.215 $Y2=1.47
r54 11 20 1.72866 $w=2.98e-07 $l=4.5e-08 $layer=LI1_cond $X=3.445 $Y=1.505
+ $X2=3.4 $Y2=1.505
r55 7 17 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.25 $Y=2.165
+ $X2=3.25 $Y2=1.635
r56 3 16 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.155 $Y=0.445
+ $X2=3.155 $Y2=1.305
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%B1 3 7 9 10 11 16
c29 16 0 1.22353e-19 $X=3.67 $Y=1.16
c30 9 0 1.41684e-20 $X=3.905 $Y=0.85
r31 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.815
+ $Y=1.16 $X2=3.815 $Y2=1.16
r32 16 18 23.9349 $w=2.92e-07 $l=1.45e-07 $layer=POLY_cond $X=3.67 $Y=1.16
+ $X2=3.815 $Y2=1.16
r33 10 11 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=3.86 $Y=1.19
+ $X2=3.86 $Y2=1.53
r34 10 19 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=3.86 $Y=1.19 $X2=3.86
+ $Y2=1.16
r35 9 19 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=3.86 $Y=0.85 $X2=3.86
+ $Y2=1.16
r36 5 16 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r37 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.67 $Y=1.325 $X2=3.67
+ $Y2=2.165
r38 1 16 15.6815 $w=2.92e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.67 $Y2=1.16
r39 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%VPWR 1 2 3 12 16 18 21 23 28 35 36 44 47 50
+ 58
c62 12 0 1.85041e-19 $X=1.115 $Y=2.32
r63 50 53 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.27 $Y=1.64
+ $X2=0.27 $Y2=2.32
r64 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r65 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 36 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r67 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 33 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.625 $Y=2.72
+ $X2=3.5 $Y2=2.72
r69 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.625 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 32 48 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.45 $Y2=2.72
r71 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 29 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.115 $Y2=2.72
r74 29 31 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.61 $Y2=2.72
r75 28 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.375 $Y=2.72
+ $X2=3.5 $Y2=2.72
r76 28 31 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=3.375 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 27 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r78 27 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r79 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 23 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=2.72
+ $X2=1.115 $Y2=2.72
r82 23 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.95 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 21 58 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=2.72
+ $X2=0.23 $Y2=2.72
r84 18 53 14.7307 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=2.32
r85 18 24 3.40825 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.177 $Y=2.72
+ $X2=0.355 $Y2=2.72
r86 18 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r87 14 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=2.635
+ $X2=3.5 $Y2=2.72
r88 14 16 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.5 $Y=2.635
+ $X2=3.5 $Y2=2.34
r89 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.635
+ $X2=1.115 $Y2=2.72
r90 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.115 $Y=2.635
+ $X2=1.115 $Y2=2.32
r91 3 16 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=1.845 $X2=3.46 $Y2=2.34
r92 2 12 600 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.485 $X2=1.115 $Y2=2.32
r93 1 53 400 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=2.32
r94 1 50 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%X 1 2 10 11 12 13 14 15 24
r23 14 15 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.652 $Y=1.87
+ $X2=0.652 $Y2=2.21
r24 14 24 4.97132 $w=2.53e-07 $l=1.1e-07 $layer=LI1_cond $X=0.652 $Y=1.87
+ $X2=0.652 $Y2=1.76
r25 11 24 4.88094 $w=2.53e-07 $l=1.08e-07 $layer=LI1_cond $X=0.652 $Y=1.652
+ $X2=0.652 $Y2=1.76
r26 11 12 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=0.652 $Y=1.652
+ $X2=0.652 $Y2=1.525
r27 10 12 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.61 $Y=0.81
+ $X2=0.61 $Y2=1.525
r28 9 13 7.81853 $w=2.53e-07 $l=1.73e-07 $layer=LI1_cond $X=0.652 $Y=0.683
+ $X2=0.652 $Y2=0.51
r29 9 10 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=0.652 $Y=0.683
+ $X2=0.652 $Y2=0.81
r30 2 24 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=1.485 $X2=0.695 $Y2=1.76
r31 1 13 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.695 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%A_574_369# 1 2 8 9 10 13 16
c29 9 0 1.64941e-19 $X=3.795 $Y=1.92
r30 11 13 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.88 $Y=2.005
+ $X2=3.88 $Y2=2.275
r31 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.795 $Y=1.92
+ $X2=3.88 $Y2=2.005
r32 9 10 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.795 $Y=1.92
+ $X2=3.205 $Y2=1.92
r33 8 16 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.12 $Y=2.255
+ $X2=3.04 $Y2=2.34
r34 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.12 $Y=2.005
+ $X2=3.205 $Y2=1.92
r35 7 8 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.12 $Y=2.005 $X2=3.12
+ $Y2=2.255
r36 2 13 600 $w=1.7e-07 $l=4.929e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.845 $X2=3.88 $Y2=2.275
r37 1 16 600 $w=1.7e-07 $l=5.73738e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.845 $X2=3.04 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_2%VGND 1 2 3 4 15 17 19 21 24 26 36 47 52 58
+ 61 63 69
r63 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r64 56 58 9.85609 $w=5.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=0.2 $X2=2.69
+ $Y2=0.2
r65 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r66 54 56 0.104919 $w=5.68e-07 $l=5e-09 $layer=LI1_cond $X=2.525 $Y=0.2 $X2=2.53
+ $Y2=0.2
r67 51 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r68 50 54 9.54764 $w=5.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.07 $Y=0.2
+ $X2=2.525 $Y2=0.2
r69 50 52 8.91182 $w=5.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.07 $Y=0.2
+ $X2=1.955 $Y2=0.2
r70 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r71 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r72 40 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r73 40 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r74 39 58 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.69
+ $Y2=0
r75 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r76 36 60 5.33421 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=3.605 $Y=0 $X2=3.872
+ $Y2=0
r77 36 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.605 $Y=0 $X2=3.45
+ $Y2=0
r78 35 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r79 35 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r80 34 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.955
+ $Y2=0
r81 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r82 32 47 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.38 $Y=0 $X2=1.165
+ $Y2=0
r83 32 34 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.38 $Y=0 $X2=1.61
+ $Y2=0
r84 30 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r85 30 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r86 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r87 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.69
+ $Y2=0
r88 26 47 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.165
+ $Y2=0
r89 26 29 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.69
+ $Y2=0
r90 24 69 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=0 $X2=0.23
+ $Y2=0
r91 21 63 13.9075 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r92 21 27 3.40825 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.177 $Y=0 $X2=0.355
+ $Y2=0
r93 21 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r94 17 60 3.0367 $w=4e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.872 $Y2=0
r95 17 19 9.93982 $w=3.98e-07 $l=3.45e-07 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0.43
r96 13 47 1.67165 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0
r97 13 15 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0.445
r98 4 19 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.785 $Y2=0.43
r99 3 54 91 $w=1.7e-07 $l=6.17009e-07 $layer=licon1_NDIFF $count=2 $X=1.985
+ $Y=0.235 $X2=2.525 $Y2=0.4
r100 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.115 $Y2=0.445
r101 1 63 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__and3b_1.pxi.spice
* Created: Thu Aug 27 14:07:56 2020
* 
x_PM_SKY130_FD_SC_HD__AND3B_1%A_N N_A_N_c_66_n N_A_N_M1008_g N_A_N_M1004_g
+ N_A_N_c_72_n A_N A_N A_N N_A_N_c_68_n N_A_N_c_69_n
+ PM_SKY130_FD_SC_HD__AND3B_1%A_N
x_PM_SKY130_FD_SC_HD__AND3B_1%A_109_93# N_A_109_93#_M1008_d N_A_109_93#_M1004_d
+ N_A_109_93#_M1003_g N_A_109_93#_M1005_g N_A_109_93#_c_92_n N_A_109_93#_c_93_n
+ N_A_109_93#_c_94_n N_A_109_93#_c_95_n PM_SKY130_FD_SC_HD__AND3B_1%A_109_93#
x_PM_SKY130_FD_SC_HD__AND3B_1%B N_B_M1006_g N_B_M1000_g N_B_c_136_n B
+ N_B_c_139_n PM_SKY130_FD_SC_HD__AND3B_1%B
x_PM_SKY130_FD_SC_HD__AND3B_1%C N_C_M1009_g N_C_M1001_g C C N_C_c_175_n
+ PM_SKY130_FD_SC_HD__AND3B_1%C
x_PM_SKY130_FD_SC_HD__AND3B_1%A_209_311# N_A_209_311#_M1005_s
+ N_A_209_311#_M1003_s N_A_209_311#_M1000_d N_A_209_311#_M1002_g
+ N_A_209_311#_M1007_g N_A_209_311#_c_225_n N_A_209_311#_c_219_n
+ N_A_209_311#_c_226_n N_A_209_311#_c_227_n N_A_209_311#_c_220_n
+ N_A_209_311#_c_229_n N_A_209_311#_c_230_n N_A_209_311#_c_221_n
+ N_A_209_311#_c_222_n N_A_209_311#_c_223_n
+ PM_SKY130_FD_SC_HD__AND3B_1%A_209_311#
x_PM_SKY130_FD_SC_HD__AND3B_1%VPWR N_VPWR_M1004_s N_VPWR_M1003_d N_VPWR_M1001_d
+ N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_321_n VPWR
+ N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_305_n N_VPWR_c_313_n
+ N_VPWR_c_314_n PM_SKY130_FD_SC_HD__AND3B_1%VPWR
x_PM_SKY130_FD_SC_HD__AND3B_1%X N_X_M1002_d N_X_M1007_d N_X_c_361_n N_X_c_358_n
+ N_X_c_359_n X X N_X_c_363_n PM_SKY130_FD_SC_HD__AND3B_1%X
x_PM_SKY130_FD_SC_HD__AND3B_1%VGND N_VGND_M1008_s N_VGND_M1009_d N_VGND_c_376_n
+ N_VGND_c_377_n N_VGND_c_378_n VGND N_VGND_c_379_n N_VGND_c_380_n
+ N_VGND_c_381_n N_VGND_c_382_n PM_SKY130_FD_SC_HD__AND3B_1%VGND
cc_1 VNB N_A_N_c_66_n 0.00932119f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.478
cc_2 VNB A_N 0.00882809f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_68_n 0.0325929f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_4 VNB N_A_N_c_69_n 0.021365f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=0.995
cc_5 VNB N_A_109_93#_M1005_g 0.0319859f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.785
cc_6 VNB N_A_109_93#_c_92_n 0.017805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_109_93#_c_93_n 0.0013167f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_8 VNB N_A_109_93#_c_94_n 0.0134771f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_9 VNB N_A_109_93#_c_95_n 0.0337288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_M1006_g 0.0249958f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_11 VNB N_B_M1000_g 0.00462445f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_12 VNB N_B_c_136_n 0.0115371f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.695
cc_13 VNB N_C_M1009_g 0.0261825f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB C 2.32476e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB C 0.0107497f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.695
cc_16 VNB N_C_c_175_n 0.0195606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_209_311#_c_219_n 0.00550334f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_18 VNB N_A_209_311#_c_220_n 0.00502922f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_209_311#_c_221_n 0.00368314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_209_311#_c_222_n 0.0230746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_209_311#_c_223_n 0.0207919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_305_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_358_n 0.0251358f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.695
cc_24 VNB N_X_c_359_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_25 VNB X 0.0136214f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.785
cc_26 VNB N_VGND_c_376_n 0.0099134f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_27 VNB N_VGND_c_377_n 0.0388434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_378_n 0.00317442f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.785
cc_29 VNB N_VGND_c_379_n 0.0534217f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_30 VNB N_VGND_c_380_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_381_n 0.206426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_382_n 0.00507625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A_N_c_66_n 0.016988f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.478
cc_34 VPB N_A_N_M1004_g 0.0422708f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_35 VPB N_A_N_c_72_n 0.0294939f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.695
cc_36 VPB A_N 0.0279341f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_37 VPB N_A_109_93#_M1003_g 0.0261578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_109_93#_c_93_n 0.0164308f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.16
cc_39 VPB N_A_109_93#_c_95_n 0.00815218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_B_M1000_g 0.0221455f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_41 VPB B 0.00941122f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_42 VPB N_B_c_139_n 0.0418573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_C_M1001_g 0.0204691f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_44 VPB N_C_c_175_n 0.00424946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_209_311#_M1007_g 0.0241986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_209_311#_c_225_n 0.00385633f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_47 VPB N_A_209_311#_c_226_n 0.00323619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_209_311#_c_227_n 0.00369523f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.87
cc_49 VPB N_A_209_311#_c_220_n 0.0011546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_209_311#_c_229_n 0.00697372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_209_311#_c_230_n 0.00553659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_209_311#_c_221_n 0.00122273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_209_311#_c_222_n 0.005118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_306_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.695
cc_55 VPB N_VPWR_c_307_n 0.0186681f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_56 VPB N_VPWR_c_308_n 0.0049827f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_57 VPB N_VPWR_c_309_n 0.0527465f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_310_n 0.0212745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_311_n 0.0177135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_305_n 0.0563135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_313_n 0.00142003f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_314_n 0.00411068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_X_c_361_n 0.00524127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_358_n 0.0183929f $X=-0.19 $Y=1.305 $X2=0.327 $Y2=1.695
cc_65 VPB N_X_c_363_n 0.0218575f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 A_N N_A_109_93#_c_92_n 0.014326f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_N_c_69_n N_A_109_93#_c_92_n 0.0169183f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_68 N_A_N_c_66_n N_A_109_93#_c_93_n 0.0212293f $X=0.327 $Y=1.478 $X2=0 $Y2=0
cc_69 A_N N_A_109_93#_c_93_n 0.0533628f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_N_c_68_n N_A_109_93#_c_95_n 0.00567702f $X=0.26 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_N_c_69_n N_A_209_311#_c_219_n 0.00474782f $X=0.327 $Y=0.995 $X2=0
+ $Y2=0
cc_72 N_A_N_M1004_g N_VPWR_c_307_n 0.00320628f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_73 N_A_N_c_72_n N_VPWR_c_307_n 0.00101412f $X=0.327 $Y=1.695 $X2=0 $Y2=0
cc_74 A_N N_VPWR_c_307_n 0.0227749f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_N_M1004_g N_VPWR_c_309_n 0.00844098f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_76 N_A_N_M1004_g N_VPWR_c_305_n 0.0120826f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_77 A_N N_VPWR_c_305_n 0.00409195f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_78 A_N N_VGND_c_377_n 0.0231087f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_N_c_68_n N_VGND_c_377_n 0.0069709f $X=0.26 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_N_c_69_n N_VGND_c_377_n 0.00710775f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_N_c_69_n N_VGND_c_379_n 0.00483902f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_N_c_69_n N_VGND_c_381_n 0.00512902f $X=0.327 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_109_93#_M1005_g N_B_M1006_g 0.0330906f $X=1.405 $Y=0.475 $X2=0 $Y2=0
cc_84 N_A_109_93#_M1003_g N_B_M1000_g 0.0211871f $X=1.38 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_109_93#_c_95_n N_B_M1000_g 0.00639148f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_109_93#_c_95_n N_B_c_136_n 0.0330906f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_109_93#_c_93_n N_A_209_311#_c_225_n 0.0222277f $X=0.68 $Y=2.26 $X2=0
+ $Y2=0
cc_88 N_A_109_93#_M1005_g N_A_209_311#_c_219_n 0.0131224f $X=1.405 $Y=0.475
+ $X2=0 $Y2=0
cc_89 N_A_109_93#_c_92_n N_A_209_311#_c_219_n 0.0071667f $X=0.68 $Y=1.245 $X2=0
+ $Y2=0
cc_90 N_A_109_93#_c_94_n N_A_209_311#_c_219_n 0.0124117f $X=1.195 $Y=1.16 $X2=0
+ $Y2=0
cc_91 N_A_109_93#_c_95_n N_A_209_311#_c_219_n 0.00498369f $X=1.405 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_A_109_93#_M1003_g N_A_209_311#_c_226_n 0.0143457f $X=1.38 $Y=1.765 $X2=0
+ $Y2=0
cc_93 N_A_109_93#_c_94_n N_A_209_311#_c_226_n 0.00915944f $X=1.195 $Y=1.16 $X2=0
+ $Y2=0
cc_94 N_A_109_93#_c_95_n N_A_209_311#_c_226_n 0.00234152f $X=1.405 $Y=1.16 $X2=0
+ $Y2=0
cc_95 N_A_109_93#_c_93_n N_A_209_311#_c_227_n 0.0112734f $X=0.68 $Y=2.26 $X2=0
+ $Y2=0
cc_96 N_A_109_93#_c_94_n N_A_209_311#_c_227_n 0.0196457f $X=1.195 $Y=1.16 $X2=0
+ $Y2=0
cc_97 N_A_109_93#_c_95_n N_A_209_311#_c_227_n 0.0049356f $X=1.405 $Y=1.16 $X2=0
+ $Y2=0
cc_98 N_A_109_93#_M1003_g N_A_209_311#_c_220_n 0.00238678f $X=1.38 $Y=1.765
+ $X2=0 $Y2=0
cc_99 N_A_109_93#_M1005_g N_A_209_311#_c_220_n 0.0140084f $X=1.405 $Y=0.475
+ $X2=0 $Y2=0
cc_100 N_A_109_93#_c_94_n N_A_209_311#_c_220_n 0.020412f $X=1.195 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_109_93#_M1003_g N_VPWR_c_321_n 0.00256209f $X=1.38 $Y=1.765 $X2=0
+ $Y2=0
cc_102 N_A_109_93#_M1003_g N_VPWR_c_309_n 0.00483317f $X=1.38 $Y=1.765 $X2=0
+ $Y2=0
cc_103 N_A_109_93#_c_93_n N_VPWR_c_309_n 0.0330845f $X=0.68 $Y=2.26 $X2=0 $Y2=0
cc_104 N_A_109_93#_M1004_d N_VPWR_c_305_n 0.00529506f $X=0.545 $Y=2.065 $X2=0
+ $Y2=0
cc_105 N_A_109_93#_c_93_n N_VPWR_c_305_n 0.00646998f $X=0.68 $Y=2.26 $X2=0 $Y2=0
cc_106 N_A_109_93#_M1003_g N_VPWR_c_313_n 0.00567892f $X=1.38 $Y=1.765 $X2=0
+ $Y2=0
cc_107 N_A_109_93#_c_93_n N_VPWR_c_313_n 0.00428127f $X=0.68 $Y=2.26 $X2=0 $Y2=0
cc_108 N_A_109_93#_c_92_n N_VGND_c_377_n 0.0166146f $X=0.68 $Y=1.245 $X2=0 $Y2=0
cc_109 N_A_109_93#_M1005_g N_VGND_c_379_n 0.00347765f $X=1.405 $Y=0.475 $X2=0
+ $Y2=0
cc_110 N_A_109_93#_c_92_n N_VGND_c_379_n 0.00841481f $X=0.68 $Y=1.245 $X2=0
+ $Y2=0
cc_111 N_A_109_93#_M1005_g N_VGND_c_381_n 0.0059338f $X=1.405 $Y=0.475 $X2=0
+ $Y2=0
cc_112 N_A_109_93#_c_92_n N_VGND_c_381_n 0.0109761f $X=0.68 $Y=1.245 $X2=0 $Y2=0
cc_113 N_B_M1006_g N_C_M1009_g 0.0416192f $X=1.765 $Y=0.475 $X2=0 $Y2=0
cc_114 N_B_M1000_g N_C_M1001_g 0.0127087f $X=1.8 $Y=1.765 $X2=0 $Y2=0
cc_115 B N_C_M1001_g 0.00197753f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_116 N_B_M1006_g C 0.00410621f $X=1.765 $Y=0.475 $X2=0 $Y2=0
cc_117 N_B_c_136_n C 0.00141844f $X=1.782 $Y=1.2 $X2=0 $Y2=0
cc_118 N_B_c_136_n N_C_c_175_n 0.017487f $X=1.782 $Y=1.2 $X2=0 $Y2=0
cc_119 N_B_c_139_n N_A_209_311#_M1007_g 0.00222866f $X=1.875 $Y=2.3 $X2=0 $Y2=0
cc_120 N_B_M1006_g N_A_209_311#_c_219_n 0.00808008f $X=1.765 $Y=0.475 $X2=0
+ $Y2=0
cc_121 N_B_M1006_g N_A_209_311#_c_220_n 0.0096969f $X=1.765 $Y=0.475 $X2=0 $Y2=0
cc_122 N_B_M1000_g N_A_209_311#_c_220_n 0.00631839f $X=1.8 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B_c_136_n N_A_209_311#_c_220_n 0.00498235f $X=1.782 $Y=1.2 $X2=0 $Y2=0
cc_124 B N_A_209_311#_c_229_n 0.00347271f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_125 N_B_M1000_g N_A_209_311#_c_230_n 0.0129761f $X=1.8 $Y=1.765 $X2=0 $Y2=0
cc_126 B N_A_209_311#_c_230_n 0.0179395f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_127 N_B_c_139_n N_A_209_311#_c_230_n 5.9549e-19 $X=1.875 $Y=2.3 $X2=0 $Y2=0
cc_128 N_B_M1000_g N_VPWR_c_308_n 8.70935e-19 $X=1.8 $Y=1.765 $X2=0 $Y2=0
cc_129 B N_VPWR_c_308_n 0.0277106f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_130 N_B_c_139_n N_VPWR_c_308_n 0.001313f $X=1.875 $Y=2.3 $X2=0 $Y2=0
cc_131 N_B_M1000_g N_VPWR_c_321_n 0.0037226f $X=1.8 $Y=1.765 $X2=0 $Y2=0
cc_132 N_B_c_139_n N_VPWR_c_309_n 0.00672592f $X=1.875 $Y=2.3 $X2=0 $Y2=0
cc_133 B N_VPWR_c_310_n 0.0314336f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_134 N_B_c_139_n N_VPWR_c_310_n 0.00611913f $X=1.875 $Y=2.3 $X2=0 $Y2=0
cc_135 B N_VPWR_c_305_n 0.0169635f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_136 N_B_c_139_n N_VPWR_c_305_n 0.00863692f $X=1.875 $Y=2.3 $X2=0 $Y2=0
cc_137 N_B_M1000_g N_VPWR_c_313_n 0.00672592f $X=1.8 $Y=1.765 $X2=0 $Y2=0
cc_138 B N_VPWR_c_313_n 0.0288891f $X=1.985 $Y=2.125 $X2=0 $Y2=0
cc_139 N_B_M1006_g N_VGND_c_379_n 0.00382191f $X=1.765 $Y=0.475 $X2=0 $Y2=0
cc_140 N_B_M1006_g N_VGND_c_381_n 0.00577482f $X=1.765 $Y=0.475 $X2=0 $Y2=0
cc_141 N_C_M1001_g N_A_209_311#_M1007_g 0.026318f $X=2.275 $Y=1.695 $X2=0 $Y2=0
cc_142 N_C_M1009_g N_A_209_311#_c_219_n 2.65899e-19 $X=2.17 $Y=0.475 $X2=0 $Y2=0
cc_143 C N_A_209_311#_c_219_n 0.0210672f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_144 N_C_M1009_g N_A_209_311#_c_220_n 6.64342e-19 $X=2.17 $Y=0.475 $X2=0 $Y2=0
cc_145 N_C_M1001_g N_A_209_311#_c_220_n 5.35136e-19 $X=2.275 $Y=1.695 $X2=0
+ $Y2=0
cc_146 C N_A_209_311#_c_220_n 0.0523822f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_147 N_C_c_175_n N_A_209_311#_c_220_n 4.85299e-19 $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_148 N_C_M1001_g N_A_209_311#_c_229_n 0.0169633f $X=2.275 $Y=1.695 $X2=0 $Y2=0
cc_149 C N_A_209_311#_c_229_n 0.0145969f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_150 N_C_c_175_n N_A_209_311#_c_229_n 3.77498e-19 $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_151 N_C_M1001_g N_A_209_311#_c_230_n 0.00182091f $X=2.275 $Y=1.695 $X2=0
+ $Y2=0
cc_152 C N_A_209_311#_c_230_n 0.0187467f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_153 N_C_c_175_n N_A_209_311#_c_230_n 0.00309114f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_154 N_C_M1001_g N_A_209_311#_c_221_n 0.00209955f $X=2.275 $Y=1.695 $X2=0
+ $Y2=0
cc_155 C N_A_209_311#_c_221_n 0.020603f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_156 N_C_c_175_n N_A_209_311#_c_221_n 0.00238051f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_157 C N_A_209_311#_c_222_n 8.36739e-19 $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_158 N_C_c_175_n N_A_209_311#_c_222_n 0.0211349f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_159 N_C_M1009_g N_A_209_311#_c_223_n 0.015251f $X=2.17 $Y=0.475 $X2=0 $Y2=0
cc_160 C N_A_209_311#_c_223_n 6.12497e-19 $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_161 C N_A_209_311#_c_223_n 0.00275588f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_162 N_C_M1001_g N_VPWR_c_321_n 2.74587e-19 $X=2.275 $Y=1.695 $X2=0 $Y2=0
cc_163 N_C_M1001_g N_VPWR_c_310_n 0.00189602f $X=2.275 $Y=1.695 $X2=0 $Y2=0
cc_164 N_C_M1001_g N_VPWR_c_305_n 0.00236577f $X=2.275 $Y=1.695 $X2=0 $Y2=0
cc_165 C N_X_c_358_n 0.00874933f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_166 N_C_M1009_g N_VGND_c_378_n 0.00582287f $X=2.17 $Y=0.475 $X2=0 $Y2=0
cc_167 C N_VGND_c_378_n 0.0164905f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_168 C N_VGND_c_378_n 0.00148069f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_169 N_C_M1009_g N_VGND_c_379_n 0.00374894f $X=2.17 $Y=0.475 $X2=0 $Y2=0
cc_170 C N_VGND_c_379_n 0.00888859f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_171 C N_VGND_c_379_n 0.00302635f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_172 N_C_M1009_g N_VGND_c_381_n 0.00557291f $X=2.17 $Y=0.475 $X2=0 $Y2=0
cc_173 C N_VGND_c_381_n 0.00701514f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_174 C N_VGND_c_381_n 0.00509342f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_175 C A_368_53# 0.00371508f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_176 N_A_209_311#_c_226_n N_VPWR_M1003_d 5.00837e-19 $X=1.56 $Y=1.51 $X2=0
+ $Y2=0
cc_177 N_A_209_311#_c_230_n N_VPWR_M1003_d 0.0011981f $X=2.207 $Y=1.657 $X2=0
+ $Y2=0
cc_178 N_A_209_311#_c_229_n N_VPWR_M1001_d 0.00275705f $X=2.565 $Y=1.657 $X2=0
+ $Y2=0
cc_179 N_A_209_311#_M1007_g N_VPWR_c_308_n 0.00549229f $X=2.75 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_209_311#_c_229_n N_VPWR_c_308_n 0.0136834f $X=2.565 $Y=1.657 $X2=0
+ $Y2=0
cc_181 N_A_209_311#_c_226_n N_VPWR_c_321_n 0.00549589f $X=1.56 $Y=1.51 $X2=0
+ $Y2=0
cc_182 N_A_209_311#_c_230_n N_VPWR_c_321_n 0.0195825f $X=2.207 $Y=1.657 $X2=0
+ $Y2=0
cc_183 N_A_209_311#_c_225_n N_VPWR_c_309_n 0.0215377f $X=1.17 $Y=1.76 $X2=0
+ $Y2=0
cc_184 N_A_209_311#_c_226_n N_VPWR_c_309_n 0.00511706f $X=1.56 $Y=1.51 $X2=0
+ $Y2=0
cc_185 N_A_209_311#_M1007_g N_VPWR_c_311_n 0.00585385f $X=2.75 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_209_311#_M1007_g N_VPWR_c_305_n 0.0123821f $X=2.75 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_209_311#_c_225_n N_VPWR_c_305_n 9.89565e-19 $X=1.17 $Y=1.76 $X2=0
+ $Y2=0
cc_188 N_A_209_311#_c_229_n N_VPWR_c_305_n 0.00854634f $X=2.565 $Y=1.657 $X2=0
+ $Y2=0
cc_189 N_A_209_311#_M1007_g N_X_c_358_n 0.00837276f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_209_311#_c_229_n N_X_c_358_n 0.0226631f $X=2.565 $Y=1.657 $X2=0 $Y2=0
cc_191 N_A_209_311#_c_221_n N_X_c_358_n 0.0313758f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_209_311#_c_222_n N_X_c_358_n 0.00753248f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_209_311#_c_223_n N_X_c_358_n 0.00624157f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_209_311#_c_221_n N_VGND_c_378_n 0.00432911f $X=2.71 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_209_311#_c_222_n N_VGND_c_378_n 4.32142e-19 $X=2.71 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_209_311#_c_223_n N_VGND_c_378_n 0.0103745f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_209_311#_c_219_n N_VGND_c_379_n 0.0355665f $X=1.56 $Y=0.437 $X2=0
+ $Y2=0
cc_198 N_A_209_311#_c_223_n N_VGND_c_380_n 0.0046653f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_209_311#_c_219_n N_VGND_c_381_n 0.0278067f $X=1.56 $Y=0.437 $X2=0
+ $Y2=0
cc_200 N_A_209_311#_c_223_n N_VGND_c_381_n 0.00895857f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_209_311#_c_219_n A_296_53# 0.00191292f $X=1.56 $Y=0.437 $X2=-0.19
+ $Y2=-0.24
cc_202 N_A_209_311#_c_220_n A_296_53# 0.00132529f $X=1.687 $Y=1.425 $X2=-0.19
+ $Y2=-0.24
cc_203 N_VPWR_c_305_n N_X_M1007_d 0.00335098f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_204 N_VPWR_c_311_n N_X_c_363_n 0.0185457f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_205 N_VPWR_c_305_n N_X_c_363_n 0.0105168f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_206 X N_VGND_c_380_n 0.0178555f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_207 N_X_M1002_d N_VGND_c_381_n 0.00387172f $X=2.825 $Y=0.235 $X2=0 $Y2=0
cc_208 X N_VGND_c_381_n 0.00990557f $X=2.9 $Y=0.425 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__xor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
M1000 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=1.4144e+12p ps=1.289e+07u
M1001 a_608_49# B a_1135_365# VNB nshort w=640000u l=150000u
+  ad=5.401e+11p pd=4.32e+06u as=3.828e+11p ps=3.78e+06u
M1002 a_480_297# C VPWR VPB phighvt w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=0p ps=0u
M1003 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1402_49# a_1031_297# a_608_49# VNB nshort w=420000u l=150000u
+  ad=5.517e+11p pd=4.37e+06u as=0p ps=0u
M1005 a_1031_297# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.526e+11p pd=2.52e+06u as=0p ps=0u
M1006 a_1402_49# a_1135_365# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.0424e+12p ps=9.75e+06u
M1007 a_79_21# C a_608_49# VNB nshort w=640000u l=150000u
+  ad=2.56e+11p pd=2.08e+06u as=0p ps=0u
M1008 a_602_325# B a_1402_49# VNB nshort w=640000u l=150000u
+  ad=5.9845e+11p pd=4.47e+06u as=0p ps=0u
M1009 a_1135_365# a_1031_297# a_608_49# VPB phighvt w=840000u l=150000u
+  ad=6.966e+11p pd=5.24e+06u as=7.326e+11p ps=5.14e+06u
M1010 a_79_21# C a_602_325# VPB phighvt w=840000u l=150000u
+  ad=3.192e+11p pd=2.44e+06u as=7.088e+11p ps=5.1e+06u
M1011 a_608_49# B a_1402_49# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=7.52e+11p ps=5.57e+06u
M1012 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.51e+11p ps=3.68e+06u
M1013 VPWR A a_1135_365# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1402_49# a_1031_297# a_602_325# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1402_49# a_1135_365# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_79_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A a_1135_365# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_602_325# B a_1135_365# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_480_297# C VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1022 a_1135_365# a_1031_297# a_602_325# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_79_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_608_49# a_480_297# a_79_21# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_602_325# a_480_297# a_79_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1031_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.653e+11p pd=1.82e+06u as=0p ps=0u
.ends


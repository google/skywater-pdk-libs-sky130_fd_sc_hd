* File: sky130_fd_sc_hd__lpflow_isobufsrc_16.spice
* Created: Tue Sep  1 19:12:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_isobufsrc_16.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_isobufsrc_16  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1038 N_VGND_M1038_d N_A_M1038_g N_A_143_297#_M1038_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75015.2 A=0.0975 P=1.6 MULT=1
MM1043 N_VGND_M1043_d N_A_M1043_g N_A_143_297#_M1038_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75014.8 A=0.0975 P=1.6 MULT=1
MM1049 N_VGND_M1043_d N_A_M1049_g N_A_143_297#_M1049_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75014.4 A=0.0975 P=1.6 MULT=1
MM1064 N_VGND_M1064_d N_A_M1064_g N_A_143_297#_M1049_s VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.08775 PD=1.26 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75014 A=0.0975 P=1.6 MULT=1
MM1002 N_X_M1002_d N_A_143_297#_M1002_g N_VGND_M1064_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.19825 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.2
+ SB=75013.2 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1002_d N_A_143_297#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75012.8 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_143_297#_M1007_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75012.4 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1007_d N_A_143_297#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75011.9 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1010_d N_A_143_297#_M1010_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.9
+ SB=75011.5 A=0.0975 P=1.6 MULT=1
MM1015 N_X_M1010_d N_A_143_297#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.3
+ SB=75011.1 A=0.0975 P=1.6 MULT=1
MM1016 N_X_M1016_d N_A_143_297#_M1016_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.7
+ SB=75010.7 A=0.0975 P=1.6 MULT=1
MM1021 N_X_M1016_d N_A_143_297#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.1
+ SB=75010.3 A=0.0975 P=1.6 MULT=1
MM1022 N_X_M1022_d N_A_143_297#_M1022_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.6
+ SB=75009.8 A=0.0975 P=1.6 MULT=1
MM1027 N_X_M1022_d N_A_143_297#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006
+ SB=75009.4 A=0.0975 P=1.6 MULT=1
MM1028 N_X_M1028_d N_A_143_297#_M1028_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.4
+ SB=75009 A=0.0975 P=1.6 MULT=1
MM1055 N_X_M1028_d N_A_143_297#_M1055_g N_VGND_M1055_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.8
+ SB=75008.6 A=0.0975 P=1.6 MULT=1
MM1062 N_X_M1062_d N_A_143_297#_M1062_g N_VGND_M1055_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.2
+ SB=75008.2 A=0.0975 P=1.6 MULT=1
MM1065 N_X_M1062_d N_A_143_297#_M1065_g N_VGND_M1065_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75007.7
+ SB=75007.7 A=0.0975 P=1.6 MULT=1
MM1067 N_X_M1067_d N_A_143_297#_M1067_g N_VGND_M1065_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.1
+ SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1068 N_X_M1067_d N_A_143_297#_M1068_g N_VGND_M1068_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.5
+ SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1018 N_X_M1018_d N_SLEEP_M1018_g N_VGND_M1068_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75008.9
+ SB=75006.5 A=0.0975 P=1.6 MULT=1
MM1029 N_X_M1018_d N_SLEEP_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009.3
+ SB=75006.1 A=0.0975 P=1.6 MULT=1
MM1030 N_X_M1030_d N_SLEEP_M1030_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75009.8
+ SB=75005.6 A=0.0975 P=1.6 MULT=1
MM1033 N_X_M1030_d N_SLEEP_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75010.2
+ SB=75005.2 A=0.0975 P=1.6 MULT=1
MM1035 N_X_M1035_d N_SLEEP_M1035_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75010.6
+ SB=75004.8 A=0.0975 P=1.6 MULT=1
MM1041 N_X_M1035_d N_SLEEP_M1041_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75011
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1042 N_X_M1042_d N_SLEEP_M1042_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75011.4
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1044 N_X_M1042_d N_SLEEP_M1044_g N_VGND_M1044_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75011.9
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1045 N_X_M1045_d N_SLEEP_M1045_g N_VGND_M1044_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75012.3
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1046 N_X_M1045_d N_SLEEP_M1046_g N_VGND_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75012.7
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1051 N_X_M1051_d N_SLEEP_M1051_g N_VGND_M1046_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75013.1
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1052 N_X_M1051_d N_SLEEP_M1052_g N_VGND_M1052_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75013.5
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1056 N_X_M1056_d N_SLEEP_M1056_g N_VGND_M1052_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75014
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1058 N_X_M1056_d N_SLEEP_M1058_g N_VGND_M1058_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75014.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1063 N_X_M1063_d N_SLEEP_M1063_g N_VGND_M1058_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75014.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1066 N_X_M1063_d N_SLEEP_M1066_g N_VGND_M1066_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75015.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1025 N_A_143_297#_M1025_d N_A_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1036 N_A_143_297#_M1025_d N_A_M1036_g N_VPWR_M1036_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1047 N_A_143_297#_M1047_d N_A_M1047_g N_VPWR_M1036_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1059 N_A_143_297#_M1047_d N_A_M1059_g N_VPWR_M1059_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_143_297#_M1000_g N_A_505_297#_M1000_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75013.2 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1000_d N_A_143_297#_M1001_g N_A_505_297#_M1001_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75012.8 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_143_297#_M1004_g N_A_505_297#_M1001_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75012.4 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1004_d N_A_143_297#_M1005_g N_A_505_297#_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.5 SB=75012 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_143_297#_M1009_g N_A_505_297#_M1005_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75011.5 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1009_d N_A_143_297#_M1011_g N_A_505_297#_M1011_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75011.1 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A_143_297#_M1019_g N_A_505_297#_M1011_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.7 SB=75010.7 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1019_d N_A_143_297#_M1020_g N_A_505_297#_M1020_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.1 SB=75010.3 A=0.15 P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_A_143_297#_M1023_g N_A_505_297#_M1020_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.6 SB=75009.9 A=0.15 P=2.3 MULT=1
MM1031 N_VPWR_M1023_d N_A_143_297#_M1031_g N_A_505_297#_M1031_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75004 SB=75009.4 A=0.15 P=2.3 MULT=1
MM1032 N_VPWR_M1032_d N_A_143_297#_M1032_g N_A_505_297#_M1031_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75004.4 SB=75009 A=0.15 P=2.3 MULT=1
MM1039 N_VPWR_M1032_d N_A_143_297#_M1039_g N_A_505_297#_M1039_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75004.8 SB=75008.6 A=0.15 P=2.3 MULT=1
MM1048 N_VPWR_M1048_d N_A_143_297#_M1048_g N_A_505_297#_M1039_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75005.2 SB=75008.2 A=0.15 P=2.3 MULT=1
MM1053 N_VPWR_M1048_d N_A_143_297#_M1053_g N_A_505_297#_M1053_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75005.7 SB=75007.8 A=0.15 P=2.3 MULT=1
MM1057 N_VPWR_M1057_d N_A_143_297#_M1057_g N_A_505_297#_M1053_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75006.1 SB=75007.3 A=0.15 P=2.3 MULT=1
MM1060 N_VPWR_M1057_d N_A_143_297#_M1060_g N_A_505_297#_M1060_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75006.5 SB=75006.9 A=0.15 P=2.3 MULT=1
MM1006 N_A_505_297#_M1060_s N_SLEEP_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.9
+ SB=75006.5 A=0.15 P=2.3 MULT=1
MM1012 N_A_505_297#_M1012_d N_SLEEP_M1012_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.3
+ SB=75006.1 A=0.15 P=2.3 MULT=1
MM1013 N_A_505_297#_M1012_d N_SLEEP_M1013_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75007.8
+ SB=75005.7 A=0.15 P=2.3 MULT=1
MM1014 N_A_505_297#_M1014_d N_SLEEP_M1014_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.2
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1017 N_A_505_297#_M1014_d N_SLEEP_M1017_g N_X_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75008.6
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1024 N_A_505_297#_M1024_d N_SLEEP_M1024_g N_X_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1026 N_A_505_297#_M1024_d N_SLEEP_M1026_g N_X_M1026_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.4
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1034 N_A_505_297#_M1034_d N_SLEEP_M1034_g N_X_M1026_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75009.9
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1037 N_A_505_297#_M1034_d N_SLEEP_M1037_g N_X_M1037_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75010.3
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1040 N_A_505_297#_M1040_d N_SLEEP_M1040_g N_X_M1037_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75010.7
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1050 N_A_505_297#_M1040_d N_SLEEP_M1050_g N_X_M1050_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75011.1
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1054 N_A_505_297#_M1054_d N_SLEEP_M1054_g N_X_M1050_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75011.5
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1061 N_A_505_297#_M1054_d N_SLEEP_M1061_g N_X_M1061_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75012
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1069 N_A_505_297#_M1069_d N_SLEEP_M1069_g N_X_M1061_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75012.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1070 N_A_505_297#_M1069_d N_SLEEP_M1070_g N_X_M1070_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75012.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1071 N_A_505_297#_M1071_d N_SLEEP_M1071_g N_X_M1070_s VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.135 PD=2.54 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75013.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX72_noxref VNB VPB NWDIODE A=27.1887 P=37.09
*
.include "sky130_fd_sc_hd__lpflow_isobufsrc_16.pxi.spice"
*
.ends
*
*
